
module topcell ( clk, ctr, rst, ai, gi, bi, po );
  input [32:1] ai;
  input [32:1] gi;
  input [32:1] bi;
  output [1:32] po;
  input clk, ctr, rst;
  wire   po1, ctro1, po2, ctro2, po3, ctro3, po4, ctro4, po5, ctro5, po6,
         ctro6, \pe1/bq[1] , \pe1/bq[2] , \pe1/bq[3] , \pe1/bq[4] ,
         \pe1/bq[5] , \pe1/bq[6] , \pe1/bq[7] , \pe1/bq[8] , \pe1/bq[9] ,
         \pe1/bq[10] , \pe1/bq[11] , \pe1/bq[12] , \pe1/bq[13] , \pe1/bq[14] ,
         \pe1/bq[15] , \pe1/bq[16] , \pe1/bq[17] , \pe1/bq[18] , \pe1/bq[19] ,
         \pe1/bq[20] , \pe1/bq[21] , \pe1/bq[22] , \pe1/bq[23] , \pe1/bq[24] ,
         \pe1/bq[25] , \pe1/bq[26] , \pe1/bq[27] , \pe1/bq[28] , \pe1/bq[29] ,
         \pe1/bq[30] , \pe1/bq[31] , \pe1/bq[32] , \pe1/ctrq , \pe2/ti_1 ,
         \pe2/ti_1t , \pe2/bq[1] , \pe2/bq[2] , \pe2/bq[3] , \pe2/bq[4] ,
         \pe2/bq[5] , \pe2/bq[6] , \pe2/bq[7] , \pe2/bq[8] , \pe2/bq[9] ,
         \pe2/bq[10] , \pe2/bq[11] , \pe2/bq[12] , \pe2/bq[13] , \pe2/bq[14] ,
         \pe2/bq[15] , \pe2/bq[16] , \pe2/bq[17] , \pe2/bq[18] , \pe2/bq[19] ,
         \pe2/bq[20] , \pe2/bq[21] , \pe2/bq[22] , \pe2/bq[23] , \pe2/bq[24] ,
         \pe2/bq[25] , \pe2/bq[26] , \pe2/bq[27] , \pe2/bq[28] , \pe2/bq[29] ,
         \pe2/bq[30] , \pe2/bq[31] , \pe2/bq[32] , \pe2/ctrq , \pe2/pq ,
         \pe3/ti_1 , \pe3/ti_1t , \pe3/bq[1] , \pe3/bq[2] , \pe3/bq[3] ,
         \pe3/bq[4] , \pe3/bq[5] , \pe3/bq[6] , \pe3/bq[7] , \pe3/bq[8] ,
         \pe3/bq[9] , \pe3/bq[10] , \pe3/bq[11] , \pe3/bq[12] , \pe3/bq[13] ,
         \pe3/bq[14] , \pe3/bq[15] , \pe3/bq[16] , \pe3/bq[17] , \pe3/bq[18] ,
         \pe3/bq[19] , \pe3/bq[20] , \pe3/bq[21] , \pe3/bq[22] , \pe3/bq[23] ,
         \pe3/bq[24] , \pe3/bq[25] , \pe3/bq[26] , \pe3/bq[27] , \pe3/bq[28] ,
         \pe3/bq[29] , \pe3/bq[30] , \pe3/bq[31] , \pe3/bq[32] , \pe3/bqt[3] ,
         \pe3/ctrq , \pe3/pq , \pe4/ti_1 , \pe4/ti_1t , \pe4/bq[1] ,
         \pe4/bq[2] , \pe4/bq[3] , \pe4/bq[4] , \pe4/bq[5] , \pe4/bq[6] ,
         \pe4/bq[7] , \pe4/bq[8] , \pe4/bq[9] , \pe4/bq[10] , \pe4/bq[11] ,
         \pe4/bq[12] , \pe4/bq[13] , \pe4/bq[14] , \pe4/bq[15] , \pe4/bq[16] ,
         \pe4/bq[17] , \pe4/bq[18] , \pe4/bq[19] , \pe4/bq[20] , \pe4/bq[21] ,
         \pe4/bq[22] , \pe4/bq[23] , \pe4/bq[24] , \pe4/bq[25] , \pe4/bq[26] ,
         \pe4/bq[27] , \pe4/bq[28] , \pe4/bq[29] , \pe4/bq[30] , \pe4/bq[31] ,
         \pe4/bq[32] , \pe4/ctrq , \pe4/pq , \pe5/ti_1 , \pe5/ti_1t ,
         \pe5/bq[1] , \pe5/bq[2] , \pe5/bq[3] , \pe5/bq[4] , \pe5/bq[5] ,
         \pe5/bq[6] , \pe5/bq[7] , \pe5/bq[8] , \pe5/bq[9] , \pe5/bq[10] ,
         \pe5/bq[11] , \pe5/bq[12] , \pe5/bq[13] , \pe5/bq[14] , \pe5/bq[15] ,
         \pe5/bq[16] , \pe5/bq[17] , \pe5/bq[18] , \pe5/bq[19] , \pe5/bq[20] ,
         \pe5/bq[21] , \pe5/bq[22] , \pe5/bq[23] , \pe5/bq[24] , \pe5/bq[25] ,
         \pe5/bq[26] , \pe5/bq[27] , \pe5/bq[28] , \pe5/bq[29] , \pe5/bq[30] ,
         \pe5/bq[31] , \pe5/bq[32] , \pe5/ctrq , \pe5/pq , \pe6/ti_1 ,
         \pe6/ti_1t , \pe6/bq[1] , \pe6/bq[2] , \pe6/bq[3] , \pe6/bq[4] ,
         \pe6/bq[5] , \pe6/bq[6] , \pe6/bq[7] , \pe6/bq[8] , \pe6/bq[9] ,
         \pe6/bq[10] , \pe6/bq[11] , \pe6/bq[12] , \pe6/bq[13] , \pe6/bq[14] ,
         \pe6/bq[15] , \pe6/bq[16] , \pe6/bq[17] , \pe6/bq[18] , \pe6/bq[19] ,
         \pe6/bq[20] , \pe6/bq[21] , \pe6/bq[22] , \pe6/bq[23] , \pe6/bq[24] ,
         \pe6/bq[25] , \pe6/bq[26] , \pe6/bq[27] , \pe6/bq[28] , \pe6/bq[29] ,
         \pe6/bq[30] , \pe6/bq[31] , \pe6/bq[32] , \pe6/ctrq , \pe6/pq ,
         n25137, n25138, n25139, n25140, n25141, n25142, n25143, n25144,
         n25145, n25146, n25147, n25148, n25149, n25150, n25151, n25152,
         n25153, n25154, n25155, n25156, n25157, n25158, n25159, n25160,
         n25161, n25162, n25163, n25164, n25165, n25166, n25167, n25168,
         n25169, n25170, n25171, n25172, n25173, n25174, n25175, n25176,
         n25177, n25178, n25179, n25180, n25181, n25182, n25183, n25184,
         n25185, n25186, n25187, n25188, n25189, n25190, n25191, n25192,
         n25193, n25194, n25195, n25196, n25197, n25198, n25199, n25200,
         n25201, n25202, n25203, n25204, n25205, n25206, n25207, n25208,
         n25209, n25210, n25211, n25212, n25213, n25214, n25215, n25216,
         n25217, n25218, n25219, n25220, n25221, n25222, n25223, n25224,
         n25225, n25226, n25227, n25228, n25229, n25230, n25231, n25232,
         n25233, n25234, n25235, n25236, n25237, n25238, n25239, n25240,
         n25241, n25242, n25243, n25244, n25245, n25246, n25247, n25248,
         n25249, n25250, n25251, n25252, n25253, n25254, n25255, n25256,
         n25257, n25258, n25259, n25260, n25261, n25262, n25263, n25264,
         n25265, n25266, n25267, n25268, n25269, n25270, n25271, n25272,
         n25273, n25274, n25275, n25276, n25277, n25278, n25279, n25280,
         n25281, n25282, n25283, n25284, n25285, n25286, n25287, n25288,
         n25289, n25290, n25291, n25292, n25293, n25294, n25295, n25296,
         n25297, n25298, n25299, n25300, n25301, n25302, n25303, n25304,
         n25305, n25306, n25307, n25308, n25309, n25310, n25311, n25312,
         n25313, n25314, n25315, n25316, n25317, n25318, n25319, n25320,
         n25321, n25322, n25323, n25324, n25325, n25326, n25327, n25328,
         n25329, n25330, n25331, n25332, n25333, n25334, n25335, n25336,
         n25337, n25338, n25339, n25340, n25341, n25342, n25343, n25344,
         n25345, n25346, n25347, n25348, n25349, n25350, n25351, n25352,
         n25353, n25354, n25355, n25356, n25357, n25358, n25359, n25360,
         n25361, n25362, n25363, n25364, n25365, n25366, n25367, n25368,
         n25369, n25370, n25371, n25372, n25373, n25374, n25375, n25376,
         n25377, n25378, n25379, n25380, n25381, n25382, n25383, n25384,
         n25385, n25386, n25387, n25388, n25389, n25390, n25391, n25392,
         n25393, n25394, n25395, n25396, n25397, n25398, n25399, n25400,
         n25401, n25402, n25403, n25404, n25405, n25406, n25407, n25408,
         n25409, n25410, n25411, n25412, n25413, n25414, n25415, n25416,
         n25417, n25418, n25419, n25420, n25421, n25422, n25423, n25424,
         n25425, n25426, n25427, n25428, n25429, n25430, n25431, n25432,
         n25433, n25434, n25435, n25436, n25437, n25438, n25439, n25440,
         n25441, n25442, n25443, n25444, n25445, n25446, n25447, n25448,
         n25449, n25450, n25451, n25452, n25453, n25454, n25455, n25456,
         n25457, n25458, n25459, n25460, n25461, n25462, n25463, n25464,
         n25465, n25466, n25467, n25468, n25469, n25470, n25471, n25472,
         n25473, n25474, n25475, n25476, n25477, n25478, n25479, n25480,
         n25481, n25482, n25483, n25484, n25485, n25486, n25487, n25488,
         n25489, n25490, n25491, n25492, n25493, n25494, n25495, n25496,
         n25497, n25498, n25499, n25500, n25501, n25502, n25503, n25504,
         n25505, n25506, n25507, n25508, n25509, n25510, n25511, n25512,
         n25513, n25514, n25515, n25516, n25517, n25518, n25519, n25520,
         n25521, n25522, n25523, n25524, n25525, n25526, n25527, n25528,
         n25529, n25530, n25531, n25532, n25533, n25534, n25535, n25536,
         n25537, n25538, n25539, n25540, n25541, n25542, n25543, n25544,
         n25545, n25546, n25547, n25548, n25549, n25550, n25551, n25552,
         n25553, n25554, n25555, n25556, n25557, n25558, n25559, n25560,
         n25561, n25562, n25563, n25564, n25565, n25566, n25567, n25568,
         n25569, n25570, n25571, n25572, n25573, n25574, n25575, n25576,
         n25577, n25578, n25579, n25580, n25581, n25582, n25583, n25584,
         n25585, n25586, n25587, n25588, n25589, n25590, n25591, n25592,
         n25593, n25594, n25595, n25596, n25597, n25598, n25599, n25600,
         n25601, n25602, n25603, n25604, n25605, n25606, n25607, n25608,
         n25609, n25610, n25611, n25612, n25613, n25614, n25615, n25616,
         n25617, n25618, n25619, n25620, n25621, n25622, n25623, n25624,
         n25625, n25626, n25627, n25628, n25629, n25630, n25631, n25632,
         n25633, n25634, n25635, n25636, n25637, n25638, n25639, n25640,
         n25641, n25642, n25643, n25644, n25645, n25646, n25647, n25648,
         n25649, n25650, n25651, n25652, n25653, n25654, n25655, n25656,
         n25657, n25658, n25659, n25660, n25661, n25662, n25663, n25664,
         n25665, n25666, n25667, n25668, n25669, n25670, n25671, n25672,
         n25673, n25674, n25675, n25676, n25677, n25678, n25679, n25680,
         n25681, n25682, n25683, n25684, n25685, n25686, n25687, n25688,
         n25689, n25690, n25691, n25692, n25693, n25694, n25695, n25696,
         n25697, n25698, n25699, n25700, n25701, n25702, n25703, n25704,
         n25705, n25706, n25707, n25708, n25709, n25710, n25711, n25712,
         n25713, n25714, n25715, n25716, n25717, n25718, n25719, n25720,
         n25721, n25722, n25723, n25724, n25725, n25726, n25727, n25728,
         n25729, n25730, n25731, n25732, n25733, n25734, n25735, n25736,
         n25737, n25738, n25739, n25740, n25741, n25742, n25743, n25744,
         n25745, n25746, n25747, n25748, n25749, n25750, n25751, n25752,
         n25753, n25754, n25755, n25756, n25757, n25758, n25759, n25760,
         n25761, n25762, n25763, n25764, n25765, n25766, n25767, n25768,
         n25769, n25770, n25771, n25772, n25773, n25774, n25775, n25776,
         n25777, n25778, n25779, n25780, n25781, n25782, n25783, n25784,
         n25785, n25786, n25787, n25788, n25789, n25790, n25791, n25792,
         n25793, n25794, n25795, n25796, n25797, n25798, n25799, n25800,
         n25801, n25802, n25803, n25804, n25805, n25806, n25807, n25808,
         n25809, n25810, n25811, n25812, n25813, n25814, n25815, n25816,
         n25817, n25818, n25819, n25820, n25821, n25822, n25823, n25824,
         n25825, n25826, n25827, n25828, n25829, n25830, n25831, n25832,
         n25833, n25834, n25835, n25836, n25837, n25838, n25839, n25840,
         n25841, n25842, n25843, n25844, n25845, n25846, n25847, n25848,
         n25849, n25850, n25851, n25852, n25853, n25854, n25855, n25856,
         n25857, n25858, n25859, n25860, n25861, n25862, n25863, n25864,
         n25865, n25866, n25867, n25868, n25869, n25870, n25871, n25872,
         n25873, n25874, n25875, n25876, n25877, n25878, n25879, n25880,
         n25881, n25882, n25883, n25884, n25885, n25886, n25887, n25888,
         n25889, n25890, n25891, n25892, n25893, n25894, n25895, n25896,
         n25897, n25898, n25899, n25900, n25901, n25902, n25903, n25904,
         n25905, n25906, n25907, n25908, n25909, n25910, n25911, n25912,
         n25913, n25914, n25915, n25916, n25917, n25918, n25919, n25920,
         n25921, n25922, n25923, n25924, n25925, n25926, n25927, n25928,
         n25929, n25930, n25931, n25932, n25933, n25934, n25935, n25936,
         n25937, n25938, n25939, n25940, n25941, n25942, n25943, n25944,
         n25945, n25946, n25947, n25948, n25949, n25950, n25951, n25952,
         n25953, n25954, n25955, n25956, n25957, n25958, n25959, n25960,
         n25961, n25962, n25963, n25964, n25965, n25966, n25967, n25968,
         n25969, n25970, n25971, n25972, n25973, n25974, n25975, n25976,
         n25977, n25978, n25979, n25980, n25981, n25982, n25983, n25984,
         n25985, n25986, n25987, n25988, n25989, n25990, n25991, n25992,
         n25993, n25994, n25995, n25996, n25997, n25998, n25999, n26000,
         n26001, n26002, n26003, n26004, n26005, n26006, n26007, n26008,
         n26009, n26010, n26011, n26012, n26013, n26014, n26015, n26016,
         n26017, n26018, n26019, n26020, n26021, n26022, n26023, n26024,
         n26025, n26026, n26027, n26028, n26029, n26030, n26031, n26032,
         n26033, n26034, n26035, n26036, n26037, n26038, n26039, n26040,
         n26041, n26042, n26043, n26044, n26045, n26046, n26047, n26048,
         n26049, n26050, n26051, n26052, n26053, n26054, n26055, n26056,
         n26057, n26058, n26059, n26060, n26061, n26062, n26063, n26064,
         n26065, n26066, n26067, n26068, n26069, n26070, n26071, n26072,
         n26073, n26074, n26075, n26076, n26077, n26078, n26079, n26080,
         n26081, n26082, n26083, n26084, n26085, n26086, n26087, n26088,
         n26089, n26090, n26091, n26092, n26093, n26094, n26095, n26096,
         n26097, n26098, n26099, n26100, n26101, n26102, n26103, n26104,
         n26105, n26106, n26107, n26108, n26109, n26110, n26111, n26112,
         n26113, n26114, n26115, n26116, n26117, n26118, n26119, n26120,
         n26121, n26122, n26123, n26124, n26125, n26126, n26127, n26128,
         n26129, n26130, n26131, n26132, n26133, n26134, n26135, n26136,
         n26137, n26138, n26139, n26140, n26141, n26142, n26143, n26144,
         n26145, n26146, n26147, n26148, n26149, n26150, n26151, n26152,
         n26153, n26154, n26155, n26156, n26157, n26158, n26159, n26160,
         n26161, n26162, n26163, n26164, n26165, n26166, n26167, n26168,
         n26169, n26170, n26171, n26172, n26173, n26174, n26175, n26176,
         n26177, n26178, n26179, n26180, n26181, n26182, n26183, n26184,
         n26185, n26186, n26187, n26188, n26189, n26190, n26191, n26192,
         n26193, n26194, n26195, n26196, n26197, n26198, n26199, n26200,
         n26201, n26202, n26203, n26204, n26205, n26206, n26207, n26208,
         n26209, n26210, n26211, n26212, n26213, n26214, n26215, n26216,
         n26217, n26218, n26219, n26220, n26221, n26222, n26223, n26224,
         n26225, n26226, n26227, n26228, n26229, n26230, n26231, n26232,
         n26233, n26234, n26235, n26236, n26237, n26238, n26239, n26240,
         n26241, n26242, n26243, n26244, n26245, n26246, n26247, n26248,
         n26249, n26250, n26251, n26252, n26253, n26254, n26255, n26256,
         n26257, n26258, n26259, n26260, n26261, n26262, n26263, n26264,
         n26265, n26266, n26267, n26268, n26269, n26270, n26271, n26272,
         n26273, n26274, n26275, n26276, n26277, n26278, n26279, n26280,
         n26281, n26282, n26283, n26284, n26285, n26286, n26287, n26288,
         n26289, n26290, n26291, n26292, n26293, n26294, n26295, n26296,
         n26297, n26298, n26299, n26300, n26301, n26302, n26303, n26304,
         n26305, n26306, n26307, n26308, n26309, n26310, n26311, n26312,
         n26313, n26314, n26315, n26316, n26317, n26318, n26319, n26320,
         n26321, n26322, n26323, n26324, n26325, n26326, n26327, n26328,
         n26329, n26330, n26331, n26332, n26333, n26334, n26335, n26336,
         n26337, n26338, n26339, n26340, n26341, n26342, n26343, n26344,
         n26345, n26346, n26347, n26348, n26349, n26350, n26351, n26352,
         n26353, n26354, n26355, n26356, n26357, n26358, n26359, n26360,
         n26361, n26362, n26363, n26364, n26365, n26366, n26367, n26368,
         n26369, n26370, n26371, n26372, n26373, n26374, n26375, n26376,
         n26377, n26378, n26379, n26380, n26381, n26382, n26383, n26384,
         n26385, n26386, n26387, n26388, n26389, n26390, n26391, n26392,
         n26393, n26394, n26395, n26396, n26397, n26398, n26399, n26400,
         n26401, n26402, n26403, n26404, n26405, n26406, n26407, n26408,
         n26409, n26410, n26411, n26412, n26413, n26414, n26415, n26416,
         n26417, n26418, n26419, n26420, n26421, n26422, n26423, n26424,
         n26425, n26426, n26427, n26428, n26429, n26430, n26431, n26432,
         n26433, n26434, n26435, n26436, n26437, n26438, n26439, n26440,
         n26441, n26442, n26443, n26444, n26445, n26446, n26447, n26448,
         n26449, n26450, n26451, n26452, n26453, n26454, n26455, n26456,
         n26457, n26458, n26459, n26460, n26461, n26462, n26463, n26464,
         n26465, n26466, n26467, n26468, n26469, n26470, n26471, n26472,
         n26473, n26474, n26475, n26476, n26477, n26478, n26479, n26480,
         n26481, n26482, n26483, n26484, n26485, n26486, n26487, n26488,
         n26489, n26490, n26491, n26492, n26493, n26494, n26495, n26496,
         n26497, n26498, n26499, n26500, n26501, n26502, n26503, n26504,
         n26505, n26506, n26507, n26508, n26509, n26510, n26511, n26512,
         n26513, n26514, n26515, n26516, n26517, n26518, n26519, n26520,
         n26521, n26522, n26523, n26524, n26525, n26526, n26527, n26528,
         n26529, n26530, n26531, n26532, n26533, n26534, n26535, n26536,
         n26537, n26538, n26539, n26540, n26541, n26542, n26543, n26544,
         n26545, n26546, n26547, n26548, n26549, n26550, n26551, n26552,
         n26553, n26554, n26555, n26556, n26557, n26558, n26559, n26560,
         n26561, n26562, n26563, n26564, n26565, n26566, n26567, n26568,
         n26569, n26570, n26571, n26572, n26573, n26574, n26575, n26576,
         n26577, n26578, n26579, n26580, n26581, n26582, n26583, n26584,
         n26585, n26586, n26587, n26588, n26589, n26590, n26591, n26592,
         n26593, n26594, n26595, n26596, n26597, n26598, n26599, n26600,
         n26601, n26602, n26603, n26604, n26605, n26606, n26607, n26608,
         n26609, n26610, n26611, n26612, n26613, n26614, n26615, n26616,
         n26617, n26618, n26619, n26620, n26621, n26622, n26623, n26624,
         n26625, n26626, n26627, n26628, n26629, n26630, n26631, n26632,
         n26633, n26634, n26635, n26636, n26637, n26638, n26639, n26640,
         n26641, n26642, n26643, n26644, n26645, n26646, n26647, n26648,
         n26649, n26650, n26651, n26652, n26653, n26654, n26655, n26656,
         n26657, n26658, n26659, n26660, n26661, n26662, n26663, n26664,
         n26665, n26666, n26667, n26668, n26669, n26670, n26671, n26672,
         n26673, n26674, n26675, n26676, n26677, n26678, n26679, n26680,
         n26681, n26682, n26683, n26684, n26685, n26686, n26687, n26688,
         n26689, n26690, n26691, n26692, n26693, n26694, n26695, n26696,
         n26697, n26698, n26699, n26700, n26701, n26702, n26703, n26704,
         n26705, n26706, n26707, n26708, n26709, n26710, n26711, n26712,
         n26713, n26714, n26715, n26716, n26717, n26718, n26719, n26720,
         n26721, n26722, n26723, n26724, n26725, n26726, n26727, n26728,
         n26729, n26730, n26731, n26732, n26733, n26734, n26735, n26736,
         n26737, n26738, n26739, n26740, n26741, n26742, n26743, n26744,
         n26745, n26746, n26747, n26748, n26749, n26750, n26751, n26752,
         n26753, n26754, n26755, n26756, n26757, n26758, n26759, n26760,
         n26761, n26762, n26763, n26764, n26765, n26766, n26767, n26768,
         n26769, n26770, n26771, n26772, n26773, n26774, n26775, n26776,
         n26777, n26778, n26779, n26780, n26781, n26782, n26783, n26784,
         n26785, n26786, n26787, n26788, n26789, n26790, n26791, n26792,
         n26793, n26794, n26795, n26796, n26797, n26798, n26799, n26800,
         n26801, n26802, n26803, n26804, n26805, n26806, n26807, n26808,
         n26809, n26810, n26811, n26812, n26813, n26814, n26815, n26816,
         n26817, n26818, n26819, n26820, n26821, n26822, n26823, n26824,
         n26825, n26826, n26827, n26828, n26829, n26830, n26831, n26832,
         n26833, n26834, n26835, n26836, n26837, n26838, n26839, n26840,
         n26841, n26842, n26843, n26844, n26845, n26846, n26847, n26848,
         n26849, n26850, n26851, n26852, n26853, n26854, n26855, n26856,
         n26857, n26858, n26859, n26860, n26861, n26862, n26863, n26864,
         n26865, n26866, n26867, n26868, n26869, n26870, n26871, n26872,
         n26873, n26874, n26875, n26876, n26877, n26878, n26879, n26880,
         n26881, n26882, n26883, n26884, n26885, n26886, n26887, n26888,
         n26889, n26890, n26891, n26892, n26893, n26894, n26895, n26896,
         n26897, n26898, n26899, n26900, n26901, n26902, n26903, n26904,
         n26905, n26906, n26907, n26908, n26909, n26910, n26911, n26912,
         n26913, n26914, n26915, n26916, n26917, n26918, n26919, n26920,
         n26921, n26922, n26923, n26924, n26925, n26926, n26927, n26928,
         n26929, n26930, n26931, n26932, n26933, n26934, n26935, n26936,
         n26937, n26938, n26939, n26940, n26941, n26942, n26943, n26944,
         n26945, n26946, n26947, n26948, n26949, n26950, n26951, n26952,
         n26953, n26954, n26955, n26956, n26957, n26958, n26959, n26960,
         n26961, n26962, n26963, n26964, n26965, n26966, n26967, n26968,
         n26969, n26970, n26971, n26972, n26973, n26974, n26975, n26976,
         n26977, n26978, n26979, n26980, n26981, n26982, n26983, n26984,
         n26985, n26986, n26987, n26988, n26989, n26990, n26991, n26992,
         n26993, n26994, n26995, n26996, n26997, n26998, n26999, n27000,
         n27001, n27002, n27003, n27004, n27005, n27006, n27007, n27008,
         n27009, n27010, n27011, n27012, n27013, n27014, n27015, n27016,
         n27017, n27018, n27019, n27020, n27021, n27022, n27023, n27024,
         n27025, n27026, n27027, n27028, n27029, n27030, n27031, n27032,
         n27033, n27034, n27035, n27036, n27037, n27038, n27039, n27040,
         n27041, n27042, n27043, n27044, n27045, n27046, n27047, n27048,
         n27049, n27050, n27051, n27052, n27053, n27054, n27055, n27056,
         n27057, n27058, n27059, n27060, n27061, n27062, n27063, n27064,
         n27065, n27066, n27067, n27068, n27069, n27070, n27071, n27072,
         n27073, n27074, n27075, n27076, n27077, n27078, n27079, n27080,
         n27081, n27082, n27083, n27084, n27085, n27086, n27087, n27088,
         n27089, n27090, n27091, n27092, n27093, n27094, n27095, n27096,
         n27097, n27098, n27099, n27100, n27101, n27102, n27103, n27104,
         n27105, n27106, n27107, n27108, n27109, n27110, n27111, n27112,
         n27113, n27114, n27115, n27116, n27117, n27118, n27119, n27120,
         n27121, n27122, n27123, n27124, n27125, n27126, n27127, n27128,
         n27129, n27130, n27131, n27132, n27133, n27134, n27135, n27136,
         n27137, n27138, n27139, n27140, n27141, n27142, n27143, n27144,
         n27145, n27146, n27147, n27148, n27149, n27150, n27151, n27152,
         n27153, n27154, n27155, n27156, n27157, n27158, n27159, n27160,
         n27161, n27162, n27163, n27164, n27165, n27166, n27167, n27168,
         n27169, n27170, n27171, n27172, n27173, n27174, n27175, n27176,
         n27177, n27178, n27179, n27180, n27181, n27182, n27183, n27184,
         n27185, n27186, n27187, n27188, n27189, n27190, n27191, n27192,
         n27193, n27194, n27195, n27196, n27197, n27198, n27199, n27200,
         n27201, n27202, n27203, n27204, n27205, n27206, n27207, n27208,
         n27209, n27210, n27211, n27212, n27213, n27214, n27215, n27216,
         n27217, n27218, n27219, n27220, n27221, n27222, n27223, n27224,
         n27225, n27226, n27227, n27228, n27229, n27230, n27231, n27232,
         n27233, n27234, n27235, n27236, n27237, n27238, n27239, n27240,
         n27241, n27242, n27243, n27244, n27245, n27246, n27247, n27248,
         n27249, n27250, n27251, n27252, n27253, n27254, n27255, n27256,
         n27257, n27258, n27259, n27260, n27261, n27262, n27263, n27264,
         n27265, n27266, n27267, n27268, n27269, n27270, n27271, n27272,
         n27273, n27274, n27275, n27276, n27277, n27278, n27279, n27280,
         n27281, n27282, n27283, n27284, n27285, n27286, n27287, n27288,
         n27289, n27290, n27291, n27292, n27293, n27294, n27295, n27296,
         n27297, n27298, n27299, n27300, n27301, n27302, n27303, n27304,
         n27305, n27306, n27307, n27308, n27309, n27310, n27311, n27312,
         n27313, n27314, n27315, n27316, n27317, n27318, n27319, n27320,
         n27321, n27322, n27323, n27324, n27325, n27326, n27327, n27328,
         n27329, n27330, n27331, n27332, n27333, n27334, n27335, n27336,
         n27337, n27338, n27339, n27340, n27341, n27342, n27343, n27344,
         n27345, n27346, n27347, n27348, n27349, n27350, n27351, n27352,
         n27353, n27354, n27355, n27356, n27357, n27358, n27359, n27360,
         n27361, n27362, n27363, n27364, n27365, n27366, n27367, n27368,
         n27369, n27370, n27371, n27372, n27373, n27374, n27375, n27376,
         n27377, n27378, n27379, n27380, n27381, n27382, n27383, n27384,
         n27385, n27386, n27387, n27388, n27389, n27390, n27391, n27392,
         n27393, n27394, n27395, n27396, n27397, n27398, n27399, n27400,
         n27401, n27402, n27403, n27404, n27405, n27406, n27407, n27408,
         n27409, n27410, n27411, n27412, n27413, n27414, n27415, n27416,
         n27417, n27418, n27419, n27420, n27421, n27422, n27423, n27424,
         n27425, n27426, n27427, n27428, n27429, n27430, n27431, n27432,
         n27433, n27434, n27435, n27436, n27437, n27438, n27439, n27440,
         n27441, n27442, n27443, n27444, n27445, n27446, n27447, n27448,
         n27449, n27450, n27451, n27452, n27453, n27454, n27455, n27456,
         n27457, n27458, n27459, n27460, n27461, n27462, n27463, n27464,
         n27465, n27466, n27467, n27468, n27469, n27470, n27471, n27472,
         n27473, n27474, n27475, n27476, n27477, n27478, n27479, n27480,
         n27481, n27482, n27483, n27484, n27485, n27486, n27487, n27488,
         n27489, n27490, n27491, n27492, n27493, n27494, n27495, n27496,
         n27497, n27498, n27499, n27500, n27501, n27502, n27503, n27504,
         n27505, n27506, n27507, n27508, n27509, n27510, n27511, n27512,
         n27513, n27514, n27515, n27516, n27517, n27518, n27519, n27520,
         n27521, n27522, n27523, n27524, n27525, n27526, n27527, n27528,
         n27529, n27530, n27531, n27532, n27533, n27534, n27535, n27536,
         n27537, n27538, n27539, n27540, n27541, n27542, n27543, n27544,
         n27545, n27546, n27547, n27548, n27549, n27550, n27551, n27552,
         n27553, n27554, n27555, n27556, n27557, n27558, n27559, n27560,
         n27561, n27562, n27563, n27564, n27565, n27566, n27567, n27568,
         n27569, n27570, n27571, n27572, n27573, n27574, n27575, n27576,
         n27577, n27578, n27579, n27580, n27581, n27582, n27583, n27584,
         n27585, n27586, n27587, n27588, n27589, n27590, n27591, n27592,
         n27593, n27594, n27595, n27596, n27597, n27598, n27599, n27600,
         n27601, n27602, n27603, n27604, n27605, n27606, n27607, n27608,
         n27609, n27610, n27611, n27612, n27613, n27614, n27615, n27616,
         n27617, n27618, n27619, n27620, n27621, n27622, n27623, n27624,
         n27625, n27626, n27627, n27628, n27629, n27630, n27631, n27632,
         n27633, n27634, n27635, n27636, n27637, n27638, n27639, n27640,
         n27641, n27642, n27643, n27644, n27645, n27646, n27647, n27648,
         n27649, n27650, n27651, n27652, n27653, n27654, n27655, n27656,
         n27657, n27658, n27659, n27660, n27661, n27662, n27663, n27664,
         n27665, n27666, n27667, n27668, n27669, n27670, n27671, n27672,
         n27673, n27674, n27675, n27676, n27677, n27678, n27679, n27680,
         n27681, n27682, n27683, n27684, n27685, n27686, n27687, n27688,
         n27689, n27690, n27691, n27692, n27693, n27694, n27695, n27696,
         n27697, n27698, n27699, n27700, n27701, n27702, n27703, n27704,
         n27705, n27706, n27707, n27708, n27709, n27710, n27711, n27712,
         n27713, n27714, n27715, n27716, n27717, n27718, n27719, n27720,
         n27721, n27722, n27723, n27724, n27725, n27726, n27727, n27728,
         n27729, n27730, n27731, n27732, n27733, n27734, n27735, n27736,
         n27737, n27738, n27739, n27740, n27741, n27742, n27743, n27744,
         n27745, n27746, n27747, n27748, n27749, n27750, n27751, n27752,
         n27753, n27754, n27755, n27756, n27757, n27758, n27759, n27760,
         n27761, n27762, n27763, n27764, n27765, n27766, n27767, n27768,
         n27769, n27770, n27771, n27772, n27773, n27774, n27775, n27776,
         n27777, n27778, n27779, n27780, n27781, n27782, n27783, n27784,
         n27785, n27786, n27787, n27788, n27789, n27790, n27791, n27792,
         n27793, n27794, n27795, n27796, n27797, n27798, n27799, n27800,
         n27801, n27802, n27803, n27804, n27805, n27806, n27807, n27808,
         n27809, n27810, n27811, n27812, n27813, n27814, n27815, n27816,
         n27817, n27818, n27819, n27820, n27821, n27822, n27823, n27824,
         n27825, n27826, n27827, n27828, n27829, n27830, n27831, n27832,
         n27833, n27834, n27835, n27836, n27837, n27838, n27839, n27840,
         n27841, n27842, n27843, n27844, n27845, n27846, n27847, n27848,
         n27849, n27850, n27851, n27852, n27853, n27854, n27855, n27856,
         n27857, n27858, n27859, n27860, n27861, n27862, n27863, n27864,
         n27865, n27866, n27867, n27868, n27869, n27870, n27871, n27872,
         n27873, n27874, n27875, n27876, n27877, n27878, n27879, n27880,
         n27881, n27882, n27883, n27884, n27885, n27886, n27887, n27888,
         n27889, n27890, n27891, n27892, n27893, n27894, n27895, n27896,
         n27897, n27898, n27899, n27900, n27901, n27902, n27903, n27904,
         n27905, n27906, n27907, n27908, n27909, n27910, n27911, n27912,
         n27913, n27914, n27915, n27916, n27917, n27918, n27919, n27920,
         n27921, n27922, n27923, n27924, n27925, n27926, n27927, n27928,
         n27929, n27930, n27931, n27932, n27933, n27934, n27935, n27936,
         n27937, n27938, n27939, n27940, n27941, n27942, n27943, n27944,
         n27945, n27946, n27947, n27948, n27949, n27950, n27951, n27952,
         n27953, n27954, n27955, n27956, n27957, n27958, n27959, n27960,
         n27961, n27962, n27963, n27964, n27965, n27966, n27967, n27968,
         n27969, n27970, n27971, n27972, n27973, n27974, n27975, n27976,
         n27977, n27978, n27979, n27980, n27981, n27982, n27983, n27984,
         n27985, n27986, n27987, n27988, n27989, n27990, n27991, n27992,
         n27993, n27994, n27995, n27996, n27997, n27998, n27999, n28000,
         n28001, n28002, n28003, n28004, n28005, n28006, n28007, n28008,
         n28009, n28010, n28011, n28012, n28013, n28014, n28015, n28016,
         n28017, n28018, n28019, n28020, n28021, n28022, n28023, n28024,
         n28025, n28026, n28027, n28028, n28029, n28030, n28031, n28032,
         n28033, n28034, n28035, n28036, n28037, n28038, n28039, n28040,
         n28041, n28042, n28043, n28044, n28045, n28046, n28047, n28048,
         n28049, n28050, n28051, n28052, n28053, n28054, n28055, n28056,
         n28057, n28058, n28059, n28060, n28061, n28062, n28063, n28064,
         n28065, n28066, n28067, n28068, n28069, n28070, n28071, n28072,
         n28073, n28074, n28075, n28076, n28077, n28078, n28079, n28080,
         n28081, n28082, n28083, n28084, n28085, n28086, n28087, n28088,
         n28089, n28090, n28091, n28092, n28093, n28094, n28095, n28096,
         n28097, n28098, n28099, n28100, n28101, n28102, n28103, n28104,
         n28105, n28106, n28107, n28108, n28109, n28110, n28111, n28112,
         n28113, n28114, n28115, n28116, n28117, n28118, n28119, n28120,
         n28121, n28122, n28123, n28124, n28125, n28126, n28127, n28128,
         n28129, n28130, n28131, n28132, n28133, n28134, n28135, n28136,
         n28137, n28138, n28139, n28140, n28141, n28142, n28143, n28144,
         n28145, n28146, n28147, n28148, n28149, n28150, n28151, n28152,
         n28153, n28154, n28155, n28156, n28157, n28158, n28159, n28160,
         n28161, n28162, n28163, n28164, n28165, n28166, n28167, n28168,
         n28169, n28170, n28171, n28172, n28173, n28174, n28175, n28176,
         n28177, n28178, n28179, n28180, n28181, n28182, n28183, n28184,
         n28185, n28186, n28187, n28188, n28189, n28190, n28191, n28192,
         n28193, n28194, n28195, n28196, n28197, n28198, n28199, n28200,
         n28201, n28202, n28203, n28204, n28205, n28206, n28207, n28208,
         n28209, n28210, n28211, n28212, n28213, n28214, n28215, n28216,
         n28217, n28218, n28219, n28220, n28221, n28222, n28223, n28224,
         n28225, n28226, n28227, n28228, n28229, n28230, n28231, n28232,
         n28233, n28234, n28235, n28236, n28237, n28238, n28239, n28240,
         n28241, n28242, n28243, n28244, n28245, n28246, n28247, n28248,
         n28249, n28250, n28251, n28252, n28253, n28254, n28255, n28256,
         n28257, n28258, n28259, n28260, n28261, n28262, n28263, n28264,
         n28265, n28266, n28267, n28268, n28269, n28270, n28271, n28272,
         n28273, n28274, n28275, n28276, n28277, n28278, n28279, n28280,
         n28281, n28282, n28283, n28284, n28285, n28286, n28287, n28288,
         n28289, n28290, n28291, n28292, n28293, n28294, n28295, n28296,
         n28297, n28298, n28299, n28300, n28301, n28302, n28303, n28304,
         n28305, n28306, n28307, n28308, n28309, n28310, n28311, n28312,
         n28313, n28314, n28315, n28316, n28317, n28318, n28319, n28320,
         n28321, n28322, n28323, n28324, n28325, n28326, n28327, n28328,
         n28329, n28330, n28331, n28332, n28333, n28334, n28335, n28336,
         n28337, n28338, n28339, n28340, n28341, n28342, n28343, n28344,
         n28345, n28346, n28347, n28348, n28349, n28350, n28351, n28352,
         n28353, n28354, n28355, n28356, n28357, n28358, n28359, n28360,
         n28361, n28362, n28363, n28364, n28365, n28366, n28367, n28368,
         n28369, n28370, n28371, n28372, n28373, n28374, n28375, n28376,
         n28377, n28378, n28379, n28380, n28381, n28382, n28383, n28384,
         n28385, n28386, n28387, n28388, n28389, n28390, n28391, n28392,
         n28393, n28394, n28395, n28396, n28397, n28398, n28399, n28400,
         n28401, n28402, n28403, n28404, n28405, n28406, n28407, n28408,
         n28409, n28410, n28411, n28412, n28413, n28414, n28415, n28416,
         n28417, n28418, n28419, n28420, n28421, n28422, n28423, n28424,
         n28425, n28426, n28427, n28428, n28429, n28430, n28431, n28432,
         n28433, n28434, n28435, n28436, n28437, n28438, n28439, n28440,
         n28441, n28442, n28443, n28444, n28445, n28446, n28447, n28448,
         n28449, n28450, n28451, n28452, n28453, n28454, n28455, n28456,
         n28457, n28458, n28459, n28460, n28461, n28462, n28463, n28464,
         n28465, n28466, n28467, n28468, n28469, n28470, n28471, n28472,
         n28473, n28474, n28475, n28476, n28477, n28478, n28479, n28480,
         n28481, n28482, n28483, n28484, n28485, n28486, n28487, n28488,
         n28489, n28490, n28491, n28492, n28493, n28494, n28495, n28496,
         n28497, n28498, n28499, n28500, n28501, n28502, n28503, n28504,
         n28505, n28506, n28507, n28508, n28509, n28510, n28511, n28512,
         n28513, n28514, n28515, n28516, n28517, n28518, n28519, n28520,
         n28521, n28522, n28523, n28524, n28525, n28526, n28527, n28528,
         n28529, n28530, n28531, n28532, n28533, n28534, n28535, n28536,
         n28537, n28538, n28539, n28540, n28541, n28542, n28543, n28544,
         n28545, n28546, n28547, n28548, n28549, n28550, n28551, n28552,
         n28553, n28554, n28555, n28556, n28557, n28558, n28559, n28560,
         n28561, n28562, n28563, n28564, n28565, n28566, n28567, n28568,
         n28569, n28570, n28571, n28572, n28573, n28574, n28575, n28576,
         n28577, n28578, n28579, n28580, n28581, n28582, n28583, n28584,
         n28585, n28586, n28587, n28588, n28589, n28590, n28591, n28592,
         n28593, n28594, n28595, n28596, n28597, n28598, n28599, n28600,
         n28601, n28602, n28603, n28604, n28605, n28606, n28607, n28608,
         n28609, n28610, n28611, n28612, n28613, n28614, n28615, n28616,
         n28617, n28618, n28619, n28620, n28621, n28622, n28623, n28624,
         n28625, n28626, n28627, n28628, n28629, n28630, n28631, n28632,
         n28633, n28634, n28635, n28636, n28637, n28638, n28639, n28640,
         n28641, n28642, n28643, n28644, n28645, n28646, n28647, n28648,
         n28649, n28650, n28651, n28652, n28653, n28654, n28655, n28656,
         n28657, n28658, n28659, n28660, n28661, n28662, n28663, n28664,
         n28665, n28666, n28667, n28668, n28669, n28670, n28671, n28672,
         n28673, n28674, n28675, n28676, n28677, n28678, n28679, n28680,
         n28681, n28682, n28683, n28684, n28685, n28686, n28687, n28688,
         n28689, n28690, n28691, n28692, n28693, n28694, n28695, n28696,
         n28697, n28698, n28699, n28700, n28701, n28702, n28703, n28704,
         n28705, n28706, n28707, n28708, n28709, n28710, n28711, n28712,
         n28713, n28714, n28715, n28716, n28717, n28718, n28719, n28720,
         n28721, n28722, n28723, n28724, n28725, n28726, n28727, n28728,
         n28729, n28730, n28731, n28732, n28733, n28734, n28735, n28736,
         n28737, n28738, n28739, n28740, n28741, n28742, n28743, n28744,
         n28745, n28746, n28747, n28748, n28749, n28750, n28751, n28752,
         n28753, n28754, n28755, n28756, n28757, n28758, n28759, n28760,
         n28761, n28762, n28763, n28764, n28765, n28766, n28767, n28768,
         n28769, n28770, n28771, n28772, n28773, n28774, n28775, n28776,
         n28777, n28778, n28779, n28780, n28781, n28782, n28783, n28784,
         n28785, n28786, n28787, n28788, n28789, n28790, n28791, n28792,
         n28793, n28794, n28795, n28796, n28797, n28798, n28799, n28800,
         n28801, n28802, n28803, n28804, n28805, n28806, n28807, n28808,
         n28809, n28810, n28811, n28812, n28813, n28814, n28815, n28816,
         n28817, n28818, n28819, n28820, n28821, n28822, n28823, n28824,
         n28825, n28826, n28827, n28828, n28829, n28830, n28831, n28832,
         n28833, n28834, n28835, n28836, n28837, n28838, n28839, n28840,
         n28841, n28842, n28843, n28844, n28845, n28846, n28847, n28848,
         n28849, n28850, n28851, n28852, n28853, n28854, n28855, n28856,
         n28857, n28858, n28859, n28860, n28861, n28862, n28863, n28864,
         n28865, n28866, n28867, n28868, n28869, n28870, n28871, n28872,
         n28873, n28874, n28875, n28876, n28877, n28878, n28879, n28880,
         n28881, n28882, n28883, n28884, n28885, n28886, n28887, n28888,
         n28889, n28890, n28891, n28892, n28893, n28894, n28895, n28896,
         n28897, n28898, n28899, n28900, n28901, n28902, n28903, n28904,
         n28905, n28906, n28907, n28908, n28909, n28910, n28911, n28912,
         n28913, n28914, n28915, n28916, n28917, n28918, n28919, n28920,
         n28921, n28922, n28923, n28924, n28925, n28926, n28927, n28928,
         n28929, n28930, n28931, n28932, n28933, n28934, n28935, n28936,
         n28937, n28938, n28939, n28940, n28941, n28942, n28943, n28944,
         n28945, n28946, n28947, n28948, n28949, n28950, n28951, n28952,
         n28953, n28954, n28955, n28956, n28957, n28958, n28959, n28960,
         n28961, n28962, n28963, n28964, n28965, n28966, n28967, n28968,
         n28969, n28970, n28971, n28972, n28973, n28974, n28975, n28976,
         n28977, n28978, n28979, n28980, n28981, n28982, n28983, n28984,
         n28985, n28986, n28987, n28988, n28989, n28990, n28991, n28992,
         n28993, n28994, n28995, n28996, n28997, n28998, n28999, n29000,
         n29001, n29002, n29003, n29004, n29005, n29006, n29007, n29008,
         n29009, n29010, n29011, n29012, n29013, n29014, n29015, n29016,
         n29017, n29018, n29019, n29020, n29021, n29022, n29023, n29024,
         n29025, n29026, n29027, n29028, n29029, n29030, n29031, n29032,
         n29033, n29034, n29035, n29036, n29037, n29038, n29039, n29040,
         n29041, n29042, n29043, n29044, n29045, n29046, n29047, n29048,
         n29049, n29050, n29051, n29052, n29053, n29054, n29055, n29056,
         n29057, n29058, n29059, n29060, n29061, n29062, n29063, n29064,
         n29065, n29066, n29067, n29068, n29069, n29070, n29071, n29072,
         n29073, n29074, n29075, n29076, n29077, n29078, n29079, n29080,
         n29081, n29082, n29083, n29084, n29085, n29086, n29087, n29088,
         n29089, n29090, n29091, n29092, n29093, n29094, n29095, n29096,
         n29097, n29098, n29099, n29100, n29101, n29102, n29103, n29104,
         n29105, n29106, n29107, n29108, n29109, n29110, n29111, n29112,
         n29113, n29114, n29115, n29116, n29117, n29118, n29119, n29120,
         n29121, n29122, n29123, n29124, n29125, n29126, n29127, n29128,
         n29129, n29130, n29131, n29132, n29133, n29134, n29135, n29136,
         n29137, n29138, n29139, n29140, n29141, n29142, n29143, n29144,
         n29145, n29146, n29147, n29148, n29149, n29150, n29151, n29152,
         n29153, n29154, n29155, n29156, n29157, n29158, n29159, n29160,
         n29161, n29162, n29163, n29164, n29165, n29166, n29167, n29168,
         n29169, n29170, n29171, n29172, n29173, n29174, n29175, n29176,
         n29177, n29178, n29179, n29180, n29181, n29182, n29183, n29184,
         n29185, n29186, n29187, n29188, n29189, n29190, n29191, n29192,
         n29193, n29194, n29195, n29196, n29197, n29198, n29199, n29200,
         n29201, n29202, n29203, n29204, n29205, n29206, n29207, n29208,
         n29209, n29210, n29211, n29212, n29213, n29214, n29215, n29216,
         n29217, n29218, n29219, n29220, n29221, n29222, n29223, n29224,
         n29225, n29226, n29227, n29228, n29229, n29230, n29231, n29232,
         n29233, n29234, n29235, n29236, n29237, n29238, n29239, n29240,
         n29241, n29242, n29243, n29244, n29245, n29246, n29247, n29248,
         n29249, n29250, n29251, n29252, n29253, n29254, n29255, n29256,
         n29257, n29258, n29259, n29260, n29261, n29262, n29263, n29264,
         n29265, n29266, n29267, n29268, n29269, n29270, n29271, n29272,
         n29273, n29274, n29275, n29276, n29277, n29278, n29279, n29280,
         n29281, n29282, n29283, n29284, n29285, n29286, n29287, n29288,
         n29289, n29290, n29291, n29292, n29293, n29294, n29295, n29296,
         n29297, n29298, n29299, n29300, n29301, n29302, n29303, n29304,
         n29305, n29306, n29307, n29308, n29309, n29310, n29311, n29312,
         n29313, n29314, n29315, n29316, n29317, n29318, n29319, n29320,
         n29321, n29322, n29323, n29324, n29325, n29326, n29327, n29328,
         n29329, n29330, n29331, n29332, n29333, n29334, n29335, n29336,
         n29337, n29338, n29339, n29340, n29341, n29342, n29343, n29344,
         n29345, n29346, n29347, n29348, n29349, n29350, n29351, n29352,
         n29353, n29354, n29355, n29356, n29357, n29358, n29359, n29360,
         n29361, n29362, n29363, n29364, n29365, n29366, n29367, n29368,
         n29369, n29370, n29371, n29372, n29373, n29374, n29375, n29376,
         n29377, n29378, n29379, n29380, n29381, n29382, n29383, n29384,
         n29385, n29386, n29387, n29388, n29389, n29390, n29391, n29392,
         n29393, n29394, n29395, n29396, n29397, n29398, n29399, n29400,
         n29401, n29402, n29403, n29404, n29405, n29406, n29407, n29408,
         n29409, n29410, n29411, n29412, n29413, n29414, n29415, n29416,
         n29417, n29418, n29419, n29420, n29421, n29422, n29423, n29424,
         n29425, n29426, n29427, n29428, n29429, n29430, n29431, n29432,
         n29433, n29434, n29435, n29436, n29437, n29438, n29439, n29440,
         n29441, n29442, n29443, n29444, n29445, n29446, n29447, n29448,
         n29449, n29450, n29451, n29452, n29453, n29454, n29455, n29456,
         n29457, n29458, n29459, n29460, n29461, n29462, n29463, n29464,
         n29465, n29466, n29467, n29468, n29469, n29470, n29471, n29472,
         n29473, n29474, n29475, n29476, n29477, n29478, n29479, n29480,
         n29481, n29482, n29483, n29484, n29485, n29486, n29487, n29488,
         n29489, n29490, n29491, n29492, n29493, n29494, n29495, n29496,
         n29497, n29498, n29499, n29500, n29501, n29502, n29503, n29504,
         n29505, n29506, n29507, n29508, n29509, n29510, n29511, n29512,
         n29513, n29514, n29515, n29516, n29517, n29518, n29519, n29520,
         n29521, n29522, n29523, n29524, n29525, n29526, n29527, n29528,
         n29529, n29530, n29531, n29532, n29533, n29534, n29535, n29536,
         n29537, n29538, n29539, n29540, n29541, n29542, n29543, n29544,
         n29545, n29546, n29547, n29548, n29549, n29550, n29551, n29552,
         n29553, n29554, n29555, n29556, n29557, n29558, n29559, n29560,
         n29561, n29562, n29563, n29564, n29565, n29566, n29567, n29568,
         n29569, n29570, n29571, n29572, n29573, n29574, n29575, n29576,
         n29577, n29578, n29579, n29580, n29581, n29582, n29583, n29584,
         n29585, n29586, n29587, n29588, n29589, n29590, n29591, n29592,
         n29593, n29594, n29595, n29596, n29597, n29598, n29599, n29600,
         n29601, n29602, n29603, n29604, n29605, n29606, n29607, n29608,
         n29609, n29610, n29611, n29612, n29613, n29614, n29615, n29616,
         n29617, n29618, n29619, n29620, n29621, n29622, n29623, n29624,
         n29625, n29626, n29627, n29628, n29629, n29630, n29631, n29632,
         n29633, n29634, n29635, n29636, n29637, n29638, n29639, n29640,
         n29641, n29642, n29643, n29644, n29645, n29646, n29647, n29648,
         n29649, n29650, n29651, n29652, n29653, n29654, n29655, n29656,
         n29657, n29658, n29659, n29660, n29661, n29662, n29663, n29664,
         n29665, n29666, n29667, n29668, n29669, n29670, n29671, n29672,
         n29673, n29674, n29675, n29676, n29677, n29678, n29679, n29680,
         n29681, n29682, n29683, n29684, n29685, n29686, n29687, n29688,
         n29689, n29690, n29691, n29692, n29693, n29694, n29695, n29696,
         n29697, n29698, n29699, n29700, n29701, n29702, n29703, n29704,
         n29705, n29706, n29707, n29708, n29709, n29710, n29711, n29712,
         n29713, n29714, n29715, n29716, n29717, n29718, n29719, n29720,
         n29721, n29722, n29723, n29724, n29725, n29726, n29727, n29728,
         n29729, n29730, n29731, n29732, n29733, n29734, n29735, n29736,
         n29737, n29738, n29739, n29740, n29741, n29742, n29743, n29744,
         n29745, n29746, n29747, n29748, n29749, n29750, n29751, n29752,
         n29753, n29754, n29755, n29756, n29757, n29758, n29759, n29760,
         n29761, n29762, n29763, n29764, n29765, n29766, n29767, n29768,
         n29769, n29770, n29771, n29772, n29773, n29774, n29775, n29776,
         n29777, n29778, n29779, n29780, n29781, n29782, n29783, n29784,
         n29785, n29786, n29787, n29788, n29789, n29790, n29791, n29792,
         n29793, n29794, n29795, n29796, n29797, n29798, n29799, n29800,
         n29801, n29802, n29803, n29804, n29805, n29806, n29807, n29808,
         n29809, n29810, n29811, n29812, n29813, n29814, n29815, n29816,
         n29817, n29818, n29819, n29820, n29821, n29822, n29823, n29824,
         n29825, n29826, n29827, n29828, n29829, n29830, n29831, n29832,
         n29833, n29834, n29835, n29836, n29837, n29838, n29839, n29840,
         n29841, n29842, n29843, n29844, n29845, n29846, n29847, n29848,
         n29849, n29850, n29851, n29852, n29853, n29854, n29855, n29856,
         n29857, n29858, n29859, n29860, n29861, n29862, n29863, n29864,
         n29865, n29866, n29867, n29868, n29869, n29870, n29871, n29872,
         n29873, n29874, n29875, n29876, n29877, n29878, n29879, n29880,
         n29881, n29882, n29883, n29884, n29885, n29886, n29887, n29888,
         n29889, n29890, n29891, n29892, n29893, n29894, n29895, n29896,
         n29897, n29898, n29899, n29900, n29901, n29902, n29903, n29904,
         n29905, n29906, n29907, n29908, n29909, n29910, n29911, n29912,
         n29913, n29914, n29915, n29916, n29917, n29918, n29919, n29920,
         n29921, n29922, n29923, n29924, n29925, n29926, n29927, n29928,
         n29929, n29930, n29931, n29932, n29933, n29934, n29935, n29936,
         n29937, n29938, n29939, n29940, n29941, n29942, n29943, n29944,
         n29945, n29946, n29947, n29948, n29949, n29950, n29951, n29952,
         n29953, n29954, n29955, n29956, n29957, n29958, n29959, n29960,
         n29961, n29962, n29963, n29964, n29965, n29966, n29967, n29968,
         n29969, n29970, n29971, n29972, n29973, n29974, n29975, n29976,
         n29977, n29978, n29979, n29980, n29981, n29982, n29983, n29984,
         n29985, n29986, n29987, n29988, n29989, n29990, n29991, n29992,
         n29993, n29994, n29995, n29996, n29997, n29998, n29999, n30000,
         n30001, n30002, n30003, n30004, n30005, n30006, n30007, n30008,
         n30009, n30010, n30011, n30012, n30013, n30014, n30015, n30016,
         n30017, n30018, n30019, n30020, n30021, n30022, n30023, n30024,
         n30025, n30026, n30027, n30028, n30029, n30030, n30031, n30032,
         n30033, n30034, n30035, n30036, n30037, n30038, n30039, n30040,
         n30041, n30042, n30043, n30044, n30045, n30046, n30047, n30048,
         n30049, n30050, n30051, n30052, n30053, n30054, n30055, n30056,
         n30057, n30058, n30059, n30060, n30061, n30062, n30063, n30064,
         n30065, n30066, n30067, n30068, n30069, n30070, n30071, n30072,
         n30073, n30074, n30075, n30076, n30077, n30078, n30079, n30080,
         n30081, n30082, n30083, n30084, n30085, n30086, n30087, n30088,
         n30089, n30090, n30091, n30092, n30093, n30094, n30095, n30096,
         n30097, n30098, n30099, n30100, n30101, n30102, n30103, n30104,
         n30105, n30106, n30107, n30108, n30109, n30110, n30111, n30112,
         n30113, n30114, n30115, n30116, n30117, n30118, n30119, n30120,
         n30121, n30122, n30123, n30124, n30125, n30126, n30127, n30128,
         n30129, n30130, n30131, n30132, n30133, n30134, n30135, n30136,
         n30137, n30138, n30139, n30140, n30141, n30142, n30143, n30144,
         n30145, n30146, n30147, n30148, n30149, n30150, n30151, n30152,
         n30153, n30154, n30155, n30156, n30157, n30158, n30159, n30160,
         n30161, n30162, n30163, n30164, n30165, n30166, n30167, n30168,
         n30169, n30170, n30171, n30172, n30173, n30174, n30175, n30176,
         n30177, n30178, n30179, n30180, n30181, n30182, n30183, n30184,
         n30185, n30186, n30187, n30188, n30189, n30190, n30191, n30192,
         n30193, n30194, n30195, n30196, n30197, n30198, n30199, n30200,
         n30201, n30202, n30203, n30204, n30205, n30206, n30207, n30208,
         n30209, n30210, n30211, n30212, n30213, n30214, n30215, n30216,
         n30217, n30218, n30219, n30220, n30221, n30222, n30223, n30224,
         n30225, n30226, n30227, n30228, n30229, n30230, n30231, n30232,
         n30233, n30234, n30235, n30236, n30237, n30238, n30239, n30240,
         n30241, n30242, n30243, n30244, n30245, n30246, n30247, n30248,
         n30249, n30250, n30251, n30252, n30253, n30254, n30255, n30256,
         n30257, n30258, n30259, n30260, n30261, n30262, n30263, n30264,
         n30265, n30266, n30267, n30268, n30269, n30270, n30271, n30272,
         n30273, n30274, n30275, n30276, n30277, n30278, n30279, n30280,
         n30281, n30282, n30283, n30284, n30285, n30286, n30287, n30288,
         n30289, n30290, n30291, n30292, n30293, n30294, n30295, n30296,
         n30297, n30298, n30299, n30300, n30301, n30302, n30303, n30304,
         n30305, n30306, n30307, n30308, n30309, n30310, n30311, n30312,
         n30313, n30314, n30315, n30316, n30317, n30318, n30319, n30320,
         n30321, n30322, n30323, n30324, n30325, n30326, n30327, n30328,
         n30329, n30330, n30331, n30332, n30333, n30334, n30335, n30336,
         n30337, n30338, n30339, n30340, n30341, n30342, n30343, n30344,
         n30345, n30346, n30347, n30348, n30349, n30350, n30351, n30352,
         n30353, n30354, n30355, n30356, n30357, n30358, n30359, n30360,
         n30361, n30362, n30363, n30364, n30365, n30366, n30367, n30368,
         n30369, n30370, n30371, n30372, n30373, n30374, n30375, n30376,
         n30377, n30378, n30379, n30380, n30381, n30382, n30383, n30384,
         n30385, n30386, n30387, n30388, n30389, n30390, n30391, n30392,
         n30393, n30394, n30395, n30396, n30397, n30398, n30399, n30400,
         n30401, n30402, n30403, n30404, n30405, n30406, n30407, n30408,
         n30409, n30410, n30411, n30412, n30413, n30414, n30415, n30416,
         n30417, n30418, n30419, n30420, n30421, n30422, n30423, n30424,
         n30425, n30426, n30427, n30428, n30429, n30430, n30431, n30432,
         n30433, n30434, n30435, n30436, n30437, n30438, n30439, n30440,
         n30441, n30442, n30443, n30444, n30445, n30446, n30447, n30448,
         n30449, n30450, n30451, n30452, n30453, n30454, n30455, n30456,
         n30457, n30458, n30459, n30460, n30461, n30462, n30463, n30464,
         n30465, n30466, n30467, n30468, n30469, n30470, n30471, n30472,
         n30473, n30474, n30475, n30476, n30477, n30478, n30479, n30480,
         n30481, n30482, n30483, n30484, n30485, n30486, n30487, n30488,
         n30489, n30490, n30491, n30492, n30493, n30494, n30495, n30496,
         n30497, n30498, n30499, n30500, n30501, n30502, n30503, n30504,
         n30505, n30506, n30507, n30508, n30509, n30510, n30511, n30512,
         n30513, n30514, n30515, n30516, n30517, n30518, n30519, n30520,
         n30521, n30522, n30523, n30524, n30525, n30526, n30527, n30528,
         n30529, n30530, n30531, n30532, n30533, n30534, n30535, n30536,
         n30537, n30538, n30539, n30540, n30541, n30542, n30543, n30544,
         n30545, n30546, n30547, n30548, n30549, n30550, n30551, n30552,
         n30553, n30554, n30555, n30556, n30557, n30558, n30559, n30560,
         n30561, n30562, n30563, n30564, n30565, n30566, n30567, n30568,
         n30569, n30570, n30571, n30572, n30573, n30574, n30575, n30576,
         n30577, n30578, n30579, n30580, n30581, n30582, n30583, n30584,
         n30585, n30586, n30587, n30588, n30589, n30590, n30591, n30592,
         n30593, n30594, n30595, n30596, n30597, n30598, n30599, n30600,
         n30601, n30602, n30603, n30604, n30605, n30606, n30607, n30608,
         n30609, n30610, n30611, n30612, n30613, n30614, n30615, n30616,
         n30617, n30618, n30619, n30620, n30621, n30622, n30623, n30624,
         n30625, n30626, n30627, n30628, n30629, n30630, n30631, n30632,
         n30633, n30634, n30635, n30636, n30637, n30638, n30639, n30640,
         n30641, n30642, n30643, n30644, n30645, n30646, n30647, n30648,
         n30649, n30650, n30651, n30652, n30653, n30654, n30655, n30656,
         n30657, n30658, n30659, n30660, n30661, n30662, n30663, n30664,
         n30665, n30666, n30667, n30668, n30669, n30670, n30671, n30672,
         n30673, n30674, n30675, n30676, n30677, n30678, n30679, n30680,
         n30681, n30682, n30683, n30684, n30685, n30686, n30687, n30688,
         n30689, n30690, n30691, n30692, n30693, n30694, n30695, n30696,
         n30697, n30698, n30699, n30700, n30701, n30702, n30703, n30704,
         n30705, n30706, n30707, n30708, n30709, n30710, n30711, n30712,
         n30713, n30714, n30715, n30716, n30717, n30718, n30719, n30720,
         n30721, n30722, n30723, n30724, n30725, n30726, n30727, n30728,
         n30729, n30730, n30731, n30732, n30733, n30734, n30735, n30736,
         n30737, n30738, n30739, n30740, n30741, n30742, n30743, n30744,
         n30745, n30746, n30747, n30748, n30749, n30750, n30751, n30752,
         n30753, n30754, n30755, n30756, n30757, n30758, n30759, n30760,
         n30761, n30762, n30763, n30764, n30765, n30766, n30767, n30768,
         n30769, n30770, n30771, n30772, n30773, n30774, n30775, n30776,
         n30777, n30778, n30779, n30780, n30781, n30782, n30783, n30784,
         n30785, n30786, n30787, n30788, n30789, n30790, n30791, n30792,
         n30793, n30794, n30795, n30796, n30797, n30798, n30799, n30800,
         n30801, n30802, n30803, n30804, n30805, n30806, n30807, n30808,
         n30809, n30810, n30811, n30812, n30813, n30814, n30815, n30816,
         n30817, n30818, n30819, n30820, n30821, n30822, n30823, n30824,
         n30825, n30826, n30827, n30828, n30829, n30830, n30831, n30832,
         n30833, n30834, n30835, n30836, n30837, n30838, n30839, n30840,
         n30841, n30842, n30843, n30844, n30845, n30846, n30847, n30848,
         n30849, n30850, n30851, n30852, n30853, n30854, n30855, n30856,
         n30857, n30858, n30859, n30860, n30861, n30862, n30863, n30864,
         n30865, n30866, n30867, n30868, n30869, n30870, n30871, n30872,
         n30873, n30874, n30875, n30876, n30877, n30878, n30879, n30880,
         n30881, n30882, n30883, n30884, n30885, n30886, n30887, n30888,
         n30889, n30890, n30891, n30892, n30893, n30894, n30895, n30896,
         n30897, n30898, n30899, n30900, n30901, n30902, n30903, n30904,
         n30905, n30906, n30907, n30908, n30909, n30910, n30911, n30912,
         n30913, n30914, n30915, n30916, n30917, n30918, n30919, n30920,
         n30921, n30922, n30923, n30924, n30925, n30926, n30927, n30928,
         n30929, n30930, n30931, n30932, n30933, n30934, n30935, n30936,
         n30937, n30938, n30939, n30940, n30941, n30942, n30943, n30944,
         n30945, n30946, n30947, n30948, n30949, n30950, n30951, n30952,
         n30953, n30954, n30955, n30956, n30957, n30958, n30959, n30960,
         n30961, n30962, n30963, n30964, n30965, n30966, n30967, n30968,
         n30969, n30970, n30971, n30972, n30973, n30974, n30975, n30976,
         n30977, n30978, n30979, n30980, n30981, n30982, n30983, n30984,
         n30985, n30986, n30987, n30988, n30989, n30990, n30991, n30992,
         n30993, n30994, n30995, n30996, n30997, n30998, n30999, n31000,
         n31001, n31002, n31003, n31004, n31005, n31006, n31007, n31008,
         n31009, n31010, n31011, n31012, n31013, n31014, n31015, n31016,
         n31017, n31018, n31019, n31020, n31021, n31022, n31023, n31024,
         n31025, n31026, n31027, n31028, n31029, n31030, n31031, n31032,
         n31033, n31034, n31035, n31036, n31037, n31038, n31039, n31040,
         n31041, n31042, n31043, n31044, n31045, n31046, n31047, n31048,
         n31049, n31050, n31051, n31052, n31053, n31054, n31055, n31056,
         n31057, n31058, n31059, n31060, n31061, n31062, n31063, n31064,
         n31065, n31066, n31067, n31068, n31069, n31070, n31071, n31072,
         n31073, n31074, n31075, n31076, n31077, n31078, n31079, n31080,
         n31081, n31082, n31083, n31084, n31085, n31086, n31087, n31088,
         n31089, n31090, n31091, n31092, n31093, n31094, n31095, n31096,
         n31097, n31098, n31099, n31100, n31101, n31102, n31103, n31104,
         n31105, n31106, n31107, n31108, n31109, n31110, n31111, n31112,
         n31113, n31114, n31115, n31116, n31117, n31118, n31119, n31120,
         n31121, n31122, n31123, n31124, n31125, n31126, n31127, n31128,
         n31129, n31130, n31131, n31132, n31133, n31134, n31135, n31136,
         n31137, n31138, n31139, n31140, n31141, n31142, n31143, n31144,
         n31145, n31146, n31147, n31148, n31149, n31150, n31151, n31152,
         n31153, n31154, n31155, n31156, n31157, n31158, n31159, n31160,
         n31161, n31162, n31163, n31164, n31165, n31166, n31167, n31168,
         n31169, n31170, n31171, n31172, n31173, n31174, n31175, n31176,
         n31177, n31178, n31179, n31180, n31181, n31182, n31183, n31184,
         n31185, n31186, n31187, n31188, n31189, n31190, n31191, n31192,
         n31193, n31194, n31195, n31196, n31197, n31198, n31199, n31200,
         n31201, n31202, n31203, n31204, n31205, n31206, n31207, n31208,
         n31209, n31210, n31211, n31212, n31213, n31214, n31215, n31216,
         n31217, n31218, n31219, n31220, n31221, n31222, n31223, n31224,
         n31225, n31226, n31227, n31228, n31229, n31230, n31231, n31232,
         n31233, n31234, n31235, n31236, n31237, n31238, n31239, n31240,
         n31241, n31242, n31243, n31244, n31245, n31246, n31247, n31248,
         n31249, n31250, n31251, n31252, n31253, n31254, n31255, n31256,
         n31257, n31258, n31259, n31260, n31261, n31262, n31263, n31264,
         n31265, n31266, n31267, n31268, n31269, n31270, n31271, n31272,
         n31273, n31274, n31275, n31276, n31277, n31278, n31279, n31280,
         n31281, n31282, n31283, n31284, n31285, n31286, n31287, n31288,
         n31289, n31290, n31291, n31292, n31293, n31294, n31295, n31296,
         n31297, n31298, n31299, n31300, n31301, n31302, n31303, n31304,
         n31305, n31306, n31307, n31308, n31309, n31310, n31311, n31312,
         n31313, n31314, n31315, n31316, n31317, n31318, n31319, n31320,
         n31321, n31322, n31323, n31324, n31325, n31326, n31327, n31328,
         n31329, n31330, n31331, n31332, n31333, n31334, n31335, n31336,
         n31337, n31338, n31339, n31340, n31341, n31342, n31343, n31344,
         n31345, n31346, n31347, n31348, n31349, n31350, n31351, n31352,
         n31353, n31354, n31355, n31356, n31357, n31358, n31359, n31360,
         n31361, n31362, n31363, n31364, n31365, n31366, n31367, n31368,
         n31369, n31370, n31371, n31372, n31373, n31374, n31375, n31376,
         n31377, n31378, n31379, n31380, n31381, n31382, n31383, n31384,
         n31385, n31386, n31387, n31388, n31389, n31390, n31391, n31392,
         n31393, n31394, n31395, n31396, n31397, n31398, n31399, n31400,
         n31401, n31402, n31403, n31404, n31405, n31406, n31407, n31408,
         n31409, n31410, n31411, n31412, n31413, n31414, n31415, n31416,
         n31417, n31418, n31419, n31420, n31421, n31422, n31423, n31424,
         n31425, n31426, n31427, n31428, n31429, n31430, n31431, n31432,
         n31433, n31434, n31435, n31436, n31437, n31438, n31439, n31440,
         n31441, n31442, n31443, n31444, n31445, n31446, n31447, n31448,
         n31449, n31450, n31451, n31452, n31453, n31454, n31455, n31456,
         n31457, n31458, n31459, n31460, n31461, n31462, n31463, n31464,
         n31465, n31466, n31467, n31468, n31469, n31470, n31471, n31472,
         n31473, n31474, n31475, n31476, n31477, n31478, n31479, n31480,
         n31481, n31482, n31483, n31484, n31485, n31486, n31487, n31488,
         n31489, n31490, n31491, n31492, n31493, n31494, n31495, n31496,
         n31497, n31498, n31499, n31500, n31501, n31502, n31503, n31504,
         n31505, n31506, n31507, n31508, n31509, n31510, n31511, n31512,
         n31513, n31514, n31515, n31516, n31517, n31518, n31519, n31520,
         n31521, n31522, n31523, n31524, n31525, n31526, n31527, n31528,
         n31529, n31530, n31531, n31532, n31533, n31534, n31535, n31536,
         n31537, n31538, n31539, n31540, n31541, n31542, n31543, n31544,
         n31545, n31546, n31547, n31548, n31549, n31550, n31551, n31552,
         n31553, n31554, n31555, n31556, n31557, n31558, n31559, n31560,
         n31561, n31562, n31563, n31564, n31565, n31566, n31567, n31568,
         n31569, n31570, n31571, n31572, n31573, n31574, n31575, n31576,
         n31577, n31578, n31579, n31580, n31581, n31582, n31583, n31584,
         n31585, n31586, n31587, n31588, n31589, n31590, n31591, n31592,
         n31593, n31594, n31595, n31596, n31597, n31598, n31599, n31600,
         n31601, n31602, n31603, n31604, n31605, n31606, n31607, n31608,
         n31609, n31610, n31611, n31612, n31613, n31614, n31615, n31616,
         n31617, n31618, n31619, n31620, n31621, n31622, n31623, n31624,
         n31625, n31626, n31627, n31628, n31629, n31630, n31631, n31632,
         n31633, n31634, n31635, n31636, n31637, n31638, n31639, n31640,
         n31641, n31642, n31643, n31644, n31645, n31646, n31647, n31648,
         n31649, n31650, n31651, n31652, n31653, n31654, n31655, n31656,
         n31657, n31658, n31659, n31660, n31661, n31662, n31663, n31664,
         n31665, n31666, n31667, n31668, n31669, n31670, n31671, n31672,
         n31673, n31674, n31675, n31676, n31677, n31678, n31679, n31680,
         n31681, n31682, n31683, n31684, n31685, n31686, n31687, n31688,
         n31689, n31690, n31691, n31692, n31693, n31694, n31695, n31696,
         n31697, n31698, n31699, n31700, n31701, n31702, n31703, n31704,
         n31705, n31706, n31707, n31708, n31709, n31710, n31711, n31712,
         n31713, n31714, n31715, n31716, n31717, n31718, n31719, n31720,
         n31721, n31722, n31723, n31724, n31725, n31726, n31727, n31728,
         n31729, n31730, n31731, n31732, n31733, n31734, n31735, n31736,
         n31737, n31738, n31739, n31740, n31741, n31742, n31743, n31744,
         n31745, n31746, n31747, n31748, n31749, n31750, n31751, n31752,
         n31753, n31754, n31755, n31756, n31757, n31758, n31759, n31760,
         n31761, n31762, n31763, n31764, n31765, n31766, n31767, n31768,
         n31769, n31770, n31771, n31772, n31773, n31774, n31775, n31776,
         n31777, n31778, n31779, n31780, n31781, n31782, n31783, n31784,
         n31785, n31786, n31787, n31788, n31789, n31790, n31791, n31792,
         n31793, n31794, n31795, n31796, n31797, n31798, n31799, n31800,
         n31801, n31802, n31803, n31804, n31805, n31806, n31807, n31808,
         n31809, n31810, n31811, n31812, n31813, n31814, n31815, n31816,
         n31817, n31818, n31819, n31820, n31821, n31822, n31823, n31824,
         n31825, n31826, n31827, n31828, n31829, n31830, n31831, n31832,
         n31833, n31834, n31835, n31836, n31837, n31838, n31839, n31840,
         n31841, n31842, n31843, n31844, n31845, n31846, n31847, n31848,
         n31849, n31850, n31851, n31852, n31853, n31854, n31855, n31856,
         n31857, n31858, n31859, n31860, n31861, n31862, n31863, n31864,
         n31865, n31866, n31867, n31868, n31869, n31870, n31871, n31872,
         n31873, n31874, n31875, n31876, n31877, n31878, n31879, n31880,
         n31881, n31882, n31883, n31884, n31885, n31886, n31887, n31888,
         n31889, n31890, n31891, n31892, n31893, n31894, n31895, n31896,
         n31897, n31898, n31899, n31900, n31901, n31902, n31903, n31904,
         n31905, n31906, n31907, n31908, n31909, n31910, n31911, n31912,
         n31913, n31914, n31915, n31916, n31917, n31918, n31919, n31920,
         n31921, n31922, n31923, n31924, n31925, n31926, n31927, n31928,
         n31929, n31930, n31931, n31932, n31933, n31934, n31935, n31936,
         n31937, n31938, n31939, n31940, n31941, n31942, n31943, n31944,
         n31945, n31946, n31947, n31948, n31949, n31950, n31951, n31952,
         n31953, n31954, n31955, n31956, n31957, n31958, n31959, n31960,
         n31961, n31962, n31963, n31964, n31965, n31966, n31967, n31968,
         n31969, n31970, n31971, n31972, n31973, n31974, n31975, n31976,
         n31977, n31978, n31979, n31980, n31981, n31982, n31983, n31984,
         n31985, n31986, n31987, n31988, n31989, n31990, n31991, n31992,
         n31993, n31994, n31995, n31996, n31997, n31998, n31999, n32000,
         n32001, n32002, n32003, n32004, n32005, n32006, n32007, n32008,
         n32009, n32010, n32011, n32012, n32013, n32014, n32015, n32016,
         n32017, n32018, n32019, n32020, n32021, n32022, n32023, n32024,
         n32025, n32026, n32027, n32028, n32029, n32030, n32031, n32032,
         n32033, n32034, n32035, n32036, n32037, n32038, n32039, n32040,
         n32041, n32042, n32043, n32044, n32045, n32046, n32047, n32048,
         n32049, n32050, n32051, n32052, n32053, n32054, n32055, n32056,
         n32057, n32058, n32059, n32060, n32061, n32062, n32063, n32064,
         n32065, n32066, n32067, n32068, n32069, n32070, n32071, n32072,
         n32073, n32074, n32075, n32076, n32077, n32078, n32079, n32080,
         n32081, n32082, n32083, n32084, n32085, n32086, n32087, n32088,
         n32089, n32090, n32091, n32092, n32093, n32094, n32095, n32096,
         n32097, n32098, n32099, n32100, n32101, n32102, n32103, n32104,
         n32105, n32106, n32107, n32108, n32109, n32110, n32111, n32112,
         n32113, n32114, n32115, n32116, n32117, n32118, n32119, n32120,
         n32121, n32122, n32123, n32124, n32125, n32126, n32127, n32128,
         n32129, n32130, n32131, n32132, n32133, n32134, n32135, n32136,
         n32137, n32138, n32139, n32140, n32141, n32142, n32143, n32144,
         n32145, n32146, n32147, n32148, n32149, n32150, n32151, n32152,
         n32153, n32154, n32155, n32156, n32157, n32158, n32159, n32160,
         n32161, n32162, n32163, n32164, n32165, n32166, n32167, n32168,
         n32169, n32170, n32171, n32172, n32173, n32174, n32175, n32176,
         n32177, n32178, n32179, n32180, n32181, n32182, n32183, n32184,
         n32185, n32186, n32187, n32188, n32189, n32190, n32191, n32192,
         n32193, n32194, n32195, n32196, n32197, n32198, n32199, n32200,
         n32201, n32202, n32203, n32204, n32205, n32206, n32207, n32208,
         n32209, n32210, n32211, n32212, n32213, n32214, n32215, n32216,
         n32217, n32218, n32219, n32220, n32221, n32222, n32223, n32224,
         n32225, n32226, n32227, n32228, n32229, n32230, n32231, n32232,
         n32233, n32234, n32235, n32236, n32237, n32238, n32239, n32240,
         n32241, n32242, n32243, n32244, n32245, n32246, n32247, n32248,
         n32249, n32250, n32251, n32252, n32253, n32254, n32255, n32256,
         n32257, n32258, n32259, n32260, n32261, n32262, n32263, n32264,
         n32265, n32266, n32267, n32268, n32269, n32270, n32271, n32272,
         n32273, n32274, n32275, n32276, n32277, n32278, n32279, n32280,
         n32281, n32282, n32283, n32284, n32285, n32286, n32287, n32288,
         n32289, n32290, n32291, n32292, n32293, n32294, n32295, n32296,
         n32297, n32298, n32299, n32300, n32301, n32302, n32303, n32304,
         n32305, n32306, n32307, n32308, n32309, n32310, n32311, n32312,
         n32313, n32314, n32315, n32316, n32317, n32318, n32319, n32320,
         n32321, n32322, n32323, n32324, n32325, n32326, n32327, n32328,
         n32329, n32330, n32331, n32332, n32333, n32334, n32335, n32336,
         n32337, n32338, n32339, n32340, n32341, n32342, n32343, n32344,
         n32345, n32346, n32347, n32348, n32349, n32350, n32351, n32352,
         n32353, n32354, n32355, n32356, n32357, n32358, n32359, n32360,
         n32361, n32362, n32363, n32364, n32365, n32366, n32367, n32368,
         n32369, n32370, n32371, n32372, n32373, n32374, n32375, n32376,
         n32377, n32378, n32379, n32380, n32381, n32382, n32383, n32384,
         n32385, n32386, n32387, n32388, n32389, n32390, n32391, n32392,
         n32393, n32394, n32395, n32396, n32397, n32398, n32399, n32400,
         n32401, n32402, n32403, n32404, n32405, n32406, n32407, n32408,
         n32409, n32410, n32411, n32412, n32413, n32414, n32415, n32416,
         n32417, n32418, n32419, n32420, n32421, n32422, n32423, n32424,
         n32425, n32426, n32427, n32428, n32429, n32430, n32431, n32432,
         n32433, n32434, n32435, n32436, n32437, n32438, n32439, n32440,
         n32441, n32442, n32443, n32444, n32445, n32446, n32447, n32448,
         n32449, n32450, n32451, n32452, n32453, n32454, n32455, n32456,
         n32457, n32458, n32459, n32460, n32461, n32462, n32463, n32464,
         n32465, n32466, n32467, n32468, n32469, n32470, n32471, n32472,
         n32473, n32474, n32475, n32476, n32477, n32478, n32479, n32480,
         n32481, n32482, n32483, n32484, n32485, n32486, n32487, n32488,
         n32489, n32490, n32491, n32492, n32493, n32494, n32495, n32496,
         n32497, n32498, n32499, n32500, n32501, n32502, n32503, n32504,
         n32505, n32506, n32507, n32508, n32509, n32510, n32511, n32512,
         n32513, n32514, n32515, n32516, n32517, n32518, n32519, n32520,
         n32521, n32522, n32523, n32524, n32525, n32526, n32527, n32528,
         n32529, n32530, n32531, n32532, n32533, n32534, n32535, n32536,
         n32537, n32538, n32539, n32540, n32541, n32542, n32543, n32544,
         n32545, n32546, n32547, n32548, n32549, n32550, n32551, n32552,
         n32553, n32554, n32555, n32556, n32557, n32558, n32559, n32560,
         n32561, n32562, n32563, n32564, n32565, n32566, n32567, n32568,
         n32569, n32570, n32571, n32572, n32573, n32574, n32575, n32576,
         n32577, n32578, n32579, n32580, n32581, n32582, n32583, n32584,
         n32585, n32586, n32587, n32588, n32589, n32590, n32591, n32592,
         n32593, n32594, n32595, n32596, n32597, n32598, n32599, n32600,
         n32601, n32602, n32603, n32604, n32605, n32606, n32607, n32608,
         n32609, n32610, n32611, n32612, n32613, n32614, n32615, n32616,
         n32617, n32618, n32619, n32620, n32621, n32622, n32623, n32624,
         n32625, n32626, n32627, n32628, n32629, n32630, n32631, n32632,
         n32633, n32634, n32635, n32636, n32637, n32638, n32639, n32640,
         n32641, n32642, n32643, n32644, n32645, n32646, n32647, n32648,
         n32649, n32650, n32651, n32652, n32653, n32654, n32655, n32656,
         n32657, n32658, n32659, n32660, n32661, n32662, n32663, n32664,
         n32665, n32666, n32667, n32668, n32669, n32670, n32671, n32672,
         n32673, n32674, n32675, n32676, n32677, n32678, n32679, n32680,
         n32681, n32682, n32683, n32684, n32685, n32686, n32687, n32688,
         n32689, n32690, n32691, n32692, n32693, n32694, n32695, n32696,
         n32697, n32698, n32699, n32700, n32701, n32702, n32703, n32704,
         n32705, n32706, n32707, n32708, n32709, n32710, n32711, n32712,
         n32713, n32714, n32715, n32716, n32717, n32718, n32719, n32720,
         n32721, n32722, n32723, n32724, n32725, n32726, n32727, n32728,
         n32729, n32730, n32731, n32732, n32733, n32734, n32735, n32736,
         n32737, n32738, n32739, n32740, n32741, n32742, n32743, n32744,
         n32745, n32746, n32747, n32748, n32749, n32750, n32751, n32752,
         n32753, n32754, n32755, n32756, n32757, n32758, n32759, n32760,
         n32761, n32762, n32763, n32764, n32765, n32766, n32767, n32768,
         n32769, n32770, n32771, n32772, n32773, n32774, n32775, n32776,
         n32777, n32778, n32779, n32780, n32781, n32782, n32783, n32784,
         n32785, n32786, n32787, n32788, n32789, n32790, n32791, n32792,
         n32793, n32794, n32795, n32796, n32797, n32798, n32799, n32800,
         n32801, n32802, n32803, n32804, n32805, n32806, n32807, n32808,
         n32809, n32810, n32811, n32812, n32813, n32814, n32815, n32816,
         n32817, n32818, n32819, n32820, n32821, n32822, n32823, n32824,
         n32825, n32826, n32827, n32828, n32829, n32830, n32831, n32832,
         n32833, n32834, n32835, n32836, n32837, n32838, n32839, n32840,
         n32841, n32842, n32843, n32844, n32845, n32846, n32847, n32848,
         n32849, n32850, n32851, n32852, n32853, n32854, n32855, n32856,
         n32857, n32858, n32859, n32860, n32861, n32862, n32863, n32864,
         n32865, n32866, n32867, n32868, n32869, n32870, n32871, n32872,
         n32873, n32874, n32875, n32876, n32877, n32878, n32879, n32880,
         n32881, n32882, n32883, n32884, n32885, n32886, n32887, n32888,
         n32889, n32890, n32891, n32892, n32893, n32894, n32895, n32896,
         n32897, n32898, n32899, n32900, n32901, n32902, n32903, n32904,
         n32905, n32906, n32907, n32908, n32909, n32910, n32911, n32912,
         n32913, n32914, n32915, n32916, n32917, n32918, n32919, n32920,
         n32921, n32922, n32923, n32924, n32925, n32926, n32927, n32928,
         n32929, n32930, n32931, n32932, n32933, n32934, n32935, n32936,
         n32937, n32938, n32939, n32940, n32941, n32942, n32943, n32944,
         n32945, n32946, n32947, n32948, n32949, n32950, n32951, n32952,
         n32953, n32954, n32955, n32956, n32957, n32958, n32959, n32960,
         n32961, n32962, n32963, n32964, n32965, n32966, n32967, n32968,
         n32969, n32970, n32971, n32972, n32973, n32974, n32975, n32976,
         n32977, n32978, n32979, n32980, n32981, n32982, n32983, n32984,
         n32985, n32986, n32987, n32988, n32989, n32990, n32991, n32992,
         n32993, n32994, n32995, n32996, n32997, n32998, n32999, n33000,
         n33001, n33002, n33003, n33004, n33005, n33006, n33007, n33008,
         n33009, n33010, n33011, n33012, n33013, n33014, n33015, n33016,
         n33017, n33018, n33019, n33020, n33021, n33022, n33023, n33024,
         n33025, n33026, n33027, n33028, n33029, n33030, n33031, n33032,
         n33033, n33034, n33035, n33036, n33037, n33038, n33039, n33040,
         n33041, n33042, n33043, n33044, n33045, n33046, n33047, n33048,
         n33049, n33050, n33051, n33052, n33053, n33054, n33055, n33056,
         n33057, n33058, n33059, n33060, n33061, n33062, n33063, n33064,
         n33065, n33066, n33067, n33068, n33069, n33070, n33071, n33072,
         n33073, n33074, n33075, n33076, n33077, n33078, n33079, n33080,
         n33081, n33082, n33083, n33084, n33085, n33086, n33087, n33088,
         n33089, n33090, n33091, n33092, n33093, n33094, n33095, n33096,
         n33097, n33098, n33099, n33100, n33101, n33102, n33103, n33104,
         n33105, n33106, n33107, n33108, n33109, n33110, n33111, n33112,
         n33113, n33114, n33115, n33116, n33117, n33118, n33119, n33120,
         n33121, n33122, n33123, n33124, n33125, n33126, n33127, n33128,
         n33129, n33130, n33131, n33132, n33133, n33134, n33135, n33136,
         n33137, n33138, n33139, n33140, n33141, n33142, n33143, n33144,
         n33145, n33146, n33147, n33148, n33149, n33150, n33151, n33152,
         n33153, n33154, n33155, n33156, n33157, n33158, n33159, n33160,
         n33161, n33162, n33163, n33164, n33165, n33166, n33167, n33168,
         n33169, n33170, n33171, n33172, n33173, n33174, n33175, n33176,
         n33177, n33178, n33179, n33180, n33181, n33182, n33183, n33184,
         n33185, n33186, n33187, n33188, n33189, n33190, n33191, n33192,
         n33193, n33194, n33195, n33196, n33197, n33198, n33199, n33200,
         n33201, n33202, n33203, n33204, n33205, n33206, n33207, n33208,
         n33209, n33210, n33211, n33212, n33213, n33214, n33215, n33216,
         n33217, n33218, n33219, n33220, n33221, n33222, n33223, n33224,
         n33225, n33226, n33227, n33228, n33229, n33230, n33231, n33232,
         n33233, n33234, n33235, n33236, n33237, n33238, n33239, n33240,
         n33241, n33242, n33243, n33244, n33245, n33246, n33247, n33248,
         n33249, n33250, n33251, n33252, n33253, n33254, n33255, n33256,
         n33257, n33258, n33259, n33260, n33261, n33262, n33263, n33264,
         n33265, n33266, n33267, n33268, n33269, n33270, n33271, n33272,
         n33273, n33274, n33275, n33276, n33277, n33278, n33279, n33280,
         n33281, n33282, n33283, n33284, n33285, n33286, n33287, n33288,
         n33289, n33290, n33291, n33292, n33293, n33294, n33295, n33296,
         n33297, n33298, n33299, n33300, n33301, n33302, n33303, n33304,
         n33305, n33306, n33307, n33308, n33309, n33310, n33311, n33312,
         n33313, n33314, n33315, n33316, n33317, n33318, n33319, n33320,
         n33321, n33322, n33323, n33324, n33325, n33326, n33327, n33328,
         n33329, n33330, n33331, n33332, n33333, n33334, n33335, n33336,
         n33337, n33338, n33339, n33340, n33341, n33342, n33343, n33344,
         n33345, n33346, n33347, n33348, n33349, n33350, n33351, n33352,
         n33353, n33354, n33355, n33356, n33357, n33358, n33359, n33360,
         n33361, n33362, n33363, n33364, n33365, n33366, n33367, n33368,
         n33369, n33370, n33371, n33372, n33373, n33374, n33375, n33376,
         n33377, n33378, n33379, n33380, n33381, n33382, n33383, n33384,
         n33385, n33386, n33387, n33388, n33389, n33390, n33391, n33392,
         n33393, n33394, n33395, n33396, n33397, n33398, n33399, n33400,
         n33401, n33402, n33403, n33404, n33405, n33406, n33407, n33408,
         n33409, n33410, n33411, n33412, n33413, n33414, n33415, n33416,
         n33417, n33418, n33419, n33420, n33421, n33422, n33423, n33424,
         n33425, n33426, n33427, n33428, n33429, n33430, n33431, n33432,
         n33433, n33434, n33435, n33436, n33437, n33438, n33439, n33440,
         n33441, n33442, n33443, n33444, n33445, n33446, n33447, n33448,
         n33449, n33450, n33451, n33452, n33453, n33454, n33455, n33456,
         n33457, n33458, n33459, n33460, n33461, n33462, n33463, n33464,
         n33465, n33466, n33467, n33468, n33469, n33470, n33471, n33472,
         n33473, n33474, n33475, n33476, n33477, n33478, n33479, n33480,
         n33481, n33482, n33483, n33484, n33485, n33486, n33487, n33488,
         n33489, n33490, n33491, n33492, n33493, n33494, n33495, n33496,
         n33497, n33498, n33499, n33500, n33501, n33502, n33503, n33504,
         n33505, n33506, n33507, n33508, n33509, n33510, n33511, n33512,
         n33513, n33514, n33515, n33516, n33517, n33518, n33519, n33520,
         n33521, n33522, n33523, n33524, n33525, n33526, n33527, n33528,
         n33529, n33530, n33531, n33532, n33533, n33534, n33535, n33536,
         n33537, n33538, n33539, n33540, n33541, n33542, n33543, n33544,
         n33545, n33546, n33547, n33548, n33549, n33550, n33551, n33552,
         n33553, n33554, n33555, n33556, n33557, n33558, n33559, n33560,
         n33561, n33562, n33563, n33564, n33565, n33566, n33567, n33568,
         n33569, n33570, n33571, n33572, n33573, n33574, n33575, n33576,
         n33577, n33578, n33579, n33580, n33581, n33582, n33583, n33584,
         n33585, n33586, n33587, n33588, n33589, n33590, n33591, n33592,
         n33593, n33594, n33595, n33596, n33597, n33598, n33599, n33600,
         n33601, n33602, n33603, n33604, n33605, n33606, n33607, n33608,
         n33609, n33610, n33611, n33612, n33613, n33614, n33615, n33616,
         n33617, n33618, n33619, n33620, n33621, n33622, n33623, n33624,
         n33625, n33626, n33627, n33628, n33629, n33630, n33631, n33632,
         n33633, n33634, n33635, n33636, n33637, n33638, n33639, n33640,
         n33641, n33642, n33643, n33644, n33645, n33646, n33647, n33648,
         n33649, n33650, n33651, n33652, n33653, n33654, n33655, n33656,
         n33657, n33658, n33659, n33660, n33661, n33662, n33663, n33664,
         n33665, n33666, n33667, n33668, n33669, n33670, n33671, n33672,
         n33673, n33674, n33675, n33676, n33677, n33678, n33679, n33680,
         n33681, n33682, n33683, n33684, n33685, n33686, n33687, n33688,
         n33689, n33690, n33691, n33692, n33693, n33694, n33695, n33696,
         n33697, n33698, n33699, n33700, n33701, n33702, n33703, n33704,
         n33705, n33706, n33707, n33708, n33709, n33710, n33711, n33712,
         n33713, n33714, n33715, n33716, n33717, n33718, n33719, n33720,
         n33721, n33722, n33723, n33724, n33725, n33726, n33727, n33728,
         n33729, n33730, n33731, n33732, n33733, n33734, n33735, n33736,
         n33737, n33738, n33739, n33740, n33741, n33742, n33743, n33744,
         n33745, n33746, n33747, n33748, n33749, n33750, n33751, n33752,
         n33753, n33754, n33755, n33756, n33757, n33758, n33759, n33760,
         n33761, n33762, n33763, n33764, n33765, n33766, n33767, n33768,
         n33769, n33770, n33771, n33772, n33773, n33774, n33775, n33776,
         n33777, n33778, n33779, n33780, n33781, n33782, n33783, n33784,
         n33785, n33786, n33787, n33788, n33789, n33790, n33791, n33792,
         n33793, n33794, n33795, n33796, n33797, n33798, n33799, n33800,
         n33801, n33802, n33803, n33804, n33805, n33806, n33807, n33808,
         n33809, n33810, n33811, n33812, n33813, n33814, n33815, n33816,
         n33817, n33818, n33819, n33820, n33821, n33822, n33823, n33824,
         n33825, n33826, n33827, n33828, n33829, n33830, n33831, n33832,
         n33833, n33834, n33835, n33836, n33837, n33838, n33839, n33840,
         n33841, n33842, n33843, n33844, n33845, n33846, n33847, n33848,
         n33849, n33850, n33851, n33852, n33853, n33854, n33855, n33856,
         n33857, n33858, n33859, n33860, n33861, n33862, n33863, n33864,
         n33865, n33866, n33867, n33868, n33869, n33870, n33871, n33872,
         n33873, n33874, n33875, n33876, n33877, n33878, n33879, n33880,
         n33881, n33882, n33883, n33884, n33885, n33886, n33887, n33888,
         n33889, n33890, n33891, n33892, n33893, n33894, n33895, n33896,
         n33897, n33898, n33899, n33900, n33901, n33902, n33903, n33904,
         n33905, n33906, n33907, n33908, n33909, n33910, n33911, n33912,
         n33913, n33914, n33915, n33916, n33917, n33918, n33919, n33920,
         n33921, n33922, n33923, n33924, n33925, n33926, n33927, n33928,
         n33929, n33930, n33931, n33932, n33933, n33934, n33935, n33936,
         n33937, n33938, n33939, n33940, n33941, n33942, n33943, n33944,
         n33945, n33946, n33947, n33948, n33949, n33950, n33951, n33952,
         n33953, n33954, n33955, n33956, n33957, n33958, n33959, n33960,
         n33961, n33962, n33963, n33964, n33965, n33966, n33967, n33968,
         n33969, n33970, n33971, n33972, n33973, n33974, n33975, n33976,
         n33977, n33978, n33979, n33980, n33981, n33982, n33983, n33984,
         n33985, n33986, n33987, n33988, n33989, n33990, n33991, n33992,
         n33993, n33994, n33995, n33996, n33997, n33998, n33999, n34000,
         n34001, n34002, n34003, n34004, n34005, n34006, n34007, n34008,
         n34009, n34010, n34011, n34012, n34013, n34014, n34015, n34016,
         n34017, n34018, n34019, n34020, n34021, n34022, n34023, n34024,
         n34025, n34026, n34027, n34028, n34029, n34030, n34031, n34032,
         n34033, n34034, n34035, n34036, n34037, n34038, n34039, n34040,
         n34041, n34042, n34043, n34044, n34045, n34046, n34047, n34048,
         n34049, n34050, n34051, n34052, n34053, n34054, n34055, n34056,
         n34057, n34058, n34059, n34060, n34061, n34062, n34063, n34064,
         n34065, n34066, n34067, n34068, n34069, n34070, n34071, n34072,
         n34073, n34074, n34075, n34076, n34077, n34078, n34079, n34080,
         n34081, n34082, n34083, n34084, n34085, n34086, n34087, n34088,
         n34089, n34090, n34091, n34092, n34093, n34094, n34095, n34096,
         n34097, n34098, n34099, n34100, n34101, n34102, n34103, n34104,
         n34105, n34106, n34107, n34108, n34109, n34110, n34111, n34112,
         n34113, n34114, n34115, n34116, n34117, n34118, n34119, n34120,
         n34121, n34122, n34123, n34124, n34125, n34126, n34127, n34128,
         n34129, n34130, n34131, n34132, n34133, n34134, n34135, n34136,
         n34137, n34138, n34139, n34140, n34141, n34142, n34143, n34144,
         n34145, n34146, n34147, n34148, n34149, n34150, n34151, n34152,
         n34153, n34154, n34155, n34156, n34157, n34158, n34159, n34160,
         n34161, n34162, n34163, n34164, n34165, n34166, n34167, n34168,
         n34169, n34170, n34171, n34172, n34173, n34174, n34175, n34176,
         n34177, n34178, n34179, n34180, n34181, n34182, n34183, n34184,
         n34185, n34186, n34187, n34188, n34189, n34190, n34191, n34192,
         n34193, n34194, n34195, n34196, n34197, n34198, n34199, n34200,
         n34201, n34202, n34203, n34204, n34205, n34206, n34207, n34208,
         n34209, n34210, n34211, n34212, n34213, n34214, n34215, n34216,
         n34217, n34218, n34219, n34220, n34221, n34222, n34223, n34224,
         n34225, n34226, n34227, n34228, n34229, n34230, n34231, n34232,
         n34233, n34234, n34235, n34236, n34237, n34238, n34239, n34240,
         n34241, n34242, n34243, n34244, n34245, n34246, n34247, n34248,
         n34249, n34250, n34251, n34252, n34253, n34254, n34255, n34256,
         n34257, n34258, n34259, n34260, n34261, n34262, n34263, n34264,
         n34265, n34266, n34267, n34268, n34269, n34270, n34271, n34272,
         n34273, n34274, n34275, n34276, n34277, n34278, n34279, n34280,
         n34281, n34282, n34283, n34284, n34285, n34286, n34287, n34288,
         n34289, n34290, n34291, n34292, n34293, n34294, n34295, n34296,
         n34297, n34298, n34299, n34300, n34301, n34302, n34303, n34304,
         n34305, n34306, n34307, n34308, n34309, n34310, n34311, n34312,
         n34313, n34314, n34315, n34316, n34317, n34318, n34319, n34320,
         n34321, n34322, n34323, n34324, n34325, n34326, n34327, n34328,
         n34329, n34330, n34331, n34332, n34333, n34334, n34335, n34336,
         n34337, n34338, n34339, n34340, n34341, n34342, n34343, n34344,
         n34345, n34346, n34347, n34348, n34349, n34350, n34351, n34352,
         n34353, n34354, n34355, n34356, n34357, n34358, n34359, n34360,
         n34361, n34362, n34363, n34364, n34365, n34366, n34367, n34368,
         n34369, n34370, n34371, n34372, n34373, n34374, n34375, n34376,
         n34377, n34378, n34379, n34380, n34381, n34382, n34383, n34384,
         n34385, n34386, n34387, n34388, n34389, n34390, n34391, n34392,
         n34393, n34394, n34395, n34396, n34397, n34398, n34399, n34400,
         n34401, n34402, n34403, n34404, n34405, n34406, n34407, n34408,
         n34409, n34410, n34411, n34412, n34413, n34414, n34415, n34416,
         n34417, n34418, n34419, n34420, n34421, n34422, n34423, n34424,
         n34425, n34426, n34427, n34428, n34429, n34430, n34431, n34432,
         n34433, n34434, n34435, n34436, n34437, n34438, n34439, n34440,
         n34441, n34442, n34443, n34444, n34445, n34446, n34447, n34448,
         n34449, n34450, n34451, n34452, n34453, n34454, n34455, n34456,
         n34457, n34458, n34459, n34460, n34461, n34462, n34463, n34464,
         n34465, n34466, n34467, n34468, n34469, n34470, n34471, n34472,
         n34473, n34474, n34475, n34476, n34477, n34478, n34479, n34480,
         n34481, n34482, n34483, n34484, n34485, n34486, n34487, n34488,
         n34489, n34490, n34491, n34492, n34493, n34494, n34495, n34496,
         n34497, n34498, n34499, n34500, n34501, n34502, n34503, n34504,
         n34505, n34506, n34507, n34508, n34509, n34510, n34511, n34512,
         n34513, n34514, n34515, n34516, n34517, n34518, n34519, n34520,
         n34521, n34522, n34523, n34524, n34525, n34526, n34527, n34528,
         n34529, n34530, n34531, n34532, n34533, n34534, n34535, n34536,
         n34537, n34538, n34539, n34540, n34541, n34542, n34543, n34544,
         n34545, n34546, n34547, n34548, n34549, n34550, n34551, n34552,
         n34553, n34554, n34555, n34556, n34557, n34558, n34559, n34560,
         n34561, n34562, n34563, n34564, n34565, n34566, n34567, n34568,
         n34569, n34570, n34571, n34572, n34573, n34574, n34575, n34576,
         n34577, n34578, n34579, n34580, n34581, n34582, n34583, n34584,
         n34585, n34586, n34587, n34588, n34589, n34590, n34591, n34592,
         n34593, n34594, n34595, n34596, n34597, n34598, n34599, n34600,
         n34601, n34602, n34603, n34604, n34605, n34606, n34607, n34608,
         n34609, n34610, n34611, n34612, n34613, n34614, n34615, n34616,
         n34617, n34618, n34619, n34620, n34621, n34622, n34623, n34624,
         n34625, n34626, n34627, n34628, n34629, n34630, n34631, n34632,
         n34633, n34634, n34635, n34636, n34637, n34638, n34639, n34640,
         n34641, n34642, n34643, n34644, n34645, n34646, n34647, n34648,
         n34649, n34650, n34651, n34652, n34653, n34654, n34655, n34656,
         n34657, n34658, n34659, n34660, n34661, n34662, n34663, n34664,
         n34665, n34666, n34667, n34668, n34669, n34670, n34671, n34672,
         n34673, n34674, n34675, n34676, n34677, n34678, n34679, n34680,
         n34681, n34682, n34683, n34684, n34685, n34686, n34687, n34688,
         n34689, n34690, n34691, n34692, n34693, n34694, n34695, n34696,
         n34697, n34698, n34699, n34700, n34701, n34702, n34703, n34704,
         n34705, n34706, n34707, n34708, n34709, n34710, n34711, n34712,
         n34713, n34714, n34715, n34716, n34717, n34718, n34719, n34720,
         n34721, n34722, n34723, n34724, n34725, n34726, n34727, n34728,
         n34729, n34730, n34731, n34732, n34733, n34734, n34735, n34736,
         n34737, n34738, n34739, n34740, n34741, n34742, n34743, n34744,
         n34745, n34746, n34747, n34748, n34749, n34750, n34751, n34752,
         n34753, n34754, n34755, n34756, n34757, n34758, n34759, n34760,
         n34761, n34762, n34763, n34764, n34765, n34766, n34767, n34768,
         n34769, n34770, n34771, n34772, n34773, n34774, n34775, n34776,
         n34777, n34778, n34779, n34780, n34781, n34782, n34783, n34784,
         n34785, n34786, n34787, n34788, n34789, n34790, n34791, n34792,
         n34793, n34794, n34795, n34796, n34797, n34798, n34799, n34800,
         n34801, n34802, n34803, n34804, n34805, n34806, n34807, n34808,
         n34809, n34810, n34811, n34812, n34813, n34814, n34815, n34816,
         n34817, n34818, n34819, n34820, n34821, n34822, n34823, n34824,
         n34825, n34826, n34827, n34828, n34829, n34830, n34831, n34832,
         n34833, n34834, n34835, n34836, n34837, n34838, n34839, n34840,
         n34841, n34842, n34843, n34844, n34845, n34846, n34847, n34848,
         n34849, n34850, n34851, n34852, n34853, n34854, n34855, n34856,
         n34857, n34858, n34859, n34860, n34861, n34862, n34863, n34864,
         n34865, n34866, n34867, n34868, n34869, n34870, n34871, n34872,
         n34873, n34874, n34875, n34876, n34877, n34878, n34879, n34880,
         n34881, n34882, n34883, n34884, n34885, n34886, n34887, n34888,
         n34889, n34890, n34891, n34892, n34893, n34894, n34895, n34896,
         n34897, n34898, n34899, n34900, n34901, n34902, n34903, n34904,
         n34905, n34906, n34907, n34908, n34909, n34910, n34911, n34912,
         n34913, n34914, n34915, n34916, n34917, n34918, n34919, n34920,
         n34921, n34922, n34923, n34924, n34925, n34926, n34927, n34928,
         n34929, n34930, n34931, n34932, n34933, n34934, n34935, n34936,
         n34937, n34938, n34939, n34940, n34941, n34942, n34943, n34944,
         n34945, n34946, n34947, n34948, n34949, n34950, n34951, n34952,
         n34953, n34954, n34955, n34956, n34957, n34958, n34959, n34960,
         n34961, n34962, n34963, n34964, n34965, n34966, n34967, n34968,
         n34969, n34970, n34971, n34972, n34973, n34974, n34975, n34976,
         n34977, n34978, n34979, n34980, n34981, n34982, n34983, n34984,
         n34985, n34986, n34987, n34988, n34989, n34990, n34991, n34992,
         n34993, n34994, n34995, n34996, n34997, n34998, n34999, n35000,
         n35001, n35002, n35003, n35004, n35005, n35006, n35007, n35008,
         n35009, n35010, n35011, n35012, n35013, n35014, n35015, n35016,
         n35017, n35018, n35019, n35020, n35021, n35022, n35023, n35024,
         n35025, n35026, n35027, n35028, n35029, n35030, n35031, n35032,
         n35033, n35034, n35035, n35036, n35037, n35038, n35039, n35040,
         n35041, n35042, n35043, n35044, n35045, n35046, n35047, n35048,
         n35049, n35050, n35051, n35052, n35053, n35054, n35055, n35056,
         n35057, n35058, n35059, n35060, n35061, n35062, n35063, n35064,
         n35065, n35066, n35067, n35068, n35069, n35070, n35071, n35072,
         n35073, n35074, n35075, n35076, n35077, n35078, n35079, n35080,
         n35081, n35082, n35083, n35084, n35085, n35086, n35087, n35088,
         n35089, n35090, n35091, n35092, n35093, n35094, n35095, n35096,
         n35097, n35098, n35099, n35100, n35101, n35102, n35103, n35104,
         n35105, n35106, n35107, n35108, n35109, n35110, n35111, n35112,
         n35113, n35114, n35115, n35116, n35117, n35118, n35119, n35120,
         n35121, n35122, n35123, n35124, n35125, n35126, n35127, n35128,
         n35129, n35130, n35131, n35132, n35133, n35134, n35135, n35136,
         n35137, n35138, n35139, n35140, n35141, n35142, n35143, n35144,
         n35145, n35146, n35147, n35148, n35149, n35150, n35151, n35152,
         n35153, n35154, n35155, n35156, n35157, n35158, n35159, n35160,
         n35161, n35162, n35163, n35164, n35165, n35166, n35167, n35168,
         n35169, n35170, n35171, n35172, n35173, n35174, n35175, n35176,
         n35177, n35178, n35179, n35180, n35181, n35182, n35183, n35184,
         n35185, n35186, n35187, n35188, n35189, n35190, n35191, n35192,
         n35193, n35194, n35195, n35196, n35197, n35198, n35199, n35200,
         n35201, n35202, n35203, n35204, n35205, n35206, n35207, n35208,
         n35209, n35210, n35211, n35212, n35213, n35214, n35215, n35216,
         n35217, n35218, n35219, n35220, n35221, n35222, n35223, n35224,
         n35225, n35226, n35227, n35228, n35229, n35230, n35231, n35232,
         n35233, n35234, n35235, n35236, n35237, n35238, n35239, n35240,
         n35241, n35242, n35243, n35244, n35245, n35246, n35247, n35248,
         n35249, n35250, n35251, n35252, n35253, n35254, n35255, n35256,
         n35257, n35258, n35259, n35260, n35261, n35262, n35263, n35264,
         n35265, n35266, n35267, n35268, n35269, n35270, n35271, n35272,
         n35273, n35274, n35275, n35276, n35277, n35278, n35279, n35280,
         n35281, n35282, n35283, n35284, n35285, n35286, n35287, n35288,
         n35289, n35290, n35291, n35292, n35293, n35294, n35295, n35296,
         n35297, n35298, n35299, n35300, n35301, n35302, n35303, n35304,
         n35305, n35306, n35307, n35308, n35309, n35310, n35311, n35312,
         n35313, n35314, n35315, n35316, n35317, n35318, n35319, n35320,
         n35321, n35322, n35323, n35324, n35325, n35326, n35327, n35328,
         n35329, n35330, n35331, n35332, n35333, n35334, n35335, n35336,
         n35337, n35338, n35339, n35340, n35341, n35342, n35343, n35344,
         n35345, n35346, n35347, n35348, n35349, n35350, n35351, n35352,
         n35353, n35354, n35355, n35356, n35357, n35358, n35359, n35360,
         n35361, n35362, n35363, n35364, n35365, n35366, n35367, n35368,
         n35369, n35370, n35371, n35372, n35373, n35374, n35375, n35376,
         n35377, n35378, n35379, n35380, n35381, n35382, n35383, n35384,
         n35385, n35386, n35387, n35388, n35389, n35390, n35391, n35392,
         n35393, n35394, n35395, n35396, n35397, n35398, n35399, n35400,
         n35401, n35402, n35403, n35404, n35405, n35406, n35407, n35408,
         n35409, n35410, n35411, n35412, n35413, n35414, n35415, n35416,
         n35417, n35418, n35419, n35420, n35421, n35422, n35423, n35424,
         n35425, n35426, n35427, n35428, n35429, n35430, n35431, n35432,
         n35433, n35434, n35435, n35436, n35437, n35438, n35439, n35440,
         n35441, n35442, n35443, n35444, n35445, n35446, n35447, n35448,
         n35449, n35450, n35451, n35452, n35453, n35454, n35455, n35456,
         n35457, n35458, n35459, n35460, n35461, n35462, n35463, n35464,
         n35465, n35466, n35467, n35468, n35469, n35470, n35471, n35472,
         n35473, n35474, n35475, n35476, n35477, n35478, n35479, n35480,
         n35481, n35482, n35483, n35484, n35485, n35486, n35487, n35488,
         n35489, n35490, n35491, n35492, n35493, n35494, n35495, n35496,
         n35497, n35498, n35499, n35500, n35501, n35502, n35503, n35504,
         n35505, n35506, n35507, n35508, n35509, n35510, n35511, n35512,
         n35513, n35514, n35515, n35516, n35517, n35518, n35519, n35520,
         n35521, n35522, n35523, n35524, n35525, n35526, n35527, n35528,
         n35529, n35530, n35531, n35532, n35533, n35534, n35535, n35536,
         n35537, n35538, n35539, n35540, n35541, n35542, n35543, n35544,
         n35545, n35546, n35547, n35548, n35549, n35550, n35551, n35552,
         n35553, n35554, n35555, n35556, n35557, n35558, n35559, n35560,
         n35561, n35562, n35563, n35564, n35565, n35566, n35567, n35568,
         n35569, n35570, n35571, n35572, n35573, n35574, n35575, n35576,
         n35577, n35578, n35579, n35580, n35581, n35582, n35583, n35584,
         n35585, n35586, n35587, n35588, n35589, n35590, n35591, n35592,
         n35593, n35594, n35595, n35596, n35597, n35598, n35599, n35600,
         n35601, n35602, n35603, n35604, n35605, n35606, n35607, n35608,
         n35609, n35610, n35611, n35612, n35613, n35614, n35615, n35616,
         n35617, n35618, n35619, n35620, n35621, n35622, n35623, n35624,
         n35625, n35626, n35627, n35628, n35629, n35630, n35631, n35632,
         n35633, n35634, n35635, n35636, n35637, n35638, n35639, n35640,
         n35641, n35642, n35643, n35644, n35645, n35646, n35647, n35648,
         n35649, n35650, n35651, n35652, n35653, n35654, n35655, n35656,
         n35657, n35658, n35659, n35660, n35661, n35662, n35663, n35664,
         n35665, n35666, n35667, n35668, n35669, n35670, n35671, n35672,
         n35673, n35674, n35675, n35676, n35677, n35678, n35679, n35680,
         n35681, n35682, n35683, n35684, n35685, n35686, n35687, n35688,
         n35689, n35690, n35691, n35692, n35693, n35694, n35695, n35696,
         n35697, n35698, n35699, n35700, n35701, n35702, n35703, n35704,
         n35705, n35706, n35707, n35708, n35709, n35710, n35711, n35712,
         n35713, n35714, n35715, n35716, n35717, n35718, n35719, n35720,
         n35721, n35722, n35723, n35724, n35725, n35726, n35727, n35728,
         n35729, n35730, n35731, n35732, n35733, n35734, n35735, n35736,
         n35737, n35738, n35739, n35740, n35741, n35742, n35743, n35744,
         n35745, n35746, n35747, n35748, n35749, n35750, n35751, n35752,
         n35753, n35754, n35755, n35756, n35757, n35758, n35759, n35760,
         n35761, n35762, n35763, n35764, n35765, n35766, n35767, n35768,
         n35769, n35770, n35771, n35772, n35773, n35774, n35775, n35776,
         n35777, n35778, n35779, n35780, n35781, n35782, n35783, n35784,
         n35785, n35786, n35787, n35788, n35789, n35790, n35791, n35792,
         n35793, n35794, n35795, n35796, n35797, n35798, n35799, n35800,
         n35801, n35802, n35803, n35804, n35805, n35806, n35807, n35808,
         n35809, n35810, n35811, n35812, n35813, n35814, n35815, n35816,
         n35817, n35818, n35819, n35820, n35821, n35822, n35823, n35824,
         n35825, n35826, n35827, n35828, n35829, n35830, n35831, n35832,
         n35833, n35834, n35835, n35836, n35837, n35838, n35839, n35840,
         n35841, n35842, n35843, n35844, n35845, n35846, n35847, n35848,
         n35849, n35850, n35851, n35852, n35853, n35854, n35855, n35856,
         n35857, n35858, n35859, n35860, n35861, n35862, n35863, n35864,
         n35865, n35866, n35867, n35868, n35869, n35870, n35871, n35872,
         n35873, n35874, n35875, n35876, n35877, n35878, n35879, n35880,
         n35881, n35882, n35883, n35884, n35885, n35886, n35887, n35888,
         n35889, n35890, n35891, n35892, n35893, n35894, n35895, n35896,
         n35897, n35898, n35899, n35900, n35901, n35902, n35903, n35904,
         n35905, n35906, n35907, n35908, n35909, n35910, n35911, n35912,
         n35913, n35914, n35915, n35916, n35917, n35918, n35919, n35920,
         n35921, n35922, n35923, n35924, n35925, n35926, n35927, n35928,
         n35929, n35930, n35931, n35932, n35933, n35934, n35935, n35936,
         n35937, n35938, n35939, n35940, n35941, n35942, n35943, n35944,
         n35945, n35946, n35947, n35948, n35949, n35950, n35951, n35952,
         n35953, n35954, n35955, n35956, n35957, n35958, n35959, n35960,
         n35961, n35962, n35963, n35964, n35965, n35966, n35967, n35968,
         n35969, n35970, n35971, n35972, n35973, n35974, n35975, n35976,
         n35977, n35978, n35979, n35980, n35981, n35982, n35983, n35984,
         n35985, n35986, n35987, n35988, n35989, n35990, n35991, n35992,
         n35993, n35994, n35995, n35996, n35997, n35998, n35999, n36000,
         n36001, n36002, n36003, n36004, n36005, n36006, n36007, n36008,
         n36009, n36010, n36011, n36012, n36013, n36014, n36015, n36016,
         n36017, n36018, n36019, n36020, n36021, n36022, n36023, n36024,
         n36025, n36026, n36027, n36028, n36029, n36030, n36031, n36032,
         n36033, n36034, n36035, n36036, n36037, n36038, n36039, n36040,
         n36041, n36042, n36043, n36044, n36045, n36046, n36047, n36048,
         n36049, n36050, n36051, n36052, n36053, n36054, n36055, n36056,
         n36057, n36058, n36059, n36060, n36061, n36062, n36063, n36064,
         n36065, n36066, n36067, n36068, n36069, n36070, n36071, n36072,
         n36073, n36074, n36075, n36076, n36077, n36078, n36079, n36080,
         n36081, n36082, n36083, n36084, n36085, n36086, n36087, n36088,
         n36089, n36090, n36091, n36092, n36093, n36094, n36095, n36096,
         n36097, n36098, n36099, n36100, n36101, n36102, n36103, n36104,
         n36105, n36106, n36107, n36108, n36109, n36110, n36111, n36112,
         n36113, n36114, n36115, n36116, n36117, n36118, n36119, n36120,
         n36121, n36122, n36123, n36124, n36125, n36126, n36127, n36128,
         n36129, n36130, n36131, n36132, n36133, n36134, n36135, n36136,
         n36137, n36138, n36139, n36140, n36141, n36142, n36143, n36144,
         n36145, n36146, n36147, n36148, n36149, n36150, n36151, n36152,
         n36153, n36154, n36155, n36156, n36157, n36158, n36159, n36160,
         n36161, n36162, n36163, n36164, n36165, n36166, n36167, n36168,
         n36169, n36170, n36171, n36172, n36173, n36174, n36175, n36176,
         n36177, n36178, n36179, n36180, n36181, n36182, n36183, n36184,
         n36185, n36186, n36187, n36188, n36189, n36190, n36191, n36192,
         n36193, n36194, n36195, n36196, n36197, n36198, n36199, n36200,
         n36201, n36202, n36203, n36204, n36205, n36206, n36207, n36208,
         n36209, n36210, n36211, n36212, n36213, n36214, n36215, n36216,
         n36217, n36218, n36219, n36220, n36221, n36222, n36223, n36224,
         n36225, n36226, n36227, n36228, n36229, n36230, n36231, n36232,
         n36233, n36234, n36235, n36236, n36237, n36238, n36239, n36240,
         n36241, n36242, n36243, n36244, n36245, n36246, n36247, n36248,
         n36249, n36250, n36251, n36252, n36253, n36254, n36255, n36256,
         n36257, n36258, n36259, n36260, n36261, n36262, n36263, n36264,
         n36265, n36266, n36267, n36268, n36269, n36270, n36271, n36272,
         n36273, n36274, n36275, n36276, n36277, n36278, n36279, n36280,
         n36281, n36282, n36283, n36284, n36285, n36286, n36287, n36288,
         n36289, n36290, n36291, n36292, n36293, n36294, n36295, n36296,
         n36297, n36298, n36299, n36300, n36301, n36302, n36303, n36304,
         n36305, n36306, n36307, n36308, n36309, n36310, n36311, n36312,
         n36313, n36314, n36315, n36316, n36317, n36318, n36319, n36320,
         n36321, n36322, n36323, n36324, n36325, n36326, n36327, n36328,
         n36329, n36330, n36331, n36332, n36333, n36334, n36335, n36336,
         n36337, n36338, n36339, n36340, n36341, n36342, n36343, n36344,
         n36345, n36346, n36347, n36348, n36349, n36350, n36351, n36352,
         n36353, n36354, n36355, n36356, n36357, n36358, n36359, n36360,
         n36361, n36362, n36363, n36364, n36365, n36366, n36367, n36368,
         n36369, n36370, n36371, n36372, n36373, n36374, n36375, n36376,
         n36377, n36378, n36379, n36380, n36381, n36382, n36383, n36384,
         n36385, n36386, n36387, n36388, n36389, n36390, n36391, n36392,
         n36393, n36394, n36395, n36396, n36397, n36398, n36399, n36400,
         n36401, n36402, n36403, n36404, n36405, n36406, n36407, n36408,
         n36409, n36410, n36411, n36412, n36413, n36414, n36415, n36416,
         n36417, n36418, n36419, n36420, n36421, n36422, n36423, n36424,
         n36425, n36426, n36427, n36428, n36429, n36430, n36431, n36432,
         n36433, n36434, n36435, n36436, n36437, n36438, n36439, n36440,
         n36441, n36442, n36443, n36444, n36445, n36446, n36447, n36448,
         n36449, n36450, n36451, n36452, n36453, n36454, n36455, n36456,
         n36457, n36458, n36459, n36460, n36461, n36462, n36463, n36464,
         n36465, n36466, n36467, n36468, n36469, n36470, n36471, n36472,
         n36473, n36474, n36475, n36476, n36477, n36478, n36479, n36480,
         n36481, n36482, n36483, n36484, n36485, n36486, n36487, n36488,
         n36489, n36490, n36491, n36492, n36493, n36494, n36495, n36496,
         n36497, n36498, n36499, n36500, n36501, n36502, n36503, n36504,
         n36505, n36506, n36507, n36508, n36509, n36510, n36511, n36512,
         n36513, n36514, n36515, n36516, n36517, n36518, n36519, n36520,
         n36521, n36522, n36523, n36524, n36525, n36526, n36527, n36528,
         n36529, n36530, n36531, n36532, n36533, n36534, n36535, n36536,
         n36537, n36538, n36539, n36540, n36541, n36542, n36543, n36544,
         n36545, n36546, n36547, n36548, n36549, n36550, n36551, n36552,
         n36553, n36554, n36555, n36556, n36557, n36558, n36559, n36560,
         n36561, n36562, n36563, n36564, n36565, n36566, n36567, n36568,
         n36569, n36570, n36571, n36572, n36573, n36574, n36575, n36576,
         n36577, n36578, n36579, n36580, n36581, n36582, n36583, n36584,
         n36585, n36586, n36587, n36588, n36589, n36590, n36591, n36592,
         n36593, n36594, n36595, n36596, n36597, n36598, n36599, n36600,
         n36601, n36602, n36603, n36604, n36605, n36606, n36607, n36608,
         n36609, n36610, n36611, n36612, n36613, n36614, n36615, n36616,
         n36617, n36618, n36619, n36620, n36621, n36622, n36623, n36624,
         n36625, n36626, n36627, n36628, n36629, n36630, n36631, n36632,
         n36633, n36634, n36635, n36636, n36637, n36638, n36639, n36640,
         n36641, n36642, n36643, n36644, n36645, n36646, n36647, n36648,
         n36649, n36650, n36651, n36652, n36653, n36654, n36655, n36656,
         n36657, n36658, n36659, n36660, n36661, n36662, n36663, n36664,
         n36665, n36666, n36667, n36668, n36669, n36670, n36671, n36672,
         n36673, n36674, n36675, n36676, n36677, n36678, n36679, n36680,
         n36681, n36682, n36683, n36684, n36685, n36686, n36687, n36688,
         n36689, n36690, n36691, n36692, n36693, n36694, n36695, n36696,
         n36697, n36698, n36699, n36700, n36701, n36702, n36703, n36704,
         n36705, n36706, n36707, n36708, n36709, n36710, n36711, n36712,
         n36713, n36714, n36715, n36716, n36717, n36718, n36719, n36720,
         n36721, n36722, n36723, n36724, n36725, n36726, n36727, n36728,
         n36729, n36730, n36731, n36732, n36733, n36734, n36735, n36736,
         n36737, n36738, n36739, n36740, n36741, n36742, n36743, n36744,
         n36745, n36746, n36747, n36748, n36749, n36750, n36751, n36752,
         n36753, n36754, n36755, n36756, n36757, n36758, n36759, n36760,
         n36761, n36762, n36763, n36764, n36765, n36766, n36767, n36768,
         n36769, n36770, n36771, n36772, n36773, n36774, n36775, n36776,
         n36777, n36778, n36779, n36780, n36781, n36782, n36783, n36784,
         n36785, n36786, n36787, n36788, n36789, n36790, n36791, n36792,
         n36793, n36794, n36795, n36796, n36797, n36798, n36799, n36800,
         n36801, n36802, n36803, n36804, n36805, n36806, n36807, n36808,
         n36809, n36810, n36811, n36812, n36813, n36814, n36815, n36816,
         n36817, n36818, n36819, n36820, n36821, n36822, n36823, n36824,
         n36825, n36826, n36827, n36828, n36829, n36830, n36831, n36832,
         n36833, n36834, n36835, n36836, n36837, n36838, n36839, n36840,
         n36841, n36842, n36843, n36844, n36845, n36846, n36847, n36848,
         n36849, n36850, n36851, n36852, n36853, n36854, n36855, n36856,
         n36857, n36858, n36859, n36860, n36861, n36862, n36863, n36864,
         n36865, n36866, n36867, n36868, n36869, n36870, n36871, n36872,
         n36873, n36874, n36875, n36876, n36877, n36878, n36879, n36880,
         n36881, n36882, n36883, n36884, n36885, n36886, n36887, n36888,
         n36889, n36890, n36891, n36892, n36893, n36894, n36895, n36896,
         n36897, n36898, n36899, n36900, n36901, n36902, n36903, n36904,
         n36905, n36906, n36907, n36908, n36909, n36910, n36911, n36912,
         n36913, n36914, n36915, n36916, n36917, n36918, n36919, n36920,
         n36921, n36922, n36923, n36924, n36925, n36926, n36927, n36928,
         n36929, n36930, n36931, n36932, n36933, n36934, n36935, n36936,
         n36937, n36938, n36939, n36940, n36941, n36942, n36943, n36944,
         n36945, n36946, n36947, n36948, n36949, n36950, n36951, n36952,
         n36953, n36954, n36955, n36956, n36957, n36958, n36959, n36960,
         n36961, n36962, n36963, n36964, n36965, n36966, n36967, n36968,
         n36969, n36970, n36971, n36972, n36973, n36974, n36975, n36976,
         n36977, n36978, n36979, n36980, n36981, n36982, n36983, n36984,
         n36985, n36986, n36987, n36988, n36989, n36990, n36991, n36992,
         n36993, n36994, n36995, n36996, n36997, n36998, n36999, n37000,
         n37001, n37002, n37003, n37004, n37005, n37006, n37007, n37008,
         n37009, n37010, n37011, n37012, n37013, n37014, n37015, n37016,
         n37017, n37018, n37019, n37020, n37021, n37022, n37023, n37024,
         n37025, n37026, n37027, n37028, n37029, n37030, n37031, n37032,
         n37033, n37034, n37035, n37036, n37037, n37038, n37039, n37040,
         n37041, n37042, n37043, n37044, n37045, n37046, n37047, n37048,
         n37049, n37050, n37051, n37052, n37053, n37054, n37055, n37056,
         n37057, n37058, n37059, n37060, n37061, n37062, n37063, n37064,
         n37065, n37066, n37067, n37068, n37069, n37070, n37071, n37072,
         n37073, n37074, n37075, n37076, n37077, n37078, n37079, n37080,
         n37081, n37082, n37083, n37084, n37085, n37086, n37087, n37088,
         n37089, n37090, n37091, n37092, n37093, n37094, n37095, n37096,
         n37097, n37098, n37099, n37100, n37101, n37102, n37103, n37104,
         n37105, n37106, n37107, n37108, n37109, n37110, n37111, n37112,
         n37113, n37114, n37115, n37116, n37117, n37118, n37119, n37120,
         n37121, n37122, n37123, n37124, n37125, n37126, n37127, n37128,
         n37129, n37130, n37131, n37132, n37133, n37134, n37135, n37136,
         n37137, n37138, n37139, n37140, n37141, n37142, n37143, n37144,
         n37145, n37146, n37147, n37148, n37149, n37150, n37151, n37152,
         n37153, n37154, n37155, n37156, n37157, n37158, n37159, n37160,
         n37161, n37162, n37163, n37164, n37165, n37166, n37167, n37168,
         n37169, n37170, n37171, n37172, n37173, n37174, n37175, n37176,
         n37177, n37178, n37179, n37180, n37181, n37182, n37183, n37184,
         n37185, n37186, n37187, n37188, n37189, n37190, n37191, n37192,
         n37193, n37194, n37195, n37196, n37197, n37198, n37199, n37200,
         n37201, n37202, n37203, n37204, n37205, n37206, n37207, n37208,
         n37209, n37210, n37211, n37212, n37213, n37214, n37215, n37216,
         n37217, n37218, n37219, n37220, n37221, n37222, n37223, n37224,
         n37225, n37226, n37227, n37228, n37229, n37230, n37231, n37232,
         n37233, n37234, n37235, n37236, n37237, n37238, n37239, n37240,
         n37241, n37242, n37243, n37244, n37245, n37246, n37247, n37248,
         n37249, n37250, n37251, n37252, n37253, n37254, n37255, n37256,
         n37257, n37258, n37259, n37260, n37261, n37262, n37263, n37264,
         n37265, n37266, n37267, n37268, n37269, n37270, n37271, n37272,
         n37273, n37274, n37275, n37276, n37277, n37278, n37279, n37280,
         n37281, n37282, n37283, n37284, n37285, n37286, n37287, n37288,
         n37289, n37290, n37291, n37292, n37293, n37294, n37295, n37296,
         n37297, n37298, n37299, n37300, n37301, n37302, n37303, n37304,
         n37305, n37306, n37307, n37308, n37309, n37310, n37311, n37312,
         n37313, n37314, n37315, n37316, n37317, n37318, n37319, n37320,
         n37321, n37322, n37323, n37324, n37325, n37326, n37327, n37328,
         n37329, n37330, n37331, n37332, n37333, n37334, n37335, n37336,
         n37337, n37338, n37339, n37340, n37341, n37342, n37343, n37344,
         n37345, n37346, n37347, n37348, n37349, n37350, n37351, n37352,
         n37353, n37354, n37355, n37356, n37357, n37358, n37359, n37360,
         n37361, n37362, n37363, n37364, n37365, n37366, n37367, n37368,
         n37369, n37370, n37371, n37372, n37373, n37374, n37375, n37376,
         n37377, n37378, n37379, n37380, n37381, n37382, n37383, n37384,
         n37385, n37386, n37387, n37388, n37389, n37390, n37391, n37392,
         n37393, n37394, n37395, n37396, n37397, n37398, n37399, n37400,
         n37401, n37402, n37403, n37404, n37405, n37406, n37407, n37408,
         n37409, n37410, n37411, n37412, n37413, n37414, n37415, n37416,
         n37417, n37418, n37419, n37420, n37421, n37422, n37423, n37424,
         n37425, n37426, n37427, n37428, n37429, n37430, n37431, n37432,
         n37433, n37434, n37435, n37436, n37437, n37438, n37439, n37440,
         n37441, n37442, n37443, n37444, n37445, n37446, n37447, n37448,
         n37449, n37450, n37451, n37452, n37453, n37454, n37455, n37456,
         n37457, n37458, n37459, n37460, n37461, n37462, n37463, n37464,
         n37465, n37466, n37467, n37468, n37469, n37470, n37471, n37472,
         n37473, n37474, n37475, n37476, n37477, n37478, n37479, n37480,
         n37481, n37482, n37483, n37484, n37485, n37486, n37487, n37488,
         n37489, n37490, n37491, n37492, n37493, n37494, n37495, n37496,
         n37497, n37498, n37499, n37500, n37501, n37502, n37503, n37504,
         n37505, n37506, n37507, n37508, n37509, n37510, n37511, n37512,
         n37513, n37514, n37515, n37516, n37517, n37518, n37519, n37520,
         n37521, n37522, n37523, n37524, n37525, n37526, n37527, n37528,
         n37529, n37530, n37531, n37532, n37533, n37534, n37535, n37536,
         n37537, n37538, n37539, n37540, n37541, n37542, n37543, n37544,
         n37545, n37546, n37547, n37548, n37549, n37550, n37551, n37552,
         n37553, n37554, n37555, n37556, n37557, n37558, n37559, n37560,
         n37561, n37562, n37563, n37564, n37565, n37566, n37567, n37568,
         n37569, n37570, n37571, n37572, n37573, n37574, n37575, n37576,
         n37577, n37578, n37579, n37580, n37581, n37582, n37583, n37584,
         n37585, n37586, n37587, n37588, n37589, n37590, n37591, n37592,
         n37593, n37594, n37595, n37596, n37597, n37598, n37599, n37600,
         n37601, n37602, n37603, n37604, n37605, n37606, n37607, n37608,
         n37609, n37610, n37611, n37612, n37613, n37614, n37615, n37616,
         n37617, n37618, n37619, n37620, n37621, n37622, n37623, n37624,
         n37625, n37626, n37627, n37628, n37629, n37630, n37631, n37632,
         n37633, n37634, n37635, n37636, n37637, n37638, n37639, n37640,
         n37641, n37642, n37643, n37644, n37645, n37646, n37647, n37648,
         n37649, n37650, n37651, n37652, n37653, n37654, n37655, n37656,
         n37657, n37658, n37659, n37660, n37661, n37662, n37663, n37664,
         n37665, n37666, n37667, n37668, n37669, n37670, n37671, n37672,
         n37673, n37674, n37675, n37676, n37677, n37678, n37679, n37680,
         n37681, n37682, n37683, n37684, n37685, n37686, n37687, n37688,
         n37689, n37690, n37691, n37692, n37693, n37694, n37695, n37696,
         n37697, n37698, n37699, n37700, n37701, n37702, n37703, n37704,
         n37705, n37706, n37707, n37708, n37709, n37710, n37711, n37712,
         n37713, n37714, n37715, n37716, n37717, n37718, n37719, n37720,
         n37721, n37722, n37723, n37724, n37725, n37726, n37727, n37728,
         n37729, n37730, n37731, n37732, n37733, n37734, n37735, n37736,
         n37737, n37738, n37739, n37740, n37741, n37742, n37743, n37744,
         n37745, n37746, n37747, n37748, n37749, n37750, n37751, n37752,
         n37753, n37754, n37755, n37756, n37757, n37758, n37759, n37760,
         n37761, n37762, n37763, n37764, n37765, n37766, n37767, n37768,
         n37769, n37770, n37771, n37772, n37773, n37774, n37775, n37776,
         n37777, n37778, n37779, n37780, n37781, n37782, n37783, n37784,
         n37785, n37786, n37787, n37788, n37789, n37790, n37791, n37792,
         n37793, n37794, n37795, n37796, n37797, n37798, n37799, n37800,
         n37801, n37802, n37803, n37804, n37805, n37806, n37807, n37808,
         n37809, n37810, n37811, n37812, n37813, n37814, n37815, n37816,
         n37817, n37818, n37819, n37820, n37821, n37822, n37823, n37824,
         n37825, n37826, n37827, n37828, n37829, n37830, n37831, n37832,
         n37833, n37834, n37835, n37836, n37837, n37838, n37839, n37840,
         n37841, n37842, n37843, n37844, n37845, n37846, n37847, n37848,
         n37849, n37850, n37851, n37852, n37853, n37854, n37855, n37856,
         n37857, n37858, n37859, n37860, n37861, n37862, n37863, n37864,
         n37865, n37866, n37867, n37868, n37869, n37870, n37871, n37872,
         n37873, n37874, n37875, n37876, n37877, n37878, n37879, n37880,
         n37881, n37882, n37883, n37884, n37885, n37886, n37887, n37888,
         n37889, n37890, n37891, n37892, n37893, n37894, n37895, n37896,
         n37897, n37898, n37899, n37900, n37901, n37902, n37903, n37904,
         n37905, n37906, n37907, n37908, n37909, n37910, n37911, n37912,
         n37913, n37914, n37915, n37916, n37917, n37918, n37919, n37920,
         n37921, n37922, n37923, n37924, n37925, n37926, n37927, n37928,
         n37929, n37930, n37931, n37932, n37933, n37934, n37935, n37936,
         n37937, n37938, n37939, n37940, n37941, n37942, n37943, n37944,
         n37945, n37946, n37947, n37948, n37949, n37950, n37951, n37952,
         n37953, n37954, n37955, n37956, n37957, n37958, n37959, n37960,
         n37961, n37962, n37963, n37964, n37965, n37966, n37967, n37968,
         n37969, n37970, n37971, n37972, n37973, n37974, n37975, n37976,
         n37977, n37978, n37979, n37980, n37981, n37982, n37983, n37984,
         n37985, n37986, n37987, n37988, n37989, n37990, n37991, n37992,
         n37993, n37994, n37995, n37996, n37997, n37998, n37999, n38000,
         n38001, n38002, n38003, n38004, n38005, n38006, n38007, n38008,
         n38009, n38010, n38011, n38012, n38013, n38014, n38015, n38016,
         n38017, n38018, n38019, n38020, n38021, n38022, n38023, n38024,
         n38025, n38026, n38027, n38028, n38029, n38030, n38031, n38032,
         n38033, n38034, n38035, n38036, n38037, n38038, n38039, n38040,
         n38041, n38042, n38043, n38044, n38045, n38046, n38047, n38048,
         n38049, n38050, n38051, n38052, n38053, n38054, n38055, n38056,
         n38057, n38058, n38059, n38060, n38061, n38062, n38063, n38064,
         n38065, n38066, n38067, n38068, n38069, n38070, n38071, n38072,
         n38073, n38074, n38075, n38076, n38077, n38078, n38079, n38080,
         n38081, n38082, n38083, n38084, n38085, n38086, n38087, n38088,
         n38089, n38090, n38091, n38092, n38093, n38094, n38095, n38096,
         n38097, n38098, n38099, n38100, n38101, n38102, n38103, n38104,
         n38105, n38106, n38107, n38108, n38109, n38110, n38111, n38112,
         n38113, n38114, n38115, n38116, n38117, n38118, n38119, n38120,
         n38121, n38122, n38123, n38124, n38125, n38126, n38127, n38128,
         n38129, n38130, n38131, n38132, n38133, n38134, n38135, n38136,
         n38137, n38138, n38139, n38140, n38141, n38142, n38143, n38144,
         n38145, n38146, n38147, n38148, n38149, n38150, n38151, n38152,
         n38153, n38154, n38155, n38156, n38157, n38158, n38159, n38160,
         n38161, n38162, n38163, n38164, n38165, n38166, n38167, n38168,
         n38169, n38170, n38171, n38172, n38173, n38174, n38175, n38176,
         n38177, n38178, n38179, n38180, n38181, n38182, n38183, n38184,
         n38185, n38186, n38187, n38188, n38189, n38190, n38191, n38192,
         n38193, n38194, n38195, n38196, n38197, n38198, n38199, n38200,
         n38201, n38202, n38203, n38204, n38205, n38206, n38207, n38208,
         n38209, n38210, n38211, n38212, n38213, n38214, n38215, n38216,
         n38217, n38218, n38219, n38220, n38221, n38222, n38223, n38224,
         n38225, n38226, n38227, n38228, n38229, n38230, n38231, n38232,
         n38233, n38234, n38235, n38236, n38237, n38238, n38239, n38240,
         n38241, n38242, n38243, n38244, n38245, n38246, n38247, n38248,
         n38249, n38250, n38251, n38252, n38253, n38254, n38255, n38256,
         n38257, n38258, n38259, n38260, n38261, n38262, n38263, n38264,
         n38265, n38266, n38267, n38268, n38269, n38270, n38271, n38272,
         n38273, n38274, n38275, n38276, n38277, n38278, n38279, n38280,
         n38281, n38282, n38283, n38284, n38285, n38286, n38287, n38288,
         n38289, n38290, n38291, n38292, n38293, n38294, n38295, n38296,
         n38297, n38298, n38299, n38300, n38301, n38302, n38303, n38304,
         n38305, n38306, n38307, n38308, n38309, n38310, n38311, n38312,
         n38313, n38314, n38315, n38316, n38317, n38318, n38319, n38320,
         n38321, n38322, n38323, n38324, n38325, n38326, n38327, n38328,
         n38329, n38330, n38331, n38332, n38333, n38334, n38335, n38336,
         n38337, n38338, n38339, n38340, n38341, n38342, n38343, n38344,
         n38345, n38346, n38347, n38348, n38349, n38350, n38351, n38352,
         n38353, n38354, n38355, n38356, n38357, n38358, n38359, n38360,
         n38361, n38362, n38363, n38364, n38365, n38366, n38367, n38368,
         n38369, n38370, n38371, n38372, n38373, n38374, n38375, n38376,
         n38377, n38378, n38379, n38380, n38381, n38382, n38383, n38384,
         n38385, n38386, n38387, n38388, n38389, n38390, n38391, n38392,
         n38393, n38394, n38395, n38396, n38397, n38398, n38399, n38400,
         n38401, n38402, n38403, n38404, n38405, n38406, n38407, n38408,
         n38409, n38410, n38411, n38412, n38413, n38414, n38415, n38416,
         n38417, n38418, n38419, n38420, n38421, n38422, n38423, n38424,
         n38425, n38426, n38427, n38428, n38429, n38430, n38431, n38432,
         n38433, n38434, n38435, n38436, n38437, n38438, n38439, n38440,
         n38441, n38442, n38443, n38444, n38445, n38446, n38447, n38448,
         n38449, n38450, n38451, n38452, n38453, n38454, n38455, n38456,
         n38457, n38458, n38459, n38460, n38461, n38462, n38463, n38464,
         n38465, n38466, n38467, n38468, n38469, n38470, n38471, n38472,
         n38473, n38474, n38475, n38476, n38477, n38478, n38479, n38480,
         n38481, n38482, n38483, n38484, n38485, n38486, n38487, n38488,
         n38489, n38490, n38491, n38492, n38493, n38494, n38495, n38496,
         n38497, n38498, n38499, n38500, n38501, n38502, n38503, n38504,
         n38505, n38506, n38507, n38508, n38509, n38510, n38511, n38512,
         n38513, n38514, n38515, n38516, n38517, n38518, n38519, n38520,
         n38521, n38522, n38523, n38524, n38525, n38526, n38527, n38528,
         n38529, n38530, n38531, n38532, n38533, n38534, n38535, n38536,
         n38537, n38538, n38539, n38540, n38541, n38542, n38543, n38544,
         n38545, n38546, n38547, n38548, n38549, n38550, n38551, n38552,
         n38553, n38554, n38555, n38556, n38557, n38558, n38559, n38560,
         n38561, n38562, n38563, n38564, n38565, n38566, n38567, n38568,
         n38569, n38570, n38571, n38572, n38573, n38574, n38575, n38576,
         n38577, n38578, n38579, n38580, n38581, n38582, n38583, n38584,
         n38585, n38586, n38587, n38588, n38589, n38590, n38591, n38592,
         n38593, n38594, n38595, n38596, n38597, n38598, n38599, n38600,
         n38601, n38602, n38603, n38604, n38605, n38606, n38607, n38608,
         n38609, n38610, n38611, n38612, n38613, n38614, n38615, n38616,
         n38617, n38618, n38619, n38620, n38621, n38622, n38623, n38624,
         n38625, n38626, n38627, n38628, n38629, n38630, n38631, n38632,
         n38633, n38634, n38635, n38636, n38637, n38638, n38639, n38640,
         n38641, n38642, n38643, n38644, n38645, n38646, n38647, n38648,
         n38649, n38650, n38651, n38652, n38653, n38654, n38655, n38656,
         n38657, n38658, n38659, n38660, n38661, n38662, n38663, n38664,
         n38665, n38666, n38667, n38668, n38669, n38670, n38671, n38672,
         n38673, n38674, n38675, n38676, n38677, n38678, n38679, n38680,
         n38681, n38682, n38683, n38684, n38685, n38686, n38687, n38688,
         n38689, n38690, n38691, n38692, n38693, n38694, n38695, n38696,
         n38697, n38698, n38699, n38700, n38701, n38702, n38703, n38704,
         n38705, n38706, n38707, n38708, n38709, n38710, n38711, n38712,
         n38713, n38714, n38715, n38716, n38717, n38718, n38719, n38720,
         n38721, n38722, n38723, n38724, n38725, n38726, n38727, n38728,
         n38729, n38730, n38731, n38732, n38733, n38734, n38735, n38736,
         n38737, n38738, n38739, n38740, n38741, n38742, n38743, n38744,
         n38745, n38746, n38747, n38748, n38749, n38750, n38751, n38752,
         n38753, n38754, n38755, n38756, n38757, n38758, n38759, n38760,
         n38761, n38762, n38763, n38764, n38765, n38766, n38767, n38768,
         n38769, n38770, n38771, n38772, n38773, n38774, n38775, n38776,
         n38777, n38778, n38779, n38780, n38781, n38782, n38783, n38784,
         n38785, n38786, n38787, n38788, n38789, n38790, n38791, n38792,
         n38793, n38794, n38795, n38796, n38797, n38798, n38799, n38800,
         n38801, n38802, n38803, n38804, n38805, n38806, n38807, n38808,
         n38809, n38810, n38811, n38812, n38813, n38814, n38815, n38816,
         n38817, n38818, n38819, n38820, n38821, n38822, n38823, n38824,
         n38825, n38826, n38827, n38828, n38829, n38830, n38831, n38832,
         n38833, n38834, n38835, n38836, n38837, n38838, n38839, n38840,
         n38841, n38842, n38843, n38844, n38845, n38846, n38847, n38848,
         n38849, n38850, n38851, n38852, n38853, n38854, n38855, n38856,
         n38857, n38858, n38859, n38860, n38861, n38862, n38863, n38864,
         n38865, n38866, n38867, n38868, n38869, n38870, n38871, n38872,
         n38873, n38874, n38875, n38876, n38877, n38878, n38879, n38880,
         n38881, n38882, n38883, n38884, n38885, n38886, n38887, n38888,
         n38889, n38890, n38891, n38892, n38893, n38894, n38895, n38896,
         n38897, n38898, n38899, n38900, n38901, n38902, n38903, n38904,
         n38905, n38906, n38907, n38908, n38909, n38910, n38911, n38912,
         n38913, n38914, n38915, n38916, n38917, n38918, n38919, n38920,
         n38921, n38922, n38923, n38924, n38925, n38926, n38927, n38928,
         n38929, n38930, n38931, n38932, n38933, n38934, n38935, n38936,
         n38937, n38938, n38939, n38940, n38941, n38942, n38943, n38944,
         n38945, n38946, n38947, n38948, n38949, n38950, n38951, n38952,
         n38953, n38954, n38955, n38956, n38957, n38958, n38959, n38960,
         n38961, n38962, n38963, n38964, n38965, n38966, n38967, n38968,
         n38969, n38970, n38971, n38972, n38973, n38974, n38975, n38976,
         n38977, n38978, n38979, n38980, n38981, n38982, n38983, n38984,
         n38985, n38986, n38987, n38988, n38989, n38990, n38991, n38992,
         n38993, n38994, n38995, n38996, n38997, n38998, n38999, n39000,
         n39001, n39002, n39003, n39004, n39005, n39006, n39007, n39008,
         n39009, n39010, n39011, n39012, n39013, n39014, n39015, n39016,
         n39017, n39018, n39019, n39020, n39021, n39022, n39023, n39024,
         n39025, n39026, n39027, n39028, n39029, n39030, n39031, n39032,
         n39033, n39034, n39035, n39036, n39037, n39038, n39039, n39040,
         n39041, n39042, n39043, n39044, n39045, n39046, n39047, n39048,
         n39049, n39050, n39051, n39052, n39053, n39054, n39055, n39056,
         n39057, n39058, n39059, n39060, n39061, n39062, n39063, n39064,
         n39065, n39066, n39067, n39068, n39069, n39070, n39071, n39072,
         n39073, n39074, n39075, n39076, n39077, n39078, n39079, n39080,
         n39081, n39082, n39083, n39084, n39085, n39086, n39087, n39088,
         n39089, n39090, n39091, n39092, n39093, n39094, n39095, n39096,
         n39097, n39098, n39099, n39100, n39101, n39102, n39103, n39104,
         n39105, n39106, n39107, n39108, n39109, n39110, n39111, n39112,
         n39113, n39114, n39115, n39116, n39117, n39118, n39119, n39120,
         n39121, n39122, n39123, n39124, n39125, n39126, n39127, n39128,
         n39129, n39130, n39131, n39132, n39133, n39134, n39135, n39136,
         n39137, n39138, n39139, n39140, n39141, n39142, n39143, n39144,
         n39145, n39146, n39147, n39148, n39149, n39150, n39151, n39152,
         n39153, n39154, n39155, n39156, n39157, n39158, n39159, n39160,
         n39161, n39162, n39163, n39164, n39165, n39166, n39167, n39168,
         n39169, n39170, n39171, n39172, n39173, n39174, n39175, n39176,
         n39177, n39178, n39179, n39180, n39181, n39182, n39183, n39184,
         n39185, n39186, n39187, n39188, n39189, n39190, n39191, n39192,
         n39193, n39194, n39195, n39196, n39197, n39198, n39199, n39200,
         n39201, n39202, n39203, n39204, n39205, n39206, n39207, n39208,
         n39209, n39210, n39211, n39212, n39213, n39214, n39215, n39216,
         n39217, n39218, n39219, n39220, n39221, n39222, n39223, n39224,
         n39225, n39226, n39227, n39228, n39229, n39230, n39231, n39232,
         n39233, n39234, n39235, n39236, n39237, n39238, n39239, n39240,
         n39241, n39242, n39243, n39244, n39245, n39246, n39247, n39248,
         n39249, n39250, n39251, n39252, n39253, n39254, n39255, n39256,
         n39257, n39258, n39259, n39260, n39261, n39262, n39263, n39264,
         n39265, n39266, n39267, n39268, n39269, n39270, n39271, n39272,
         n39273, n39274, n39275, n39276, n39277, n39278, n39279, n39280,
         n39281, n39282, n39283, n39284, n39285, n39286, n39287, n39288,
         n39289, n39290, n39291, n39292, n39293, n39294, n39295, n39296,
         n39297, n39298, n39299, n39300, n39301, n39302, n39303, n39304,
         n39305, n39306, n39307, n39308, n39309, n39310, n39311, n39312,
         n39313, n39314, n39315, n39316, n39317, n39318, n39319, n39320,
         n39321, n39322, n39323, n39324, n39325, n39326, n39327, n39328,
         n39329, n39330, n39331, n39332, n39333, n39334, n39335, n39336,
         n39337, n39338, n39339, n39340, n39341, n39342, n39343, n39344,
         n39345, n39346, n39347, n39348, n39349, n39350, n39351, n39352,
         n39353, n39354, n39355, n39356, n39357, n39358, n39359, n39360,
         n39361, n39362, n39363, n39364, n39365, n39366, n39367, n39368,
         n39369, n39370, n39371, n39372, n39373, n39374, n39375, n39376,
         n39377, n39378, n39379, n39380, n39381, n39382, n39383, n39384,
         n39385, n39386, n39387, n39388, n39389, n39390, n39391, n39392,
         n39393, n39394, n39395, n39396, n39397, n39398, n39399, n39400,
         n39401, n39402, n39403, n39404, n39405, n39406, n39407, n39408,
         n39409, n39410, n39411, n39412, n39413, n39414, n39415, n39416,
         n39417, n39418, n39419, n39420, n39421, n39422, n39423, n39424,
         n39425, n39426, n39427, n39428, n39429, n39430, n39431, n39432,
         n39433, n39434, n39435, n39436, n39437, n39438, n39439, n39440,
         n39441, n39442, n39443, n39444, n39445, n39446, n39447, n39448,
         n39449, n39450, n39451, n39452, n39453, n39454, n39455, n39456,
         n39457, n39458, n39459, n39460, n39461, n39462, n39463, n39464,
         n39465, n39466, n39467, n39468, n39469, n39470, n39471, n39472,
         n39473, n39474, n39475, n39476, n39477, n39478, n39479, n39480,
         n39481, n39482, n39483, n39484, n39485, n39486, n39487, n39488,
         n39489, n39490, n39491, n39492, n39493, n39494, n39495, n39496,
         n39497, n39498, n39499, n39500, n39501, n39502, n39503, n39504,
         n39505, n39506, n39507, n39508, n39509, n39510, n39511, n39512,
         n39513, n39514, n39515, n39516, n39517, n39518, n39519, n39520,
         n39521, n39522, n39523, n39524, n39525, n39526, n39527, n39528,
         n39529, n39530, n39531, n39532, n39533, n39534, n39535, n39536,
         n39537, n39538, n39539, n39540, n39541, n39542, n39543, n39544,
         n39545, n39546, n39547, n39548, n39549, n39550, n39551, n39552,
         n39553, n39554, n39555, n39556, n39557, n39558, n39559, n39560,
         n39561, n39562, n39563, n39564, n39565, n39566, n39567, n39568,
         n39569, n39570, n39571, n39572, n39573, n39574, n39575, n39576,
         n39577, n39578, n39579, n39580, n39581, n39582, n39583, n39584,
         n39585, n39586, n39587, n39588, n39589, n39590, n39591, n39592,
         n39593, n39594, n39595, n39596, n39597, n39598, n39599, n39600,
         n39601, n39602, n39603, n39604, n39605, n39606, n39607, n39608,
         n39609, n39610, n39611, n39612, n39613, n39614, n39615, n39616,
         n39617, n39618, n39619, n39620, n39621, n39622, n39623, n39624,
         n39625, n39626, n39627, n39628, n39629, n39630, n39631, n39632,
         n39633, n39634, n39635, n39636, n39637, n39638, n39639, n39640,
         n39641, n39642, n39643, n39644, n39645, n39646, n39647, n39648,
         n39649, n39650, n39651, n39652, n39653, n39654, n39655, n39656,
         n39657, n39658, n39659, n39660, n39661, n39662, n39663, n39664,
         n39665, n39666, n39667, n39668, n39669, n39670, n39671, n39672,
         n39673, n39674, n39675, n39676, n39677, n39678, n39679, n39680,
         n39681, n39682, n39683, n39684, n39685, n39686, n39687, n39688,
         n39689, n39690, n39691, n39692, n39693, n39694, n39695, n39696,
         n39697, n39698, n39699, n39700, n39701, n39702, n39703, n39704,
         n39705, n39706, n39707, n39708, n39709, n39710, n39711, n39712,
         n39713, n39714, n39715, n39716, n39717, n39718, n39719, n39720,
         n39721, n39722, n39723, n39724, n39725, n39726, n39727, n39728,
         n39729, n39730, n39731, n39732, n39733, n39734, n39735, n39736,
         n39737, n39738, n39739, n39740, n39741, n39742, n39743, n39744,
         n39745, n39746, n39747, n39748, n39749, n39750, n39751, n39752,
         n39753, n39754, n39755, n39756, n39757, n39758, n39759, n39760,
         n39761, n39762, n39763, n39764, n39765, n39766, n39767, n39768,
         n39769, n39770, n39771, n39772, n39773, n39774, n39775, n39776,
         n39777, n39778, n39779, n39780, n39781, n39782, n39783, n39784,
         n39785, n39786, n39787, n39788, n39789, n39790, n39791, n39792,
         n39793, n39794, n39795, n39796, n39797, n39798, n39799, n39800,
         n39801, n39802, n39803, n39804, n39805, n39806, n39807, n39808,
         n39809, n39810, n39811, n39812, n39813, n39814, n39815, n39816,
         n39817, n39818, n39819, n39820, n39821, n39822, n39823, n39824,
         n39825, n39826, n39827, n39828, n39829, n39830, n39831, n39832,
         n39833, n39834, n39835, n39836, n39837, n39838, n39839, n39840,
         n39841, n39842, n39843, n39844, n39845, n39846, n39847, n39848,
         n39849, n39850, n39851, n39852, n39853, n39854, n39855, n39856,
         n39857, n39858, n39859, n39860, n39861, n39862, n39863, n39864,
         n39865, n39866, n39867, n39868, n39869, n39870, n39871, n39872,
         n39873, n39874, n39875, n39876, n39877, n39878, n39879, n39880,
         n39881, n39882, n39883, n39884, n39885, n39886, n39887, n39888,
         n39889, n39890, n39891, n39892, n39893, n39894, n39895, n39896,
         n39897, n39898, n39899, n39900, n39901, n39902, n39903, n39904,
         n39905, n39906, n39907, n39908, n39909, n39910, n39911, n39912,
         n39913, n39914, n39915, n39916, n39917, n39918, n39919, n39920,
         n39921, n39922, n39923, n39924, n39925, n39926, n39927, n39928,
         n39929, n39930, n39931, n39932, n39933, n39934, n39935, n39936,
         n39937, n39938, n39939, n39940, n39941, n39942, n39943, n39944,
         n39945, n39946, n39947, n39948, n39949, n39950, n39951, n39952,
         n39953, n39954, n39955, n39956, n39957, n39958, n39959, n39960,
         n39961, n39962, n39963, n39964, n39965, n39966, n39967, n39968,
         n39969, n39970, n39971, n39972, n39973, n39974, n39975, n39976,
         n39977, n39978, n39979, n39980, n39981, n39982, n39983, n39984,
         n39985, n39986, n39987, n39988, n39989, n39990, n39991, n39992,
         n39993, n39994, n39995, n39996, n39997, n39998, n39999, n40000,
         n40001, n40002, n40003, n40004, n40005, n40006, n40007, n40008,
         n40009, n40010, n40011, n40012, n40013, n40014, n40015, n40016,
         n40017, n40018, n40019, n40020, n40021, n40022, n40023, n40024,
         n40025, n40026, n40027, n40028, n40029, n40030, n40031, n40032,
         n40033, n40034, n40035, n40036, n40037, n40038, n40039, n40040,
         n40041, n40042, n40043, n40044, n40045, n40046, n40047, n40048,
         n40049, n40050, n40051, n40052, n40053, n40054, n40055, n40056,
         n40057, n40058, n40059, n40060, n40061, n40062, n40063, n40064,
         n40065, n40066, n40067, n40068, n40069, n40070, n40071, n40072,
         n40073, n40074, n40075, n40076, n40077, n40078, n40079, n40080,
         n40081, n40082, n40083, n40084, n40085, n40086, n40087, n40088,
         n40089, n40090, n40091, n40092, n40093, n40094, n40095, n40096,
         n40097, n40098, n40099, n40100, n40101, n40102, n40103, n40104,
         n40105, n40106, n40107, n40108, n40109, n40110, n40111, n40112,
         n40113, n40114, n40115, n40116, n40117, n40118, n40119, n40120,
         n40121, n40122, n40123, n40124, n40125, n40126, n40127, n40128,
         n40129, n40130, n40131, n40132, n40133, n40134, n40135, n40136,
         n40137, n40138, n40139, n40140, n40141, n40142, n40143, n40144,
         n40145, n40146, n40147, n40148, n40149, n40150, n40151, n40152,
         n40153, n40154, n40155, n40156, n40157, n40158, n40159, n40160,
         n40161, n40162, n40163, n40164, n40165, n40166, n40167, n40168,
         n40169, n40170, n40171, n40172, n40173, n40174, n40175, n40176,
         n40177, n40178, n40179, n40180, n40181, n40182, n40183, n40184,
         n40185, n40186, n40187, n40188, n40189, n40190, n40191, n40192,
         n40193, n40194, n40195, n40196, n40197, n40198, n40199, n40200,
         n40201, n40202, n40203, n40204, n40205, n40206, n40207, n40208,
         n40209, n40210, n40211, n40212, n40213, n40214, n40215, n40216,
         n40217, n40218, n40219, n40220, n40221, n40222, n40223, n40224,
         n40225, n40226, n40227, n40228, n40229, n40230, n40231, n40232,
         n40233, n40234, n40235, n40236, n40237, n40238, n40239, n40240,
         n40241, n40242, n40243, n40244, n40245, n40246, n40247, n40248,
         n40249, n40250, n40251, n40252, n40253, n40254, n40255, n40256,
         n40257, n40258, n40259, n40260, n40261, n40262, n40263, n40264,
         n40265, n40266, n40267, n40268, n40269, n40270, n40271, n40272,
         n40273, n40274, n40275, n40276, n40277, n40278, n40279, n40280,
         n40281, n40282, n40283, n40284, n40285, n40286, n40287, n40288,
         n40289, n40290, n40291, n40292, n40293, n40294, n40295, n40296,
         n40297, n40298, n40299, n40300, n40301, n40302, n40303, n40304,
         n40305, n40306, n40307, n40308, n40309, n40310, n40311, n40312,
         n40313, n40314, n40315, n40316, n40317, n40318, n40319, n40320,
         n40321, n40322, n40323, n40324, n40325, n40326, n40327, n40328,
         n40329, n40330, n40331, n40332, n40333, n40334, n40335, n40336,
         n40337, n40338, n40339, n40340, n40341, n40342, n40343, n40344,
         n40345, n40346, n40347, n40348, n40349, n40350, n40351, n40352,
         n40353, n40354, n40355, n40356, n40357, n40358, n40359, n40360,
         n40361, n40362, n40363, n40364, n40365, n40366, n40367, n40368,
         n40369, n40370, n40371, n40372, n40373, n40374, n40375, n40376,
         n40377, n40378, n40379, n40380, n40381, n40382, n40383, n40384,
         n40385, n40386, n40387, n40388, n40389, n40390, n40391, n40392,
         n40393, n40394, n40395, n40396, n40397, n40398, n40399, n40400,
         n40401, n40402, n40403, n40404, n40405, n40406, n40407, n40408,
         n40409, n40410, n40411, n40412, n40413, n40414, n40415, n40416,
         n40417, n40418, n40419, n40420, n40421, n40422, n40423, n40424,
         n40425, n40426, n40427, n40428, n40429, n40430, n40431, n40432,
         n40433, n40434, n40435, n40436, n40437, n40438, n40439, n40440,
         n40441, n40442, n40443, n40444, n40445, n40446, n40447, n40448,
         n40449, n40450, n40451, n40452, n40453, n40454, n40455, n40456,
         n40457, n40458, n40459, n40460, n40461, n40462, n40463, n40464,
         n40465, n40466, n40467, n40468, n40469, n40470, n40471, n40472,
         n40473, n40474, n40475, n40476, n40477, n40478, n40479, n40480,
         n40481, n40482, n40483, n40484, n40485, n40486, n40487, n40488,
         n40489, n40490, n40491, n40492, n40493, n40494, n40495, n40496,
         n40497, n40498, n40499, n40500, n40501, n40502, n40503, n40504,
         n40505, n40506, n40507, n40508, n40509, n40510, n40511, n40512,
         n40513, n40514, n40515, n40516, n40517, n40518, n40519, n40520,
         n40521, n40522, n40523, n40524, n40525, n40526, n40527, n40528,
         n40529, n40530, n40531, n40532, n40533, n40534, n40535, n40536,
         n40537, n40538, n40539, n40540, n40541, n40542, n40543, n40544,
         n40545, n40546, n40547, n40548, n40549, n40550, n40551, n40552,
         n40553, n40554, n40555, n40556, n40557, n40558, n40559, n40560,
         n40561, n40562, n40563, n40564, n40565, n40566, n40567, n40568,
         n40569, n40570, n40571, n40572, n40573, n40574, n40575, n40576,
         n40577, n40578, n40579, n40580, n40581, n40582, n40583, n40584,
         n40585, n40586, n40587, n40588, n40589, n40590, n40591, n40592,
         n40593, n40594, n40595, n40596, n40597, n40598, n40599, n40600,
         n40601, n40602, n40603, n40604, n40605, n40606, n40607, n40608,
         n40609, n40610, n40611, n40612, n40613, n40614, n40615, n40616,
         n40617, n40618, n40619, n40620, n40621, n40622, n40623, n40624,
         n40625, n40626, n40627, n40628, n40629, n40630, n40631, n40632,
         n40633, n40634, n40635, n40636, n40637, n40638, n40639, n40640,
         n40641, n40642, n40643, n40644, n40645, n40646, n40647, n40648,
         n40649, n40650, n40651, n40652, n40653, n40654, n40655, n40656,
         n40657, n40658, n40659, n40660, n40661, n40662, n40663, n40664,
         n40665, n40666, n40667, n40668, n40669, n40670, n40671, n40672,
         n40673, n40674, n40675, n40676, n40677, n40678, n40679, n40680,
         n40681, n40682, n40683, n40684, n40685, n40686, n40687, n40688,
         n40689, n40690, n40691, n40692, n40693, n40694, n40695, n40696,
         n40697, n40698, n40699, n40700, n40701, n40702, n40703, n40704,
         n40705, n40706, n40707, n40708, n40709, n40710, n40711, n40712,
         n40713, n40714, n40715, n40716, n40717, n40718, n40719, n40720,
         n40721, n40722, n40723, n40724, n40725, n40726, n40727, n40728,
         n40729, n40730, n40731, n40732, n40733, n40734, n40735, n40736,
         n40737, n40738, n40739, n40740, n40741, n40742, n40743, n40744,
         n40745, n40746, n40747, n40748, n40749, n40750, n40751, n40752,
         n40753, n40754, n40755, n40756, n40757, n40758, n40759, n40760,
         n40761, n40762, n40763, n40764, n40765, n40766, n40767, n40768,
         n40769, n40770, n40771, n40772, n40773, n40774, n40775, n40776,
         n40777, n40778, n40779, n40780, n40781, n40782, n40783, n40784,
         n40785, n40786, n40787, n40788, n40789, n40790, n40791, n40792,
         n40793, n40794, n40795, n40796, n40797, n40798, n40799, n40800,
         n40801, n40802, n40803, n40804, n40805, n40806, n40807, n40808,
         n40809, n40810, n40811, n40812, n40813, n40814, n40815, n40816,
         n40817, n40818, n40819, n40820, n40821, n40822, n40823, n40824,
         n40825, n40826, n40827, n40828, n40829, n40830, n40831, n40832,
         n40833, n40834, n40835, n40836, n40837, n40838, n40839, n40840,
         n40841, n40842, n40843, n40844, n40845, n40846, n40847, n40848,
         n40849, n40850, n40851, n40852, n40853, n40854, n40855, n40856,
         n40857, n40858, n40859, n40860, n40861, n40862, n40863, n40864,
         n40865, n40866, n40867, n40868, n40869, n40870, n40871, n40872,
         n40873, n40874, n40875, n40876, n40877, n40878, n40879, n40880,
         n40881, n40882, n40883, n40884, n40885, n40886, n40887, n40888,
         n40889, n40890, n40891, n40892, n40893, n40894, n40895, n40896,
         n40897, n40898, n40899, n40900, n40901, n40902, n40903, n40904,
         n40905, n40906, n40907, n40908, n40909, n40910, n40911, n40912,
         n40913, n40914, n40915, n40916, n40917, n40918, n40919, n40920,
         n40921, n40922, n40923, n40924, n40925, n40926, n40927, n40928,
         n40929, n40930, n40931, n40932, n40933, n40934, n40935, n40936,
         n40937, n40938, n40939, n40940, n40941, n40942, n40943, n40944,
         n40945, n40946, n40947, n40948, n40949, n40950, n40951, n40952,
         n40953, n40954, n40955, n40956, n40957, n40958, n40959, n40960,
         n40961, n40962, n40963, n40964, n40965, n40966, n40967, n40968,
         n40969, n40970, n40971, n40972, n40973, n40974, n40975, n40976,
         n40977, n40978, n40979, n40980, n40981, n40982, n40983, n40984,
         n40985, n40986, n40987, n40988, n40989, n40990, n40991, n40992,
         n40993, n40994, n40995, n40996, n40997, n40998, n40999, n41000,
         n41001, n41002, n41003, n41004, n41005, n41006, n41007, n41008,
         n41009, n41010, n41011, n41012, n41013, n41014, n41015, n41016,
         n41017, n41018, n41019, n41020, n41021, n41022, n41023, n41024,
         n41025, n41026, n41027, n41028, n41029, n41030, n41031, n41032,
         n41033, n41034, n41035, n41036, n41037, n41038, n41039, n41040,
         n41041, n41042, n41043, n41044, n41045, n41046, n41047, n41048,
         n41049, n41050, n41051, n41052, n41053, n41054, n41055, n41056,
         n41057, n41058, n41059, n41060, n41061, n41062, n41063, n41064,
         n41065, n41066, n41067, n41068, n41069, n41070, n41071, n41072,
         n41073, n41074, n41075, n41076, n41077, n41078, n41079, n41080,
         n41081, n41082, n41083, n41084, n41085, n41086, n41087, n41088,
         n41089, n41090, n41091, n41092, n41093, n41094, n41095, n41096,
         n41097, n41098, n41099, n41100, n41101, n41102, n41103, n41104,
         n41105, n41106, n41107, n41108, n41109, n41110, n41111, n41112,
         n41113, n41114, n41115, n41116, n41117, n41118, n41119, n41120,
         n41121, n41122, n41123, n41124, n41125, n41126, n41127, n41128,
         n41129, n41130, n41131, n41132, n41133, n41134, n41135, n41136,
         n41137, n41138, n41139, n41140, n41141, n41142, n41143, n41144,
         n41145, n41146, n41147, n41148, n41149, n41150, n41151, n41152,
         n41153, n41154, n41155, n41156, n41157, n41158, n41159, n41160,
         n41161, n41162, n41163, n41164, n41165, n41166, n41167, n41168,
         n41169, n41170, n41171, n41172, n41173, n41174, n41175, n41176,
         n41177, n41178, n41179, n41180, n41181, n41182, n41183, n41184,
         n41185, n41186, n41187, n41188, n41189, n41190, n41191, n41192,
         n41193, n41194, n41195, n41196, n41197, n41198, n41199, n41200,
         n41201, n41202, n41203, n41204, n41205, n41206, n41207, n41208,
         n41209, n41210, n41211, n41212, n41213, n41214, n41215, n41216,
         n41217, n41218, n41219, n41220, n41221, n41222, n41223, n41224,
         n41225, n41226, n41227, n41228, n41229, n41230, n41231, n41232,
         n41233, n41234, n41235, n41236, n41237, n41238, n41239, n41240,
         n41241, n41242, n41243, n41244, n41245, n41246, n41247, n41248,
         n41249, n41250, n41251, n41252, n41253, n41254, n41255, n41256,
         n41257, n41258, n41259, n41260, n41261, n41262, n41263, n41264,
         n41265, n41266, n41267, n41268, n41269, n41270, n41271, n41272,
         n41273, n41274, n41275, n41276, n41277, n41278, n41279, n41280,
         n41281, n41282, n41283, n41284, n41285, n41286, n41287, n41288,
         n41289, n41290, n41291, n41292, n41293, n41294, n41295, n41296,
         n41297, n41298, n41299, n41300, n41301, n41302, n41303, n41304,
         n41305, n41306, n41307, n41308, n41309, n41310, n41311, n41312,
         n41313, n41314, n41315, n41316, n41317, n41318, n41319, n41320,
         n41321, n41322, n41323, n41324, n41325, n41326, n41327, n41328,
         n41329, n41330, n41331, n41332, n41333, n41334, n41335, n41336,
         n41337, n41338, n41339, n41340, n41341, n41342, n41343, n41344,
         n41345, n41346, n41347, n41348, n41349, n41350, n41351, n41352,
         n41353, n41354, n41355, n41356, n41357, n41358, n41359, n41360,
         n41361, n41362, n41363, n41364, n41365, n41366, n41367, n41368,
         n41369, n41370, n41371, n41372, n41373, n41374, n41375, n41376,
         n41377, n41378, n41379, n41380, n41381, n41382, n41383, n41384,
         n41385, n41386, n41387, n41388, n41389, n41390, n41391, n41392,
         n41393, n41394, n41395, n41396, n41397, n41398, n41399, n41400,
         n41401, n41402, n41403, n41404, n41405, n41406, n41407, n41408,
         n41409, n41410, n41411, n41412, n41413, n41414, n41415, n41416,
         n41417, n41418, n41419, n41420, n41421, n41422, n41423, n41424,
         n41425, n41426, n41427, n41428, n41429, n41430, n41431, n41432,
         n41433, n41434, n41435, n41436, n41437, n41438, n41439, n41440,
         n41441, n41442, n41443, n41444, n41445, n41446, n41447, n41448,
         n41449, n41450, n41451, n41452, n41453, n41454, n41455, n41456,
         n41457, n41458, n41459, n41460, n41461, n41462, n41463, n41464,
         n41465, n41466, n41467, n41468, n41469, n41470, n41471, n41472,
         n41473, n41474, n41475, n41476, n41477, n41478, n41479, n41480,
         n41481, n41482, n41483, n41484, n41485, n41486, n41487, n41488,
         n41489, n41490, n41491, n41492, n41493, n41494, n41495, n41496,
         n41497, n41498, n41499, n41500, n41501, n41502, n41503, n41504,
         n41505, n41506, n41507, n41508, n41509, n41510, n41511, n41512,
         n41513, n41514, n41515, n41516, n41517, n41518, n41519, n41520,
         n41521, n41522, n41523, n41524, n41525, n41526, n41527, n41528,
         n41529, n41530, n41531, n41532, n41533, n41534, n41535, n41536,
         n41537, n41538, n41539, n41540, n41541, n41542, n41543, n41544,
         n41545, n41546, n41547, n41548, n41549, n41550, n41551, n41552,
         n41553, n41554, n41555, n41556, n41557, n41558, n41559, n41560,
         n41561, n41562, n41563, n41564, n41565, n41566, n41567, n41568,
         n41569, n41570, n41571, n41572, n41573, n41574, n41575, n41576,
         n41577, n41578, n41579, n41580, n41581, n41582, n41583, n41584,
         n41585, n41586, n41587, n41588, n41589, n41590, n41591, n41592,
         n41593, n41594, n41595, n41596, n41597, n41598, n41599, n41600,
         n41601, n41602, n41603, n41604, n41605, n41606, n41607, n41608,
         n41609, n41610, n41611, n41612, n41613, n41614, n41615, n41616,
         n41617, n41618, n41619, n41620, n41621, n41622, n41623, n41624,
         n41625, n41626, n41627, n41628, n41629, n41630, n41631, n41632,
         n41633, n41634, n41635, n41636, n41637, n41638, n41639, n41640,
         n41641, n41642, n41643, n41644, n41645, n41646, n41647, n41648,
         n41649, n41650, n41651, n41652, n41653, n41654, n41655, n41656,
         n41657, n41658, n41659, n41660, n41661, n41662, n41663, n41664,
         n41665, n41666, n41667, n41668, n41669, n41670, n41671, n41672,
         n41673, n41674, n41675, n41676, n41677, n41678, n41679, n41680,
         n41681, n41682, n41683, n41684, n41685, n41686, n41687, n41688,
         n41689, n41690, n41691, n41692, n41693, n41694, n41695, n41696,
         n41697, n41698, n41699, n41700, n41701, n41702, n41703, n41704,
         n41705, n41706, n41707, n41708, n41709, n41710, n41711, n41712,
         n41713, n41714, n41715, n41716, n41717, n41718, n41719, n41720,
         n41721, n41722, n41723, n41724, n41725, n41726, n41727, n41728,
         n41729, n41730, n41731, n41732, n41733, n41734, n41735, n41736,
         n41737, n41738, n41739, n41740, n41741, n41742, n41743, n41744,
         n41745, n41746, n41747, n41748, n41749, n41750, n41751, n41752,
         n41753, n41754, n41755, n41756, n41757, n41758, n41759, n41760,
         n41761, n41762, n41763, n41764, n41765, n41766, n41767, n41768,
         n41769, n41770, n41771, n41772, n41773, n41774, n41775, n41776,
         n41777, n41778, n41779, n41780, n41781, n41782, n41783, n41784,
         n41785, n41786, n41787, n41788, n41789, n41790, n41791, n41792,
         n41793, n41794, n41795, n41796, n41797, n41798, n41799, n41800,
         n41801, n41802, n41803, n41804, n41805, n41806, n41807, n41808,
         n41809, n41810, n41811, n41812, n41813, n41814, n41815, n41816,
         n41817, n41818, n41819, n41820, n41821, n41822, n41823, n41824,
         n41825, n41826, n41827, n41828, n41829, n41830, n41831, n41832,
         n41833, n41834, n41835, n41836, n41837, n41838, n41839, n41840,
         n41841, n41842, n41843, n41844, n41845, n41846, n41847, n41848,
         n41849, n41850, n41851, n41852, n41853, n41854, n41855, n41856,
         n41857, n41858, n41859, n41860, n41861, n41862, n41863, n41864,
         n41865, n41866, n41867, n41868, n41869, n41870, n41871, n41872,
         n41873, n41874, n41875, n41876, n41877, n41878, n41879, n41880,
         n41881, n41882, n41883, n41884, n41885, n41886, n41887, n41888,
         n41889, n41890, n41891, n41892, n41893, n41894, n41895, n41896,
         n41897, n41898, n41899, n41900, n41901, n41902, n41903, n41904,
         n41905, n41906, n41907, n41908, n41909, n41910, n41911, n41912,
         n41913, n41914, n41915, n41916, n41917, n41918, n41919, n41920,
         n41921, n41922, n41923, n41924, n41925, n41926, n41927, n41928,
         n41929, n41930, n41931, n41932, n41933, n41934, n41935, n41936,
         n41937, n41938, n41939, n41940, n41941, n41942, n41943, n41944,
         n41945, n41946, n41947, n41948, n41949, n41950, n41951, n41952,
         n41953, n41954, n41955, n41956, n41957, n41958, n41959, n41960,
         n41961, n41962, n41963, n41964, n41965, n41966, n41967, n41968,
         n41969, n41970, n41971, n41972, n41973, n41974, n41975, n41976,
         n41977, n41978, n41979, n41980, n41981, n41982, n41983, n41984,
         n41985, n41986, n41987, n41988, n41989, n41990, n41991, n41992,
         n41993, n41994, n41995, n41996, n41997, n41998, n41999, n42000,
         n42001, n42002, n42003, n42004, n42005, n42006, n42007, n42008,
         n42009, n42010, n42011, n42012, n42013, n42014, n42015, n42016,
         n42017, n42018, n42019, n42020, n42021, n42022, n42023, n42024,
         n42025, n42026, n42027, n42028, n42029, n42030, n42031, n42032,
         n42033, n42034, n42035, n42036, n42037, n42038, n42039, n42040,
         n42041, n42042, n42043, n42044, n42045, n42046, n42047, n42048,
         n42049, n42050, n42051, n42052, n42053, n42054, n42055, n42056,
         n42057, n42058, n42059, n42060, n42061, n42062, n42063, n42064,
         n42065, n42066, n42067, n42068, n42069, n42070, n42071, n42072,
         n42073, n42074, n42075, n42076, n42077, n42078, n42079, n42080,
         n42081, n42082, n42083, n42084, n42085, n42086, n42087, n42088,
         n42089, n42090, n42091, n42092, n42093, n42094, n42095, n42096,
         n42097, n42098, n42099, n42100, n42101, n42102, n42103, n42104,
         n42105, n42106, n42107, n42108, n42109, n42110, n42111, n42112,
         n42113, n42114, n42115, n42116, n42117, n42118, n42119, n42120,
         n42121, n42122, n42123, n42124, n42125, n42126, n42127, n42128,
         n42129, n42130, n42131, n42132, n42133, n42134, n42135, n42136,
         n42137, n42138, n42139, n42140, n42141, n42142, n42143, n42144,
         n42145, n42146, n42147, n42148, n42149, n42150, n42151, n42152,
         n42153, n42154, n42155, n42156, n42157, n42158, n42159, n42160,
         n42161, n42162, n42163, n42164, n42165, n42166, n42167, n42168,
         n42169, n42170, n42171, n42172, n42173, n42174, n42175, n42176,
         n42177, n42178, n42179, n42180, n42181, n42182, n42183, n42184,
         n42185, n42186, n42187, n42188, n42189, n42190, n42191, n42192,
         n42193, n42194, n42195, n42196, n42197, n42198, n42199, n42200,
         n42201, n42202, n42203, n42204, n42205, n42206, n42207, n42208,
         n42209, n42210, n42211, n42212, n42213, n42214, n42215, n42216,
         n42217, n42218, n42219, n42220, n42221, n42222, n42223, n42224,
         n42225, n42226, n42227, n42228, n42229, n42230, n42231, n42232,
         n42233, n42234, n42235, n42236, n42237, n42238, n42239, n42240,
         n42241, n42242, n42243, n42244, n42245, n42246, n42247, n42248,
         n42249, n42250, n42251, n42252, n42253, n42254, n42255, n42256,
         n42257, n42258, n42259, n42260, n42261, n42262, n42263, n42264,
         n42265, n42266, n42267, n42268, n42269, n42270, n42271, n42272,
         n42273, n42274, n42275, n42276, n42277, n42278, n42279, n42280,
         n42281, n42282, n42283, n42284, n42285, n42286, n42287, n42288,
         n42289, n42290, n42291, n42292, n42293, n42294, n42295, n42296,
         n42297, n42298, n42299, n42300, n42301, n42302, n42303, n42304,
         n42305, n42306, n42307, n42308, n42309, n42310, n42311, n42312,
         n42313, n42314, n42315, n42316, n42317, n42318, n42319, n42320,
         n42321, n42322, n42323, n42324, n42325, n42326, n42327, n42328,
         n42329, n42330, n42331, n42332, n42333, n42334, n42335, n42336,
         n42337, n42338, n42339, n42340, n42341, n42342, n42343, n42344,
         n42345, n42346, n42347, n42348, n42349, n42350, n42351, n42352,
         n42353, n42354, n42355, n42356, n42357, n42358, n42359, n42360,
         n42361, n42362, n42363, n42364, n42365, n42366, n42367, n42368,
         n42369, n42370, n42371, n42372, n42373, n42374, n42375, n42376,
         n42377, n42378, n42379, n42380, n42381, n42382, n42383, n42384,
         n42385, n42386, n42387, n42388, n42389, n42390, n42391, n42392,
         n42393, n42394, n42395, n42396, n42397, n42398, n42399, n42400,
         n42401, n42402, n42403, n42404, n42405, n42406, n42407, n42408,
         n42409, n42410, n42411, n42412, n42413, n42414, n42415, n42416,
         n42417, n42418, n42419, n42420, n42421, n42422, n42423, n42424,
         n42425, n42426, n42427, n42428, n42429, n42430, n42431, n42432,
         n42433, n42434, n42435, n42436, n42437, n42438, n42439, n42440,
         n42441, n42442, n42443, n42444, n42445, n42446, n42447, n42448,
         n42449, n42450, n42451, n42452, n42453, n42454, n42455, n42456,
         n42457, n42458, n42459, n42460, n42461, n42462, n42463, n42464,
         n42465, n42466, n42467, n42468, n42469, n42470, n42471, n42472,
         n42473, n42474, n42475, n42476, n42477, n42478, n42479, n42480,
         n42481, n42482, n42483, n42484, n42485, n42486, n42487, n42488,
         n42489, n42490, n42491, n42492, n42493, n42494, n42495, n42496,
         n42497, n42498, n42499, n42500, n42501, n42502, n42503, n42504,
         n42505, n42506, n42507, n42508, n42509, n42510, n42511, n42512,
         n42513, n42514, n42515, n42516, n42517, n42518, n42519, n42520,
         n42521, n42522, n42523, n42524, n42525, n42526, n42527, n42528,
         n42529, n42530, n42531, n42532, n42533, n42534, n42535, n42536,
         n42537, n42538, n42539, n42540, n42541, n42542, n42543, n42544,
         n42545, n42546, n42547, n42548, n42549, n42550, n42551, n42552,
         n42553, n42554, n42555, n42556, n42557, n42558, n42559, n42560,
         n42561, n42562, n42563, n42564, n42565, n42566, n42567, n42568,
         n42569, n42570, n42571, n42572, n42573, n42574, n42575, n42576,
         n42577, n42578, n42579, n42580, n42581, n42582, n42583, n42584,
         n42585, n42586, n42587, n42588, n42589, n42590, n42591, n42592,
         n42593, n42594, n42595, n42596, n42597, n42598, n42599, n42600,
         n42601, n42602, n42603, n42604, n42605, n42606, n42607, n42608,
         n42609, n42610, n42611, n42612, n42613, n42614, n42615, n42616,
         n42617, n42618, n42619, n42620, n42621, n42622, n42623, n42624,
         n42625, n42626, n42627, n42628, n42629, n42630, n42631, n42632,
         n42633, n42634, n42635, n42636, n42637, n42638, n42639, n42640,
         n42641, n42642, n42643, n42644, n42645, n42646, n42647, n42648,
         n42649, n42650, n42651, n42652, n42653, n42654, n42655, n42656,
         n42657, n42658, n42659, n42660, n42661, n42662, n42663, n42664,
         n42665, n42666, n42667, n42668, n42669, n42670, n42671, n42672,
         n42673, n42674, n42675, n42676, n42677, n42678, n42679, n42680,
         n42681, n42682, n42683, n42684, n42685, n42686, n42687, n42688,
         n42689, n42690, n42691, n42692, n42693, n42694, n42695, n42696,
         n42697, n42698, n42699, n42700, n42701, n42702, n42703, n42704,
         n42705, n42706, n42707, n42708, n42709, n42710, n42711, n42712,
         n42713, n42714, n42715, n42716, n42717, n42718, n42719, n42720,
         n42721, n42722, n42723, n42724, n42725, n42726, n42727, n42728,
         n42729, n42730, n42731, n42732, n42733, n42734, n42735, n42736,
         n42737, n42738, n42739, n42740, n42741, n42742, n42743, n42744,
         n42745, n42746, n42747, n42748, n42749, n42750, n42751, n42752,
         n42753, n42754, n42755, n42756, n42757, n42758, n42759, n42760,
         n42761, n42762, n42763, n42764, n42765, n42766, n42767, n42768,
         n42769, n42770, n42771, n42772, n42773, n42774, n42775, n42776,
         n42777, n42778, n42779, n42780, n42781, n42782, n42783, n42784,
         n42785, n42786, n42787, n42788, n42789, n42790, n42791, n42792,
         n42793, n42794, n42795, n42796, n42797, n42798, n42799, n42800,
         n42801, n42802, n42803, n42804, n42805, n42806, n42807, n42808,
         n42809, n42810, n42811, n42812, n42813, n42814, n42815, n42816,
         n42817, n42818, n42819, n42820, n42821, n42822, n42823, n42824,
         n42825, n42826, n42827, n42828, n42829, n42830, n42831, n42832,
         n42833, n42834, n42835, n42836, n42837, n42838, n42839, n42840,
         n42841, n42842, n42843, n42844, n42845, n42846, n42847, n42848,
         n42849, n42850, n42851, n42852, n42853, n42854, n42855, n42856,
         n42857, n42858, n42859, n42860, n42861, n42862, n42863, n42864,
         n42865, n42866, n42867, n42868, n42869, n42870, n42871, n42872,
         n42873, n42874, n42875, n42876, n42877, n42878, n42879, n42880,
         n42881, n42882, n42883, n42884, n42885, n42886, n42887, n42888,
         n42889, n42890, n42891, n42892, n42893, n42894, n42895, n42896,
         n42897, n42898, n42899, n42900, n42901, n42902, n42903, n42904,
         n42905, n42906, n42907, n42908, n42909, n42910, n42911, n42912,
         n42913, n42914, n42915, n42916, n42917, n42918, n42919, n42920,
         n42921, n42922, n42923, n42924, n42925, n42926, n42927, n42928,
         n42929, n42930, n42931, n42932, n42933, n42934, n42935, n42936,
         n42937, n42938, n42939, n42940, n42941, n42942, n42943, n42944,
         n42945, n42946, n42947, n42948, n42949, n42950, n42951, n42952,
         n42953, n42954, n42955, n42956, n42957, n42958, n42959, n42960,
         n42961, n42962, n42963, n42964, n42965, n42966, n42967, n42968,
         n42969, n42970, n42971, n42972, n42973, n42974, n42975, n42976,
         n42977, n42978, n42979, n42980, n42981, n42982, n42983, n42984,
         n42985, n42986, n42987, n42988, n42989, n42990, n42991, n42992,
         n42993, n42994, n42995, n42996, n42997, n42998, n42999, n43000,
         n43001, n43002, n43003, n43004, n43005, n43006, n43007, n43008,
         n43009, n43010, n43011, n43012, n43013, n43014, n43015, n43016,
         n43017, n43018, n43019, n43020, n43021, n43022, n43023, n43024,
         n43025, n43026, n43027, n43028, n43029, n43030, n43031, n43032,
         n43033, n43034, n43035, n43036, n43037, n43038, n43039, n43040,
         n43041, n43042, n43043, n43044, n43045, n43046, n43047, n43048,
         n43049, n43050, n43051, n43052, n43053, n43054, n43055, n43056,
         n43057, n43058, n43059, n43060, n43061, n43062, n43063, n43064,
         n43065, n43066, n43067, n43068, n43069, n43070, n43071, n43072,
         n43073, n43074, n43075, n43076, n43077, n43078, n43079, n43080,
         n43081, n43082, n43083, n43084, n43085, n43086, n43087, n43088,
         n43089, n43090, n43091, n43092, n43093, n43094, n43095, n43096,
         n43097, n43098, n43099, n43100, n43101, n43102, n43103, n43104,
         n43105, n43106, n43107, n43108, n43109, n43110, n43111, n43112,
         n43113, n43114, n43115, n43116, n43117, n43118, n43119, n43120,
         n43121, n43122, n43123, n43124, n43125, n43126, n43127, n43128,
         n43129, n43130, n43131, n43132, n43133, n43134, n43135, n43136,
         n43137, n43138, n43139, n43140, n43141, n43142, n43143, n43144,
         n43145, n43146, n43147, n43148, n43149, n43150, n43151, n43152,
         n43153, n43154, n43155, n43156, n43157, n43158, n43159, n43160,
         n43161, n43162, n43163, n43164, n43165, n43166, n43167, n43168,
         n43169, n43170, n43171, n43172, n43173, n43174, n43175, n43176,
         n43177, n43178, n43179, n43180, n43181, n43182, n43183, n43184,
         n43185, n43186, n43187, n43188, n43189, n43190, n43191, n43192,
         n43193, n43194, n43195, n43196, n43197, n43198, n43199, n43200,
         n43201, n43202, n43203, n43204, n43205, n43206, n43207, n43208,
         n43209, n43210, n43211, n43212, n43213, n43214, n43215, n43216,
         n43217, n43218, n43219, n43220, n43221, n43222, n43223, n43224,
         n43225, n43226, n43227, n43228, n43229, n43230, n43231, n43232,
         n43233, n43234, n43235, n43236, n43237, n43238, n43239, n43240,
         n43241, n43242, n43243, n43244, n43245, n43246, n43247, n43248,
         n43249, n43250, n43251, n43252, n43253, n43254, n43255, n43256,
         n43257, n43258, n43259, n43260, n43261, n43262, n43263, n43264,
         n43265, n43266, n43267, n43268, n43269, n43270, n43271, n43272,
         n43273, n43274, n43275, n43276, n43277, n43278, n43279, n43280,
         n43281, n43282, n43283, n43284, n43285, n43286, n43287, n43288,
         n43289, n43290, n43291, n43292, n43293, n43294, n43295, n43296,
         n43297, n43298, n43299, n43300, n43301, n43302, n43303, n43304,
         n43305, n43306, n43307, n43308, n43309, n43310, n43311, n43312,
         n43313, n43314, n43315, n43316, n43317, n43318, n43319, n43320,
         n43321, n43322, n43323, n43324, n43325, n43326, n43327, n43328,
         n43329, n43330, n43331, n43332, n43333, n43334, n43335, n43336,
         n43337, n43338, n43339, n43340, n43341, n43342, n43343, n43344,
         n43345, n43346, n43347, n43348, n43349, n43350, n43351, n43352,
         n43353, n43354, n43355, n43356, n43357, n43358, n43359, n43360,
         n43361, n43362, n43363, n43364, n43365, n43366, n43367, n43368,
         n43369, n43370, n43371, n43372, n43373, n43374, n43375, n43376,
         n43377, n43378, n43379, n43380, n43381, n43382, n43383, n43384,
         n43385, n43386, n43387, n43388, n43389, n43390, n43391, n43392,
         n43393, n43394, n43395, n43396, n43397, n43398, n43399, n43400,
         n43401, n43402, n43403, n43404, n43405, n43406, n43407, n43408,
         n43409, n43410, n43411, n43412, n43413, n43414, n43415, n43416,
         n43417, n43418, n43419, n43420, n43421, n43422, n43423, n43424,
         n43425, n43426, n43427, n43428, n43429, n43430, n43431, n43432,
         n43433, n43434, n43435, n43436, n43437, n43438, n43439, n43440,
         n43441, n43442, n43443, n43444, n43445, n43446, n43447, n43448,
         n43449, n43450, n43451, n43452, n43453, n43454, n43455, n43456,
         n43457, n43458, n43459, n43460, n43461, n43462, n43463, n43464,
         n43465, n43466, n43467, n43468, n43469, n43470, n43471, n43472,
         n43473, n43474, n43475, n43476, n43477, n43478, n43479, n43480,
         n43481, n43482, n43483, n43484, n43485, n43486, n43487, n43488,
         n43489, n43490, n43491, n43492, n43493, n43494, n43495, n43496,
         n43497, n43498, n43499, n43500, n43501, n43502, n43503, n43504,
         n43505, n43506, n43507, n43508, n43509, n43510, n43511, n43512,
         n43513, n43514, n43515, n43516, n43517, n43518, n43519, n43520,
         n43521, n43522, n43523, n43524, n43525, n43526, n43527, n43528,
         n43529, n43530, n43531, n43532, n43533, n43534, n43535, n43536,
         n43537, n43538, n43539, n43540, n43541, n43542, n43543, n43544,
         n43545, n43546, n43547, n43548, n43549, n43550, n43551, n43552,
         n43553, n43554, n43555, n43556, n43557, n43558, n43559, n43560,
         n43561, n43562, n43563, n43564, n43565, n43566, n43567, n43568,
         n43569, n43570, n43571, n43572, n43573, n43574, n43575, n43576,
         n43577, n43578, n43579, n43580, n43581, n43582, n43583, n43584,
         n43585, n43586, n43587, n43588, n43589, n43590, n43591, n43592,
         n43593, n43594, n43595, n43596, n43597, n43598, n43599, n43600,
         n43601, n43602, n43603, n43604, n43605, n43606, n43607, n43608,
         n43609, n43610, n43611, n43612, n43613, n43614, n43615, n43616,
         n43617, n43618, n43619, n43620, n43621, n43622, n43623, n43624,
         n43625, n43626, n43627, n43628, n43629, n43630, n43631, n43632,
         n43633, n43634, n43635, n43636, n43637, n43638, n43639, n43640,
         n43641, n43642, n43643, n43644, n43645, n43646, n43647, n43648,
         n43649, n43650, n43651, n43652, n43653, n43654, n43655, n43656,
         n43657, n43658, n43659, n43660, n43661, n43662, n43663, n43664,
         n43665, n43666, n43667, n43668, n43669, n43670, n43671, n43672,
         n43673, n43674, n43675, n43676, n43677, n43678, n43679, n43680,
         n43681, n43682, n43683, n43684, n43685, n43686, n43687, n43688,
         n43689, n43690, n43691, n43692, n43693, n43694, n43695, n43696,
         n43697, n43698, n43699, n43700, n43701, n43702, n43703, n43704,
         n43705, n43706, n43707, n43708, n43709, n43710, n43711, n43712,
         n43713, n43714, n43715, n43716, n43717, n43718, n43719, n43720,
         n43721, n43722, n43723, n43724, n43725, n43726, n43727, n43728,
         n43729, n43730, n43731, n43732, n43733, n43734, n43735, n43736,
         n43737, n43738, n43739, n43740, n43741, n43742, n43743, n43744,
         n43745, n43746, n43747, n43748, n43749, n43750, n43751, n43752,
         n43753, n43754, n43755, n43756, n43757, n43758, n43759, n43760,
         n43761, n43762, n43763, n43764, n43765, n43766, n43767, n43768,
         n43769, n43770, n43771, n43772, n43773, n43774, n43775, n43776,
         n43777, n43778, n43779, n43780, n43781, n43782, n43783, n43784,
         n43785, n43786, n43787, n43788, n43789, n43790, n43791, n43792,
         n43793, n43794, n43795, n43796, n43797, n43798, n43799, n43800,
         n43801, n43802, n43803, n43804, n43805, n43806, n43807, n43808,
         n43809, n43810, n43811, n43812, n43813, n43814, n43815, n43816,
         n43817, n43818, n43819, n43820, n43821, n43822, n43823, n43824,
         n43825, n43826, n43827, n43828, n43829, n43830, n43831, n43832,
         n43833, n43834, n43835, n43836, n43837, n43838, n43839, n43840,
         n43841, n43842, n43843, n43844, n43845, n43846, n43847, n43848,
         n43849, n43850, n43851, n43852, n43853, n43854, n43855, n43856,
         n43857, n43858, n43859, n43860, n43861, n43862, n43863, n43864,
         n43865, n43866, n43867, n43868, n43869, n43870, n43871, n43872,
         n43873, n43874, n43875, n43876, n43877, n43878, n43879, n43880,
         n43881, n43882, n43883, n43884, n43885, n43886, n43887, n43888,
         n43889, n43890, n43891, n43892, n43893, n43894, n43895, n43896,
         n43897, n43898, n43899, n43900, n43901, n43902, n43903, n43904,
         n43905, n43906, n43907, n43908, n43909, n43910, n43911, n43912,
         n43913, n43914, n43915, n43916, n43917, n43918, n43919, n43920,
         n43921, n43922, n43923, n43924, n43925, n43926, n43927, n43928,
         n43929, n43930, n43931, n43932, n43933, n43934, n43935, n43936,
         n43937, n43938, n43939, n43940, n43941, n43942, n43943, n43944,
         n43945, n43946, n43947, n43948, n43949, n43950, n43951, n43952,
         n43953, n43954, n43955, n43956, n43957, n43958, n43959, n43960,
         n43961, n43962, n43963, n43964, n43965, n43966, n43967, n43968,
         n43969, n43970, n43971, n43972, n43973, n43974, n43975, n43976,
         n43977, n43978, n43979, n43980, n43981, n43982, n43983, n43984,
         n43985, n43986, n43987, n43988, n43989, n43990, n43991, n43992,
         n43993, n43994, n43995, n43996, n43997, n43998, n43999, n44000,
         n44001, n44002, n44003, n44004, n44005, n44006, n44007, n44008,
         n44009, n44010, n44011, n44012, n44013, n44014, n44015, n44016,
         n44017, n44018, n44019, n44020, n44021, n44022, n44023, n44024,
         n44025, n44026, n44027, n44028, n44029, n44030, n44031, n44032,
         n44033, n44034, n44035, n44036, n44037, n44038, n44039, n44040,
         n44041, n44042, n44043, n44044, n44045, n44046, n44047, n44048,
         n44049, n44050, n44051, n44052, n44053, n44054, n44055, n44056,
         n44057, n44058, n44059, n44060, n44061, n44062, n44063, n44064,
         n44065, n44066, n44067, n44068, n44069, n44070, n44071, n44072,
         n44073, n44074, n44075, n44076, n44077, n44078, n44079, n44080,
         n44081, n44082, n44083, n44084, n44085, n44086, n44087, n44088,
         n44089, n44090, n44091, n44092, n44093, n44094, n44095, n44096,
         n44097, n44098, n44099, n44100, n44101, n44102, n44103, n44104,
         n44105, n44106, n44107, n44108, n44109, n44110, n44111, n44112,
         n44113, n44114, n44115, n44116, n44117, n44118, n44119, n44120,
         n44121, n44122, n44123, n44124, n44125, n44126, n44127, n44128,
         n44129, n44130, n44131, n44132, n44133, n44134, n44135, n44136,
         n44137, n44138, n44139, n44140, n44141, n44142, n44143, n44144,
         n44145, n44146, n44147, n44148, n44149, n44150, n44151, n44152,
         n44153, n44154, n44155, n44156, n44157, n44158, n44159, n44160,
         n44161, n44162, n44163, n44164, n44165, n44166, n44167, n44168,
         n44169, n44170, n44171, n44172, n44173, n44174, n44175, n44176,
         n44177, n44178, n44179, n44180, n44181, n44182, n44183, n44184,
         n44185, n44186, n44187, n44188, n44189, n44190, n44191, n44192,
         n44193, n44194, n44195, n44196, n44197, n44198, n44199, n44200,
         n44201, n44202, n44203, n44204, n44205, n44206, n44207, n44208,
         n44209, n44210, n44211, n44212, n44213, n44214, n44215, n44216,
         n44217, n44218, n44219, n44220, n44221, n44222, n44223, n44224,
         n44225, n44226, n44227, n44228, n44229, n44230, n44231, n44232,
         n44233, n44234, n44235, n44236, n44237, n44238, n44239, n44240,
         n44241, n44242, n44243, n44244, n44245, n44246, n44247, n44248,
         n44249, n44250, n44251, n44252, n44253, n44254, n44255, n44256,
         n44257, n44258, n44259, n44260, n44261, n44262, n44263, n44264,
         n44265, n44266, n44267, n44268, n44269, n44270, n44271, n44272,
         n44273, n44274, n44275, n44276, n44277, n44278, n44279, n44280,
         n44281, n44282, n44283, n44284, n44285, n44286, n44287, n44288,
         n44289, n44290, n44291, n44292, n44293, n44294, n44295, n44296,
         n44297, n44298, n44299, n44300, n44301, n44302, n44303, n44304,
         n44305, n44306, n44307, n44308, n44309, n44310, n44311, n44312,
         n44313, n44314, n44315, n44316, n44317, n44318, n44319, n44320,
         n44321, n44322, n44323, n44324, n44325, n44326, n44327, n44328,
         n44329, n44330, n44331, n44332, n44333, n44334, n44335, n44336,
         n44337, n44338, n44339, n44340, n44341, n44342, n44343, n44344,
         n44345, n44346, n44347, n44348, n44349, n44350, n44351, n44352,
         n44353, n44354, n44355, n44356, n44357, n44358, n44359, n44360,
         n44361, n44362, n44363, n44364, n44365, n44366, n44367, n44368,
         n44369, n44370, n44371, n44372, n44373, n44374, n44375, n44376,
         n44377, n44378, n44379, n44380, n44381, n44382, n44383, n44384,
         n44385, n44386, n44387, n44388, n44389, n44390, n44391, n44392,
         n44393, n44394, n44395, n44396, n44397, n44398, n44399, n44400,
         n44401, n44402, n44403, n44404, n44405, n44406, n44407, n44408,
         n44409, n44410, n44411, n44412, n44413, n44414, n44415, n44416,
         n44417, n44418, n44419, n44420, n44421, n44422, n44423, n44424,
         n44425, n44426, n44427, n44428, n44429, n44430, n44431, n44432,
         n44433, n44434, n44435, n44436, n44437, n44438, n44439, n44440,
         n44441, n44442, n44443, n44444, n44445, n44446, n44447, n44448,
         n44449, n44450, n44451, n44452, n44453, n44454, n44455, n44456,
         n44457, n44458, n44459, n44460, n44461, n44462, n44463, n44464,
         n44465, n44466, n44467, n44468, n44469, n44470, n44471, n44472,
         n44473, n44474, n44475, n44476, n44477, n44478, n44479, n44480,
         n44481, n44482, n44483, n44484, n44485, n44486, n44487, n44488,
         n44489, n44490, n44491, n44492, n44493, n44494, n44495, n44496,
         n44497, n44498, n44499, n44500, n44501, n44502, n44503, n44504,
         n44505, n44506, n44507, n44508, n44509, n44510, n44511, n44512,
         n44513, n44514, n44515, n44516, n44517, n44518, n44519, n44520,
         n44521, n44522, n44523, n44524, n44525, n44526, n44527, n44528,
         n44529, n44530, n44531, n44532, n44533, n44534, n44535, n44536,
         n44537, n44538, n44539, n44540, n44541, n44542, n44543, n44544,
         n44545, n44546, n44547, n44548, n44549, n44550, n44551, n44552,
         n44553, n44554, n44555, n44556, n44557, n44558, n44559, n44560,
         n44561, n44562, n44563, n44564, n44565, n44566, n44567, n44568,
         n44569, n44570, n44571, n44572, n44573, n44574, n44575, n44576,
         n44577, n44578, n44579, n44580, n44581, n44582, n44583, n44584,
         n44585, n44586, n44587, n44588, n44589, n44590, n44591, n44592,
         n44593, n44594, n44595, n44596, n44597, n44598, n44599, n44600,
         n44601, n44602, n44603, n44604, n44605, n44606, n44607, n44608,
         n44609, n44610, n44611, n44612, n44613, n44614, n44615, n44616,
         n44617, n44618, n44619, n44620, n44621, n44622, n44623, n44624,
         n44625, n44626, n44627, n44628, n44629, n44630, n44631, n44632,
         n44633, n44634, n44635, n44636, n44637, n44638, n44639, n44640,
         n44641, n44642, n44643, n44644, n44645, n44646, n44647, n44648,
         n44649, n44650, n44651, n44652, n44653, n44654, n44655, n44656,
         n44657, n44658, n44659, n44660, n44661, n44662, n44663, n44664,
         n44665, n44666, n44667, n44668, n44669, n44670, n44671, n44672,
         n44673, n44674, n44675, n44676, n44677, n44678, n44679, n44680,
         n44681, n44682, n44683, n44684, n44685, n44686, n44687, n44688,
         n44689, n44690, n44691, n44692, n44693, n44694, n44695, n44696,
         n44697, n44698, n44699, n44700, n44701, n44702, n44703, n44704,
         n44705, n44706, n44707, n44708, n44709, n44710, n44711, n44712,
         n44713, n44714, n44715, n44716, n44717, n44718, n44719, n44720,
         n44721, n44722, n44723, n44724, n44725, n44726, n44727, n44728,
         n44729, n44730, n44731, n44732, n44733, n44734, n44735, n44736,
         n44737, n44738, n44739, n44740, n44741, n44742, n44743, n44744,
         n44745, n44746, n44747, n44748, n44749, n44750, n44751, n44752,
         n44753, n44754, n44755, n44756, n44757, n44758, n44759, n44760,
         n44761, n44762, n44763, n44764, n44765, n44766, n44767, n44768,
         n44769, n44770, n44771, n44772, n44773, n44774, n44775, n44776,
         n44777, n44778, n44779, n44780, n44781, n44782, n44783, n44784,
         n44785, n44786, n44787, n44788, n44789, n44790, n44791, n44792,
         n44793, n44794, n44795, n44796, n44797, n44798, n44799, n44800,
         n44801, n44802, n44803, n44804, n44805, n44806, n44807, n44808,
         n44809, n44810, n44811, n44812, n44813, n44814, n44815, n44816,
         n44817, n44818, n44819, n44820, n44821, n44822, n44823, n44824,
         n44825, n44826, n44827, n44828, n44829, n44830, n44831, n44832,
         n44833, n44834, n44835, n44836, n44837, n44838, n44839, n44840,
         n44841, n44842, n44843, n44844, n44845, n44846, n44847, n44848,
         n44849, n44850, n44851, n44852, n44853, n44854, n44855, n44856,
         n44857, n44858, n44859, n44860, n44861, n44862, n44863, n44864,
         n44865, n44866, n44867, n44868, n44869, n44870, n44871, n44872,
         n44873, n44874, n44875, n44876, n44877, n44878, n44879, n44880,
         n44881, n44882, n44883, n44884, n44885, n44886, n44887, n44888,
         n44889, n44890, n44891, n44892, n44893, n44894, n44895, n44896,
         n44897, n44898, n44899, n44900, n44901, n44902, n44903, n44904,
         n44905, n44906, n44907, n44908, n44909, n44910, n44911, n44912,
         n44913, n44914, n44915, n44916, n44917, n44918, n44919, n44920,
         n44921, n44922, n44923, n44924, n44925, n44926, n44927, n44928,
         n44929, n44930, n44931, n44932, n44933, n44934, n44935, n44936,
         n44937, n44938, n44939, n44940, n44941, n44942, n44943, n44944,
         n44945, n44946, n44947, n44948, n44949, n44950, n44951, n44952,
         n44953, n44954, n44955, n44956, n44957, n44958, n44959, n44960,
         n44961, n44962, n44963, n44964, n44965, n44966, n44967, n44968,
         n44969, n44970, n44971, n44972, n44973, n44974, n44975, n44976,
         n44977, n44978, n44979, n44980, n44981, n44982, n44983, n44984,
         n44985, n44986, n44987, n44988, n44989, n44990, n44991, n44992,
         n44993, n44994, n44995, n44996, n44997, n44998, n44999, n45000,
         n45001, n45002, n45003, n45004, n45005, n45006, n45007, n45008,
         n45009, n45010, n45011, n45012, n45013, n45014, n45015, n45016,
         n45017, n45018, n45019, n45020, n45021, n45022, n45023, n45024,
         n45025, n45026, n45027, n45028, n45029, n45030, n45031, n45032,
         n45033, n45034, n45035, n45036, n45037, n45038, n45039, n45040,
         n45041, n45042, n45043, n45044, n45045, n45046, n45047, n45048,
         n45049, n45050, n45051, n45052, n45053, n45054, n45055, n45056,
         n45057, n45058, n45059, n45060, n45061, n45062, n45063, n45064,
         n45065, n45066, n45067, n45068, n45069, n45070, n45071, n45072,
         n45073, n45074, n45075, n45076, n45077, n45078, n45079, n45080,
         n45081, n45082, n45083, n45084, n45085, n45086, n45087, n45088,
         n45089, n45090, n45091, n45092, n45093, n45094, n45095, n45096,
         n45097, n45098, n45099, n45100, n45101, n45102, n45103, n45104,
         n45105, n45106, n45107, n45108, n45109, n45110, n45111, n45112,
         n45113, n45114, n45115, n45116, n45117, n45118, n45119, n45120,
         n45121, n45122, n45123, n45124, n45125, n45126, n45127, n45128,
         n45129, n45130, n45131, n45132, n45133, n45134, n45135, n45136,
         n45137, n45138, n45139, n45140, n45141, n45142, n45143, n45144,
         n45145, n45146, n45147, n45148, n45149, n45150, n45151, n45152,
         n45153, n45154, n45155, n45156, n45157, n45158, n45159, n45160,
         n45161, n45162, n45163, n45164, n45165, n45166, n45167, n45168,
         n45169, n45170, n45171, n45172, n45173, n45174, n45175, n45176,
         n45177, n45178, n45179, n45180, n45181, n45182, n45183, n45184,
         n45185, n45186, n45187, n45188, n45189, n45190, n45191, n45192,
         n45193, n45194, n45195, n45196, n45197, n45198, n45199, n45200,
         n45201, n45202, n45203, n45204, n45205, n45206, n45207, n45208,
         n45209, n45210, n45211, n45212, n45213, n45214, n45215, n45216,
         n45217, n45218, n45219, n45220, n45221, n45222, n45223, n45224,
         n45225, n45226, n45227, n45228, n45229, n45230, n45231, n45232,
         n45233, n45234, n45235, n45236, n45237, n45238, n45239, n45240,
         n45241, n45242, n45243, n45244, n45245, n45246, n45247, n45248,
         n45249, n45250, n45251, n45252, n45253, n45254, n45255, n45256,
         n45257, n45258, n45259, n45260, n45261, n45262, n45263, n45264,
         n45265, n45266, n45267, n45268, n45269, n45270, n45271, n45272,
         n45273, n45274, n45275, n45276, n45277, n45278, n45279, n45280,
         n45281, n45282, n45283, n45284, n45285, n45286, n45287, n45288,
         n45289, n45290, n45291, n45292, n45293, n45294, n45295, n45296,
         n45297, n45298, n45299, n45300, n45301, n45302, n45303, n45304,
         n45305, n45306, n45307, n45308, n45309, n45310, n45311, n45312,
         n45313, n45314, n45315, n45316, n45317, n45318, n45319, n45320,
         n45321, n45322, n45323, n45324, n45325, n45326, n45327, n45328,
         n45329, n45330, n45331, n45332, n45333, n45334, n45335, n45336,
         n45337, n45338, n45339, n45340, n45341, n45342, n45343, n45344,
         n45345, n45346, n45347, n45348, n45349, n45350, n45351, n45352,
         n45353, n45354, n45355, n45356, n45357, n45358, n45359, n45360,
         n45361, n45362, n45363, n45364, n45365, n45366, n45367, n45368,
         n45369, n45370, n45371, n45372, n45373, n45374, n45375, n45376,
         n45377, n45378, n45379, n45380, n45381, n45382, n45383, n45384,
         n45385, n45386, n45387, n45388, n45389, n45390, n45391, n45392,
         n45393, n45394, n45395, n45396, n45397, n45398, n45399, n45400,
         n45401, n45402, n45403, n45404, n45405, n45406, n45407, n45408,
         n45409, n45410, n45411, n45412, n45413, n45414, n45415, n45416,
         n45417, n45418, n45419, n45420, n45421, n45422, n45423, n45424,
         n45425, n45426, n45427, n45428, n45429, n45430, n45431, n45432,
         n45433, n45434, n45435, n45436, n45437, n45438, n45439, n45440,
         n45441, n45442, n45443, n45444, n45445, n45446, n45447, n45448,
         n45449, n45450, n45451, n45452, n45453, n45454, n45455, n45456,
         n45457, n45458, n45459, n45460, n45461, n45462, n45463, n45464,
         n45465, n45466, n45467, n45468, n45469, n45470, n45471, n45472,
         n45473, n45474, n45475, n45476, n45477, n45478, n45479, n45480,
         n45481, n45482, n45483, n45484, n45485, n45486, n45487, n45488,
         n45489, n45490, n45491, n45492, n45493, n45494, n45495, n45496,
         n45497, n45498, n45499, n45500, n45501, n45502, n45503, n45504,
         n45505, n45506, n45507, n45508, n45509, n45510, n45511, n45512,
         n45513, n45514, n45515, n45516, n45517, n45518, n45519, n45520,
         n45521, n45522, n45523, n45524, n45525, n45526, n45527, n45528,
         n45529, n45530, n45531, n45532, n45533, n45534, n45535, n45536,
         n45537, n45538, n45539, n45540, n45541, n45542, n45543, n45544,
         n45545, n45546, n45547, n45548, n45549, n45550, n45551, n45552,
         n45553, n45554, n45555, n45556, n45557, n45558, n45559, n45560,
         n45561, n45562, n45563, n45564, n45565, n45566, n45567, n45568,
         n45569, n45570, n45571, n45572, n45573, n45574, n45575, n45576,
         n45577, n45578, n45579, n45580, n45581, n45582, n45583, n45584,
         n45585, n45586, n45587, n45588, n45589, n45590, n45591, n45592,
         n45593, n45594, n45595, n45596, n45597, n45598, n45599, n45600,
         n45601, n45602, n45603, n45604, n45605, n45606, n45607, n45608,
         n45609, n45610, n45611, n45612, n45613, n45614, n45615, n45616,
         n45617, n45618, n45619, n45620, n45621, n45622, n45623, n45624,
         n45625, n45626, n45627, n45628, n45629, n45630, n45631, n45632,
         n45633, n45634, n45635, n45636, n45637, n45638, n45639, n45640,
         n45641, n45642, n45643, n45644, n45645, n45646, n45647, n45648,
         n45649, n45650, n45651, n45652, n45653, n45654, n45655, n45656,
         n45657, n45658, n45659, n45660, n45661, n45662, n45663, n45664,
         n45665, n45666, n45667, n45668, n45669, n45670, n45671, n45672,
         n45673, n45674, n45675, n45676, n45677, n45678, n45679, n45680,
         n45681, n45682, n45683, n45684, n45685, n45686, n45687, n45688,
         n45689, n45690, n45691, n45692, n45693, n45694, n45695, n45696,
         n45697, n45698, n45699, n45700, n45701, n45702, n45703, n45704,
         n45705, n45706, n45707, n45708, n45709, n45710, n45711, n45712,
         n45713, n45714, n45715, n45716, n45717, n45718, n45719, n45720,
         n45721, n45722, n45723, n45724, n45725, n45726, n45727, n45728,
         n45729, n45730, n45731, n45732, n45733, n45734, n45735, n45736,
         n45737, n45738, n45739, n45740, n45741, n45742, n45743, n45744,
         n45745, n45746, n45747, n45748, n45749, n45750, n45751, n45752,
         n45753, n45754, n45755, n45756, n45757, n45758, n45759, n45760,
         n45761, n45762, n45763, n45764, n45765, n45766, n45767, n45768,
         n45769, n45770, n45771, n45772, n45773, n45774, n45775, n45776,
         n45777, n45778, n45779, n45780, n45781, n45782, n45783, n45784,
         n45785, n45786, n45787, n45788, n45789, n45790, n45791, n45792,
         n45793, n45794, n45795, n45796, n45797, n45798, n45799, n45800,
         n45801, n45802, n45803, n45804, n45805, n45806, n45807, n45808,
         n45809, n45810, n45811, n45812, n45813, n45814, n45815, n45816,
         n45817, n45818, n45819, n45820, n45821, n45822, n45823, n45824,
         n45825, n45826, n45827, n45828, n45829, n45830, n45831, n45832,
         n45833, n45834, n45835, n45836, n45837, n45838, n45839, n45840,
         n45841, n45842, n45843, n45844, n45845, n45846, n45847, n45848,
         n45849, n45850, n45851, n45852, n45853, n45854, n45855, n45856,
         n45857, n45858, n45859, n45860, n45861, n45862, n45863, n45864,
         n45865, n45866, n45867, n45868, n45869, n45870, n45871, n45872,
         n45873, n45874, n45875, n45876, n45877, n45878, n45879, n45880,
         n45881, n45882, n45883, n45884, n45885, n45886, n45887, n45888,
         n45889, n45890, n45891, n45892, n45893, n45894, n45895, n45896,
         n45897, n45898, n45899, n45900, n45901, n45902, n45903, n45904,
         n45905, n45906, n45907, n45908, n45909, n45910, n45911, n45912,
         n45913, n45914, n45915, n45916, n45917, n45918, n45919, n45920,
         n45921, n45922, n45923, n45924, n45925, n45926, n45927, n45928,
         n45929, n45930, n45931, n45932, n45933, n45934, n45935, n45936,
         n45937, n45938, n45939, n45940, n45941, n45942, n45943, n45944,
         n45945, n45946, n45947, n45948, n45949, n45950, n45951, n45952,
         n45953, n45954, n45955, n45956, n45957, n45958, n45959, n45960,
         n45961, n45962, n45963, n45964, n45965, n45966, n45967, n45968,
         n45969, n45970, n45971, n45972, n45973, n45974, n45975, n45976,
         n45977, n45978, n45979, n45980, n45981, n45982, n45983, n45984,
         n45985, n45986, n45987, n45988, n45989, n45990, n45991, n45992,
         n45993, n45994, n45995, n45996, n45997, n45998, n45999, n46000,
         n46001, n46002, n46003, n46004, n46005, n46006, n46007, n46008,
         n46009, n46010, n46011, n46012, n46013, n46014, n46015, n46016,
         n46017, n46018, n46019, n46020, n46021, n46022, n46023, n46024,
         n46025, n46026, n46027, n46028, n46029, n46030, n46031, n46032,
         n46033, n46034, n46035, n46036, n46037, n46038, n46039, n46040,
         n46041, n46042, n46043, n46044, n46045, n46046, n46047, n46048,
         n46049, n46050, n46051, n46052, n46053, n46054, n46055, n46056,
         n46057, n46058, n46059, n46060, n46061, n46062, n46063, n46064,
         n46065, n46066, n46067, n46068, n46069, n46070, n46071, n46072,
         n46073, n46074, n46075, n46076, n46077, n46078, n46079, n46080,
         n46081, n46082, n46083, n46084, n46085, n46086, n46087, n46088,
         n46089, n46090, n46091, n46092, n46093, n46094, n46095, n46096,
         n46097, n46098, n46099, n46100, n46101, n46102, n46103, n46104,
         n46105, n46106, n46107, n46108, n46109, n46110, n46111, n46112,
         n46113, n46114, n46115, n46116, n46117, n46118, n46119, n46120,
         n46121, n46122, n46123, n46124, n46125, n46126, n46127, n46128,
         n46129, n46130, n46131, n46132, n46133, n46134, n46135, n46136,
         n46137, n46138, n46139, n46140, n46141, n46142, n46143, n46144,
         n46145, n46146, n46147, n46148, n46149, n46150, n46151, n46152,
         n46153, n46154, n46155, n46156, n46157, n46158, n46159, n46160,
         n46161, n46162, n46163, n46164, n46165, n46166, n46167, n46168,
         n46169, n46170, n46171, n46172, n46173, n46174, n46175, n46176,
         n46177, n46178, n46179, n46180, n46181, n46182, n46183, n46184,
         n46185, n46186, n46187, n46188, n46189, n46190, n46191, n46192,
         n46193, n46194, n46195, n46196, n46197, n46198, n46199, n46200,
         n46201, n46202, n46203, n46204, n46205, n46206, n46207, n46208,
         n46209, n46210, n46211, n46212, n46213, n46214, n46215, n46216,
         n46217, n46218, n46219, n46220, n46221, n46222, n46223, n46224,
         n46225, n46226, n46227, n46228, n46229, n46230, n46231, n46232,
         n46233, n46234, n46235, n46236, n46237, n46238, n46239, n46240,
         n46241, n46242, n46243, n46244, n46245, n46246, n46247, n46248,
         n46249, n46250, n46251, n46252, n46253, n46254, n46255, n46256,
         n46257, n46258, n46259, n46260, n46261, n46262, n46263, n46264,
         n46265, n46266, n46267, n46268, n46269, n46270, n46271, n46272,
         n46273, n46274, n46275, n46276, n46277, n46278, n46279, n46280,
         n46281, n46282, n46283, n46284, n46285, n46286, n46287, n46288,
         n46289, n46290, n46291, n46292, n46293, n46294, n46295, n46296,
         n46297, n46298, n46299, n46300, n46301, n46302, n46303, n46304,
         n46305, n46306, n46307, n46308, n46309, n46310, n46311, n46312,
         n46313, n46314, n46315, n46316, n46317, n46318, n46319, n46320,
         n46321, n46322, n46323, n46324, n46325, n46326, n46327, n46328,
         n46329, n46330, n46331, n46332, n46333, n46334, n46335, n46336,
         n46337, n46338, n46339, n46340, n46341, n46342, n46343, n46344,
         n46345, n46346, n46347, n46348, n46349, n46350, n46351, n46352,
         n46353, n46354, n46355, n46356, n46357, n46358, n46359, n46360,
         n46361, n46362, n46363, n46364, n46365, n46366, n46367, n46368,
         n46369, n46370, n46371, n46372, n46373, n46374, n46375, n46376,
         n46377, n46378, n46379, n46380, n46381, n46382, n46383, n46384,
         n46385, n46386, n46387, n46388, n46389, n46390, n46391, n46392,
         n46393, n46394, n46395, n46396, n46397, n46398, n46399, n46400,
         n46401, n46402, n46403, n46404, n46405, n46406, n46407, n46408,
         n46409, n46410, n46411, n46412, n46413, n46414, n46415, n46416,
         n46417, n46418, n46419, n46420, n46421, n46422, n46423, n46424,
         n46425, n46426, n46427, n46428, n46429, n46430, n46431, n46432,
         n46433, n46434, n46435, n46436, n46437, n46438, n46439, n46440,
         n46441, n46442, n46443, n46444, n46445, n46446, n46447, n46448,
         n46449, n46450, n46451, n46452, n46453, n46454, n46455, n46456,
         n46457, n46458, n46459, n46460, n46461, n46462, n46463, n46464,
         n46465, n46466, n46467, n46468, n46469, n46470, n46471, n46472,
         n46473, n46474, n46475, n46476, n46477, n46478, n46479, n46480,
         n46481, n46482, n46483, n46484, n46485, n46486, n46487, n46488,
         n46489, n46490, n46491, n46492, n46493, n46494, n46495, n46496,
         n46497, n46498, n46499, n46500, n46501, n46502, n46503, n46504,
         n46505, n46506, n46507, n46508, n46509, n46510, n46511, n46512,
         n46513, n46514, n46515, n46516, n46517, n46518, n46519, n46520,
         n46521, n46522, n46523, n46524, n46525, n46526, n46527, n46528,
         n46529, n46530, n46531, n46532, n46533, n46534, n46535, n46536,
         n46537, n46538, n46539, n46540, n46541, n46542, n46543, n46544,
         n46545, n46546, n46547, n46548, n46549, n46550, n46551, n46552,
         n46553, n46554, n46555, n46556, n46557, n46558, n46559, n46560,
         n46561, n46562, n46563, n46564, n46565, n46566, n46567, n46568,
         n46569, n46570, n46571, n46572, n46573, n46574, n46575, n46576,
         n46577, n46578, n46579, n46580, n46581, n46582, n46583, n46584,
         n46585, n46586, n46587, n46588, n46589, n46590, n46591, n46592,
         n46593, n46594, n46595, n46596, n46597, n46598, n46599, n46600,
         n46601, n46602, n46603, n46604, n46605, n46606, n46607, n46608,
         n46609, n46610, n46611, n46612, n46613, n46614, n46615, n46616,
         n46617, n46618, n46619, n46620, n46621, n46622, n46623, n46624,
         n46625, n46626, n46627, n46628, n46629, n46630, n46631, n46632,
         n46633, n46634, n46635, n46636, n46637, n46638, n46639, n46640,
         n46641, n46642, n46643, n46644, n46645, n46646, n46647, n46648,
         n46649, n46650, n46651, n46652, n46653, n46654, n46655, n46656,
         n46657, n46658, n46659, n46660, n46661, n46662, n46663, n46664,
         n46665, n46666, n46667, n46668, n46669, n46670, n46671, n46672,
         n46673, n46674, n46675, n46676, n46677, n46678, n46679, n46680,
         n46681, n46682, n46683, n46684, n46685, n46686, n46687, n46688,
         n46689, n46690, n46691, n46692, n46693, n46694, n46695, n46696,
         n46697, n46698, n46699, n46700, n46701, n46702, n46703, n46704,
         n46705, n46706, n46707, n46708, n46709, n46710, n46711, n46712,
         n46713, n46714, n46715, n46716, n46717, n46718, n46719, n46720,
         n46721, n46722, n46723, n46724, n46725, n46726, n46727, n46728,
         n46729, n46730, n46731, n46732, n46733, n46734, n46735, n46736,
         n46737, n46738, n46739, n46740, n46741, n46742, n46743, n46744,
         n46745, n46746, n46747, n46748, n46749, n46750, n46751, n46752,
         n46753, n46754, n46755, n46756, n46757, n46758, n46759, n46760,
         n46761, n46762, n46763, n46764, n46765, n46766, n46767, n46768,
         n46769, n46770, n46771, n46772, n46773, n46774, n46775, n46776,
         n46777, n46778, n46779, n46780, n46781, n46782, n46783, n46784,
         n46785, n46786, n46787, n46788, n46789, n46790, n46791, n46792,
         n46793, n46794, n46795, n46796, n46797, n46798, n46799, n46800,
         n46801, n46802, n46803, n46804, n46805, n46806, n46807, n46808,
         n46809, n46810, n46811, n46812, n46813, n46814, n46815, n46816,
         n46817, n46818, n46819, n46820, n46821, n46822, n46823, n46824,
         n46825, n46826, n46827, n46828, n46829, n46830, n46831, n46832,
         n46833, n46834, n46835, n46836, n46837, n46838, n46839, n46840,
         n46841, n46842, n46843, n46844, n46845, n46846, n46847, n46848,
         n46849, n46850, n46851, n46852, n46853, n46854, n46855, n46856,
         n46857, n46858, n46859, n46860, n46861, n46862, n46863, n46864,
         n46865, n46866, n46867, n46868, n46869, n46870, n46871, n46872,
         n46873, n46874, n46875, n46876, n46877, n46878, n46879, n46880,
         n46881, n46882, n46883, n46884, n46885, n46886, n46887, n46888,
         n46889, n46890, n46891, n46892, n46893, n46894, n46895, n46896,
         n46897, n46898, n46899, n46900, n46901, n46902, n46903, n46904,
         n46905, n46906, n46907, n46908, n46909, n46910, n46911, n46912,
         n46913, n46914, n46915, n46916, n46917, n46918, n46919, n46920,
         n46921, n46922, n46923, n46924, n46925, n46926, n46927, n46928,
         n46929, n46930, n46931, n46932, n46933, n46934, n46935, n46936,
         n46937, n46938, n46939, n46940, n46941, n46942, n46943, n46944,
         n46945, n46946, n46947, n46948, n46949, n46950, n46951, n46952,
         n46953, n46954, n46955, n46956, n46957, n46958, n46959, n46960,
         n46961, n46962, n46963, n46964, n46965, n46966, n46967, n46968,
         n46969, n46970, n46971, n46972, n46973, n46974, n46975, n46976,
         n46977, n46978, n46979, n46980, n46981, n46982, n46983, n46984,
         n46985, n46986, n46987, n46988, n46989, n46990, n46991, n46992,
         n46993, n46994, n46995, n46996, n46997, n46998, n46999, n47000,
         n47001, n47002, n47003, n47004, n47005, n47006, n47007, n47008,
         n47009, n47010, n47011, n47012, n47013, n47014, n47015, n47016,
         n47017, n47018, n47019, n47020, n47021, n47022, n47023, n47024,
         n47025, n47026, n47027, n47028, n47029, n47030, n47031, n47032,
         n47033, n47034, n47035, n47036, n47037, n47038, n47039, n47040,
         n47041, n47042, n47043, n47044, n47045, n47046, n47047, n47048,
         n47049, n47050, n47051, n47052, n47053, n47054, n47055, n47056,
         n47057, n47058, n47059, n47060, n47061, n47062, n47063, n47064,
         n47065, n47066, n47067, n47068, n47069, n47070, n47071, n47072,
         n47073, n47074, n47075, n47076, n47077, n47078, n47079, n47080,
         n47081, n47082, n47083, n47084, n47085, n47086, n47087, n47088,
         n47089, n47090, n47091, n47092, n47093, n47094, n47095, n47096,
         n47097, n47098, n47099, n47100, n47101, n47102, n47103, n47104,
         n47105, n47106, n47107, n47108, n47109, n47110, n47111, n47112,
         n47113, n47114, n47115, n47116, n47117, n47118, n47119, n47120,
         n47121, n47122, n47123, n47124, n47125, n47126, n47127, n47128,
         n47129, n47130, n47131, n47132, n47133, n47134, n47135, n47136,
         n47137, n47138, n47139, n47140, n47141, n47142, n47143, n47144,
         n47145, n47146, n47147, n47148, n47149, n47150, n47151, n47152,
         n47153, n47154, n47155, n47156, n47157, n47158, n47159, n47160,
         n47161, n47162, n47163, n47164, n47165, n47166, n47167, n47168,
         n47169, n47170, n47171, n47172, n47173, n47174, n47175, n47176,
         n47177, n47178, n47179, n47180, n47181, n47182, n47183, n47184,
         n47185, n47186, n47187, n47188, n47189, n47190, n47191, n47192,
         n47193, n47194, n47195, n47196, n47197, n47198, n47199, n47200,
         n47201, n47202, n47203, n47204, n47205, n47206, n47207, n47208,
         n47209, n47210, n47211, n47212, n47213, n47214, n47215, n47216,
         n47217, n47218, n47219, n47220, n47221, n47222, n47223, n47224,
         n47225, n47226, n47227, n47228, n47229, n47230, n47231, n47232,
         n47233, n47234, n47235, n47236, n47237, n47238, n47239, n47240,
         n47241, n47242, n47243, n47244, n47245, n47246, n47247, n47248,
         n47249, n47250, n47251, n47252, n47253, n47254, n47255, n47256,
         n47257, n47258, n47259, n47260, n47261, n47262, n47263, n47264,
         n47265, n47266, n47267, n47268, n47269, n47270, n47271, n47272,
         n47273, n47274, n47275, n47276, n47277, n47278, n47279, n47280,
         n47281, n47282, n47283, n47284, n47285, n47286, n47287, n47288,
         n47289, n47290, n47291, n47292, n47293, n47294, n47295, n47296,
         n47297, n47298, n47299, n47300, n47301, n47302, n47303, n47304,
         n47305, n47306, n47307, n47308, n47309, n47310, n47311, n47312,
         n47313, n47314, n47315, n47316, n47317, n47318, n47319, n47320,
         n47321, n47322, n47323, n47324, n47325, n47326, n47327, n47328,
         n47329, n47330, n47331, n47332, n47333, n47334, n47335, n47336,
         n47337, n47338, n47339, n47340, n47341, n47342, n47343, n47344,
         n47345, n47346, n47347, n47348, n47349, n47350, n47351, n47352,
         n47353, n47354, n47355, n47356, n47357, n47358, n47359, n47360,
         n47361, n47362, n47363, n47364, n47365, n47366, n47367, n47368,
         n47369, n47370, n47371, n47372, n47373, n47374, n47375, n47376,
         n47377, n47378, n47379, n47380, n47381, n47382, n47383, n47384,
         n47385, n47386, n47387, n47388, n47389, n47390, n47391, n47392,
         n47393, n47394, n47395, n47396, n47397, n47398, n47399, n47400,
         n47401, n47402, n47403, n47404, n47405, n47406, n47407, n47408,
         n47409, n47410, n47411, n47412, n47413, n47414, n47415, n47416,
         n47417, n47418, n47419, n47420, n47421, n47422, n47423, n47424,
         n47425, n47426, n47427, n47428, n47429, n47430, n47431, n47432,
         n47433, n47434, n47435, n47436, n47437, n47438, n47439, n47440,
         n47441, n47442, n47443, n47444, n47445, n47446, n47447, n47448,
         n47449, n47450, n47451, n47452, n47453, n47454, n47455, n47456,
         n47457, n47458, n47459, n47460, n47461, n47462, n47463, n47464,
         n47465, n47466, n47467, n47468, n47469, n47470, n47471, n47472,
         n47473, n47474, n47475, n47476, n47477, n47478, n47479, n47480,
         n47481, n47482, n47483, n47484, n47485, n47486, n47487, n47488,
         n47489, n47490, n47491, n47492, n47493, n47494, n47495, n47496,
         n47497, n47498, n47499, n47500, n47501, n47502, n47503, n47504,
         n47505, n47506, n47507, n47508, n47509, n47510, n47511, n47512,
         n47513, n47514, n47515, n47516, n47517, n47518, n47519, n47520,
         n47521, n47522, n47523, n47524, n47525, n47526, n47527, n47528,
         n47529, n47530, n47531, n47532, n47533, n47534, n47535, n47536,
         n47537, n47538, n47539, n47540, n47541, n47542, n47543, n47544,
         n47545, n47546, n47547, n47548, n47549, n47550, n47551, n47552,
         n47553, n47554, n47555, n47556, n47557, n47558, n47559, n47560,
         n47561, n47562, n47563, n47564, n47565, n47566, n47567, n47568,
         n47569, n47570, n47571, n47572, n47573, n47574, n47575, n47576,
         n47577, n47578, n47579, n47580, n47581, n47582, n47583, n47584,
         n47585, n47586, n47587, n47588, n47589, n47590, n47591, n47592,
         n47593, n47594, n47595, n47596, n47597, n47598, n47599, n47600,
         n47601, n47602, n47603, n47604, n47605, n47606, n47607, n47608,
         n47609, n47610, n47611, n47612, n47613, n47614, n47615, n47616,
         n47617, n47618, n47619, n47620, n47621, n47622, n47623, n47624,
         n47625, n47626, n47627, n47628, n47629, n47630, n47631, n47632,
         n47633, n47634, n47635, n47636, n47637, n47638, n47639, n47640,
         n47641, n47642, n47643, n47644, n47645, n47646, n47647, n47648,
         n47649, n47650, n47651, n47652, n47653, n47654, n47655, n47656,
         n47657, n47658, n47659, n47660, n47661, n47662, n47663, n47664,
         n47665, n47666, n47667, n47668, n47669, n47670, n47671, n47672,
         n47673, n47674, n47675, n47676, n47677, n47678, n47679, n47680,
         n47681, n47682, n47683, n47684, n47685, n47686, n47687, n47688,
         n47689, n47690, n47691, n47692, n47693, n47694, n47695, n47696,
         n47697, n47698, n47699, n47700, n47701, n47702, n47703, n47704,
         n47705, n47706, n47707, n47708, n47709, n47710, n47711, n47712,
         n47713, n47714, n47715, n47716, n47717, n47718, n47719, n47720,
         n47721, n47722, n47723, n47724, n47725, n47726, n47727, n47728,
         n47729, n47730, n47731, n47732, n47733, n47734, n47735, n47736,
         n47737, n47738, n47739, n47740, n47741, n47742, n47743, n47744,
         n47745, n47746, n47747, n47748, n47749, n47750, n47751, n47752,
         n47753, n47754, n47755, n47756, n47757, n47758, n47759, n47760,
         n47761, n47762, n47763, n47764, n47765, n47766, n47767, n47768,
         n47769, n47770, n47771, n47772, n47773, n47774, n47775, n47776,
         n47777, n47778, n47779, n47780, n47781, n47782, n47783, n47784,
         n47785, n47786, n47787, n47788, n47789, n47790, n47791, n47792,
         n47793, n47794, n47795, n47796, n47797, n47798, n47799, n47800,
         n47801, n47802, n47803, n47804, n47805, n47806, n47807, n47808,
         n47809, n47810, n47811, n47812, n47813, n47814, n47815, n47816,
         n47817, n47818, n47819, n47820, n47821, n47822, n47823, n47824,
         n47825, n47826, n47827, n47828, n47829, n47830, n47831, n47832,
         n47833, n47834, n47835, n47836, n47837, n47838, n47839, n47840,
         n47841, n47842, n47843, n47844, n47845, n47846, n47847, n47848,
         n47849, n47850, n47851, n47852, n47853, n47854, n47855, n47856,
         n47857, n47858, n47859, n47860, n47861, n47862, n47863, n47864,
         n47865, n47866, n47867, n47868, n47869, n47870, n47871, n47872,
         n47873, n47874, n47875, n47876, n47877, n47878, n47879, n47880,
         n47881, n47882, n47883, n47884, n47885, n47886, n47887, n47888,
         n47889, n47890, n47891, n47892, n47893, n47894, n47895, n47896,
         n47897, n47898, n47899, n47900, n47901, n47902, n47903, n47904,
         n47905, n47906, n47907, n47908, n47909, n47910, n47911, n47912,
         n47913, n47914, n47915, n47916, n47917, n47918, n47919, n47920,
         n47921, n47922, n47923, n47924, n47925, n47926, n47927, n47928,
         n47929, n47930, n47931, n47932, n47933, n47934, n47935, n47936,
         n47937, n47938, n47939, n47940, n47941, n47942, n47943, n47944,
         n47945, n47946, n47947, n47948, n47949, n47950, n47951, n47952,
         n47953, n47954, n47955, n47956, n47957, n47958, n47959, n47960,
         n47961, n47962, n47963, n47964, n47965, n47966, n47967, n47968,
         n47969, n47970, n47971, n47972, n47973, n47974, n47975, n47976,
         n47977, n47978, n47979, n47980, n47981, n47982, n47983, n47984,
         n47985, n47986, n47987, n47988, n47989, n47990, n47991, n47992,
         n47993, n47994, n47995, n47996, n47997, n47998, n47999, n48000,
         n48001, n48002, n48003, n48004, n48005, n48006, n48007, n48008,
         n48009, n48010, n48011, n48012, n48013, n48014, n48015, n48016,
         n48017, n48018, n48019, n48020, n48021, n48022, n48023, n48024,
         n48025, n48026, n48027, n48028, n48029, n48030, n48031, n48032,
         n48033, n48034, n48035, n48036, n48037, n48038, n48039, n48040,
         n48041, n48042, n48043, n48044, n48045, n48046, n48047, n48048,
         n48049, n48050, n48051, n48052, n48053, n48054, n48055, n48056,
         n48057, n48058, n48059, n48060, n48061, n48062, n48063, n48064,
         n48065, n48066, n48067, n48068, n48069, n48070, n48071, n48072,
         n48073, n48074, n48075, n48076, n48077, n48078, n48079, n48080,
         n48081, n48082, n48083, n48084, n48085, n48086, n48087, n48088,
         n48089, n48090, n48091, n48092, n48093, n48094, n48095, n48096,
         n48097, n48098, n48099, n48100, n48101, n48102, n48103, n48104,
         n48105, n48106, n48107, n48108, n48109, n48110, n48111, n48112,
         n48113, n48114, n48115, n48116, n48117, n48118, n48119, n48120,
         n48121, n48122, n48123, n48124, n48125, n48126, n48127, n48128,
         n48129, n48130, n48131, n48132, n48133, n48134, n48135, n48136,
         n48137, n48138, n48139, n48140, n48141, n48142, n48143, n48144,
         n48145, n48146, n48147, n48148, n48149, n48150, n48151, n48152,
         n48153, n48154, n48155, n48156, n48157, n48158, n48159, n48160,
         n48161, n48162, n48163, n48164, n48165, n48166, n48167, n48168,
         n48169, n48170, n48171, n48172, n48173, n48174, n48175, n48176,
         n48177, n48178, n48179, n48180, n48181, n48182, n48183, n48184,
         n48185, n48186, n48187, n48188, n48189, n48190, n48191, n48192,
         n48193, n48194, n48195, n48196, n48197, n48198, n48199, n48200,
         n48201, n48202, n48203, n48204, n48205, n48206, n48207, n48208,
         n48209, n48210, n48211, n48212, n48213, n48214, n48215, n48216,
         n48217, n48218, n48219, n48220, n48221, n48222, n48223, n48224,
         n48225, n48226, n48227, n48228, n48229, n48230, n48231, n48232,
         n48233, n48234, n48235, n48236, n48237, n48238, n48239, n48240,
         n48241, n48242, n48243, n48244, n48245, n48246, n48247, n48248,
         n48249, n48250, n48251, n48252, n48253, n48254, n48255, n48256,
         n48257, n48258, n48259, n48260, n48261, n48262, n48263, n48264,
         n48265, n48266, n48267, n48268, n48269, n48270, n48271, n48272,
         n48273, n48274, n48275, n48276, n48277, n48278, n48279, n48280,
         n48281, n48282, n48283, n48284, n48285, n48286, n48287, n48288,
         n48289, n48290, n48291, n48292, n48293, n48294, n48295, n48296,
         n48297, n48298, n48299, n48300, n48301, n48302, n48303, n48304,
         n48305, n48306, n48307, n48308, n48309, n48310, n48311, n48312,
         n48313, n48314, n48315, n48316, n48317, n48318, n48319, n48320,
         n48321, n48322, n48323, n48324, n48325, n48326, n48327, n48328,
         n48329, n48330, n48331, n48332, n48333, n48334, n48335, n48336,
         n48337, n48338, n48339, n48340, n48341, n48342, n48343, n48344,
         n48345, n48346, n48347, n48348, n48349, n48350, n48351, n48352,
         n48353, n48354, n48355, n48356, n48357, n48358, n48359, n48360,
         n48361, n48362, n48363, n48364, n48365, n48366, n48367, n48368,
         n48369, n48370, n48371, n48372, n48373, n48374, n48375, n48376,
         n48377, n48378, n48379, n48380, n48381, n48382, n48383, n48384,
         n48385, n48386, n48387, n48388, n48389, n48390, n48391, n48392,
         n48393, n48394, n48395, n48396, n48397, n48398, n48399, n48400,
         n48401, n48402, n48403, n48404, n48405, n48406, n48407, n48408,
         n48409, n48410, n48411, n48412, n48413, n48414, n48415, n48416,
         n48417, n48418, n48419, n48420, n48421, n48422, n48423, n48424,
         n48425, n48426, n48427, n48428, n48429, n48430, n48431, n48432,
         n48433, n48434, n48435, n48436, n48437, n48438, n48439, n48440,
         n48441, n48442, n48443, n48444, n48445, n48446, n48447, n48448,
         n48449, n48450, n48451, n48452, n48453, n48454, n48455, n48456,
         n48457, n48458, n48459, n48460, n48461, n48462, n48463, n48464,
         n48465, n48466, n48467, n48468, n48469, n48470, n48471, n48472,
         n48473, n48474, n48475, n48476, n48477, n48478, n48479, n48480,
         n48481, n48482, n48483, n48484, n48485, n48486, n48487, n48488,
         n48489, n48490, n48491, n48492, n48493, n48494, n48495, n48496,
         n48497, n48498, n48499, n48500, n48501, n48502, n48503, n48504,
         n48505, n48506, n48507, n48508, n48509, n48510, n48511, n48512,
         n48513, n48514, n48515, n48516, n48517, n48518, n48519, n48520,
         n48521, n48522, n48523, n48524, n48525, n48526, n48527, n48528,
         n48529, n48530, n48531, n48532, n48533, n48534, n48535, n48536,
         n48537, n48538, n48539, n48540, n48541, n48542, n48543, n48544,
         n48545, n48546, n48547, n48548, n48549, n48550, n48551, n48552,
         n48553, n48554, n48555, n48556, n48557, n48558, n48559, n48560,
         n48561, n48562, n48563, n48564, n48565, n48566, n48567, n48568,
         n48569, n48570, n48571, n48572, n48573, n48574, n48575, n48576,
         n48577, n48578, n48579, n48580, n48581, n48582, n48583, n48584,
         n48585, n48586, n48587, n48588, n48589, n48590, n48591, n48592,
         n48593, n48594, n48595, n48596, n48597, n48598, n48599, n48600,
         n48601, n48602, n48603, n48604, n48605, n48606, n48607, n48608,
         n48609, n48610, n48611, n48612, n48613, n48614, n48615, n48616,
         n48617, n48618, n48619, n48620, n48621, n48622, n48623, n48624,
         n48625, n48626, n48627, n48628, n48629, n48630, n48631, n48632,
         n48633, n48634, n48635, n48636, n48637, n48638, n48639, n48640,
         n48641, n48642, n48643, n48644, n48645, n48646, n48647, n48648,
         n48649, n48650, n48651, n48652, n48653, n48654, n48655, n48656,
         n48657, n48658, n48659, n48660, n48661, n48662, n48663, n48664,
         n48665, n48666, n48667, n48668, n48669, n48670, n48671, n48672,
         n48673, n48674, n48675, n48676, n48677, n48678, n48679, n48680,
         n48681, n48682, n48683, n48684, n48685, n48686, n48687, n48688,
         n48689, n48690, n48691, n48692, n48693, n48694, n48695, n48696,
         n48697, n48698, n48699, n48700, n48701, n48702, n48703, n48704,
         n48705, n48706, n48707, n48708, n48709, n48710, n48711, n48712,
         n48713, n48714, n48715, n48716, n48717, n48718, n48719, n48720,
         n48721, n48722, n48723, n48724, n48725, n48726, n48727, n48728,
         n48729, n48730, n48731, n48732, n48733, n48734, n48735, n48736,
         n48737, n48738, n48739, n48740, n48741, n48742, n48743, n48744,
         n48745, n48746, n48747, n48748, n48749, n48750, n48751, n48752,
         n48753, n48754, n48755, n48756, n48757, n48758, n48759, n48760,
         n48761, n48762, n48763, n48764, n48765, n48766, n48767, n48768,
         n48769, n48770, n48771, n48772, n48773, n48774, n48775, n48776,
         n48777, n48778, n48779, n48780, n48781, n48782, n48783, n48784,
         n48785, n48786, n48787, n48788, n48789, n48790, n48791, n48792,
         n48793, n48794, n48795, n48796, n48797, n48798, n48799, n48800,
         n48801, n48802, n48803, n48804, n48805, n48806, n48807, n48808,
         n48809, n48810, n48811, n48812, n48813, n48814, n48815, n48816,
         n48817, n48818, n48819, n48820, n48821, n48822, n48823, n48824,
         n48825, n48826, n48827, n48828, n48829, n48830, n48831, n48832,
         n48833, n48834, n48835, n48836, n48837, n48838, n48839, n48840,
         n48841, n48842, n48843, n48844, n48845, n48846, n48847, n48848,
         n48849, n48850, n48851, n48852, n48853, n48854, n48855, n48856,
         n48857, n48858, n48859, n48860, n48861, n48862, n48863, n48864,
         n48865, n48866, n48867, n48868, n48869, n48870, n48871, n48872,
         n48873, n48874, n48875, n48876, n48877, n48878, n48879, n48880,
         n48881, n48882, n48883, n48884, n48885, n48886, n48887, n48888,
         n48889, n48890, n48891, n48892, n48893, n48894, n48895, n48896,
         n48897, n48898, n48899, n48900, n48901, n48902, n48903, n48904,
         n48905, n48906, n48907, n48908, n48909, n48910, n48911, n48912,
         n48913, n48914, n48915, n48916, n48917, n48918, n48919, n48920,
         n48921, n48922, n48923, n48924, n48925, n48926, n48927, n48928,
         n48929, n48930, n48931, n48932, n48933, n48934, n48935, n48936,
         n48937, n48938, n48939, n48940, n48941, n48942, n48943, n48944,
         n48945, n48946, n48947, n48948, n48949, n48950, n48951, n48952,
         n48953, n48954, n48955, n48956, n48957, n48958, n48959, n48960,
         n48961, n48962, n48963, n48964, n48965, n48966, n48967, n48968,
         n48969, n48970, n48971, n48972, n48973, n48974, n48975, n48976,
         n48977, n48978, n48979, n48980, n48981, n48982, n48983, n48984,
         n48985, n48986, n48987, n48988, n48989, n48990, n48991, n48992,
         n48993, n48994, n48995, n48996, n48997, n48998, n48999, n49000,
         n49001, n49002, n49003, n49004, n49005, n49006, n49007, n49008,
         n49009, n49010, n49011, n49012, n49013, n49014, n49015, n49016,
         n49017, n49018, n49019, n49020, n49021, n49022, n49023, n49024,
         n49025, n49026, n49027, n49028, n49029, n49030, n49031, n49032,
         n49033, n49034, n49035, n49036, n49037, n49038, n49039, n49040,
         n49041, n49042, n49043, n49044, n49045, n49046, n49047, n49048,
         n49049, n49050, n49051, n49052, n49053, n49054, n49055, n49056,
         n49057, n49058, n49059, n49060, n49061, n49062, n49063, n49064,
         n49065, n49066, n49067, n49068, n49069, n49070, n49071, n49072,
         n49073, n49074, n49075, n49076, n49077, n49078, n49079, n49080,
         n49081, n49082, n49083, n49084, n49085, n49086, n49087, n49088,
         n49089, n49090, n49091, n49092, n49093, n49094, n49095, n49096,
         n49097, n49098, n49099, n49100, n49101, n49102, n49103, n49104,
         n49105, n49106, n49107, n49108, n49109, n49110, n49111, n49112,
         n49113, n49114, n49115, n49116, n49117, n49118, n49119, n49120,
         n49121, n49122, n49123, n49124, n49125, n49126, n49127, n49128,
         n49129, n49130, n49131, n49132, n49133, n49134, n49135, n49136,
         n49137, n49138, n49139, n49140, n49141, n49142, n49143, n49144,
         n49145, n49146, n49147, n49148, n49149, n49150, n49151, n49152,
         n49153, n49154, n49155, n49156, n49157, n49158, n49159, n49160,
         n49161, n49162, n49163, n49164, n49165, n49166, n49167, n49168,
         n49169, n49170, n49171, n49172, n49173, n49174, n49175, n49176,
         n49177, n49178, n49179, n49180, n49181, n49182, n49183, n49184,
         n49185, n49186, n49187, n49188, n49189, n49190, n49191, n49192,
         n49193, n49194, n49195, n49196, n49197, n49198, n49199, n49200,
         n49201, n49202, n49203, n49204, n49205, n49206, n49207, n49208,
         n49209, n49210, n49211, n49212, n49213, n49214, n49215, n49216,
         n49217, n49218, n49219, n49220, n49221, n49222, n49223, n49224,
         n49225, n49226, n49227, n49228, n49229, n49230, n49231, n49232,
         n49233, n49234, n49235, n49236, n49237, n49238, n49239, n49240,
         n49241, n49242, n49243, n49244, n49245, n49246, n49247, n49248,
         n49249, n49250, n49251, n49252, n49253, n49254, n49255, n49256,
         n49257, n49258, n49259, n49260, n49261, n49262, n49263, n49264,
         n49265, n49266, n49267, n49268, n49269, n49270, n49271, n49272,
         n49273, n49274, n49275, n49276, n49277, n49278, n49279, n49280,
         n49281, n49282, n49283, n49284, n49285, n49286, n49287, n49288,
         n49289, n49290, n49291, n49292, n49293, n49294, n49295, n49296,
         n49297, n49298, n49299, n49300, n49301, n49302, n49303, n49304,
         n49305, n49306, n49307, n49308, n49309, n49310, n49311, n49312,
         n49313, n49314, n49315, n49316, n49317, n49318, n49319, n49320,
         n49321, n49322, n49323, n49324, n49325, n49326, n49327, n49328,
         n49329, n49330, n49331, n49332, n49333, n49334, n49335, n49336,
         n49337, n49338, n49339, n49340, n49341, n49342, n49343, n49344,
         n49345, n49346, n49347, n49348, n49349, n49350, n49351, n49352,
         n49353, n49354, n49355, n49356, n49357, n49358, n49359, n49360,
         n49361, n49362, n49363, n49364, n49365, n49366, n49367, n49368,
         n49369, n49370, n49371, n49372, n49373, n49374, n49375, n49376,
         n49377, n49378, n49379, n49380, n49381, n49382, n49383, n49384,
         n49385, n49386, n49387, n49388, n49389, n49390, n49391, n49392,
         n49393, n49394, n49395, n49396, n49397, n49398, n49399, n49400,
         n49401, n49402, n49403, n49404, n49405, n49406, n49407, n49408,
         n49409, n49410, n49411, n49412, n49413, n49414, n49415, n49416,
         n49417, n49418, n49419, n49420, n49421, n49422, n49423, n49424,
         n49425, n49426, n49427, n49428, n49429, n49430, n49431, n49432,
         n49433, n49434, n49435, n49436, n49437, n49438, n49439, n49440,
         n49441, n49442, n49443, n49444, n49445, n49446, n49447, n49448,
         n49449, n49450, n49451, n49452, n49453, n49454, n49455, n49456,
         n49457, n49458, n49459, n49460, n49461, n49462, n49463, n49464,
         n49465, n49466, n49467, n49468, n49469, n49470, n49471, n49472,
         n49473, n49474, n49475, n49476, n49477, n49478, n49479, n49480,
         n49481, n49482, n49483, n49484, n49485, n49486, n49487, n49488,
         n49489, n49490, n49491, n49492, n49493, n49494, n49495, n49496,
         n49497, n49498, n49499, n49500, n49501, n49502, n49503, n49504,
         n49505, n49506, n49507, n49508, n49509, n49510, n49511, n49512,
         n49513, n49514, n49515, n49516, n49517, n49518, n49519, n49520,
         n49521, n49522, n49523, n49524, n49525, n49526, n49527, n49528,
         n49529, n49530, n49531, n49532, n49533, n49534, n49535, n49536,
         n49537, n49538, n49539, n49540, n49541, n49542, n49543, n49544,
         n49545, n49546, n49547, n49548, n49549, n49550, n49551, n49552,
         n49553, n49554, n49555, n49556, n49557, n49558, n49559, n49560,
         n49561, n49562, n49563, n49564, n49565, n49566, n49567, n49568,
         n49569, n49570, n49571, n49572, n49573, n49574, n49575, n49576,
         n49577, n49578, n49579, n49580, n49581, n49582, n49583, n49584,
         n49585, n49586, n49587, n49588, n49589, n49590, n49591, n49592,
         n49593, n49594, n49595, n49596, n49597, n49598, n49599, n49600,
         n49601, n49602, n49603, n49604, n49605, n49606, n49607, n49608,
         n49609, n49610, n49611, n49612, n49613, n49614, n49615, n49616,
         n49617, n49618, n49619, n49620, n49621, n49622, n49623, n49624,
         n49625, n49626, n49627, n49628, n49629, n49630, n49631, n49632,
         n49633, n49634, n49635, n49636, n49637, n49638, n49639, n49640,
         n49641, n49642, n49643, n49644, n49645, n49646, n49647, n49648,
         n49649, n49650, n49651, n49652, n49653, n49654, n49655, n49656,
         n49657, n49658, n49659, n49660, n49661, n49662, n49663, n49664,
         n49665, n49666, n49667, n49668, n49669, n49670, n49671, n49672,
         n49673, n49674, n49675, n49676, n49677, n49678, n49679, n49680,
         n49681, n49682, n49683, n49684, n49685, n49686, n49687, n49688,
         n49689, n49690, n49691, n49692, n49693, n49694, n49695, n49696,
         n49697, n49698, n49699, n49700, n49701, n49702, n49703, n49704,
         n49705, n49706, n49707, n49708, n49709, n49710, n49711, n49712,
         n49713, n49714, n49715, n49716, n49717, n49718, n49719, n49720,
         n49721, n49722, n49723, n49724, n49725, n49726, n49727, n49728,
         n49729, n49730, n49731, n49732, n49733, n49734, n49735, n49736,
         n49737, n49738, n49739, n49740, n49741, n49742, n49743, n49744,
         n49745, n49746, n49747, n49748, n49749, n49750, n49751, n49752,
         n49753, n49754, n49755, n49756, n49757, n49758, n49759, n49760,
         n49761, n49762, n49763, n49764, n49765, n49766, n49767, n49768,
         n49769, n49770, n49771, n49772, n49773, n49774, n49775, n49776,
         n49777, n49778, n49779, n49780, n49781, n49782, n49783, n49784,
         n49785, n49786, n49787, n49788, n49789, n49790, n49791, n49792,
         n49793, n49794, n49795, n49796, n49797, n49798, n49799, n49800,
         n49801, n49802, n49803, n49804, n49805, n49806, n49807, n49808,
         n49809, n49810, n49811, n49812, n49813, n49814, n49815, n49816,
         n49817, n49818, n49819, n49820, n49821, n49822, n49823, n49824,
         n49825, n49826, n49827, n49828, n49829, n49830, n49831, n49832,
         n49833, n49834, n49835, n49836, n49837, n49838, n49839, n49840,
         n49841, n49842, n49843, n49844, n49845, n49846, n49847, n49848,
         n49849, n49850, n49851, n49852, n49853, n49854, n49855, n49856,
         n49857, n49858, n49859, n49860, n49861, n49862, n49863, n49864,
         n49865, n49866, n49867, n49868, n49869, n49870, n49871, n49872,
         n49873, n49874, n49875, n49876, n49877, n49878, n49879, n49880,
         n49881, n49882, n49883, n49884, n49885, n49886, n49887, n49888,
         n49889, n49890, n49891, n49892, n49893, n49894, n49895, n49896,
         n49897, n49898, n49899, n49900, n49901, n49902, n49903, n49904,
         n49905, n49906, n49907, n49908, n49909, n49910, n49911, n49912,
         n49913, n49914, n49915, n49916, n49917, n49918, n49919, n49920,
         n49921, n49922, n49923, n49924, n49925, n49926, n49927, n49928,
         n49929, n49930, n49931, n49932, n49933, n49934, n49935, n49936,
         n49937, n49938, n49939, n49940, n49941, n49942, n49943, n49944,
         n49945, n49946, n49947, n49948, n49949, n49950, n49951, n49952,
         n49953, n49954, n49955, n49956, n49957, n49958, n49959, n49960,
         n49961, n49962, n49963, n49964, n49965, n49966, n49967, n49968,
         n49969, n49970, n49971, n49972, n49973, n49974, n49975, n49976,
         n49977, n49978, n49979, n49980, n49981, n49982, n49983, n49984,
         n49985, n49986, n49987, n49988, n49989, n49990, n49991, n49992,
         n49993, n49994, n49995, n49996, n49997, n49998, n49999, n50000,
         n50001, n50002, n50003, n50004, n50005, n50006, n50007, n50008,
         n50009, n50010, n50011, n50012, n50013, n50014, n50015, n50016,
         n50017, n50018, n50019, n50020, n50021, n50022, n50023, n50024,
         n50025, n50026, n50027, n50028, n50029, n50030, n50031, n50032,
         n50033, n50034, n50035, n50036, n50037, n50038, n50039, n50040,
         n50041, n50042, n50043, n50044, n50045, n50046, n50047, n50048,
         n50049, n50050, n50051, n50052, n50053, n50054, n50055, n50056,
         n50057, n50058, n50059, n50060, n50061, n50062, n50063, n50064,
         n50065, n50066, n50067, n50068, n50069, n50070, n50071, n50072,
         n50073, n50074, n50075, n50076, n50077, n50078, n50079, n50080,
         n50081, n50082, n50083, n50084, n50085, n50086, n50087, n50088,
         n50089, n50090, n50091, n50092, n50093, n50094, n50095, n50096,
         n50097, n50098, n50099, n50100, n50101, n50102, n50103, n50104,
         n50105, n50106, n50107, n50108, n50109, n50110, n50111, n50112,
         n50113, n50114, n50115, n50116, n50117, n50118, n50119, n50120,
         n50121, n50122, n50123, n50124, n50125, n50126, n50127, n50128,
         n50129, n50130, n50131, n50132, n50133, n50134, n50135, n50136,
         n50137, n50138, n50139, n50140, n50141, n50142, n50143, n50144,
         n50145, n50146, n50147, n50148, n50149, n50150, n50151, n50152,
         n50153, n50154, n50155, n50156, n50157, n50158, n50159, n50160,
         n50161, n50162, n50163, n50164, n50165, n50166, n50167, n50168,
         n50169, n50170, n50171, n50172, n50173, n50174, n50175, n50176,
         n50177, n50178, n50179, n50180, n50181, n50182, n50183, n50184,
         n50185, n50186, n50187, n50188, n50189, n50190, n50191, n50192,
         n50193, n50194, n50195, n50196, n50197, n50198, n50199, n50200,
         n50201, n50202, n50203, n50204, n50205, n50206, n50207, n50208,
         n50209, n50210, n50211, n50212, n50213, n50214, n50215, n50216,
         n50217, n50218, n50219, n50220, n50221, n50222, n50223, n50224,
         n50225, n50226, n50227, n50228, n50229, n50230, n50231, n50232,
         n50233, n50234, n50235, n50236, n50237, n50238, n50239, n50240,
         n50241, n50242, n50243, n50244, n50245, n50246, n50247, n50248,
         n50249, n50250, n50251, n50252, n50253, n50254, n50255, n50256,
         n50257, n50258, n50259, n50260, n50261, n50262, n50263, n50264,
         n50265, n50266, n50267, n50268, n50269, n50270, n50271, n50272,
         n50273, n50274, n50275, n50276, n50277, n50278, n50279, n50280,
         n50281, n50282, n50283, n50284, n50285, n50286, n50287, n50288,
         n50289, n50290, n50291, n50292, n50293, n50294, n50295, n50296,
         n50297, n50298, n50299, n50300, n50301, n50302, n50303, n50304,
         n50305, n50306, n50307, n50308, n50309, n50310, n50311, n50312,
         n50313, n50314, n50315, n50316, n50317, n50318, n50319, n50320,
         n50321, n50322, n50323, n50324, n50325, n50326, n50327, n50328,
         n50329, n50330, n50331, n50332, n50333, n50334, n50335, n50336,
         n50337, n50338, n50339, n50340, n50341, n50342, n50343, n50344,
         n50345, n50346, n50347, n50348, n50349, n50350, n50351, n50352,
         n50353, n50354, n50355, n50356, n50357, n50358, n50359, n50360,
         n50361, n50362, n50363, n50364, n50365, n50366, n50367, n50368,
         n50369, n50370, n50371, n50372, n50373, n50374, n50375, n50376,
         n50377, n50378, n50379, n50380, n50381, n50382, n50383, n50384,
         n50385, n50386, n50387, n50388, n50389, n50390, n50391, n50392,
         n50393, n50394, n50395, n50396, n50397, n50398, n50399, n50400,
         n50401, n50402, n50403, n50404, n50405, n50406, n50407, n50408,
         n50409, n50410, n50411, n50412, n50413, n50414, n50415, n50416,
         n50417, n50418, n50419, n50420, n50421, n50422, n50423, n50424,
         n50425, n50426, n50427, n50428, n50429, n50430, n50431, n50432,
         n50433, n50434, n50435, n50436, n50437, n50438, n50439, n50440,
         n50441, n50442, n50443, n50444, n50445, n50446, n50447, n50448,
         n50449, n50450, n50451, n50452, n50453, n50454, n50455, n50456,
         n50457, n50458, n50459, n50460, n50461, n50462, n50463, n50464,
         n50465, n50466, n50467, n50468, n50469, n50470, n50471, n50472,
         n50473, n50474, n50475, n50476, n50477, n50478, n50479, n50480,
         n50481, n50482, n50483, n50484, n50485, n50486, n50487, n50488,
         n50489, n50490, n50491, n50492, n50493, n50494, n50495, n50496,
         n50497, n50498, n50499, n50500, n50501, n50502, n50503, n50504,
         n50505, n50506, n50507, n50508, n50509, n50510, n50511, n50512,
         n50513, n50514, n50515, n50516, n50517, n50518, n50519, n50520,
         n50521, n50522, n50523, n50524, n50525, n50526, n50527, n50528,
         n50529, n50530, n50531, n50532, n50533, n50534, n50535, n50536,
         n50537, n50538, n50539, n50540, n50541, n50542, n50543, n50544,
         n50545, n50546, n50547, n50548, n50549, n50550, n50551, n50552,
         n50553, n50554, n50555, n50556, n50557, n50558, n50559, n50560,
         n50561, n50562, n50563, n50564, n50565, n50566, n50567, n50568,
         n50569, n50570, n50571, n50572, n50573, n50574, n50575, n50576,
         n50577, n50578, n50579, n50580, n50581, n50582, n50583, n50584,
         n50585, n50586, n50587, n50588, n50589, n50590, n50591, n50592,
         n50593, n50594, n50595, n50596, n50597, n50598, n50599, n50600,
         n50601, n50602, n50603, n50604, n50605, n50606, n50607, n50608,
         n50609, n50610, n50611, n50612, n50613, n50614, n50615, n50616,
         n50617, n50618, n50619, n50620, n50621, n50622, n50623, n50624,
         n50625, n50626, n50627, n50628, n50629, n50630, n50631, n50632,
         n50633, n50634, n50635, n50636, n50637, n50638, n50639, n50640,
         n50641, n50642, n50643, n50644, n50645, n50646, n50647, n50648,
         n50649, n50650, n50651, n50652, n50653, n50654, n50655, n50656,
         n50657, n50658, n50659, n50660, n50661, n50662, n50663, n50664,
         n50665, n50666, n50667, n50668, n50669, n50670, n50671, n50672,
         n50673, n50674, n50675, n50676, n50677, n50678, n50679, n50680,
         n50681, n50682, n50683, n50684, n50685, n50686, n50687, n50688,
         n50689, n50690, n50691, n50692, n50693, n50694, n50695, n50696,
         n50697, n50698, n50699, n50700, n50701, n50702, n50703, n50704,
         n50705, n50706, n50707, n50708, n50709, n50710, n50711, n50712,
         n50713, n50714, n50715, n50716, n50717, n50718, n50719, n50720,
         n50721, n50722, n50723, n50724, n50725, n50726, n50727, n50728,
         n50729, n50730, n50731, n50732, n50733, n50734, n50735, n50736,
         n50737, n50738, n50739, n50740, n50741, n50742, n50743, n50744,
         n50745, n50746, n50747, n50748, n50749, n50750, n50751, n50752,
         n50753, n50754, n50755, n50756, n50757, n50758, n50759, n50760,
         n50761, n50762, n50763, n50764, n50765, n50766, n50767, n50768,
         n50769, n50770, n50771, n50772, n50773, n50774, n50775, n50776,
         n50777, n50778, n50779, n50780, n50781, n50782, n50783, n50784,
         n50785, n50786, n50787, n50788, n50789, n50790, n50791, n50792,
         n50793, n50794, n50795, n50796, n50797, n50798, n50799, n50800,
         n50801, n50802, n50803, n50804, n50805, n50806, n50807, n50808,
         n50809, n50810, n50811, n50812, n50813, n50814, n50815, n50816,
         n50817, n50818, n50819, n50820, n50821, n50822, n50823, n50824,
         n50825, n50826, n50827, n50828, n50829, n50830, n50831, n50832,
         n50833, n50834, n50835, n50836, n50837, n50838, n50839, n50840,
         n50841, n50842, n50843, n50844, n50845, n50846, n50847, n50848,
         n50849, n50850, n50851, n50852, n50853, n50854, n50855, n50856,
         n50857, n50858, n50859, n50860, n50861, n50862, n50863, n50864,
         n50865, n50866, n50867, n50868, n50869, n50870, n50871, n50872,
         n50873, n50874, n50875, n50876, n50877, n50878, n50879, n50880,
         n50881, n50882, n50883, n50884, n50885, n50886, n50887, n50888,
         n50889, n50890, n50891, n50892, n50893, n50894, n50895, n50896,
         n50897, n50898, n50899, n50900, n50901, n50902, n50903, n50904,
         n50905, n50906, n50907, n50908, n50909, n50910, n50911, n50912,
         n50913, n50914, n50915, n50916, n50917, n50918, n50919, n50920,
         n50921, n50922, n50923, n50924, n50925, n50926, n50927, n50928,
         n50929, n50930, n50931, n50932, n50933, n50934, n50935, n50936,
         n50937, n50938, n50939, n50940, n50941, n50942, n50943, n50944,
         n50945, n50946, n50947, n50948, n50949, n50950, n50951, n50952,
         n50953, n50954, n50955, n50956, n50957, n50958, n50959, n50960,
         n50961, n50962, n50963, n50964, n50965, n50966, n50967, n50968,
         n50969, n50970, n50971, n50972, n50973, n50974, n50975, n50976,
         n50977, n50978, n50979, n50980, n50981, n50982, n50983, n50984,
         n50985, n50986, n50987, n50988, n50989, n50990, n50991, n50992,
         n50993, n50994, n50995, n50996, n50997, n50998, n50999, n51000,
         n51001, n51002, n51003, n51004, n51005, n51006, n51007, n51008,
         n51009, n51010, n51011, n51012, n51013, n51014, n51015, n51016,
         n51017, n51018, n51019, n51020, n51021, n51022, n51023, n51024,
         n51025, n51026, n51027, n51028, n51029, n51030, n51031, n51032,
         n51033, n51034, n51035, n51036, n51037, n51038, n51039, n51040,
         n51041, n51042, n51043, n51044, n51045, n51046, n51047, n51048,
         n51049, n51050, n51051, n51052, n51053, n51054, n51055, n51056,
         n51057, n51058, n51059, n51060, n51061, n51062, n51063, n51064,
         n51065, n51066, n51067, n51068, n51069, n51070, n51071, n51072,
         n51073, n51074, n51075, n51076, n51077, n51078, n51079, n51080,
         n51081, n51082, n51083, n51084, n51085, n51086, n51087, n51088,
         n51089, n51090, n51091, n51092, n51093, n51094, n51095, n51096,
         n51097, n51098, n51099, n51100, n51101, n51102, n51103, n51104,
         n51105, n51106, n51107, n51108, n51109, n51110, n51111, n51112,
         n51113, n51114, n51115, n51116, n51117, n51118, n51119, n51120,
         n51121, n51122, n51123, n51124, n51125, n51126, n51127, n51128,
         n51129, n51130, n51131, n51132, n51133, n51134, n51135, n51136,
         n51137, n51138, n51139, n51140, n51141, n51142, n51143, n51144,
         n51145, n51146, n51147, n51148, n51149, n51150, n51151, n51152,
         n51153, n51154, n51155, n51156, n51157, n51158, n51159, n51160,
         n51161, n51162, n51163, n51164, n51165, n51166, n51167, n51168,
         n51169, n51170, n51171, n51172, n51173, n51174, n51175, n51176,
         n51177, n51178, n51179, n51180, n51181, n51182, n51183, n51184,
         n51185, n51186, n51187, n51188, n51189, n51190, n51191, n51192,
         n51193, n51194, n51195, n51196, n51197, n51198, n51199, n51200,
         n51201, n51202, n51203, n51204, n51205, n51206, n51207, n51208,
         n51209, n51210, n51211, n51212, n51213, n51214, n51215, n51216,
         n51217, n51218, n51219, n51220, n51221, n51222, n51223, n51224,
         n51225, n51226, n51227, n51228, n51229, n51230, n51231, n51232,
         n51233, n51234, n51235, n51236, n51237, n51238, n51239, n51240,
         n51241, n51242, n51243, n51244, n51245, n51246, n51247, n51248,
         n51249, n51250, n51251, n51252, n51253, n51254, n51255, n51256,
         n51257, n51258, n51259, n51260, n51261, n51262, n51263, n51264,
         n51265, n51266, n51267, n51268, n51269, n51270, n51271, n51272,
         n51273, n51274, n51275, n51276, n51277, n51278, n51279, n51280,
         n51281, n51282, n51283, n51284, n51285, n51286, n51287, n51288,
         n51289, n51290, n51291, n51292, n51293, n51294, n51295, n51296,
         n51297, n51298, n51299, n51300, n51301, n51302, n51303, n51304,
         n51305, n51306, n51307, n51308, n51309, n51310, n51311, n51312,
         n51313, n51314, n51315, n51316, n51317, n51318, n51319, n51320,
         n51321, n51322, n51323, n51324, n51325, n51326, n51327, n51328,
         n51329, n51330, n51331, n51332, n51333, n51334, n51335, n51336,
         n51337, n51338, n51339, n51340, n51341, n51342, n51343, n51344,
         n51345, n51346, n51347, n51348, n51349, n51350, n51351, n51352,
         n51353, n51354, n51355, n51356, n51357, n51358, n51359, n51360,
         n51361, n51362, n51363, n51364, n51365, n51366, n51367, n51368,
         n51369, n51370, n51371, n51372, n51373, n51374, n51375, n51376,
         n51377, n51378, n51379, n51380, n51381, n51382, n51383, n51384,
         n51385, n51386, n51387, n51388, n51389, n51390, n51391, n51392,
         n51393, n51394, n51395, n51396, n51397, n51398, n51399, n51400,
         n51401, n51402, n51403, n51404, n51405, n51406, n51407, n51408,
         n51409, n51410, n51411, n51412, n51413, n51414, n51415, n51416,
         n51417, n51418, n51419, n51420, n51421, n51422, n51423, n51424,
         n51425, n51426, n51427, n51428, n51429, n51430, n51431, n51432,
         n51433, n51434, n51435, n51436, n51437, n51438, n51439, n51440,
         n51441, n51442, n51443, n51444, n51445, n51446, n51447, n51448,
         n51449, n51450, n51451, n51452, n51453, n51454, n51455, n51456,
         n51457, n51458, n51459, n51460, n51461, n51462, n51463, n51464,
         n51465, n51466, n51467, n51468, n51469, n51470, n51471, n51472,
         n51473, n51474, n51475, n51476, n51477, n51478, n51479, n51480,
         n51481, n51482, n51483, n51484, n51485, n51486, n51487, n51488,
         n51489, n51490, n51491, n51492, n51493, n51494, n51495, n51496,
         n51497, n51498, n51499, n51500, n51501, n51502, n51503, n51504,
         n51505, n51506, n51507, n51508, n51509, n51510, n51511, n51512,
         n51513, n51514, n51515, n51516, n51517, n51518, n51519, n51520,
         n51521, n51522, n51523, n51524, n51525, n51526, n51527, n51528,
         n51529, n51530, n51531, n51532, n51533, n51534, n51535, n51536,
         n51537, n51538, n51539, n51540, n51541, n51542, n51543, n51544,
         n51545, n51546, n51547, n51548, n51549, n51550, n51551, n51552,
         n51553, n51554, n51555, n51556, n51557, n51558, n51559, n51560,
         n51561, n51562, n51563, n51564, n51565, n51566, n51567, n51568,
         n51569, n51570, n51571, n51572, n51573, n51574, n51575, n51576,
         n51577, n51578, n51579, n51580, n51581, n51582, n51583, n51584,
         n51585, n51586, n51587, n51588, n51589, n51590, n51591, n51592,
         n51593, n51594, n51595, n51596, n51597, n51598, n51599, n51600,
         n51601, n51602, n51603, n51604, n51605, n51606, n51607, n51608,
         n51609, n51610, n51611, n51612, n51613, n51614, n51615, n51616,
         n51617, n51618, n51619, n51620, n51621, n51622, n51623, n51624,
         n51625, n51626, n51627, n51628, n51629, n51630, n51631, n51632,
         n51633, n51634, n51635, n51636, n51637, n51638, n51639, n51640,
         n51641, n51642, n51643, n51644, n51645, n51646, n51647, n51648,
         n51649, n51650, n51651, n51652, n51653, n51654, n51655, n51656,
         n51657, n51658, n51659, n51660, n51661, n51662, n51663, n51664,
         n51665, n51666, n51667, n51668, n51669, n51670, n51671, n51672,
         n51673, n51674, n51675, n51676, n51677, n51678, n51679, n51680,
         n51681, n51682, n51683, n51684, n51685, n51686, n51687, n51688,
         n51689, n51690, n51691, n51692, n51693, n51694, n51695, n51696,
         n51697, n51698, n51699, n51700, n51701, n51702, n51703, n51704,
         n51705, n51706, n51707, n51708, n51709, n51710, n51711, n51712,
         n51713, n51714, n51715, n51716, n51717, n51718, n51719, n51720,
         n51721, n51722, n51723, n51724, n51725, n51726, n51727, n51728,
         n51729, n51730, n51731, n51732, n51733, n51734, n51735, n51736,
         n51737, n51738, n51739, n51740, n51741, n51742, n51743, n51744,
         n51745, n51746, n51747, n51748, n51749, n51750, n51751, n51752,
         n51753, n51754, n51755, n51756, n51757, n51758, n51759, n51760,
         n51761, n51762, n51763, n51764, n51765, n51766, n51767, n51768,
         n51769, n51770, n51771, n51772, n51773, n51774, n51775, n51776,
         n51777, n51778, n51779, n51780, n51781, n51782, n51783, n51784,
         n51785, n51786, n51787, n51788, n51789, n51790, n51791, n51792,
         n51793, n51794, n51795, n51796, n51797, n51798, n51799, n51800,
         n51801, n51802, n51803, n51804, n51805, n51806, n51807, n51808,
         n51809, n51810, n51811, n51812, n51813, n51814, n51815, n51816,
         n51817, n51818, n51819, n51820, n51821, n51822, n51823, n51824,
         n51825, n51826, n51827, n51828, n51829, n51830, n51831, n51832,
         n51833, n51834, n51835, n51836, n51837, n51838, n51839, n51840,
         n51841, n51842, n51843, n51844, n51845, n51846, n51847, n51848,
         n51849, n51850, n51851, n51852, n51853, n51854, n51855, n51856,
         n51857, n51858, n51859, n51860, n51861, n51862, n51863, n51864,
         n51865, n51866, n51867, n51868, n51869, n51870, n51871, n51872,
         n51873, n51874, n51875, n51876, n51877, n51878, n51879, n51880,
         n51881, n51882, n51883, n51884, n51885, n51886, n51887, n51888,
         n51889, n51890, n51891, n51892, n51893, n51894, n51895, n51896,
         n51897, n51898, n51899, n51900, n51901, n51902, n51903, n51904,
         n51905, n51906, n51907, n51908, n51909, n51910, n51911, n51912,
         n51913, n51914, n51915, n51916, n51917, n51918, n51919, n51920,
         n51921, n51922, n51923, n51924, n51925, n51926, n51927, n51928,
         n51929, n51930, n51931, n51932, n51933, n51934, n51935, n51936,
         n51937, n51938, n51939, n51940, n51941, n51942, n51943, n51944,
         n51945, n51946, n51947, n51948, n51949, n51950, n51951, n51952,
         n51953, n51954, n51955, n51956, n51957, n51958, n51959, n51960,
         n51961, n51962, n51963, n51964, n51965, n51966, n51967, n51968,
         n51969, n51970, n51971, n51972, n51973, n51974, n51975, n51976,
         n51977, n51978, n51979, n51980, n51981, n51982, n51983, n51984,
         n51985, n51986, n51987, n51988, n51989, n51990, n51991, n51992,
         n51993, n51994, n51995, n51996, n51997, n51998, n51999, n52000,
         n52001, n52002, n52003, n52004, n52005, n52006, n52007, n52008,
         n52009, n52010, n52011, n52012, n52013, n52014, n52015, n52016,
         n52017, n52018, n52019, n52020, n52021, n52022, n52023, n52024,
         n52025, n52026, n52027, n52028, n52029, n52030, n52031, n52032,
         n52033, n52034, n52035, n52036, n52037, n52038, n52039, n52040,
         n52041, n52042, n52043, n52044, n52045, n52046, n52047, n52048,
         n52049, n52050, n52051, n52052, n52053, n52054, n52055, n52056,
         n52057, n52058, n52059, n52060, n52061, n52062, n52063, n52064,
         n52065, n52066, n52067, n52068, n52069, n52070, n52071, n52072,
         n52073, n52074, n52075, n52076, n52077, n52078, n52079, n52080,
         n52081, n52082, n52083, n52084, n52085, n52086, n52087, n52088,
         n52089, n52090, n52091, n52092, n52093, n52094, n52095, n52096,
         n52097, n52098, n52099, n52100, n52101, n52102, n52103, n52104,
         n52105, n52106, n52107, n52108, n52109, n52110, n52111, n52112,
         n52113, n52114, n52115, n52116, n52117, n52118, n52119, n52120,
         n52121, n52122, n52123, n52124, n52125, n52126, n52127, n52128,
         n52129, n52130, n52131, n52132, n52133, n52134, n52135, n52136,
         n52137, n52138, n52139, n52140, n52141, n52142, n52143, n52144,
         n52145, n52146, n52147, n52148, n52149, n52150, n52151, n52152,
         n52153, n52154, n52155, n52156, n52157, n52158, n52159, n52160,
         n52161, n52162, n52163, n52164, n52165, n52166, n52167, n52168,
         n52169, n52170, n52171, n52172, n52173, n52174, n52175, n52176,
         n52177, n52178, n52179, n52180, n52181, n52182, n52183, n52184,
         n52185, n52186, n52187, n52188, n52189, n52190, n52191, n52192,
         n52193, n52194, n52195, n52196, n52197, n52198, n52199, n52200,
         n52201, n52202, n52203, n52204, n52205, n52206, n52207, n52208,
         n52209, n52210, n52211, n52212, n52213, n52214, n52215, n52216,
         n52217, n52218, n52219, n52220, n52221, n52222, n52223, n52224,
         n52225, n52226, n52227, n52228, n52229, n52230, n52231, n52232,
         n52233, n52234, n52235, n52236, n52237, n52238, n52239, n52240,
         n52241, n52242, n52243, n52244, n52245, n52246, n52247, n52248,
         n52249, n52250, n52251, n52252, n52253, n52254, n52255, n52256,
         n52257, n52258, n52259, n52260, n52261, n52262, n52263, n52264,
         n52265, n52266, n52267, n52268, n52269, n52270, n52271, n52272,
         n52273, n52274, n52275, n52276, n52277, n52278, n52279, n52280,
         n52281, n52282, n52283, n52284, n52285, n52286, n52287, n52288,
         n52289, n52290, n52291, n52292, n52293, n52294, n52295, n52296,
         n52297, n52298, n52299, n52300, n52301, n52302, n52303, n52304,
         n52305, n52306, n52307, n52308, n52309, n52310, n52311, n52312,
         n52313, n52314, n52315, n52316, n52317, n52318, n52319, n52320,
         n52321, n52322, n52323, n52324, n52325, n52326, n52327, n52328,
         n52329, n52330, n52331, n52332, n52333, n52334, n52335, n52336,
         n52337, n52338, n52339, n52340, n52341, n52342, n52343, n52344,
         n52345, n52346, n52347, n52348, n52349, n52350, n52351, n52352,
         n52353, n52354, n52355, n52356, n52357, n52358, n52359, n52360,
         n52361, n52362, n52363, n52364, n52365, n52366, n52367, n52368,
         n52369, n52370, n52371, n52372, n52373, n52374, n52375, n52376,
         n52377, n52378, n52379, n52380, n52381, n52382, n52383, n52384,
         n52385, n52386, n52387, n52388, n52389, n52390, n52391, n52392,
         n52393, n52394, n52395, n52396, n52397, n52398, n52399, n52400,
         n52401, n52402, n52403, n52404, n52405, n52406, n52407, n52408,
         n52409, n52410, n52411, n52412, n52413, n52414, n52415, n52416,
         n52417, n52418, n52419, n52420, n52421, n52422, n52423, n52424,
         n52425, n52426, n52427, n52428, n52429, n52430, n52431, n52432,
         n52433, n52434, n52435, n52436, n52437, n52438, n52439, n52440,
         n52441, n52442, n52443, n52444, n52445, n52446, n52447, n52448,
         n52449, n52450, n52451, n52452, n52453, n52454, n52455, n52456,
         n52457, n52458, n52459, n52460, n52461, n52462, n52463, n52464,
         n52465, n52466, n52467, n52468, n52469, n52470, n52471, n52472,
         n52473, n52474, n52475, n52476, n52477, n52478, n52479, n52480,
         n52481, n52482, n52483, n52484, n52485, n52486, n52487, n52488,
         n52489, n52490, n52491, n52492, n52493, n52494, n52495, n52496,
         n52497, n52498, n52499, n52500, n52501, n52502, n52503, n52504,
         n52505, n52506, n52507, n52508, n52509, n52510, n52511, n52512,
         n52513, n52514, n52515, n52516, n52517, n52518, n52519, n52520,
         n52521, n52522, n52523, n52524, n52525, n52526, n52527, n52528,
         n52529, n52530, n52531, n52532, n52533, n52534, n52535, n52536,
         n52537, n52538, n52539, n52540, n52541, n52542, n52543, n52544,
         n52545, n52546, n52547, n52548, n52549, n52550, n52551, n52552,
         n52553, n52554, n52555, n52556, n52557, n52558, n52559, n52560,
         n52561, n52562, n52563, n52564, n52565, n52566, n52567, n52568,
         n52569, n52570, n52571, n52572, n52573, n52574, n52575, n52576,
         n52577, n52578, n52579, n52580, n52581, n52582, n52583, n52584,
         n52585, n52586, n52587, n52588, n52589, n52590, n52591, n52592,
         n52593, n52594, n52595, n52596, n52597, n52598, n52599, n52600,
         n52601, n52602, n52603, n52604, n52605, n52606, n52607, n52608,
         n52609, n52610, n52611, n52612, n52613, n52614, n52615, n52616,
         n52617, n52618, n52619, n52620, n52621, n52622, n52623, n52624,
         n52625, n52626, n52627, n52628, n52629, n52630, n52631, n52632,
         n52633, n52634, n52635, n52636, n52637, n52638, n52639, n52640,
         n52641, n52642, n52643, n52644, n52645, n52646, n52647, n52648,
         n52649, n52650, n52651, n52652, n52653, n52654, n52655, n52656,
         n52657, n52658, n52659, n52660, n52661, n52662, n52663, n52664,
         n52665, n52666, n52667, n52668, n52669, n52670, n52671, n52672,
         n52673, n52674, n52675, n52676, n52677, n52678, n52679, n52680,
         n52681, n52682, n52683, n52684, n52685, n52686, n52687, n52688,
         n52689, n52690, n52691, n52692, n52693, n52694, n52695, n52696,
         n52697, n52698, n52699, n52700, n52701, n52702, n52703, n52704,
         n52705, n52706, n52707, n52708, n52709, n52710, n52711, n52712,
         n52713, n52714, n52715, n52716, n52717, n52718, n52719, n52720,
         n52721, n52722, n52723, n52724, n52725, n52726, n52727, n52728,
         n52729, n52730, n52731, n52732, n52733, n52734, n52735, n52736,
         n52737, n52738, n52739, n52740, n52741, n52742, n52743, n52744,
         n52745, n52746, n52747, n52748, n52749, n52750, n52751, n52752,
         n52753, n52754, n52755, n52756, n52757, n52758, n52759, n52760,
         n52761, n52762, n52763, n52764, n52765, n52766, n52767, n52768,
         n52769, n52770, n52771, n52772, n52773, n52774, n52775, n52776,
         n52777, n52778, n52779, n52780, n52781, n52782, n52783, n52784,
         n52785, n52786, n52787, n52788, n52789, n52790, n52791, n52792,
         n52793, n52794, n52795, n52796, n52797, n52798, n52799, n52800,
         n52801, n52802, n52803, n52804, n52805, n52806, n52807, n52808,
         n52809, n52810, n52811, n52812, n52813, n52814, n52815, n52816,
         n52817, n52818, n52819, n52820, n52821, n52822, n52823, n52824,
         n52825, n52826, n52827, n52828, n52829, n52830, n52831, n52832,
         n52833, n52834, n52835, n52836, n52837, n52838, n52839, n52840,
         n52841, n52842, n52843, n52844, n52845, n52846, n52847, n52848,
         n52849, n52850, n52851, n52852, n52853, n52854, n52855, n52856,
         n52857, n52858, n52859, n52860, n52861, n52862, n52863, n52864,
         n52865, n52866, n52867, n52868, n52869, n52870, n52871, n52872,
         n52873, n52874, n52875, n52876, n52877, n52878, n52879, n52880,
         n52881, n52882, n52883, n52884, n52885, n52886, n52887, n52888,
         n52889, n52890, n52891, n52892, n52893, n52894, n52895, n52896,
         n52897, n52898, n52899, n52900, n52901, n52902, n52903, n52904,
         n52905, n52906, n52907, n52908, n52909, n52910, n52911, n52912,
         n52913, n52914, n52915, n52916, n52917, n52918, n52919, n52920,
         n52921, n52922, n52923, n52924, n52925, n52926, n52927, n52928,
         n52929, n52930, n52931, n52932, n52933, n52934, n52935, n52936,
         n52937, n52938, n52939, n52940, n52941, n52942, n52943, n52944,
         n52945, n52946, n52947, n52948, n52949, n52950, n52951, n52952,
         n52953, n52954, n52955, n52956, n52957, n52958, n52959, n52960,
         n52961, n52962, n52963, n52964, n52965, n52966, n52967, n52968,
         n52969, n52970, n52971, n52972, n52973, n52974, n52975, n52976,
         n52977, n52978, n52979, n52980, n52981, n52982, n52983, n52984,
         n52985, n52986, n52987, n52988, n52989, n52990, n52991, n52992,
         n52993, n52994, n52995, n52996, n52997, n52998, n52999, n53000,
         n53001, n53002, n53003, n53004, n53005, n53006, n53007, n53008,
         n53009, n53010, n53011, n53012, n53013, n53014, n53015, n53016,
         n53017, n53018, n53019, n53020, n53021, n53022, n53023, n53024,
         n53025, n53026, n53027, n53028, n53029, n53030, n53031, n53032,
         n53033, n53034, n53035, n53036, n53037, n53038, n53039, n53040,
         n53041, n53042, n53043, n53044, n53045, n53046, n53047, n53048,
         n53049, n53050, n53051, n53052, n53053, n53054, n53055, n53056,
         n53057, n53058, n53059, n53060, n53061, n53062, n53063, n53064,
         n53065, n53066, n53067, n53068, n53069, n53070, n53071, n53072,
         n53073, n53074, n53075, n53076, n53077, n53078, n53079, n53080,
         n53081, n53082, n53083, n53084, n53085, n53086, n53087, n53088,
         n53089, n53090, n53091, n53092, n53093, n53094, n53095, n53096,
         n53097, n53098, n53099, n53100, n53101, n53102, n53103, n53104,
         n53105, n53106, n53107, n53108, n53109, n53110, n53111, n53112,
         n53113, n53114, n53115, n53116, n53117, n53118, n53119, n53120,
         n53121, n53122, n53123, n53124, n53125, n53126, n53127, n53128,
         n53129, n53130, n53131, n53132, n53133, n53134, n53135, n53136,
         n53137, n53138, n53139, n53140, n53141, n53142, n53143, n53144,
         n53145, n53146, n53147, n53148, n53149, n53150, n53151, n53152,
         n53153, n53154, n53155, n53156, n53157, n53158, n53159, n53160,
         n53161, n53162, n53163, n53164, n53165, n53166, n53167, n53168,
         n53169, n53170, n53171, n53172, n53173, n53174, n53175, n53176,
         n53177, n53178, n53179, n53180, n53181, n53182, n53183, n53184,
         n53185, n53186, n53187, n53188, n53189, n53190, n53191, n53192,
         n53193, n53194, n53195, n53196, n53197, n53198, n53199, n53200,
         n53201, n53202, n53203, n53204, n53205, n53206, n53207, n53208,
         n53209, n53210, n53211, n53212, n53213, n53214, n53215, n53216,
         n53217, n53218, n53219, n53220, n53221, n53222, n53223, n53224,
         n53225, n53226, n53227, n53228, n53229, n53230, n53231, n53232,
         n53233, n53234, n53235, n53236, n53237, n53238, n53239, n53240,
         n53241, n53242, n53243, n53244, n53245, n53246, n53247, n53248,
         n53249, n53250, n53251, n53252, n53253, n53254, n53255, n53256,
         n53257, n53258, n53259, n53260, n53261, n53262, n53263, n53264,
         n53265, n53266, n53267, n53268, n53269, n53270, n53271, n53272,
         n53273, n53274, n53275, n53276, n53277, n53278, n53279, n53280,
         n53281, n53282, n53283, n53284, n53285, n53286, n53287, n53288,
         n53289, n53290, n53291, n53292, n53293, n53294, n53295, n53296,
         n53297, n53298, n53299, n53300, n53301, n53302, n53303, n53304,
         n53305, n53306, n53307, n53308, n53309, n53310, n53311, n53312,
         n53313, n53314, n53315, n53316, n53317, n53318, n53319, n53320,
         n53321, n53322, n53323, n53324, n53325, n53326, n53327, n53328,
         n53329, n53330, n53331, n53332, n53333, n53334, n53335, n53336,
         n53337, n53338, n53339, n53340, n53341, n53342, n53343, n53344,
         n53345, n53346, n53347, n53348, n53349, n53350, n53351, n53352,
         n53353, n53354, n53355, n53356, n53357, n53358, n53359, n53360,
         n53361, n53362, n53363, n53364, n53365, n53366, n53367, n53368,
         n53369, n53370, n53371, n53372, n53373, n53374, n53375, n53376,
         n53377, n53378, n53379, n53380, n53381, n53382, n53383, n53384,
         n53385, n53386, n53387, n53388, n53389, n53390, n53391, n53392,
         n53393, n53394, n53395, n53396, n53397, n53398, n53399, n53400,
         n53401, n53402, n53403, n53404, n53405, n53406, n53407, n53408,
         n53409, n53410, n53411, n53412, n53413, n53414, n53415, n53416,
         n53417, n53418, n53419, n53420, n53421, n53422, n53423, n53424,
         n53425, n53426, n53427, n53428, n53429, n53430, n53431, n53432,
         n53433, n53434, n53435, n53436, n53437, n53438, n53439, n53440,
         n53441, n53442, n53443, n53444, n53445, n53446, n53447, n53448,
         n53449, n53450, n53451, n53452, n53453, n53454, n53455, n53456,
         n53457, n53458, n53459, n53460, n53461, n53462, n53463, n53464,
         n53465, n53466, n53467, n53468, n53469, n53470, n53471, n53472,
         n53473, n53474, n53475, n53476, n53477, n53478, n53479, n53480,
         n53481, n53482, n53483, n53484, n53485, n53486, n53487, n53488,
         n53489, n53490, n53491, n53492, n53493, n53494, n53495, n53496,
         n53497, n53498, n53499, n53500, n53501, n53502, n53503, n53504,
         n53505, n53506, n53507, n53508, n53509, n53510, n53511, n53512,
         n53513, n53514, n53515, n53516, n53517, n53518, n53519, n53520,
         n53521, n53522, n53523, n53524, n53525, n53526, n53527, n53528,
         n53529, n53530, n53531, n53532, n53533, n53534, n53535, n53536,
         n53537, n53538, n53539, n53540, n53541, n53542, n53543, n53544,
         n53545, n53546, n53547, n53548, n53549, n53550, n53551, n53552,
         n53553, n53554, n53555, n53556, n53557, n53558, n53559, n53560,
         n53561, n53562, n53563, n53564, n53565, n53566, n53567, n53568,
         n53569, n53570, n53571, n53572, n53573, n53574, n53575, n53576,
         n53577, n53578, n53579, n53580, n53581, n53582, n53583, n53584,
         n53585, n53586, n53587, n53588, n53589, n53590, n53591, n53592,
         n53593, n53594, n53595, n53596, n53597, n53598, n53599, n53600,
         n53601, n53602, n53603, n53604, n53605, n53606, n53607, n53608,
         n53609, n53610, n53611, n53612, n53613, n53614, n53615, n53616,
         n53617, n53618, n53619, n53620, n53621, n53622, n53623, n53624,
         n53625, n53626, n53627, n53628, n53629, n53630, n53631, n53632,
         n53633, n53634, n53635, n53636, n53637, n53638, n53639, n53640,
         n53641, n53642, n53643, n53644, n53645, n53646, n53647, n53648,
         n53649, n53650, n53651, n53652, n53653, n53654, n53655, n53656,
         n53657, n53658, n53659, n53660, n53661, n53662, n53663, n53664,
         n53665, n53666, n53667, n53668, n53669, n53670, n53671, n53672,
         n53673, n53674, n53675, n53676, n53677, n53678, n53679, n53680,
         n53681, n53682, n53683, n53684, n53685, n53686, n53687, n53688,
         n53689, n53690, n53691, n53692, n53693, n53694, n53695, n53696,
         n53697, n53698, n53699, n53700, n53701, n53702, n53703, n53704,
         n53705, n53706, n53707, n53708, n53709, n53710, n53711, n53712,
         n53713, n53714, n53715, n53716, n53717, n53718, n53719, n53720,
         n53721, n53722, n53723, n53724, n53725, n53726, n53727, n53728,
         n53729, n53730, n53731, n53732, n53733, n53734, n53735, n53736,
         n53737, n53738, n53739, n53740, n53741, n53742, n53743, n53744,
         n53745, n53746, n53747, n53748, n53749, n53750, n53751, n53752,
         n53753, n53754, n53755, n53756, n53757, n53758, n53759, n53760,
         n53761, n53762, n53763, n53764, n53765, n53766, n53767, n53768,
         n53769, n53770, n53771, n53772, n53773, n53774, n53775, n53776,
         n53777, n53778, n53779, n53780, n53781, n53782, n53783, n53784,
         n53785, n53786, n53787, n53788, n53789, n53790, n53791, n53792,
         n53793, n53794, n53795, n53796, n53797, n53798, n53799, n53800,
         n53801, n53802, n53803, n53804, n53805, n53806, n53807, n53808,
         n53809, n53810, n53811, n53812, n53813, n53814, n53815, n53816,
         n53817, n53818, n53819, n53820, n53821, n53822, n53823, n53824,
         n53825, n53826, n53827, n53828, n53829, n53830, n53831, n53832,
         n53833, n53834, n53835, n53836, n53837, n53838, n53839, n53840,
         n53841, n53842, n53843, n53844, n53845, n53846, n53847, n53848,
         n53849, n53850, n53851, n53852, n53853, n53854, n53855, n53856,
         n53857, n53858, n53859, n53860, n53861, n53862, n53863, n53864,
         n53865, n53866, n53867, n53868, n53869, n53870, n53871, n53872,
         n53873, n53874, n53875, n53876, n53877, n53878, n53879, n53880,
         n53881, n53882, n53883, n53884, n53885, n53886, n53887, n53888,
         n53889, n53890, n53891, n53892, n53893, n53894, n53895, n53896,
         n53897, n53898, n53899, n53900, n53901, n53902, n53903, n53904,
         n53905, n53906, n53907, n53908, n53909, n53910, n53911, n53912,
         n53913, n53914, n53915, n53916, n53917, n53918, n53919, n53920,
         n53921, n53922, n53923, n53924, n53925, n53926, n53927, n53928,
         n53929, n53930, n53931, n53932, n53933, n53934, n53935, n53936,
         n53937, n53938, n53939, n53940, n53941, n53942, n53943, n53944,
         n53945, n53946, n53947, n53948, n53949, n53950, n53951, n53952,
         n53953, n53954, n53955, n53956, n53957, n53958, n53959, n53960,
         n53961, n53962, n53963, n53964, n53965, n53966, n53967, n53968,
         n53969, n53970, n53971, n53972, n53973, n53974, n53975, n53976,
         n53977, n53978, n53979, n53980, n53981, n53982, n53983, n53984,
         n53985, n53986, n53987, n53988, n53989, n53990, n53991, n53992,
         n53993, n53994, n53995, n53996, n53997, n53998, n53999, n54000,
         n54001, n54002, n54003, n54004, n54005, n54006, n54007, n54008,
         n54009, n54010, n54011, n54012, n54013, n54014, n54015, n54016,
         n54017, n54018, n54019, n54020, n54021, n54022, n54023, n54024,
         n54025, n54026, n54027, n54028, n54029, n54030, n54031, n54032,
         n54033, n54034, n54035, n54036, n54037, n54038, n54039, n54040,
         n54041, n54042, n54043, n54044, n54045, n54046, n54047, n54048,
         n54049, n54050, n54051, n54052, n54053, n54054, n54055, n54056,
         n54057, n54058, n54059, n54060, n54061, n54062, n54063, n54064,
         n54065, n54066, n54067, n54068, n54069, n54070, n54071, n54072,
         n54073, n54074, n54075, n54076, n54077, n54078, n54079, n54080,
         n54081, n54082, n54083, n54084, n54085, n54086, n54087, n54088,
         n54089, n54090, n54091, n54092, n54093, n54094, n54095, n54096,
         n54097, n54098, n54099, n54100, n54101, n54102, n54103, n54104,
         n54105, n54106, n54107, n54108, n54109, n54110, n54111, n54112,
         n54113, n54114, n54115, n54116, n54117, n54118, n54119, n54120,
         n54121, n54122, n54123, n54124, n54125, n54126, n54127, n54128,
         n54129, n54130, n54131, n54132, n54133, n54134, n54135, n54136,
         n54137, n54138, n54139, n54140, n54141, n54142, n54143, n54144,
         n54145, n54146, n54147, n54148, n54149, n54150, n54151, n54152,
         n54153, n54154, n54155, n54156, n54157, n54158, n54159, n54160,
         n54161, n54162, n54163, n54164, n54165, n54166, n54167, n54168,
         n54169, n54170, n54171, n54172, n54173, n54174, n54175, n54176,
         n54177, n54178, n54179, n54180, n54181, n54182, n54183, n54184,
         n54185, n54186, n54187, n54188, n54189, n54190, n54191, n54192,
         n54193, n54194, n54195, n54196, n54197, n54198, n54199, n54200,
         n54201, n54202, n54203, n54204, n54205, n54206, n54207, n54208,
         n54209, n54210, n54211, n54212, n54213, n54214, n54215, n54216,
         n54217, n54218, n54219, n54220, n54221, n54222, n54223, n54224,
         n54225, n54226, n54227, n54228, n54229, n54230, n54231, n54232,
         n54233, n54234, n54235, n54236, n54237, n54238, n54239, n54240,
         n54241, n54242, n54243, n54244, n54245, n54246, n54247, n54248,
         n54249, n54250, n54251, n54252, n54253, n54254, n54255, n54256,
         n54257, n54258, n54259, n54260, n54261, n54262, n54263, n54264,
         n54265, n54266, n54267, n54268, n54269, n54270, n54271, n54272,
         n54273, n54274, n54275, n54276, n54277, n54278, n54279, n54280,
         n54281, n54282, n54283, n54284, n54285, n54286, n54287, n54288,
         n54289, n54290, n54291, n54292, n54293, n54294, n54295, n54296,
         n54297, n54298, n54299, n54300, n54301, n54302, n54303, n54304,
         n54305, n54306, n54307, n54308, n54309, n54310, n54311, n54312,
         n54313, n54314, n54315, n54316, n54317, n54318, n54319, n54320,
         n54321, n54322, n54323, n54324, n54325, n54326, n54327, n54328,
         n54329, n54330, n54331, n54332, n54333, n54334, n54335, n54336,
         n54337, n54338, n54339, n54340, n54341, n54342, n54343, n54344,
         n54345, n54346, n54347, n54348, n54349, n54350, n54351, n54352,
         n54353, n54354, n54355, n54356, n54357, n54358, n54359, n54360,
         n54361, n54362, n54363, n54364, n54365, n54366, n54367, n54368,
         n54369, n54370, n54371, n54372, n54373, n54374, n54375, n54376,
         n54377, n54378, n54379, n54380, n54381, n54382, n54383, n54384,
         n54385, n54386, n54387, n54388, n54389, n54390, n54391, n54392,
         n54393, n54394, n54395, n54396, n54397, n54398, n54399, n54400,
         n54401, n54402, n54403, n54404, n54405, n54406, n54407, n54408,
         n54409, n54410, n54411, n54412, n54413, n54414, n54415, n54416,
         n54417, n54418, n54419, n54420, n54421, n54422, n54423, n54424,
         n54425, n54426, n54427, n54428, n54429, n54430, n54431, n54432,
         n54433, n54434, n54435, n54436, n54437, n54438, n54439, n54440,
         n54441, n54442, n54443, n54444, n54445, n54446, n54447, n54448,
         n54449, n54450, n54451, n54452, n54453, n54454, n54455, n54456,
         n54457, n54458, n54459, n54460, n54461, n54462, n54463, n54464,
         n54465, n54466, n54467, n54468, n54469, n54470, n54471, n54472,
         n54473, n54474, n54475, n54476, n54477, n54478, n54479, n54480,
         n54481, n54482, n54483, n54484, n54485, n54486, n54487, n54488,
         n54489, n54490, n54491, n54492, n54493, n54494, n54495, n54496,
         n54497, n54498, n54499, n54500, n54501, n54502, n54503, n54504,
         n54505, n54506, n54507, n54508, n54509, n54510, n54511, n54512,
         n54513, n54514, n54515, n54516, n54517, n54518, n54519, n54520,
         n54521, n54522, n54523, n54524, n54525, n54526, n54527, n54528,
         n54529, n54530, n54531, n54532, n54533, n54534, n54535, n54536,
         n54537, n54538, n54539, n54540, n54541, n54542, n54543, n54544,
         n54545, n54546, n54547, n54548, n54549, n54550, n54551, n54552,
         n54553, n54554, n54555, n54556, n54557, n54558, n54559, n54560,
         n54561, n54562, n54563, n54564, n54565, n54566, n54567, n54568,
         n54569, n54570, n54571, n54572, n54573, n54574, n54575, n54576,
         n54577, n54578, n54579, n54580, n54581, n54582, n54583, n54584,
         n54585, n54586, n54587, n54588, n54589, n54590, n54591, n54592,
         n54593, n54594, n54595, n54596, n54597, n54598, n54599, n54600,
         n54601, n54602, n54603, n54604, n54605, n54606, n54607, n54608,
         n54609, n54610, n54611, n54612, n54613, n54614, n54615, n54616,
         n54617, n54618, n54619, n54620, n54621, n54622, n54623, n54624,
         n54625, n54626, n54627, n54628, n54629, n54630, n54631, n54632,
         n54633, n54634, n54635, n54636, n54637, n54638, n54639, n54640,
         n54641, n54642, n54643, n54644, n54645, n54646, n54647, n54648,
         n54649, n54650, n54651, n54652, n54653, n54654, n54655, n54656,
         n54657, n54658, n54659, n54660, n54661, n54662, n54663, n54664,
         n54665, n54666, n54667, n54668, n54669, n54670, n54671, n54672,
         n54673, n54674, n54675, n54676, n54677, n54678, n54679, n54680,
         n54681, n54682, n54683, n54684, n54685, n54686, n54687, n54688,
         n54689, n54690, n54691, n54692, n54693, n54694, n54695, n54696,
         n54697, n54698, n54699, n54700, n54701, n54702, n54703, n54704,
         n54705, n54706, n54707, n54708, n54709, n54710, n54711, n54712,
         n54713, n54714, n54715, n54716, n54717, n54718, n54719, n54720,
         n54721, n54722, n54723, n54724, n54725, n54726, n54727, n54728,
         n54729, n54730, n54731, n54732, n54733, n54734, n54735, n54736,
         n54737, n54738, n54739, n54740, n54741, n54742, n54743, n54744,
         n54745, n54746, n54747, n54748, n54749, n54750, n54751, n54752,
         n54753, n54754, n54755, n54756, n54757, n54758, n54759, n54760,
         n54761, n54762, n54763, n54764, n54765, n54766, n54767, n54768,
         n54769, n54770, n54771, n54772, n54773, n54774, n54775, n54776,
         n54777, n54778, n54779, n54780, n54781, n54782, n54783, n54784,
         n54785, n54786, n54787, n54788, n54789, n54790, n54791, n54792,
         n54793, n54794, n54795, n54796, n54797, n54798, n54799, n54800,
         n54801, n54802, n54803, n54804, n54805, n54806, n54807, n54808,
         n54809, n54810, n54811, n54812, n54813, n54814, n54815, n54816,
         n54817, n54818, n54819, n54820, n54821, n54822, n54823, n54824,
         n54825, n54826, n54827, n54828, n54829, n54830, n54831, n54832,
         n54833, n54834, n54835, n54836, n54837, n54838, n54839, n54840,
         n54841, n54842, n54843, n54844, n54845, n54846, n54847, n54848,
         n54849, n54850, n54851, n54852, n54853, n54854, n54855, n54856,
         n54857, n54858, n54859, n54860, n54861, n54862, n54863, n54864,
         n54865, n54866, n54867, n54868, n54869, n54870, n54871, n54872,
         n54873, n54874, n54875, n54876, n54877, n54878, n54879, n54880,
         n54881, n54882, n54883, n54884, n54885, n54886, n54887, n54888,
         n54889, n54890, n54891, n54892, n54893, n54894, n54895, n54896,
         n54897, n54898, n54899, n54900, n54901, n54902, n54903, n54904,
         n54905, n54906, n54907, n54908, n54909, n54910, n54911, n54912,
         n54913, n54914, n54915, n54916, n54917, n54918, n54919, n54920,
         n54921, n54922, n54923, n54924, n54925, n54926, n54927, n54928,
         n54929, n54930, n54931, n54932, n54933, n54934, n54935, n54936,
         n54937, n54938, n54939, n54940, n54941, n54942, n54943, n54944,
         n54945, n54946, n54947, n54948, n54949, n54950, n54951, n54952,
         n54953, n54954, n54955, n54956, n54957, n54958, n54959, n54960,
         n54961, n54962, n54963, n54964, n54965, n54966, n54967, n54968,
         n54969, n54970, n54971, n54972, n54973, n54974, n54975, n54976,
         n54977, n54978, n54979, n54980, n54981, n54982, n54983, n54984,
         n54985, n54986, n54987, n54988, n54989, n54990, n54991, n54992,
         n54993, n54994, n54995, n54996, n54997, n54998, n54999, n55000,
         n55001, n55002, n55003, n55004, n55005, n55006, n55007, n55008,
         n55009, n55010, n55011, n55012, n55013, n55014, n55015, n55016,
         n55017, n55018, n55019, n55020, n55021, n55022, n55023, n55024,
         n55025, n55026, n55027, n55028, n55029, n55030, n55031, n55032,
         n55033, n55034, n55035, n55036, n55037, n55038, n55039, n55040,
         n55041, n55042, n55043, n55044, n55045, n55046, n55047, n55048,
         n55049, n55050, n55051, n55052, n55053, n55054, n55055, n55056,
         n55057, n55058, n55059, n55060, n55061, n55062, n55063, n55064,
         n55065, n55066, n55067, n55068, n55069, n55070, n55071, n55072,
         n55073, n55074, n55075, n55076, n55077, n55078, n55079, n55080,
         n55081, n55082, n55083, n55084, n55085, n55086, n55087, n55088,
         n55089, n55090, n55091, n55092, n55093, n55094, n55095, n55096,
         n55097, n55098, n55099, n55100, n55101, n55102, n55103, n55104,
         n55105, n55106, n55107, n55108, n55109, n55110, n55111, n55112,
         n55113, n55114, n55115, n55116, n55117, n55118, n55119, n55120,
         n55121, n55122, n55123, n55124, n55125, n55126, n55127, n55128,
         n55129, n55130, n55131, n55132, n55133, n55134, n55135, n55136,
         n55137, n55138, n55139, n55140, n55141, n55142, n55143, n55144,
         n55145, n55146, n55147, n55148, n55149, n55150, n55151, n55152,
         n55153, n55154, n55155, n55156, n55157, n55158, n55159, n55160,
         n55161, n55162, n55163, n55164, n55165, n55166, n55167, n55168,
         n55169, n55170, n55171, n55172, n55173, n55174, n55175, n55176,
         n55177, n55178, n55179, n55180, n55181, n55182, n55183, n55184,
         n55185, n55186, n55187, n55188, n55189, n55190, n55191, n55192,
         n55193, n55194, n55195, n55196, n55197, n55198, n55199, n55200,
         n55201, n55202, n55203, n55204, n55205, n55206, n55207, n55208,
         n55209, n55210, n55211, n55212, n55213, n55214, n55215, n55216,
         n55217, n55218, n55219, n55220, n55221, n55222, n55223, n55224,
         n55225, n55226, n55227, n55228, n55229, n55230, n55231, n55232,
         n55233, n55234, n55235, n55236, n55237, n55238, n55239, n55240,
         n55241, n55242, n55243, n55244, n55245, n55246, n55247, n55248,
         n55249, n55250, n55251, n55252, n55253, n55254, n55255, n55256,
         n55257, n55258, n55259, n55260, n55261, n55262, n55263, n55264,
         n55265, n55266, n55267, n55268, n55269, n55270, n55271, n55272,
         n55273, n55274, n55275, n55276, n55277, n55278, n55279, n55280,
         n55281, n55282, n55283, n55284, n55285, n55286, n55287, n55288,
         n55289, n55290, n55291, n55292, n55293, n55294, n55295, n55296,
         n55297, n55298, n55299, n55300, n55301, n55302, n55303, n55304,
         n55305, n55306, n55307, n55308, n55309, n55310, n55311, n55312,
         n55313, n55314, n55315, n55316, n55317, n55318, n55319, n55320,
         n55321, n55322, n55323, n55324, n55325, n55326, n55327, n55328,
         n55329, n55330, n55331, n55332, n55333, n55334, n55335, n55336,
         n55337, n55338, n55339, n55340, n55341, n55342, n55343, n55344,
         n55345, n55346, n55347, n55348, n55349, n55350, n55351, n55352,
         n55353, n55354, n55355, n55356, n55357, n55358, n55359, n55360,
         n55361, n55362, n55363, n55364, n55365, n55366, n55367, n55368,
         n55369, n55370, n55371, n55372, n55373, n55374, n55375, n55376,
         n55377, n55378, n55379, n55380, n55381, n55382, n55383, n55384,
         n55385, n55386, n55387, n55388, n55389, n55390, n55391, n55392,
         n55393, n55394, n55395, n55396, n55397, n55398, n55399, n55400,
         n55401, n55402, n55403, n55404, n55405, n55406, n55407, n55408,
         n55409, n55410, n55411, n55412, n55413, n55414, n55415, n55416,
         n55417, n55418, n55419, n55420, n55421, n55422, n55423, n55424,
         n55425, n55426, n55427, n55428, n55429, n55430, n55431, n55432,
         n55433, n55434, n55435, n55436, n55437, n55438, n55439, n55440,
         n55441, n55442, n55443, n55444, n55445, n55446, n55447, n55448,
         n55449, n55450, n55451, n55452, n55453, n55454, n55455, n55456,
         n55457, n55458, n55459, n55460, n55461, n55462, n55463, n55464,
         n55465, n55466, n55467, n55468, n55469, n55470, n55471, n55472,
         n55473, n55474, n55475, n55476, n55477, n55478, n55479, n55480,
         n55481, n55482, n55483, n55484, n55485, n55486, n55487, n55488,
         n55489, n55490, n55491, n55492, n55493, n55494, n55495, n55496,
         n55497, n55498, n55499, n55500, n55501, n55502, n55503, n55504,
         n55505, n55506, n55507, n55508, n55509, n55510, n55511, n55512,
         n55513, n55514, n55515, n55516, n55517, n55518, n55519, n55520,
         n55521, n55522, n55523, n55524, n55525, n55526, n55527, n55528,
         n55529, n55530, n55531, n55532, n55533, n55534, n55535, n55536,
         n55537, n55538, n55539, n55540, n55541, n55542, n55543, n55544,
         n55545, n55546, n55547, n55548, n55549, n55550, n55551, n55552,
         n55553, n55554, n55555, n55556, n55557, n55558, n55559, n55560,
         n55561, n55562, n55563, n55564, n55565, n55566, n55567, n55568,
         n55569, n55570, n55571, n55572, n55573, n55574, n55575, n55576,
         n55577, n55578, n55579, n55580, n55581, n55582, n55583, n55584,
         n55585, n55586, n55587, n55588, n55589, n55590, n55591, n55592,
         n55593, n55594, n55595, n55596, n55597, n55598, n55599, n55600,
         n55601, n55602, n55603, n55604, n55605, n55606, n55607, n55608,
         n55609, n55610, n55611, n55612, n55613, n55614, n55615, n55616,
         n55617, n55618, n55619, n55620, n55621, n55622, n55623, n55624,
         n55625, n55626, n55627, n55628, n55629, n55630, n55631, n55632,
         n55633, n55634, n55635, n55636, n55637, n55638, n55639, n55640,
         n55641, n55642, n55643, n55644, n55645, n55646, n55647, n55648,
         n55649, n55650, n55651, n55652, n55653, n55654, n55655, n55656,
         n55657, n55658, n55659, n55660, n55661, n55662, n55663, n55664,
         n55665, n55666, n55667, n55668, n55669, n55670, n55671, n55672,
         n55673, n55674, n55675, n55676, n55677, n55678, n55679, n55680,
         n55681, n55682, n55683, n55684, n55685, n55686, n55687, n55688,
         n55689, n55690, n55691, n55692, n55693, n55694, n55695, n55696,
         n55697, n55698, n55699, n55700, n55701, n55702, n55703, n55704,
         n55705, n55706, n55707, n55708, n55709, n55710, n55711, n55712,
         n55713, n55714, n55715, n55716, n55717, n55718, n55719, n55720,
         n55721, n55722, n55723, n55724, n55725, n55726, n55727, n55728,
         n55729, n55730, n55731, n55732, n55733, n55734, n55735, n55736,
         n55737, n55738, n55739, n55740, n55741, n55742, n55743, n55744,
         n55745, n55746, n55747, n55748, n55749, n55750, n55751, n55752,
         n55753, n55754, n55755, n55756, n55757, n55758, n55759, n55760,
         n55761, n55762, n55763, n55764, n55765, n55766, n55767, n55768,
         n55769, n55770, n55771, n55772, n55773, n55774, n55775, n55776,
         n55777, n55778, n55779, n55780, n55781, n55782, n55783, n55784,
         n55785, n55786, n55787, n55788, n55789, n55790, n55791, n55792,
         n55793, n55794, n55795, n55796, n55797, n55798, n55799, n55800,
         n55801, n55802, n55803, n55804, n55805, n55806, n55807, n55808,
         n55809, n55810, n55811, n55812, n55813, n55814, n55815, n55816,
         n55817, n55818, n55819, n55820, n55821, n55822, n55823, n55824,
         n55825, n55826, n55827, n55828, n55829, n55830, n55831, n55832,
         n55833, n55834, n55835, n55836, n55837, n55838, n55839, n55840,
         n55841, n55842, n55843, n55844, n55845, n55846, n55847, n55848,
         n55849, n55850, n55851, n55852, n55853, n55854, n55855, n55856,
         n55857, n55858, n55859, n55860, n55861, n55862, n55863, n55864,
         n55865, n55866, n55867, n55868, n55869, n55870, n55871, n55872,
         n55873, n55874, n55875, n55876, n55877, n55878, n55879, n55880,
         n55881, n55882, n55883, n55884, n55885, n55886, n55887, n55888,
         n55889, n55890, n55891, n55892, n55893, n55894, n55895, n55896,
         n55897, n55898, n55899, n55900, n55901, n55902, n55903, n55904,
         n55905, n55906, n55907, n55908, n55909, n55910, n55911, n55912,
         n55913, n55914, n55915, n55916, n55917, n55918, n55919, n55920,
         n55921, n55922, n55923, n55924, n55925, n55926, n55927, n55928,
         n55929, n55930, n55931, n55932, n55933, n55934, n55935, n55936,
         n55937, n55938, n55939, n55940, n55941, n55942, n55943, n55944,
         n55945, n55946, n55947, n55948, n55949, n55950, n55951, n55952,
         n55953, n55954, n55955, n55956, n55957, n55958, n55959, n55960,
         n55961, n55962, n55963, n55964, n55965, n55966, n55967, n55968,
         n55969, n55970, n55971, n55972, n55973, n55974, n55975, n55976,
         n55977, n55978, n55979, n55980, n55981, n55982, n55983, n55984,
         n55985, n55986, n55987, n55988, n55989, n55990, n55991, n55992,
         n55993, n55994, n55995, n55996, n55997, n55998, n55999, n56000,
         n56001, n56002, n56003, n56004, n56005, n56006, n56007, n56008,
         n56009, n56010, n56011, n56012, n56013, n56014, n56015, n56016,
         n56017, n56018, n56019, n56020, n56021, n56022, n56023, n56024,
         n56025, n56026, n56027, n56028, n56029, n56030, n56031, n56032,
         n56033, n56034, n56035, n56036, n56037, n56038, n56039, n56040,
         n56041, n56042, n56043, n56044, n56045, n56046, n56047, n56048,
         n56049, n56050, n56051, n56052, n56053, n56054, n56055, n56056,
         n56057, n56058, n56059, n56060, n56061, n56062, n56063, n56064,
         n56065, n56066, n56067, n56068, n56069, n56070, n56071, n56072,
         n56073, n56074, n56075, n56076, n56077, n56078, n56079, n56080,
         n56081, n56082, n56083, n56084, n56085, n56086, n56087, n56088,
         n56089, n56090, n56091, n56092, n56093, n56094, n56095, n56096,
         n56097, n56098, n56099, n56100, n56101, n56102, n56103, n56104,
         n56105, n56106, n56107, n56108, n56109, n56110, n56111, n56112,
         n56113, n56114, n56115, n56116, n56117, n56118, n56119, n56120,
         n56121, n56122, n56123, n56124, n56125, n56126, n56127, n56128,
         n56129, n56130, n56131, n56132, n56133, n56134, n56135, n56136,
         n56137, n56138, n56139, n56140, n56141, n56142, n56143, n56144,
         n56145, n56146, n56147, n56148, n56149, n56150, n56151, n56152,
         n56153, n56154, n56155, n56156, n56157, n56158, n56159, n56160,
         n56161, n56162, n56163, n56164, n56165, n56166, n56167, n56168,
         n56169, n56170, n56171, n56172, n56173, n56174, n56175, n56176,
         n56177, n56178, n56179, n56180, n56181, n56182, n56183, n56184,
         n56185, n56186, n56187, n56188, n56189, n56190, n56191, n56192,
         n56193, n56194, n56195, n56196, n56197, n56198, n56199, n56200,
         n56201, n56202, n56203, n56204, n56205, n56206, n56207, n56208,
         n56209, n56210, n56211, n56212, n56213, n56214, n56215, n56216,
         n56217, n56218, n56219, n56220, n56221, n56222, n56223, n56224,
         n56225, n56226, n56227, n56228, n56229, n56230, n56231, n56232,
         n56233, n56234, n56235, n56236, n56237, n56238, n56239, n56240,
         n56241, n56242, n56243, n56244, n56245, n56246, n56247, n56248,
         n56249, n56250, n56251, n56252, n56253, n56254, n56255, n56256,
         n56257, n56258, n56259, n56260, n56261, n56262, n56263, n56264,
         n56265, n56266, n56267, n56268, n56269, n56270, n56271, n56272,
         n56273, n56274, n56275, n56276, n56277, n56278, n56279, n56280,
         n56281, n56282, n56283, n56284, n56285, n56286, n56287, n56288,
         n56289, n56290, n56291, n56292, n56293, n56294, n56295, n56296,
         n56297, n56298, n56299, n56300, n56301, n56302, n56303, n56304,
         n56305, n56306, n56307, n56308, n56309, n56310, n56311, n56312,
         n56313, n56314, n56315, n56316, n56317, n56318, n56319, n56320,
         n56321, n56322, n56323, n56324, n56325, n56326, n56327, n56328,
         n56329, n56330, n56331, n56332, n56333, n56334, n56335, n56336,
         n56337, n56338, n56339, n56340, n56341, n56342, n56343, n56344,
         n56345, n56346, n56347, n56348, n56349, n56350, n56351, n56352,
         n56353, n56354, n56355, n56356, n56357, n56358, n56359, n56360,
         n56361, n56362, n56363, n56364, n56365, n56366, n56367, n56368,
         n56369, n56370, n56371, n56372, n56373, n56374, n56375, n56376,
         n56377, n56378, n56379, n56380, n56381, n56382, n56383, n56384,
         n56385, n56386, n56387, n56388, n56389, n56390, n56391, n56392,
         n56393, n56394, n56395, n56396, n56397, n56398, n56399, n56400,
         n56401, n56402, n56403, n56404, n56405, n56406, n56407, n56408,
         n56409, n56410, n56411, n56412, n56413, n56414, n56415, n56416,
         n56417, n56418, n56419, n56420, n56421, n56422, n56423, n56424,
         n56425, n56426, n56427, n56428, n56429, n56430, n56431, n56432,
         n56433, n56434, n56435, n56436, n56437, n56438, n56439, n56440,
         n56441, n56442, n56443, n56444, n56445, n56446, n56447, n56448,
         n56449, n56450, n56451, n56452, n56453, n56454, n56455, n56456,
         n56457, n56458, n56459, n56460, n56461, n56462, n56463, n56464,
         n56465, n56466, n56467, n56468, n56469, n56470, n56471, n56472,
         n56473, n56474, n56475, n56476, n56477, n56478, n56479, n56480,
         n56481, n56482, n56483, n56484, n56485, n56486, n56487, n56488,
         n56489, n56490, n56491, n56492, n56493, n56494, n56495, n56496,
         n56497, n56498, n56499, n56500, n56501, n56502, n56503, n56504,
         n56505, n56506, n56507, n56508, n56509, n56510, n56511, n56512,
         n56513, n56514, n56515, n56516, n56517, n56518, n56519, n56520,
         n56521, n56522, n56523, n56524, n56525, n56526, n56527, n56528,
         n56529, n56530, n56531, n56532, n56533, n56534, n56535, n56536,
         n56537, n56538, n56539, n56540, n56541, n56542, n56543, n56544,
         n56545, n56546, n56547, n56548, n56549, n56550, n56551, n56552,
         n56553, n56554, n56555, n56556, n56557, n56558, n56559, n56560,
         n56561, n56562, n56563, n56564, n56565, n56566, n56567, n56568,
         n56569, n56570, n56571, n56572, n56573, n56574, n56575, n56576,
         n56577, n56578, n56579, n56580, n56581, n56582, n56583, n56584,
         n56585, n56586, n56587, n56588, n56589, n56590, n56591, n56592,
         n56593, n56594, n56595, n56596, n56597, n56598, n56599, n56600,
         n56601, n56602, n56603, n56604, n56605, n56606, n56607, n56608,
         n56609, n56610, n56611, n56612, n56613, n56614, n56615, n56616,
         n56617, n56618, n56619, n56620, n56621, n56622, n56623, n56624,
         n56625, n56626, n56627, n56628, n56629, n56630, n56631, n56632,
         n56633, n56634, n56635, n56636, n56637, n56638, n56639, n56640,
         n56641, n56642, n56643, n56644, n56645, n56646, n56647, n56648,
         n56649, n56650, n56651, n56652, n56653, n56654, n56655, n56656,
         n56657, n56658, n56659, n56660, n56661, n56662, n56663, n56664,
         n56665, n56666, n56667, n56668, n56669, n56670, n56671, n56672,
         n56673, n56674, n56675, n56676, n56677, n56678, n56679, n56680,
         n56681, n56682, n56683, n56684, n56685, n56686, n56687, n56688,
         n56689, n56690, n56691, n56692, n56693, n56694, n56695, n56696,
         n56697, n56698, n56699, n56700, n56701, n56702, n56703, n56704,
         n56705, n56706, n56707, n56708, n56709, n56710, n56711, n56712,
         n56713, n56714, n56715, n56716, n56717, n56718, n56719, n56720,
         n56721, n56722, n56723, n56724, n56725, n56726, n56727, n56728,
         n56729, n56730, n56731, n56732, n56733, n56734, n56735, n56736,
         n56737, n56738, n56739, n56740, n56741, n56742, n56743, n56744,
         n56745, n56746, n56747, n56748, n56749, n56750, n56751, n56752,
         n56753, n56754, n56755, n56756, n56757, n56758, n56759, n56760,
         n56761, n56762, n56763, n56764, n56765, n56766, n56767, n56768,
         n56769, n56770, n56771, n56772, n56773, n56774, n56775, n56776,
         n56777, n56778, n56779, n56780, n56781, n56782, n56783, n56784,
         n56785, n56786, n56787, n56788, n56789, n56790, n56791, n56792,
         n56793, n56794, n56795, n56796, n56797, n56798, n56799, n56800,
         n56801, n56802, n56803, n56804, n56805, n56806, n56807, n56808,
         n56809, n56810, n56811, n56812, n56813, n56814, n56815, n56816,
         n56817, n56818, n56819, n56820, n56821, n56822, n56823, n56824,
         n56825, n56826, n56827, n56828, n56829, n56830, n56831, n56832,
         n56833, n56834, n56835, n56836, n56837, n56838, n56839, n56840,
         n56841, n56842, n56843, n56844, n56845, n56846, n56847, n56848,
         n56849, n56850, n56851, n56852, n56853, n56854, n56855, n56856,
         n56857, n56858, n56859, n56860, n56861, n56862, n56863, n56864,
         n56865, n56866, n56867, n56868, n56869, n56870, n56871, n56872,
         n56873, n56874, n56875, n56876, n56877, n56878, n56879, n56880,
         n56881, n56882, n56883, n56884, n56885, n56886, n56887, n56888,
         n56889, n56890, n56891, n56892, n56893, n56894, n56895, n56896,
         n56897, n56898, n56899, n56900, n56901, n56902, n56903, n56904,
         n56905, n56906, n56907, n56908, n56909, n56910, n56911, n56912,
         n56913, n56914, n56915, n56916, n56917, n56918, n56919, n56920,
         n56921, n56922, n56923, n56924, n56925, n56926, n56927, n56928,
         n56929, n56930, n56931, n56932, n56933, n56934, n56935, n56936,
         n56937, n56938, n56939, n56940, n56941, n56942, n56943, n56944,
         n56945, n56946, n56947, n56948, n56949, n56950, n56951, n56952,
         n56953, n56954, n56955, n56956, n56957, n56958, n56959, n56960,
         n56961, n56962, n56963, n56964, n56965, n56966, n56967, n56968,
         n56969, n56970, n56971, n56972, n56973, n56974, n56975, n56976,
         n56977, n56978, n56979, n56980, n56981, n56982, n56983, n56984,
         n56985, n56986, n56987, n56988, n56989, n56990, n56991, n56992,
         n56993, n56994, n56995, n56996, n56997, n56998, n56999, n57000,
         n57001, n57002, n57003, n57004, n57005, n57006, n57007, n57008,
         n57009, n57010, n57011, n57012, n57013, n57014, n57015, n57016,
         n57017, n57018, n57019, n57020, n57021, n57022, n57023, n57024,
         n57025, n57026, n57027, n57028, n57029, n57030, n57031, n57032,
         n57033, n57034, n57035, n57036, n57037, n57038, n57039, n57040,
         n57041, n57042, n57043, n57044, n57045, n57046, n57047, n57048,
         n57049, n57050, n57051, n57052, n57053, n57054, n57055, n57056,
         n57057, n57058, n57059, n57060, n57061, n57062, n57063, n57064,
         n57065, n57066, n57067, n57068, n57069, n57070, n57071, n57072,
         n57073, n57074, n57075, n57076, n57077, n57078, n57079, n57080,
         n57081, n57082, n57083, n57084, n57085, n57086, n57087, n57088,
         n57089, n57090, n57091, n57092, n57093, n57094, n57095, n57096,
         n57097, n57098, n57099, n57100, n57101, n57102, n57103, n57104,
         n57105, n57106, n57107, n57108, n57109, n57110, n57111, n57112,
         n57113, n57114, n57115, n57116, n57117, n57118, n57119, n57120,
         n57121, n57122, n57123, n57124, n57125, n57126, n57127, n57128,
         n57129, n57130, n57131, n57132, n57133, n57134, n57135, n57136,
         n57137, n57138, n57139, n57140, n57141, n57142, n57143, n57144,
         n57145, n57146, n57147, n57148, n57149, n57150, n57151, n57152,
         n57153, n57154, n57155, n57156, n57157, n57158, n57159, n57160,
         n57161, n57162, n57163, n57164, n57165, n57166, n57167, n57168,
         n57169, n57170, n57171, n57172, n57173, n57174, n57175, n57176,
         n57177, n57178, n57179, n57180, n57181, n57182, n57183, n57184,
         n57185, n57186, n57187, n57188, n57189, n57190, n57191, n57192,
         n57193, n57194, n57195, n57196, n57197, n57198, n57199, n57200,
         n57201, n57202, n57203, n57204, n57205, n57206, n57207, n57208,
         n57209, n57210, n57211, n57212, n57213, n57214, n57215, n57216,
         n57217, n57218, n57219, n57220, n57221, n57222, n57223, n57224,
         n57225, n57226, n57227, n57228, n57229, n57230, n57231, n57232,
         n57233, n57234, n57235, n57236, n57237, n57238, n57239, n57240,
         n57241, n57242, n57243, n57244, n57245, n57246, n57247, n57248,
         n57249, n57250, n57251, n57252, n57253, n57254, n57255, n57256,
         n57257, n57258, n57259, n57260, n57261, n57262, n57263, n57264,
         n57265, n57266, n57267, n57268, n57269, n57270, n57271, n57272,
         n57273, n57274, n57275, n57276, n57277, n57278, n57279, n57280,
         n57281, n57282, n57283, n57284, n57285, n57286, n57287, n57288,
         n57289, n57290, n57291, n57292, n57293, n57294, n57295, n57296,
         n57297, n57298, n57299, n57300, n57301, n57302, n57303, n57304,
         n57305, n57306, n57307, n57308, n57309, n57310, n57311, n57312,
         n57313, n57314, n57315, n57316, n57317, n57318, n57319, n57320,
         n57321, n57322, n57323, n57324, n57325, n57326, n57327, n57328,
         n57329, n57330, n57331, n57332, n57333, n57334, n57335, n57336,
         n57337, n57338, n57339, n57340, n57341, n57342, n57343, n57344,
         n57345, n57346, n57347, n57348, n57349, n57350, n57351, n57352,
         n57353, n57354, n57355, n57356, n57357, n57358, n57359, n57360,
         n57361, n57362, n57363, n57364, n57365, n57366, n57367, n57368,
         n57369, n57370, n57371, n57372, n57373, n57374, n57375, n57376,
         n57377, n57378, n57379, n57380, n57381, n57382, n57383, n57384,
         n57385, n57386, n57387, n57388, n57389, n57390, n57391, n57392,
         n57393, n57394, n57395, n57396, n57397, n57398, n57399, n57400,
         n57401, n57402, n57403, n57404, n57405, n57406, n57407, n57408,
         n57409, n57410, n57411, n57412, n57413, n57414, n57415, n57416,
         n57417, n57418, n57419, n57420, n57421, n57422, n57423, n57424,
         n57425, n57426, n57427, n57428, n57429, n57430, n57431, n57432,
         n57433, n57434, n57435, n57436, n57437, n57438, n57439, n57440,
         n57441, n57442, n57443, n57444, n57445, n57446, n57447, n57448,
         n57449, n57450, n57451, n57452, n57453, n57454, n57455, n57456,
         n57457, n57458, n57459, n57460, n57461, n57462, n57463, n57464,
         n57465, n57466, n57467, n57468, n57469, n57470, n57471, n57472,
         n57473, n57474, n57475, n57476, n57477, n57478, n57479, n57480,
         n57481, n57482, n57483, n57484, n57485, n57486, n57487, n57488,
         n57489, n57490, n57491, n57492, n57493, n57494, n57495, n57496,
         n57497, n57498, n57499, n57500, n57501, n57502, n57503, n57504,
         n57505, n57506, n57507, n57508, n57509, n57510, n57511, n57512,
         n57513, n57514, n57515, n57516, n57517, n57518, n57519, n57520,
         n57521, n57522, n57523, n57524, n57525, n57526, n57527, n57528,
         n57529, n57530, n57531, n57532, n57533, n57534, n57535, n57536,
         n57537, n57538, n57539, n57540, n57541, n57542, n57543, n57544,
         n57545, n57546, n57547, n57548, n57549, n57550, n57551, n57552,
         n57553, n57554, n57555, n57556, n57557, n57558, n57559, n57560,
         n57561, n57562, n57563, n57564, n57565, n57566, n57567, n57568,
         n57569, n57570, n57571, n57572, n57573, n57574, n57575, n57576,
         n57577, n57578, n57579, n57580, n57581, n57582, n57583, n57584,
         n57585, n57586, n57587, n57588, n57589, n57590, n57591, n57592,
         n57593, n57594, n57595, n57596, n57597, n57598, n57599, n57600,
         n57601, n57602, n57603, n57604, n57605, n57606, n57607, n57608,
         n57609, n57610, n57611, n57612, n57613, n57614, n57615, n57616,
         n57617, n57618, n57619, n57620, n57621, n57622, n57623, n57624,
         n57625, n57626, n57627, n57628, n57629, n57630, n57631, n57632,
         n57633, n57634, n57635, n57636, n57637, n57638, n57639, n57640,
         n57641, n57642, n57643, n57644, n57645, n57646, n57647, n57648,
         n57649, n57650, n57651, n57652, n57653, n57654, n57655, n57656,
         n57657, n57658, n57659, n57660, n57661, n57662, n57663, n57664,
         n57665, n57666, n57667, n57668, n57669, n57670, n57671, n57672,
         n57673, n57674, n57675, n57676, n57677, n57678, n57679, n57680,
         n57681, n57682, n57683, n57684, n57685, n57686, n57687, n57688,
         n57689, n57690, n57691, n57692, n57693, n57694, n57695, n57696,
         n57697, n57698, n57699, n57700, n57701, n57702, n57703, n57704,
         n57705, n57706, n57707, n57708, n57709, n57710, n57711, n57712,
         n57713, n57714, n57715, n57716, n57717, n57718, n57719, n57720,
         n57721, n57722, n57723, n57724, n57725, n57726, n57727, n57728,
         n57729, n57730, n57731, n57732, n57733, n57734, n57735, n57736,
         n57737, n57738, n57739, n57740, n57741, n57742, n57743, n57744,
         n57745, n57746, n57747, n57748, n57749, n57750, n57751, n57752,
         n57753, n57754, n57755, n57756, n57757, n57758, n57759, n57760,
         n57761, n57762, n57763, n57764, n57765, n57766, n57767, n57768,
         n57769, n57770, n57771, n57772, n57773, n57774, n57775, n57776,
         n57777, n57778, n57779, n57780, n57781, n57782, n57783, n57784,
         n57785, n57786, n57787, n57788, n57789, n57790, n57791, n57792,
         n57793, n57794, n57795, n57796, n57797, n57798, n57799, n57800,
         n57801, n57802, n57803, n57804, n57805, n57806, n57807, n57808,
         n57809, n57810, n57811, n57812, n57813, n57814, n57815, n57816,
         n57817, n57818, n57819, n57820, n57821, n57822, n57823, n57824,
         n57825, n57826, n57827, n57828, n57829, n57830, n57831, n57832,
         n57833, n57834, n57835, n57836, n57837, n57838, n57839, n57840,
         n57841, n57842, n57843, n57844, n57845, n57846, n57847, n57848,
         n57849, n57850, n57851, n57852, n57853, n57854, n57855, n57856,
         n57857, n57858, n57859, n57860, n57861, n57862, n57863, n57864,
         n57865, n57866, n57867, n57868, n57869, n57870, n57871, n57872,
         n57873, n57874, n57875, n57876, n57877, n57878, n57879, n57880,
         n57881, n57882, n57883, n57884, n57885, n57886, n57887, n57888,
         n57889, n57890, n57891, n57892, n57893, n57894, n57895, n57896,
         n57897, n57898, n57899, n57900, n57901, n57902, n57903, n57904,
         n57905, n57906, n57907, n57908, n57909, n57910, n57911, n57912,
         n57913, n57914, n57915, n57916, n57917, n57918, n57919, n57920,
         n57921, n57922, n57923, n57924, n57925, n57926, n57927, n57928,
         n57929, n57930, n57931, n57932, n57933, n57934, n57935, n57936,
         n57937, n57938, n57939, n57940, n57941, n57942, n57943, n57944,
         n57945, n57946, n57947, n57948, n57949, n57950, n57951, n57952,
         n57953, n57954, n57955, n57956, n57957, n57958, n57959, n57960,
         n57961, n57962, n57963, n57964, n57965, n57966, n57967, n57968,
         n57969, n57970, n57971, n57972, n57973, n57974, n57975, n57976,
         n57977, n57978, n57979, n57980, n57981, n57982, n57983, n57984,
         n57985, n57986, n57987, n57988, n57989, n57990, n57991, n57992,
         n57993, n57994, n57995, n57996, n57997, n57998, n57999, n58000,
         n58001, n58002, n58003, n58004, n58005, n58006, n58007, n58008,
         n58009, n58010, n58011, n58012, n58013, n58014, n58015, n58016,
         n58017, n58018, n58019, n58020, n58021, n58022, n58023, n58024,
         n58025, n58026, n58027, n58028, n58029, n58030, n58031, n58032,
         n58033, n58034, n58035, n58036, n58037, n58038, n58039, n58040,
         n58041, n58042, n58043, n58044, n58045, n58046, n58047, n58048,
         n58049, n58050, n58051, n58052, n58053, n58054, n58055, n58056,
         n58057, n58058, n58059, n58060, n58061, n58062, n58063, n58064,
         n58065, n58066, n58067, n58068, n58069, n58070, n58071, n58072,
         n58073, n58074, n58075, n58076, n58077, n58078, n58079, n58080,
         n58081, n58082, n58083, n58084, n58085, n58086, n58087, n58088,
         n58089, n58090, n58091, n58092, n58093, n58094, n58095, n58096,
         n58097, n58098, n58099, n58100, n58101, n58102, n58103, n58104,
         n58105, n58106, n58107, n58108, n58109, n58110, n58111, n58112,
         n58113, n58114, n58115, n58116, n58117, n58118, n58119, n58120,
         n58121, n58122, n58123, n58124, n58125, n58126, n58127, n58128,
         n58129, n58130, n58131, n58132, n58133, n58134, n58135, n58136,
         n58137, n58138, n58139, n58140, n58141, n58142, n58143, n58144,
         n58145, n58146, n58147, n58148, n58149, n58150, n58151, n58152,
         n58153, n58154, n58155, n58156, n58157, n58158, n58159, n58160,
         n58161, n58162, n58163, n58164, n58165, n58166, n58167, n58168,
         n58169, n58170, n58171, n58172, n58173, n58174, n58175, n58176,
         n58177, n58178, n58179, n58180, n58181, n58182, n58183, n58184,
         n58185, n58186, n58187, n58188, n58189, n58190, n58191, n58192,
         n58193, n58194, n58195, n58196, n58197, n58198, n58199, n58200,
         n58201, n58202, n58203, n58204, n58205, n58206, n58207, n58208,
         n58209, n58210, n58211, n58212, n58213, n58214, n58215, n58216,
         n58217, n58218, n58219, n58220, n58221, n58222, n58223, n58224,
         n58225, n58226, n58227, n58228, n58229, n58230, n58231, n58232,
         n58233, n58234, n58235, n58236, n58237, n58238, n58239, n58240,
         n58241, n58242, n58243, n58244, n58245, n58246, n58247, n58248,
         n58249, n58250, n58251, n58252, n58253, n58254, n58255, n58256,
         n58257, n58258, n58259, n58260, n58261, n58262, n58263, n58264,
         n58265, n58266, n58267, n58268, n58269, n58270, n58271, n58272,
         n58273, n58274, n58275, n58276, n58277, n58278, n58279, n58280,
         n58281, n58282, n58283, n58284, n58285, n58286, n58287, n58288,
         n58289, n58290, n58291, n58292, n58293, n58294, n58295, n58296,
         n58297, n58298, n58299, n58300, n58301, n58302, n58303, n58304,
         n58305, n58306, n58307, n58308, n58309, n58310, n58311, n58312,
         n58313, n58314, n58315, n58316, n58317, n58318, n58319, n58320,
         n58321, n58322, n58323, n58324, n58325, n58326, n58327, n58328,
         n58329, n58330, n58331, n58332, n58333, n58334, n58335, n58336,
         n58337, n58338, n58339, n58340, n58341, n58342, n58343, n58344,
         n58345, n58346, n58347, n58348, n58349, n58350, n58351, n58352,
         n58353, n58354, n58355, n58356, n58357, n58358, n58359, n58360,
         n58361, n58362, n58363, n58364, n58365, n58366, n58367, n58368,
         n58369, n58370, n58371, n58372, n58373, n58374, n58375, n58376,
         n58377, n58378, n58379, n58380, n58381, n58382, n58383, n58384,
         n58385, n58386, n58387, n58388, n58389, n58390, n58391, n58392,
         n58393, n58394, n58395, n58396, n58397, n58398, n58399, n58400,
         n58401, n58402, n58403, n58404, n58405, n58406, n58407, n58408,
         n58409, n58410, n58411, n58412, n58413, n58414, n58415, n58416,
         n58417, n58418, n58419, n58420, n58421, n58422, n58423, n58424,
         n58425, n58426, n58427, n58428, n58429, n58430, n58431, n58432,
         n58433, n58434, n58435, n58436, n58437, n58438, n58439, n58440,
         n58441, n58442, n58443, n58444, n58445, n58446, n58447, n58448,
         n58449, n58450, n58451, n58452, n58453, n58454, n58455, n58456,
         n58457, n58458, n58459, n58460, n58461, n58462, n58463, n58464,
         n58465, n58466, n58467, n58468, n58469, n58470, n58471, n58472,
         n58473, n58474, n58475, n58476, n58477, n58478, n58479, n58480,
         n58481, n58482, n58483, n58484, n58485, n58486, n58487, n58488,
         n58489, n58490, n58491, n58492, n58493, n58494, n58495, n58496,
         n58497, n58498, n58499, n58500, n58501, n58502, n58503, n58504,
         n58505, n58506, n58507, n58508, n58509, n58510, n58511, n58512,
         n58513, n58514, n58515, n58516, n58517, n58518, n58519, n58520,
         n58521, n58522, n58523, n58524, n58525, n58526, n58527, n58528,
         n58529, n58530, n58531, n58532, n58533, n58534, n58535, n58536,
         n58537, n58538, n58539, n58540, n58541, n58542, n58543, n58544,
         n58545, n58546, n58547, n58548, n58549, n58550, n58551, n58552,
         n58553, n58554, n58555, n58556, n58557, n58558, n58559, n58560,
         n58561, n58562, n58563, n58564, n58565, n58566, n58567, n58568,
         n58569, n58570, n58571, n58572, n58573, n58574, n58575, n58576,
         n58577, n58578, n58579, n58580, n58581, n58582, n58583, n58584,
         n58585, n58586, n58587, n58588, n58589, n58590, n58591, n58592,
         n58593, n58594, n58595, n58596, n58597, n58598, n58599, n58600,
         n58601, n58602, n58603, n58604, n58605, n58606, n58607, n58608,
         n58609, n58610, n58611, n58612, n58613, n58614, n58615, n58616,
         n58617, n58618, n58619, n58620, n58621, n58622, n58623, n58624,
         n58625, n58626, n58627, n58628, n58629, n58630, n58631, n58632,
         n58633, n58634, n58635, n58636, n58637, n58638, n58639, n58640,
         n58641, n58642, n58643, n58644, n58645, n58646, n58647, n58648,
         n58649, n58650, n58651, n58652, n58653, n58654, n58655, n58656,
         n58657, n58658, n58659, n58660, n58661, n58662, n58663, n58664,
         n58665, n58666, n58667, n58668, n58669, n58670, n58671, n58672,
         n58673, n58674, n58675, n58676, n58677, n58678, n58679, n58680,
         n58681, n58682, n58683, n58684, n58685, n58686, n58687, n58688,
         n58689, n58690, n58691, n58692, n58693, n58694, n58695, n58696,
         n58697, n58698, n58699, n58700, n58701, n58702, n58703, n58704,
         n58705, n58706, n58707, n58708, n58709, n58710, n58711, n58712,
         n58713, n58714, n58715, n58716, n58717, n58718, n58719, n58720,
         n58721, n58722, n58723, n58724, n58725, n58726, n58727, n58728,
         n58729, n58730, n58731, n58732, n58733, n58734, n58735, n58736,
         n58737, n58738, n58739, n58740, n58741, n58742, n58743, n58744,
         n58745, n58746, n58747, n58748, n58749, n58750, n58751, n58752,
         n58753, n58754, n58755, n58756, n58757, n58758, n58759, n58760,
         n58761, n58762, n58763, n58764, n58765, n58766, n58767, n58768,
         n58769, n58770, n58771, n58772, n58773, n58774, n58775, n58776,
         n58777, n58778, n58779, n58780, n58781, n58782, n58783, n58784,
         n58785, n58786, n58787, n58788, n58789, n58790, n58791, n58792,
         n58793, n58794, n58795, n58796, n58797, n58798, n58799, n58800,
         n58801, n58802, n58803, n58804, n58805, n58806, n58807, n58808,
         n58809, n58810, n58811, n58812, n58813, n58814, n58815, n58816,
         n58817, n58818, n58819, n58820, n58821, n58822, n58823, n58824,
         n58825, n58826, n58827, n58828, n58829, n58830, n58831, n58832,
         n58833, n58834, n58835, n58836, n58837, n58838, n58839, n58840,
         n58841, n58842, n58843, n58844, n58845, n58846, n58847, n58848,
         n58849, n58850, n58851, n58852, n58853, n58854, n58855, n58856,
         n58857, n58858, n58859, n58860, n58861, n58862, n58863, n58864,
         n58865, n58866, n58867, n58868, n58869, n58870, n58871, n58872,
         n58873, n58874, n58875, n58876, n58877, n58878, n58879, n58880,
         n58881, n58882, n58883, n58884, n58885, n58886, n58887, n58888,
         n58889, n58890, n58891, n58892, n58893, n58894, n58895, n58896,
         n58897, n58898, n58899, n58900, n58901, n58902, n58903, n58904,
         n58905, n58906, n58907, n58908, n58909, n58910, n58911, n58912,
         n58913, n58914, n58915, n58916, n58917, n58918, n58919, n58920,
         n58921, n58922, n58923, n58924, n58925, n58926, n58927, n58928,
         n58929, n58930, n58931, n58932, n58933, n58934, n58935, n58936,
         n58937, n58938, n58939, n58940, n58941, n58942, n58943, n58944,
         n58945, n58946, n58947, n58948, n58949, n58950, n58951, n58952,
         n58953, n58954, n58955, n58956, n58957, n58958, n58959, n58960,
         n58961, n58962, n58963, n58964, n58965, n58966, n58967, n58968,
         n58969, n58970, n58971, n58972, n58973, n58974, n58975, n58976,
         n58977, n58978, n58979, n58980, n58981, n58982, n58983, n58984,
         n58985, n58986, n58987, n58988, n58989, n58990, n58991, n58992,
         n58993, n58994, n58995, n58996, n58997, n58998, n58999, n59000,
         n59001, n59002, n59003, n59004, n59005, n59006, n59007, n59008,
         n59009, n59010, n59011, n59012, n59013, n59014, n59015, n59016,
         n59017, n59018, n59019, n59020, n59021, n59022, n59023, n59024,
         n59025, n59026, n59027, n59028, n59029, n59030, n59031, n59032,
         n59033, n59034, n59035, n59036, n59037, n59038, n59039, n59040,
         n59041, n59042, n59043, n59044, n59045, n59046, n59047, n59048,
         n59049, n59050, n59051, n59052, n59053, n59054, n59055, n59056,
         n59057, n59058, n59059, n59060, n59061, n59062, n59063, n59064,
         n59065, n59066, n59067, n59068, n59069, n59070, n59071, n59072,
         n59073, n59074, n59075, n59076, n59077, n59078, n59079, n59080,
         n59081, n59082, n59083, n59084, n59085, n59086, n59087, n59088,
         n59089, n59090, n59091, n59092, n59093, n59094, n59095, n59096,
         n59097, n59098, n59099, n59100, n59101, n59102, n59103, n59104,
         n59105, n59106, n59107, n59108, n59109, n59110, n59111, n59112,
         n59113, n59114, n59115, n59116, n59117, n59118, n59119, n59120,
         n59121, n59122, n59123, n59124, n59125, n59126, n59127, n59128,
         n59129, n59130, n59131, n59132, n59133, n59134, n59135, n59136,
         n59137, n59138, n59139, n59140, n59141, n59142, n59143, n59144,
         n59145, n59146, n59147, n59148, n59149, n59150, n59151, n59152,
         n59153, n59154, n59155, n59156, n59157, n59158, n59159, n59160,
         n59161, n59162, n59163, n59164, n59165, n59166, n59167, n59168,
         n59169, n59170, n59171, n59172, n59173, n59174, n59175, n59176,
         n59177, n59178, n59179, n59180, n59181, n59182, n59183, n59184,
         n59185, n59186, n59187, n59188, n59189, n59190, n59191, n59192,
         n59193, n59194, n59195, n59196, n59197, n59198, n59199, n59200,
         n59201, n59202, n59203, n59204, n59205, n59206, n59207, n59208,
         n59209, n59210, n59211, n59212, n59213, n59214, n59215, n59216,
         n59217, n59218, n59219, n59220, n59221, n59222, n59223, n59224,
         n59225, n59226, n59227, n59228, n59229, n59230, n59231, n59232,
         n59233, n59234, n59235, n59236, n59237, n59238, n59239, n59240,
         n59241, n59242, n59243, n59244, n59245, n59246, n59247, n59248,
         n59249, n59250, n59251, n59252, n59253, n59254, n59255, n59256,
         n59257, n59258, n59259, n59260, n59261, n59262, n59263, n59264,
         n59265, n59266, n59267, n59268, n59269, n59270, n59271, n59272,
         n59273, n59274, n59275, n59276, n59277, n59278, n59279, n59280,
         n59281, n59282, n59283, n59284, n59285, n59286, n59287, n59288,
         n59289, n59290, n59291, n59292, n59293, n59294, n59295, n59296,
         n59297, n59298, n59299, n59300, n59301, n59302, n59303, n59304,
         n59305, n59306, n59307, n59308, n59309, n59310, n59311, n59312,
         n59313, n59314, n59315, n59316, n59317, n59318, n59319, n59320,
         n59321, n59322, n59323, n59324, n59325, n59326, n59327, n59328,
         n59329, n59330, n59331, n59332, n59333, n59334, n59335, n59336,
         n59337, n59338, n59339, n59340, n59341, n59343, n59344, n59345,
         n59346, n59347, n59348, n59349, n59350, n59351, n59352, n59353,
         n59354, n59355, n59356, n59357, n59358, n59359, n59360, n59361,
         n59362, n59363, n59364, n59365, n59366, n59367, n59368, n59369,
         n59370, n59371, n59372, n59373, n59374, n59375, n59376, n59377,
         n59378, n59379, n59380, n59381, n59382, n59383, n59384, n59385,
         n59386, n59387, n59388, n59389, n59390, n59391, n59392, n59393,
         n59394, n59395, n59396, n59397, n59398, n59399, n59400, n59401,
         n59402, n59403, n59404, n59405, n59406, n59407, n59408, n59409,
         n59410, n59411, n59412, n59413, n59414, n59415, n59416, n59417,
         n59418, n59419, n59420, n59421, n59422, n59423, n59424, n59425,
         n59426, n59427, n59428, n59429, n59430, n59431, n59432, n59433,
         n59434, n59435, n59436, n59437, n59438, n59439, n59440, n59441,
         n59442, n59443, n59444, n59445, n59446, n59447, n59448, n59449,
         n59450, n59451, n59452, n59453, n59454, n59455, n59456, n59457,
         n59458, n59459, n59460, n59461, n59462, n59463, n59464, n59465,
         n59466, n59467, n59468, n59469, n59470, n59471, n59472, n59473,
         n59474, n59475, n59476, n59477, n59478, n59479, n59480, n59481,
         n59482, n59483, n59484, n59485, n59486, n59487, n59488, n59489,
         n59490, n59491, n59492, n59493, n59494, n59495, n59496, n59497,
         n59498, n59499, n59500, n59501, n59502, n59503, n59504, n59505,
         n59506, n59507, n59508, n59509, n59510, n59511, n59512, n59513,
         n59514, n59515, n59516, n59517, n59518, n59519, n59520, n59521,
         n59522, n59523, n59524, n59525, n59526, n59527, n59528, n59529,
         n59530, n59531, n59532, n59533, n59534, n59535, n59536, n59537,
         n59538, n59539, n59540, n59541, n59542, n59543, n59544, n59545,
         n59546, n59547, n59548, n59549, n59550, n59551, n59552, n59553,
         n59554, n59555, n59556, n59557, n59558, n59559, n59560, n59561,
         n59562, n59563, n59564, n59565, n59566, n59567, n59568, n59569,
         n59570, n59571, n59572, n59573, n59574, n59575, n59576, n59577,
         n59578, n59579, n59580, n59581, n59582, n59583, n59584, n59585,
         n59586, n59587, n59588, n59589, n59590, n59591, n59592, n59593,
         n59594, n59595, n59596, n59597, n59598, n59599, n59600, n59601,
         n59602, n59603, n59604, n59605, n59606, n59607, n59608, n59609,
         n59610, n59611, n59612, n59613, n59614, n59615, n59616, n59617,
         n59618, n59619, n59620, n59621, n59622, n59623, n59624, n59625,
         n59626, n59627, n59628, n59629, n59630, n59631, n59632, n59633,
         n59634, n59635, n59636, n59637, n59638, n59639, n59640, n59641,
         n59642, n59643, n59644, n59645, n59646, n59647, n59648, n59649,
         n59650, n59651, n59652, n59653, n59654, n59655, n59656, n59657,
         n59658, n59659, n59660, n59661, n59662, n59663, n59664, n59665,
         n59666, n59667, n59668, n59669, n59670, n59671, n59672, n59673,
         n59674, n59675, n59676, n59677, n59678, n59679, n59680, n59681,
         n59682, n59683, n59684, n59685, n59686, n59687, n59688, n59689,
         n59690, n59691, n59692, n59693, n59694, n59695, n59696, n59697,
         n59698, n59699, n59700, n59701, n59702, n59703, n59704, n59705,
         n59706, n59707, n59708, n59709, n59710, n59711, n59712, n59713,
         n59714, n59715, n59716, n59717, n59718, n59719, n59720, n59721,
         n59722, n59723, n59724, n59725, n59726, n59727, n59728, n59729,
         n59730, n59731, n59732, n59733, n59734, n59735, n59736, n59737,
         n59738, n59739, n59740, n59741, n59742, n59743, n59744, n59745,
         n59746, n59747, n59748, n59749, n59750, n59751, n59752, n59753,
         n59754, n59755, n59756, n59757, n59758, n59759, n59760, n59761,
         n59762, n59763, n59764, n59765, n59766, n59767, n59768, n59769,
         n59770, n59771, n59772, n59773, n59774, n59775, n59776, n59777,
         n59778, n59779, n59780, n59781, n59782, n59783, n59784, n59785,
         n59786, n59787, n59788, n59789, n59790, n59791, n59792, n59793,
         n59794, n59795, n59796, n59797, n59798, n59799, n59800, n59801,
         n59802, n59803, n59804, n59805, n59806, n59807, n59808, n59809,
         n59810, n59811, n59812, n59813, n59814, n59815, n59816, n59817,
         n59818, n59819, n59820, n59821, n59822, n59823, n59824, n59825,
         n59826, n59827, n59828, n59829, n59830, n59831, n59832, n59833,
         n59834, n59835, n59836, n59837, n59838, n59839, n59840, n59841,
         n59842, n59843, n59844, n59845, n59846, n59847, n59848, n59849,
         n59850, n59851, n59852, n59853, n59854, n59855, n59856, n59857,
         n59858, n59859, n59860, n59861, n59862, n59863, n59864, n59865,
         n59866, n59867, n59868, n59869, n59870, n59871, n59872, n59873,
         n59874, n59875, n59876, n59877, n59878, n59879, n59880, n59881,
         n59882, n59883, n59884, n59885, n59886, n59887, n59888, n59889,
         n59890, n59891, n59892, n59893, n59894, n59895, n59896, n59897,
         n59898, n59899, n59900, n59901, n59902, n59903, n59904, n59905,
         n59906, n59907, n59908, n59909, n59910, n59911, n59912, n59913,
         n59914, n59915, n59916, n59917, n59918, n59919, n59920, n59921,
         n59922, n59923, n59924, n59925, n59926, n59927, n59928, n59929,
         n59930, n59931, n59932, n59933, n59934, n59935, n59936, n59937,
         n59938, n59939, n59940, n59941, n59942, n59943, n59944, n59945,
         n59946, n59947, n59948, n59949, n59950, n59951, n59952, n59953,
         n59954, n59955, n59956, n59957, n59958, n59959, n59960, n59961,
         n59962, n59963, n59964, n59965, n59966, n59967, n59968, n59969,
         n59970, n59971, n59972, n59973, n59974, n59975, n59976, n59977,
         n59978, n59979, n59980, n59981, n59982, n59983, n59984, n59985,
         n59986, n59987, n59988, n59989, n59990, n59991, n59992, n59993,
         n59994, n59995, n59996, n59997, n59998, n59999, n60000, n60001,
         n60002, n60003, n60004, n60005, n60006, n60007, n60008, n60009,
         n60010, n60011, n60012, n60013, n60014, n60015, n60016, n60017,
         n60018, n60019, n60020, n60021, n60022, n60023, n60024, n60025,
         n60026, n60027, n60028, n60029, n60030, n60031, n60032, n60033,
         n60034, n60035, n60036, n60037, n60038, n60039, n60040, n60041,
         n60042, n60043, n60044, n60045, n60046, n60047, n60048, n60049,
         n60050, n60051, n60052, n60053, n60054, n60055, n60056, n60057,
         n60058, n60059, n60060, n60061, n60062, n60063, n60064, n60065,
         n60066, n60067, n60068, n60069, n60070, n60071, n60072, n60073,
         n60074, n60075, n60076, n60077, n60078, n60079, n60080, n60081,
         n60082, n60083, n60084, n60085, n60086, n60087, n60088, n60089,
         n60090, n60091, n60092, n60093, n60094, n60095, n60096, n60097,
         n60098, n60099, n60100, n60101, n60102, n60103, n60104, n60105,
         n60106, n60107, n60108, n60109, n60110;
  wire   [32:1] ao1;
  wire   [32:1] go1;
  wire   [32:1] bo1;
  wire   [1:31] poh1;
  wire   [1:31] pov1;
  wire   [32:1] ao2;
  wire   [32:1] go2;
  wire   [32:1] bo2;
  wire   [1:31] poh2;
  wire   [1:31] pov2;
  wire   [32:1] ao3;
  wire   [32:1] go3;
  wire   [32:1] bo3;
  wire   [1:31] poh3;
  wire   [1:31] pov3;
  wire   [32:1] ao4;
  wire   [32:1] go4;
  wire   [32:1] bo4;
  wire   [1:31] poh4;
  wire   [1:31] pov4;
  wire   [32:1] ao5;
  wire   [32:1] go5;
  wire   [32:1] bo5;
  wire   [1:31] poh5;
  wire   [1:31] pov5;
  wire   [32:1] bo6;
  wire   [1:31] poh6;
  wire   [1:31] \pe1/poht ;
  wire   [32:1] \pe1/got ;
  wire   [32:1] \pe1/aot ;
  wire   [1:31] \pe1/ti_7t ;
  wire   [1:31] \pe2/poht ;
  wire   [32:1] \pe2/got ;
  wire   [32:1] \pe2/aot ;
  wire   [1:31] \pe2/ti_7t ;
  wire   [1:31] \pe2/phq ;
  wire   [1:31] \pe2/pvq ;
  wire   [1:31] \pe3/poht ;
  wire   [32:1] \pe3/got ;
  wire   [32:1] \pe3/aot ;
  wire   [1:31] \pe3/ti_7t ;
  wire   [1:31] \pe3/phq ;
  wire   [1:31] \pe3/pvq ;
  wire   [1:31] \pe4/poht ;
  wire   [32:1] \pe4/got ;
  wire   [32:1] \pe4/aot ;
  wire   [1:31] \pe4/ti_7t ;
  wire   [1:31] \pe4/phq ;
  wire   [1:31] \pe4/pvq ;
  wire   [1:31] \pe5/poht ;
  wire   [32:1] \pe5/got ;
  wire   [32:1] \pe5/aot ;
  wire   [1:31] \pe5/ti_7t ;
  wire   [1:31] \pe5/phq ;
  wire   [1:31] \pe5/pvq ;
  wire   [1:31] \pe6/poht ;
  wire   [32:1] \pe6/got ;
  wire   [32:1] \pe6/aot ;
  wire   [1:31] \pe6/ti_7t ;
  wire   [1:31] \pe6/phq ;
  wire   [1:31] \pe6/pvq ;

  DRNQHSV4 \pe1/pe1/q_reg[32]  ( .D(ai[1]), .CK(clk), .RDN(n59649), .Q(
        \pe1/aot [1]) );
  DRNQHSV4 \pe1/pe1/q_reg[30]  ( .D(ai[3]), .CK(clk), .RDN(n59447), .Q(
        \pe1/aot [3]) );
  DRNQHSV4 \pe1/pe1/q_reg[29]  ( .D(ai[4]), .CK(clk), .RDN(n59476), .Q(
        \pe1/aot [4]) );
  DRNQHSV4 \pe1/pe1/q_reg[28]  ( .D(ai[5]), .CK(clk), .RDN(n59434), .Q(
        \pe1/aot [5]) );
  DRNQHSV4 \pe1/pe1/q_reg[27]  ( .D(ai[6]), .CK(clk), .RDN(rst), .Q(
        \pe1/aot [6]) );
  DRNQHSV4 \pe1/pe1/q_reg[26]  ( .D(ai[7]), .CK(clk), .RDN(n59436), .Q(
        \pe1/aot [7]) );
  DRNQHSV4 \pe1/pe1/q_reg[25]  ( .D(ai[8]), .CK(clk), .RDN(n59424), .Q(
        \pe1/aot [8]) );
  DRNQHSV4 \pe1/pe1/q_reg[24]  ( .D(ai[9]), .CK(clk), .RDN(n59492), .Q(
        \pe1/aot [9]) );
  DRNQHSV4 \pe1/pe1/q_reg[23]  ( .D(ai[10]), .CK(clk), .RDN(n59438), .Q(
        \pe1/aot [10]) );
  DRNQHSV4 \pe1/pe1/q_reg[22]  ( .D(ai[11]), .CK(clk), .RDN(n59437), .Q(
        \pe1/aot [11]) );
  DRNQHSV4 \pe1/pe1/q_reg[21]  ( .D(ai[12]), .CK(clk), .RDN(n59429), .Q(
        \pe1/aot [12]) );
  DRNQHSV4 \pe1/pe1/q_reg[20]  ( .D(ai[13]), .CK(clk), .RDN(n59446), .Q(
        \pe1/aot [13]) );
  DRNQHSV4 \pe1/pe1/q_reg[19]  ( .D(ai[14]), .CK(clk), .RDN(n59397), .Q(
        \pe1/aot [14]) );
  DRNQHSV4 \pe1/pe1/q_reg[18]  ( .D(ai[15]), .CK(clk), .RDN(n59491), .Q(
        \pe1/aot [15]) );
  DRNQHSV4 \pe1/pe1/q_reg[17]  ( .D(ai[16]), .CK(clk), .RDN(n59424), .Q(
        \pe1/aot [16]) );
  DRNQHSV4 \pe1/pe1/q_reg[16]  ( .D(ai[17]), .CK(clk), .RDN(n59496), .Q(
        \pe1/aot [17]) );
  DRNQHSV4 \pe1/pe1/q_reg[15]  ( .D(ai[18]), .CK(clk), .RDN(n59458), .Q(
        \pe1/aot [18]) );
  DRNQHSV4 \pe1/pe1/q_reg[14]  ( .D(ai[19]), .CK(clk), .RDN(n59659), .Q(
        \pe1/aot [19]) );
  DRNQHSV4 \pe1/pe1/q_reg[13]  ( .D(ai[20]), .CK(clk), .RDN(n59496), .Q(
        \pe1/aot [20]) );
  DRNQHSV4 \pe1/pe1/q_reg[12]  ( .D(ai[21]), .CK(clk), .RDN(n59512), .Q(
        \pe1/aot [21]) );
  DRNQHSV4 \pe1/pe1/q_reg[11]  ( .D(ai[22]), .CK(clk), .RDN(n59496), .Q(
        \pe1/aot [22]) );
  DRNQHSV4 \pe1/pe1/q_reg[10]  ( .D(ai[23]), .CK(clk), .RDN(rst), .Q(
        \pe1/aot [23]) );
  DRNQHSV4 \pe1/pe1/q_reg[9]  ( .D(ai[24]), .CK(clk), .RDN(n59448), .Q(
        \pe1/aot [24]) );
  DRNQHSV4 \pe1/pe1/q_reg[8]  ( .D(ai[25]), .CK(clk), .RDN(n59425), .Q(
        \pe1/aot [25]) );
  DRNQHSV4 \pe1/pe1/q_reg[7]  ( .D(ai[26]), .CK(clk), .RDN(n59442), .Q(
        \pe1/aot [26]) );
  DRNQHSV4 \pe1/pe1/q_reg[6]  ( .D(ai[27]), .CK(clk), .RDN(n59418), .Q(
        \pe1/aot [27]) );
  DRNQHSV4 \pe1/pe1/q_reg[5]  ( .D(ai[28]), .CK(clk), .RDN(n59454), .Q(
        \pe1/aot [28]) );
  DRNQHSV4 \pe1/pe1/q_reg[4]  ( .D(ai[29]), .CK(clk), .RDN(n29733), .Q(
        \pe1/aot [29]) );
  DRNQHSV4 \pe1/pe1/q_reg[3]  ( .D(ai[30]), .CK(clk), .RDN(n59448), .Q(
        \pe1/aot [30]) );
  DRNQHSV4 \pe1/pe1/q_reg[2]  ( .D(ai[31]), .CK(clk), .RDN(n59925), .Q(
        \pe1/aot [31]) );
  DRNQHSV4 \pe1/pe1/q_reg[1]  ( .D(ai[32]), .CK(clk), .RDN(n29731), .Q(
        \pe1/aot [32]) );
  DRNQHSV4 \pe1/pe2/q_reg[32]  ( .D(gi[1]), .CK(clk), .RDN(n59494), .Q(
        \pe1/got [1]) );
  DRNQHSV4 \pe1/pe2/q_reg[31]  ( .D(gi[2]), .CK(clk), .RDN(rst), .Q(
        \pe1/got [2]) );
  DRNQHSV4 \pe1/pe2/q_reg[30]  ( .D(gi[3]), .CK(clk), .RDN(n59434), .Q(
        \pe1/got [3]) );
  DRNQHSV4 \pe1/pe2/q_reg[29]  ( .D(gi[4]), .CK(clk), .RDN(rst), .Q(
        \pe1/got [4]) );
  DRNQHSV4 \pe1/pe2/q_reg[28]  ( .D(gi[5]), .CK(clk), .RDN(n59452), .Q(
        \pe1/got [5]) );
  DRNQHSV4 \pe1/pe2/q_reg[27]  ( .D(gi[6]), .CK(clk), .RDN(rst), .Q(
        \pe1/got [6]) );
  DRNQHSV4 \pe1/pe2/q_reg[26]  ( .D(gi[7]), .CK(clk), .RDN(n59424), .Q(
        \pe1/got [7]) );
  DRNQHSV4 \pe1/pe2/q_reg[25]  ( .D(gi[8]), .CK(clk), .RDN(rst), .Q(
        \pe1/got [8]) );
  DRNQHSV4 \pe1/pe2/q_reg[24]  ( .D(gi[9]), .CK(clk), .RDN(rst), .Q(
        \pe1/got [9]) );
  DRNQHSV4 \pe1/pe2/q_reg[23]  ( .D(gi[10]), .CK(clk), .RDN(n59925), .Q(
        \pe1/got [10]) );
  DRNQHSV4 \pe1/pe2/q_reg[22]  ( .D(gi[11]), .CK(clk), .RDN(n59490), .Q(
        \pe1/got [11]) );
  DRNQHSV4 \pe1/pe2/q_reg[21]  ( .D(gi[12]), .CK(clk), .RDN(n59490), .Q(
        \pe1/got [12]) );
  DRNQHSV4 \pe1/pe2/q_reg[20]  ( .D(gi[13]), .CK(clk), .RDN(n59493), .Q(
        \pe1/got [13]) );
  DRNQHSV4 \pe1/pe2/q_reg[19]  ( .D(gi[14]), .CK(clk), .RDN(n59404), .Q(
        \pe1/got [14]) );
  DRNQHSV4 \pe1/pe2/q_reg[18]  ( .D(gi[15]), .CK(clk), .RDN(n59492), .Q(
        \pe1/got [15]) );
  DRNQHSV4 \pe1/pe2/q_reg[17]  ( .D(gi[16]), .CK(clk), .RDN(n59483), .Q(
        \pe1/got [16]) );
  DRNQHSV4 \pe1/pe2/q_reg[16]  ( .D(gi[17]), .CK(clk), .RDN(rst), .Q(
        \pe1/got [17]) );
  DRNQHSV4 \pe1/pe2/q_reg[15]  ( .D(gi[18]), .CK(clk), .RDN(n59445), .Q(
        \pe1/got [18]) );
  DRNQHSV4 \pe1/pe2/q_reg[14]  ( .D(gi[19]), .CK(clk), .RDN(n29730), .Q(
        \pe1/got [19]) );
  DRNQHSV4 \pe1/pe2/q_reg[13]  ( .D(gi[20]), .CK(clk), .RDN(n59446), .Q(
        \pe1/got [20]) );
  DRNQHSV4 \pe1/pe2/q_reg[12]  ( .D(gi[21]), .CK(clk), .RDN(n59411), .Q(
        \pe1/got [21]) );
  DRNQHSV4 \pe1/pe2/q_reg[11]  ( .D(gi[22]), .CK(clk), .RDN(n59467), .Q(
        \pe1/got [22]) );
  DRNQHSV4 \pe1/pe2/q_reg[10]  ( .D(gi[23]), .CK(clk), .RDN(n59653), .Q(
        \pe1/got [23]) );
  DRNQHSV4 \pe1/pe2/q_reg[9]  ( .D(gi[24]), .CK(clk), .RDN(n59458), .Q(
        \pe1/got [24]) );
  DRNQHSV4 \pe1/pe2/q_reg[8]  ( .D(gi[25]), .CK(clk), .RDN(n29732), .Q(
        \pe1/got [25]) );
  DRNQHSV4 \pe1/pe2/q_reg[7]  ( .D(gi[26]), .CK(clk), .RDN(n59651), .Q(
        \pe1/got [26]) );
  DRNQHSV4 \pe1/pe2/q_reg[6]  ( .D(gi[27]), .CK(clk), .RDN(n59460), .Q(
        \pe1/got [27]) );
  DRNQHSV4 \pe1/pe2/q_reg[5]  ( .D(gi[28]), .CK(clk), .RDN(rst), .Q(
        \pe1/got [28]) );
  DRNQHSV4 \pe1/pe2/q_reg[4]  ( .D(gi[29]), .CK(clk), .RDN(n59656), .Q(
        \pe1/got [29]) );
  DRNQHSV4 \pe1/pe2/q_reg[3]  ( .D(gi[30]), .CK(clk), .RDN(n59659), .Q(
        \pe1/got [30]) );
  DRNQHSV4 \pe1/pe2/q_reg[2]  ( .D(gi[31]), .CK(clk), .RDN(n29732), .Q(
        \pe1/got [31]) );
  DRNQHSV4 \pe1/pe2/q_reg[1]  ( .D(gi[32]), .CK(clk), .RDN(n59414), .Q(
        \pe1/got [32]) );
  DRNQHSV4 \pe1/pe8/q_reg  ( .D(\pe1/ctrq ), .CK(clk), .RDN(n59496), .Q(ctro1)
         );
  DRNQHSV4 \pe1/pe12/q_reg[32]  ( .D(n59718), .CK(clk), .RDN(n59397), .Q(
        \pe1/bq[1] ) );
  DRNQHSV4 \pe1/pe12/q_reg[31]  ( .D(n59719), .CK(clk), .RDN(n59493), .Q(
        \pe1/bq[2] ) );
  DRNQHSV4 \pe1/pe12/q_reg[30]  ( .D(n59720), .CK(clk), .RDN(n59463), .Q(
        \pe1/bq[3] ) );
  DRNQHSV4 \pe1/pe12/q_reg[29]  ( .D(n59717), .CK(clk), .RDN(n59461), .Q(
        \pe1/bq[4] ) );
  DRNQHSV4 \pe1/pe12/q_reg[28]  ( .D(n59715), .CK(clk), .RDN(n29730), .Q(
        \pe1/bq[5] ) );
  DRNQHSV4 \pe1/pe12/q_reg[27]  ( .D(n59714), .CK(clk), .RDN(n59478), .Q(
        \pe1/bq[6] ) );
  DRNQHSV4 \pe1/pe12/q_reg[26]  ( .D(n59716), .CK(clk), .RDN(n59510), .Q(
        \pe1/bq[7] ) );
  DRNQHSV4 \pe1/pe12/q_reg[25]  ( .D(n59711), .CK(clk), .RDN(n59510), .Q(
        \pe1/bq[8] ) );
  DRNQHSV4 \pe1/pe12/q_reg[23]  ( .D(n59713), .CK(clk), .RDN(n59480), .Q(
        \pe1/bq[10] ) );
  DRNQHSV4 \pe1/pe12/q_reg[21]  ( .D(n59709), .CK(clk), .RDN(n59656), .Q(
        \pe1/bq[12] ) );
  DRNQHSV4 \pe1/pe12/q_reg[20]  ( .D(n59707), .CK(clk), .RDN(n59474), .Q(
        \pe1/bq[13] ) );
  DRNQHSV4 \pe1/pe12/q_reg[19]  ( .D(n59708), .CK(clk), .RDN(n59510), .Q(
        \pe1/bq[14] ) );
  DRNQHSV4 \pe1/pe12/q_reg[18]  ( .D(n59706), .CK(clk), .RDN(n59455), .Q(
        \pe1/bq[15] ) );
  DRNQHSV4 \pe1/pe12/q_reg[17]  ( .D(n59705), .CK(clk), .RDN(n59463), .Q(
        \pe1/bq[16] ) );
  DRNQHSV4 \pe1/pe12/q_reg[16]  ( .D(n59703), .CK(clk), .RDN(n59396), .Q(
        \pe1/bq[17] ) );
  DRNQHSV4 \pe1/pe12/q_reg[14]  ( .D(n59702), .CK(clk), .RDN(n59659), .Q(
        \pe1/bq[19] ) );
  DRNQHSV4 \pe1/pe12/q_reg[13]  ( .D(n59701), .CK(clk), .RDN(n59433), .Q(
        \pe1/bq[20] ) );
  DRNQHSV4 \pe1/pe12/q_reg[11]  ( .D(n59700), .CK(clk), .RDN(n59492), .Q(
        \pe1/bq[22] ) );
  DRNQHSV4 \pe1/pe12/q_reg[10]  ( .D(n59698), .CK(clk), .RDN(n59436), .Q(
        \pe1/bq[23] ) );
  DRNQHSV4 \pe1/pe12/q_reg[9]  ( .D(n59696), .CK(clk), .RDN(n59512), .Q(
        \pe1/bq[24] ) );
  DRNQHSV4 \pe1/pe12/q_reg[8]  ( .D(n59697), .CK(clk), .RDN(n59450), .Q(
        \pe1/bq[25] ) );
  DRNQHSV4 \pe1/pe12/q_reg[7]  ( .D(n59695), .CK(clk), .RDN(n59431), .Q(
        \pe1/bq[26] ) );
  DRNQHSV4 \pe1/pe12/q_reg[6]  ( .D(n59694), .CK(clk), .RDN(n59512), .Q(
        \pe1/bq[27] ) );
  DRNQHSV4 \pe1/pe12/q_reg[5]  ( .D(n59689), .CK(clk), .RDN(n59491), .Q(
        \pe1/bq[28] ) );
  DRNQHSV4 \pe1/pe12/q_reg[4]  ( .D(n59693), .CK(clk), .RDN(n59413), .Q(
        \pe1/bq[29] ) );
  DRNQHSV4 \pe1/pe12/q_reg[2]  ( .D(n59690), .CK(clk), .RDN(n59659), .Q(
        \pe1/bq[31] ) );
  DRNQHSV4 \pe1/pe12/q_reg[1]  ( .D(n59692), .CK(clk), .RDN(n59439), .Q(
        \pe1/bq[32] ) );
  DRNQHSV4 \pe1/pe14/q_reg[1]  ( .D(n59675), .CK(clk), .RDN(n59472), .Q(
        \pe1/ti_7t [1]) );
  DRNQHSV4 \pe2/pe1/q_reg[32]  ( .D(ao1[1]), .CK(clk), .RDN(n59654), .Q(
        \pe2/aot [1]) );
  DRNQHSV4 \pe2/pe1/q_reg[30]  ( .D(ao1[3]), .CK(clk), .RDN(n59399), .Q(
        \pe2/aot [3]) );
  DRNQHSV4 \pe2/pe1/q_reg[29]  ( .D(ao1[4]), .CK(clk), .RDN(n59414), .Q(
        \pe2/aot [4]) );
  DRNQHSV4 \pe2/pe1/q_reg[28]  ( .D(ao1[5]), .CK(clk), .RDN(n59410), .Q(
        \pe2/aot [5]) );
  DRNQHSV4 \pe2/pe1/q_reg[27]  ( .D(ao1[6]), .CK(clk), .RDN(n59438), .Q(
        \pe2/aot [6]) );
  DRNQHSV4 \pe2/pe1/q_reg[26]  ( .D(ao1[7]), .CK(clk), .RDN(n59414), .Q(
        \pe2/aot [7]) );
  DRNQHSV4 \pe2/pe1/q_reg[25]  ( .D(ao1[8]), .CK(clk), .RDN(n59455), .Q(
        \pe2/aot [8]) );
  DRNQHSV4 \pe2/pe1/q_reg[24]  ( .D(ao1[9]), .CK(clk), .RDN(n59476), .Q(
        \pe2/aot [9]) );
  DRNQHSV4 \pe2/pe1/q_reg[23]  ( .D(ao1[10]), .CK(clk), .RDN(n59480), .Q(
        \pe2/aot [10]) );
  DRNQHSV4 \pe2/pe1/q_reg[22]  ( .D(ao1[11]), .CK(clk), .RDN(n59468), .Q(
        \pe2/aot [11]) );
  DRNQHSV4 \pe2/pe1/q_reg[21]  ( .D(ao1[12]), .CK(clk), .RDN(n59469), .Q(
        \pe2/aot [12]) );
  DRNQHSV4 \pe2/pe1/q_reg[20]  ( .D(ao1[13]), .CK(clk), .RDN(n59653), .Q(
        \pe2/aot [13]) );
  DRNQHSV4 \pe2/pe1/q_reg[19]  ( .D(ao1[14]), .CK(clk), .RDN(n59474), .Q(
        \pe2/aot [14]) );
  DRNQHSV4 \pe2/pe1/q_reg[18]  ( .D(ao1[15]), .CK(clk), .RDN(n59404), .Q(
        \pe2/aot [15]) );
  DRNQHSV4 \pe2/pe1/q_reg[17]  ( .D(ao1[16]), .CK(clk), .RDN(n59471), .Q(
        \pe2/aot [16]) );
  DRNQHSV4 \pe2/pe1/q_reg[16]  ( .D(ao1[17]), .CK(clk), .RDN(n59418), .Q(
        \pe2/aot [17]) );
  DRNQHSV4 \pe2/pe1/q_reg[15]  ( .D(ao1[18]), .CK(clk), .RDN(n59431), .Q(
        \pe2/aot [18]) );
  DRNQHSV4 \pe2/pe1/q_reg[14]  ( .D(ao1[19]), .CK(clk), .RDN(n59474), .Q(
        \pe2/aot [19]) );
  DRNQHSV4 \pe2/pe1/q_reg[13]  ( .D(ao1[20]), .CK(clk), .RDN(n29730), .Q(
        \pe2/aot [20]) );
  DRNQHSV4 \pe2/pe1/q_reg[12]  ( .D(ao1[21]), .CK(clk), .RDN(n59463), .Q(
        \pe2/aot [21]) );
  DRNQHSV4 \pe2/pe1/q_reg[11]  ( .D(ao1[22]), .CK(clk), .RDN(n59434), .Q(
        \pe2/aot [22]) );
  DRNQHSV4 \pe2/pe1/q_reg[10]  ( .D(ao1[23]), .CK(clk), .RDN(n59449), .Q(
        \pe2/aot [23]) );
  DRNQHSV4 \pe2/pe1/q_reg[9]  ( .D(ao1[24]), .CK(clk), .RDN(n59454), .Q(
        \pe2/aot [24]) );
  DRNQHSV4 \pe2/pe1/q_reg[8]  ( .D(ao1[25]), .CK(clk), .RDN(n59454), .Q(
        \pe2/aot [25]) );
  DRNQHSV4 \pe2/pe1/q_reg[7]  ( .D(ao1[26]), .CK(clk), .RDN(n59438), .Q(
        \pe2/aot [26]) );
  DRNQHSV4 \pe2/pe1/q_reg[6]  ( .D(ao1[27]), .CK(clk), .RDN(n59417), .Q(
        \pe2/aot [27]) );
  DRNQHSV4 \pe2/pe1/q_reg[5]  ( .D(ao1[28]), .CK(clk), .RDN(n59413), .Q(
        \pe2/aot [28]) );
  DRNQHSV4 \pe2/pe1/q_reg[4]  ( .D(ao1[29]), .CK(clk), .RDN(n59411), .Q(
        \pe2/aot [29]) );
  DRNQHSV4 \pe2/pe1/q_reg[3]  ( .D(ao1[30]), .CK(clk), .RDN(n59410), .Q(
        \pe2/aot [30]) );
  DRNQHSV4 \pe2/pe1/q_reg[2]  ( .D(ao1[31]), .CK(clk), .RDN(n59405), .Q(
        \pe2/aot [31]) );
  DRNQHSV4 \pe2/pe1/q_reg[1]  ( .D(ao1[32]), .CK(clk), .RDN(n59922), .Q(
        \pe2/aot [32]) );
  DRNQHSV4 \pe2/pe2/q_reg[32]  ( .D(go1[1]), .CK(clk), .RDN(n59469), .Q(
        \pe2/got [1]) );
  DRNQHSV4 \pe2/pe2/q_reg[31]  ( .D(go1[2]), .CK(clk), .RDN(n59484), .Q(
        \pe2/got [2]) );
  DRNQHSV4 \pe2/pe2/q_reg[30]  ( .D(go1[3]), .CK(clk), .RDN(n59491), .Q(
        \pe2/got [3]) );
  DRNQHSV4 \pe2/pe2/q_reg[29]  ( .D(go1[4]), .CK(clk), .RDN(n59482), .Q(
        \pe2/got [4]) );
  DRNQHSV4 \pe2/pe2/q_reg[28]  ( .D(go1[5]), .CK(clk), .RDN(n59482), .Q(
        \pe2/got [5]) );
  DRNQHSV4 \pe2/pe2/q_reg[27]  ( .D(go1[6]), .CK(clk), .RDN(n59403), .Q(
        \pe2/got [6]) );
  DRNQHSV4 \pe2/pe2/q_reg[26]  ( .D(go1[7]), .CK(clk), .RDN(n59403), .Q(
        \pe2/got [7]) );
  DRNQHSV4 \pe2/pe2/q_reg[25]  ( .D(go1[8]), .CK(clk), .RDN(n59396), .Q(
        \pe2/got [8]) );
  DRNQHSV4 \pe2/pe2/q_reg[24]  ( .D(go1[9]), .CK(clk), .RDN(n59452), .Q(
        \pe2/got [9]) );
  DRNQHSV4 \pe2/pe2/q_reg[23]  ( .D(go1[10]), .CK(clk), .RDN(n59397), .Q(
        \pe2/got [10]) );
  DRNQHSV4 \pe2/pe2/q_reg[22]  ( .D(go1[11]), .CK(clk), .RDN(n59416), .Q(
        \pe2/got [11]) );
  DRNQHSV4 \pe2/pe2/q_reg[21]  ( .D(go1[12]), .CK(clk), .RDN(n59411), .Q(
        \pe2/got [12]) );
  DRNQHSV4 \pe2/pe2/q_reg[20]  ( .D(go1[13]), .CK(clk), .RDN(n59458), .Q(
        \pe2/got [13]) );
  DRNQHSV4 \pe2/pe2/q_reg[19]  ( .D(go1[14]), .CK(clk), .RDN(n59659), .Q(
        \pe2/got [14]) );
  DRNQHSV4 \pe2/pe2/q_reg[18]  ( .D(go1[15]), .CK(clk), .RDN(n59434), .Q(
        \pe2/got [15]) );
  DRNQHSV4 \pe2/pe2/q_reg[17]  ( .D(go1[16]), .CK(clk), .RDN(n59397), .Q(
        \pe2/got [16]) );
  DRNQHSV4 \pe2/pe2/q_reg[16]  ( .D(go1[17]), .CK(clk), .RDN(n59457), .Q(
        \pe2/got [17]) );
  DRNQHSV4 \pe2/pe2/q_reg[15]  ( .D(go1[18]), .CK(clk), .RDN(n59444), .Q(
        \pe2/got [18]) );
  DRNQHSV4 \pe2/pe2/q_reg[14]  ( .D(go1[19]), .CK(clk), .RDN(n59922), .Q(
        \pe2/got [19]) );
  DRNQHSV4 \pe2/pe2/q_reg[13]  ( .D(go1[20]), .CK(clk), .RDN(n59437), .Q(
        \pe2/got [20]) );
  DRNQHSV4 \pe2/pe2/q_reg[12]  ( .D(go1[21]), .CK(clk), .RDN(n59458), .Q(
        \pe2/got [21]) );
  DRNQHSV4 \pe2/pe2/q_reg[11]  ( .D(go1[22]), .CK(clk), .RDN(n59445), .Q(
        \pe2/got [22]) );
  DRNQHSV4 \pe2/pe2/q_reg[10]  ( .D(go1[23]), .CK(clk), .RDN(n59430), .Q(
        \pe2/got [23]) );
  DRNQHSV4 \pe2/pe2/q_reg[9]  ( .D(go1[24]), .CK(clk), .RDN(n59454), .Q(
        \pe2/got [24]) );
  DRNQHSV4 \pe2/pe2/q_reg[8]  ( .D(go1[25]), .CK(clk), .RDN(n59405), .Q(
        \pe2/got [25]) );
  DRNQHSV4 \pe2/pe2/q_reg[7]  ( .D(go1[26]), .CK(clk), .RDN(n59403), .Q(
        \pe2/got [26]) );
  DRNQHSV4 \pe2/pe2/q_reg[6]  ( .D(go1[27]), .CK(clk), .RDN(n59472), .Q(
        \pe2/got [27]) );
  DRNQHSV4 \pe2/pe2/q_reg[5]  ( .D(go1[28]), .CK(clk), .RDN(n59653), .Q(
        \pe2/got [28]) );
  DRNQHSV4 \pe2/pe2/q_reg[4]  ( .D(go1[29]), .CK(clk), .RDN(n59435), .Q(
        \pe2/got [29]) );
  DRNQHSV4 \pe2/pe2/q_reg[3]  ( .D(go1[30]), .CK(clk), .RDN(n59923), .Q(
        \pe2/got [30]) );
  DRNQHSV4 \pe2/pe2/q_reg[2]  ( .D(go1[31]), .CK(clk), .RDN(n59925), .Q(
        \pe2/got [31]) );
  DRNQHSV4 \pe2/pe2/q_reg[1]  ( .D(go1[32]), .CK(clk), .RDN(n59449), .Q(
        \pe2/got [32]) );
  DRNQHSV4 \pe2/pe5/q_reg[21]  ( .D(pov1[21]), .CK(clk), .RDN(n59651), .Q(
        \pe2/pvq [21]) );
  DRNQHSV4 \pe2/pe5/q_reg[15]  ( .D(n60039), .CK(clk), .RDN(n59510), .Q(
        \pe2/pvq [15]) );
  DRNQHSV4 \pe2/pe5/q_reg[14]  ( .D(pov1[14]), .CK(clk), .RDN(n59408), .Q(
        \pe2/pvq [14]) );
  DRNQHSV4 \pe2/pe5/q_reg[12]  ( .D(pov1[12]), .CK(clk), .RDN(n59400), .Q(
        \pe2/pvq [12]) );
  DRNQHSV4 \pe2/pe5/q_reg[11]  ( .D(pov1[11]), .CK(clk), .RDN(n59463), .Q(
        \pe2/pvq [11]) );
  DRNQHSV4 \pe2/pe5/q_reg[9]  ( .D(n60017), .CK(clk), .RDN(n59449), .Q(
        \pe2/pvq [9]) );
  DRNQHSV4 \pe2/pe5/q_reg[7]  ( .D(n60065), .CK(clk), .RDN(n59925), .Q(
        \pe2/pvq [7]) );
  DRNQHSV4 \pe2/pe5/q_reg[6]  ( .D(pov1[6]), .CK(clk), .RDN(n29733), .Q(
        \pe2/pvq [6]) );
  DRNQHSV4 \pe2/pe5/q_reg[2]  ( .D(n60109), .CK(clk), .RDN(n59440), .Q(
        \pe2/pvq [2]) );
  DRNQHSV4 \pe2/pe6/q_reg[30]  ( .D(poh1[30]), .CK(clk), .RDN(n29731), .Q(
        \pe2/phq [30]) );
  DRNQHSV4 \pe2/pe6/q_reg[29]  ( .D(poh1[29]), .CK(clk), .RDN(n59397), .Q(
        \pe2/phq [29]) );
  DRNQHSV4 \pe2/pe6/q_reg[28]  ( .D(poh1[28]), .CK(clk), .RDN(n59466), .Q(
        \pe2/phq [28]) );
  DRNQHSV4 \pe2/pe6/q_reg[27]  ( .D(poh1[27]), .CK(clk), .RDN(n59510), .Q(
        \pe2/phq [27]) );
  DRNQHSV4 \pe2/pe6/q_reg[26]  ( .D(poh1[26]), .CK(clk), .RDN(n59650), .Q(
        \pe2/phq [26]) );
  DRNQHSV4 \pe2/pe6/q_reg[25]  ( .D(poh1[25]), .CK(clk), .RDN(n59650), .Q(
        \pe2/phq [25]) );
  DRNQHSV4 \pe2/pe6/q_reg[24]  ( .D(poh1[24]), .CK(clk), .RDN(n59432), .Q(
        \pe2/phq [24]) );
  DRNQHSV4 \pe2/pe6/q_reg[23]  ( .D(poh1[23]), .CK(clk), .RDN(n59402), .Q(
        \pe2/phq [23]) );
  DRNQHSV4 \pe2/pe6/q_reg[22]  ( .D(poh1[22]), .CK(clk), .RDN(n59658), .Q(
        \pe2/phq [22]) );
  DRNQHSV4 \pe2/pe6/q_reg[21]  ( .D(poh1[21]), .CK(clk), .RDN(n59448), .Q(
        \pe2/phq [21]) );
  DRNQHSV4 \pe2/pe6/q_reg[20]  ( .D(poh1[20]), .CK(clk), .RDN(n59404), .Q(
        \pe2/phq [20]) );
  DRNQHSV4 \pe2/pe6/q_reg[19]  ( .D(poh1[19]), .CK(clk), .RDN(n59439), .Q(
        \pe2/phq [19]) );
  DRNQHSV4 \pe2/pe6/q_reg[18]  ( .D(poh1[18]), .CK(clk), .RDN(n29732), .Q(
        \pe2/phq [18]) );
  DRNQHSV4 \pe2/pe6/q_reg[17]  ( .D(poh1[17]), .CK(clk), .RDN(n59459), .Q(
        \pe2/phq [17]) );
  DRNQHSV4 \pe2/pe6/q_reg[16]  ( .D(poh1[16]), .CK(clk), .RDN(n59484), .Q(
        \pe2/phq [16]) );
  DRNQHSV4 \pe2/pe6/q_reg[15]  ( .D(poh1[15]), .CK(clk), .RDN(n59479), .Q(
        \pe2/phq [15]) );
  DRNQHSV4 \pe2/pe6/q_reg[14]  ( .D(poh1[14]), .CK(clk), .RDN(n59923), .Q(
        \pe2/phq [14]) );
  DRNQHSV4 \pe2/pe6/q_reg[13]  ( .D(poh1[13]), .CK(clk), .RDN(n59453), .Q(
        \pe2/phq [13]) );
  DRNQHSV4 \pe2/pe6/q_reg[12]  ( .D(poh1[12]), .CK(clk), .RDN(n59512), .Q(
        \pe2/phq [12]) );
  DRNQHSV4 \pe2/pe6/q_reg[11]  ( .D(poh1[11]), .CK(clk), .RDN(n59510), .Q(
        \pe2/phq [11]) );
  DRNQHSV4 \pe2/pe6/q_reg[10]  ( .D(poh1[10]), .CK(clk), .RDN(n59649), .Q(
        \pe2/phq [10]) );
  DRNQHSV4 \pe2/pe6/q_reg[9]  ( .D(poh1[9]), .CK(clk), .RDN(n59502), .Q(
        \pe2/phq [9]) );
  DRNQHSV4 \pe2/pe6/q_reg[8]  ( .D(poh1[8]), .CK(clk), .RDN(n59419), .Q(
        \pe2/phq [8]) );
  DRNQHSV4 \pe2/pe6/q_reg[7]  ( .D(poh1[7]), .CK(clk), .RDN(n59424), .Q(
        \pe2/phq [7]) );
  DRNQHSV4 \pe2/pe6/q_reg[6]  ( .D(poh1[6]), .CK(clk), .RDN(n59454), .Q(
        \pe2/phq [6]) );
  DRNQHSV4 \pe2/pe6/q_reg[5]  ( .D(poh1[5]), .CK(clk), .RDN(n59407), .Q(
        \pe2/phq [5]) );
  DRNQHSV4 \pe2/pe6/q_reg[4]  ( .D(poh1[4]), .CK(clk), .RDN(n59431), .Q(
        \pe2/phq [4]) );
  DRNQHSV4 \pe2/pe6/q_reg[3]  ( .D(poh1[3]), .CK(clk), .RDN(n59656), .Q(
        \pe2/phq [3]) );
  DRNQHSV4 \pe2/pe6/q_reg[2]  ( .D(poh1[2]), .CK(clk), .RDN(n59657), .Q(
        \pe2/phq [2]) );
  DRNQHSV4 \pe2/pe6/q_reg[1]  ( .D(poh1[1]), .CK(clk), .RDN(n59456), .Q(
        \pe2/phq [1]) );
  DRNQHSV4 \pe2/pe7/q_reg  ( .D(n59999), .CK(clk), .RDN(n59923), .Q(\pe2/ctrq ) );
  DRNQHSV4 \pe2/pe8/q_reg  ( .D(n59497), .CK(clk), .RDN(n59652), .Q(ctro2) );
  DRNQHSV4 \pe2/pe12/q_reg[31]  ( .D(n59567), .CK(clk), .RDN(n59479), .Q(
        \pe2/bq[2] ) );
  DRNQHSV4 \pe2/pe12/q_reg[30]  ( .D(n59754), .CK(clk), .RDN(n29730), .Q(
        \pe2/bq[3] ) );
  DRNQHSV4 \pe2/pe12/q_reg[29]  ( .D(n59752), .CK(clk), .RDN(n59491), .Q(
        \pe2/bq[4] ) );
  DRNQHSV4 \pe2/pe12/q_reg[28]  ( .D(n59566), .CK(clk), .RDN(n59433), .Q(
        \pe2/bq[5] ) );
  DRNQHSV4 \pe2/pe12/q_reg[27]  ( .D(n59749), .CK(clk), .RDN(n59449), .Q(
        \pe2/bq[6] ) );
  DRNQHSV4 \pe2/pe12/q_reg[26]  ( .D(n59746), .CK(clk), .RDN(n59415), .Q(
        \pe2/bq[7] ) );
  DRNQHSV4 \pe2/pe12/q_reg[25]  ( .D(n59565), .CK(clk), .RDN(n59488), .Q(
        \pe2/bq[8] ) );
  DRNQHSV4 \pe2/pe12/q_reg[24]  ( .D(n59748), .CK(clk), .RDN(n59651), .Q(
        \pe2/bq[9] ) );
  DRNQHSV4 \pe2/pe12/q_reg[23]  ( .D(n59747), .CK(clk), .RDN(n59478), .Q(
        \pe2/bq[10] ) );
  DRNQHSV4 \pe2/pe12/q_reg[22]  ( .D(n59745), .CK(clk), .RDN(n29733), .Q(
        \pe2/bq[11] ) );
  DRNQHSV4 \pe2/pe12/q_reg[21]  ( .D(n59564), .CK(clk), .RDN(n59402), .Q(
        \pe2/bq[12] ) );
  DRNQHSV4 \pe2/pe12/q_reg[20]  ( .D(n59744), .CK(clk), .RDN(n59411), .Q(
        \pe2/bq[13] ) );
  DRNQHSV4 \pe2/pe12/q_reg[19]  ( .D(n59742), .CK(clk), .RDN(n59425), .Q(
        \pe2/bq[14] ) );
  DRNQHSV4 \pe2/pe12/q_reg[18]  ( .D(n59743), .CK(clk), .RDN(n59464), .Q(
        \pe2/bq[15] ) );
  DRNQHSV4 \pe2/pe12/q_reg[17]  ( .D(n59741), .CK(clk), .RDN(n59399), .Q(
        \pe2/bq[16] ) );
  DRNQHSV4 \pe2/pe12/q_reg[16]  ( .D(n59740), .CK(clk), .RDN(n59468), .Q(
        \pe2/bq[17] ) );
  DRNQHSV4 \pe2/pe12/q_reg[15]  ( .D(n59739), .CK(clk), .RDN(n59402), .Q(
        \pe2/bq[18] ) );
  DRNQHSV4 \pe2/pe12/q_reg[14]  ( .D(n59563), .CK(clk), .RDN(n59399), .Q(
        \pe2/bq[19] ) );
  DRNQHSV4 \pe2/pe12/q_reg[13]  ( .D(n59738), .CK(clk), .RDN(n59457), .Q(
        \pe2/bq[20] ) );
  DRNQHSV4 \pe2/pe12/q_reg[12]  ( .D(n59735), .CK(clk), .RDN(n59480), .Q(
        \pe2/bq[21] ) );
  DRNQHSV4 \pe2/pe12/q_reg[11]  ( .D(n59734), .CK(clk), .RDN(n59455), .Q(
        \pe2/bq[22] ) );
  DRNQHSV4 \pe2/pe12/q_reg[10]  ( .D(n59562), .CK(clk), .RDN(n59460), .Q(
        \pe2/bq[23] ) );
  DRNQHSV4 \pe2/pe12/q_reg[9]  ( .D(n59731), .CK(clk), .RDN(n59484), .Q(
        \pe2/bq[24] ) );
  DRNQHSV4 \pe2/pe12/q_reg[8]  ( .D(n59729), .CK(clk), .RDN(n29733), .Q(
        \pe2/bq[25] ) );
  DRNQHSV4 \pe2/pe12/q_reg[7]  ( .D(n59728), .CK(clk), .RDN(n59458), .Q(
        \pe2/bq[26] ) );
  DRNQHSV4 \pe2/pe12/q_reg[6]  ( .D(n59727), .CK(clk), .RDN(n59656), .Q(
        \pe2/bq[27] ) );
  DRNQHSV4 \pe2/pe12/q_reg[5]  ( .D(n59726), .CK(clk), .RDN(n59412), .Q(
        \pe2/bq[28] ) );
  DRNQHSV4 \pe2/pe12/q_reg[4]  ( .D(n59723), .CK(clk), .RDN(n59921), .Q(
        \pe2/bq[29] ) );
  DRNQHSV4 \pe2/pe12/q_reg[3]  ( .D(n59724), .CK(clk), .RDN(n59399), .Q(
        \pe2/bq[30] ) );
  DRNQHSV4 \pe2/pe12/q_reg[2]  ( .D(n59722), .CK(clk), .RDN(n59466), .Q(
        \pe2/bq[31] ) );
  DRNQHSV4 \pe2/pe12/q_reg[1]  ( .D(n59721), .CK(clk), .RDN(n59412), .Q(
        \pe2/bq[32] ) );
  DRNQHSV4 \pe2/pe13/q_reg  ( .D(\pe2/ti_1t ), .CK(clk), .RDN(n59440), .Q(
        \pe2/ti_1 ) );
  DRNQHSV4 \pe2/pe14/q_reg[3]  ( .D(n59684), .CK(clk), .RDN(n59440), .Q(
        \pe2/ti_7t [3]) );
  DRNQHSV4 \pe2/pe14/q_reg[5]  ( .D(n59679), .CK(clk), .RDN(n29731), .Q(
        \pe2/ti_7t [5]) );
  DRNQHSV4 \pe2/pe14/q_reg[7]  ( .D(n45149), .CK(clk), .RDN(n59493), .Q(
        \pe2/ti_7t [7]) );
  DRNQHSV4 \pe3/pe1/q_reg[32]  ( .D(ao2[1]), .CK(clk), .RDN(n29729), .Q(
        \pe3/aot [1]) );
  DRNQHSV4 \pe3/pe1/q_reg[31]  ( .D(ao2[2]), .CK(clk), .RDN(n59468), .Q(
        \pe3/aot [2]) );
  DRNQHSV4 \pe3/pe1/q_reg[30]  ( .D(ao2[3]), .CK(clk), .RDN(n59465), .Q(
        \pe3/aot [3]) );
  DRNQHSV4 \pe3/pe1/q_reg[29]  ( .D(ao2[4]), .CK(clk), .RDN(n59471), .Q(
        \pe3/aot [4]) );
  DRNQHSV4 \pe3/pe1/q_reg[28]  ( .D(ao2[5]), .CK(clk), .RDN(n59443), .Q(
        \pe3/aot [5]) );
  DRNQHSV4 \pe3/pe1/q_reg[27]  ( .D(ao2[6]), .CK(clk), .RDN(n59450), .Q(
        \pe3/aot [6]) );
  DRNQHSV4 \pe3/pe1/q_reg[26]  ( .D(ao2[7]), .CK(clk), .RDN(n29730), .Q(
        \pe3/aot [7]) );
  DRNQHSV4 \pe3/pe1/q_reg[25]  ( .D(ao2[8]), .CK(clk), .RDN(n59408), .Q(
        \pe3/aot [8]) );
  DRNQHSV4 \pe3/pe1/q_reg[24]  ( .D(ao2[9]), .CK(clk), .RDN(n59419), .Q(
        \pe3/aot [9]) );
  DRNQHSV4 \pe3/pe1/q_reg[23]  ( .D(ao2[10]), .CK(clk), .RDN(n59452), .Q(
        \pe3/aot [10]) );
  DRNQHSV4 \pe3/pe1/q_reg[22]  ( .D(ao2[11]), .CK(clk), .RDN(n59444), .Q(
        \pe3/aot [11]) );
  DRNQHSV4 \pe3/pe1/q_reg[21]  ( .D(ao2[12]), .CK(clk), .RDN(n59419), .Q(
        \pe3/aot [12]) );
  DRNQHSV4 \pe3/pe1/q_reg[20]  ( .D(ao2[13]), .CK(clk), .RDN(n59503), .Q(
        \pe3/aot [13]) );
  DRNQHSV4 \pe3/pe1/q_reg[19]  ( .D(ao2[14]), .CK(clk), .RDN(n59434), .Q(
        \pe3/aot [14]) );
  DRNQHSV4 \pe3/pe1/q_reg[18]  ( .D(ao2[15]), .CK(clk), .RDN(n59430), .Q(
        \pe3/aot [15]) );
  DRNQHSV4 \pe3/pe1/q_reg[17]  ( .D(ao2[16]), .CK(clk), .RDN(n59396), .Q(
        \pe3/aot [16]) );
  DRNQHSV4 \pe3/pe1/q_reg[16]  ( .D(ao2[17]), .CK(clk), .RDN(n59502), .Q(
        \pe3/aot [17]) );
  DRNQHSV4 \pe3/pe1/q_reg[15]  ( .D(ao2[18]), .CK(clk), .RDN(n59442), .Q(
        \pe3/aot [18]) );
  DRNQHSV4 \pe3/pe1/q_reg[14]  ( .D(ao2[19]), .CK(clk), .RDN(n59652), .Q(
        \pe3/aot [19]) );
  DRNQHSV4 \pe3/pe1/q_reg[13]  ( .D(ao2[20]), .CK(clk), .RDN(n59651), .Q(
        \pe3/aot [20]) );
  DRNQHSV4 \pe3/pe1/q_reg[12]  ( .D(ao2[21]), .CK(clk), .RDN(n59417), .Q(
        \pe3/aot [21]) );
  DRNQHSV4 \pe3/pe1/q_reg[11]  ( .D(ao2[22]), .CK(clk), .RDN(n59437), .Q(
        \pe3/aot [22]) );
  DRNQHSV4 \pe3/pe1/q_reg[10]  ( .D(ao2[23]), .CK(clk), .RDN(n29731), .Q(
        \pe3/aot [23]) );
  DRNQHSV4 \pe3/pe1/q_reg[9]  ( .D(ao2[24]), .CK(clk), .RDN(n59658), .Q(
        \pe3/aot [24]) );
  DRNQHSV4 \pe3/pe1/q_reg[8]  ( .D(ao2[25]), .CK(clk), .RDN(n59922), .Q(
        \pe3/aot [25]) );
  DRNQHSV4 \pe3/pe1/q_reg[7]  ( .D(ao2[26]), .CK(clk), .RDN(n59446), .Q(
        \pe3/aot [26]) );
  DRNQHSV4 \pe3/pe1/q_reg[6]  ( .D(ao2[27]), .CK(clk), .RDN(n59402), .Q(
        \pe3/aot [27]) );
  DRNQHSV4 \pe3/pe1/q_reg[5]  ( .D(ao2[28]), .CK(clk), .RDN(n59446), .Q(
        \pe3/aot [28]) );
  DRNQHSV4 \pe3/pe1/q_reg[4]  ( .D(ao2[29]), .CK(clk), .RDN(n59512), .Q(
        \pe3/aot [29]) );
  DRNQHSV4 \pe3/pe1/q_reg[3]  ( .D(ao2[30]), .CK(clk), .RDN(n59652), .Q(
        \pe3/aot [30]) );
  DRNQHSV4 \pe3/pe1/q_reg[2]  ( .D(ao2[31]), .CK(clk), .RDN(n59416), .Q(
        \pe3/aot [31]) );
  DRNQHSV4 \pe3/pe2/q_reg[32]  ( .D(go2[1]), .CK(clk), .RDN(n59652), .Q(
        \pe3/got [1]) );
  DRNQHSV4 \pe3/pe2/q_reg[31]  ( .D(go2[2]), .CK(clk), .RDN(n59418), .Q(
        \pe3/got [2]) );
  DRNQHSV4 \pe3/pe2/q_reg[30]  ( .D(go2[3]), .CK(clk), .RDN(n59461), .Q(
        \pe3/got [3]) );
  DRNQHSV4 \pe3/pe2/q_reg[29]  ( .D(go2[4]), .CK(clk), .RDN(n59925), .Q(
        \pe3/got [4]) );
  DRNQHSV4 \pe3/pe2/q_reg[28]  ( .D(go2[5]), .CK(clk), .RDN(n59503), .Q(
        \pe3/got [5]) );
  DRNQHSV4 \pe3/pe2/q_reg[27]  ( .D(go2[6]), .CK(clk), .RDN(n59450), .Q(
        \pe3/got [6]) );
  DRNQHSV4 \pe3/pe2/q_reg[26]  ( .D(go2[7]), .CK(clk), .RDN(n59652), .Q(
        \pe3/got [7]) );
  DRNQHSV4 \pe3/pe2/q_reg[25]  ( .D(go2[8]), .CK(clk), .RDN(n59652), .Q(
        \pe3/got [8]) );
  DRNQHSV4 \pe3/pe2/q_reg[24]  ( .D(go2[9]), .CK(clk), .RDN(n59425), .Q(
        \pe3/got [9]) );
  DRNQHSV4 \pe3/pe2/q_reg[23]  ( .D(go2[10]), .CK(clk), .RDN(n59488), .Q(
        \pe3/got [10]) );
  DRNQHSV4 \pe3/pe2/q_reg[22]  ( .D(go2[11]), .CK(clk), .RDN(n59425), .Q(
        \pe3/got [11]) );
  DRNQHSV4 \pe3/pe2/q_reg[21]  ( .D(go2[12]), .CK(clk), .RDN(n59443), .Q(
        \pe3/got [12]) );
  DRNQHSV4 \pe3/pe2/q_reg[20]  ( .D(go2[13]), .CK(clk), .RDN(n59658), .Q(
        \pe3/got [13]) );
  DRNQHSV4 \pe3/pe2/q_reg[19]  ( .D(go2[14]), .CK(clk), .RDN(n59482), .Q(
        \pe3/got [14]) );
  DRNQHSV4 \pe3/pe2/q_reg[18]  ( .D(go2[15]), .CK(clk), .RDN(n29731), .Q(
        \pe3/got [15]) );
  DRNQHSV4 \pe3/pe2/q_reg[17]  ( .D(go2[16]), .CK(clk), .RDN(n59490), .Q(
        \pe3/got [16]) );
  DRNQHSV4 \pe3/pe2/q_reg[16]  ( .D(go2[17]), .CK(clk), .RDN(n59488), .Q(
        \pe3/got [17]) );
  DRNQHSV4 \pe3/pe2/q_reg[15]  ( .D(go2[18]), .CK(clk), .RDN(n59461), .Q(
        \pe3/got [18]) );
  DRNQHSV4 \pe3/pe2/q_reg[14]  ( .D(go2[19]), .CK(clk), .RDN(n59431), .Q(
        \pe3/got [19]) );
  DRNQHSV4 \pe3/pe2/q_reg[13]  ( .D(go2[20]), .CK(clk), .RDN(n59462), .Q(
        \pe3/got [20]) );
  DRNQHSV4 \pe3/pe2/q_reg[12]  ( .D(go2[21]), .CK(clk), .RDN(n59474), .Q(
        \pe3/got [21]) );
  DRNQHSV4 \pe3/pe2/q_reg[11]  ( .D(go2[22]), .CK(clk), .RDN(n59431), .Q(
        \pe3/got [22]) );
  DRNQHSV4 \pe3/pe2/q_reg[10]  ( .D(go2[23]), .CK(clk), .RDN(n59433), .Q(
        \pe3/got [23]) );
  DRNQHSV4 \pe3/pe2/q_reg[9]  ( .D(go2[24]), .CK(clk), .RDN(n59455), .Q(
        \pe3/got [24]) );
  DRNQHSV4 \pe3/pe2/q_reg[8]  ( .D(go2[25]), .CK(clk), .RDN(n59446), .Q(
        \pe3/got [25]) );
  DRNQHSV4 \pe3/pe2/q_reg[7]  ( .D(go2[26]), .CK(clk), .RDN(n59472), .Q(
        \pe3/got [26]) );
  DRNQHSV4 \pe3/pe2/q_reg[6]  ( .D(go2[27]), .CK(clk), .RDN(n59416), .Q(
        \pe3/got [27]) );
  DRNQHSV4 \pe3/pe2/q_reg[5]  ( .D(go2[28]), .CK(clk), .RDN(n59402), .Q(
        \pe3/got [28]) );
  DRNQHSV4 \pe3/pe2/q_reg[4]  ( .D(go2[29]), .CK(clk), .RDN(n59450), .Q(
        \pe3/got [29]) );
  DRNQHSV4 \pe3/pe2/q_reg[3]  ( .D(go2[30]), .CK(clk), .RDN(n59922), .Q(
        \pe3/got [30]) );
  DRNQHSV4 \pe3/pe5/q_reg[24]  ( .D(n60093), .CK(clk), .RDN(n59478), .Q(
        \pe3/pvq [24]) );
  DRNQHSV4 \pe3/pe5/q_reg[23]  ( .D(n60094), .CK(clk), .RDN(n59444), .Q(
        \pe3/pvq [23]) );
  DRNQHSV4 \pe3/pe5/q_reg[21]  ( .D(n60062), .CK(clk), .RDN(n59417), .Q(
        \pe3/pvq [21]) );
  DRNQHSV4 \pe3/pe5/q_reg[19]  ( .D(n60047), .CK(clk), .RDN(n59447), .Q(
        \pe3/pvq [19]) );
  DRNQHSV4 \pe3/pe5/q_reg[18]  ( .D(n60052), .CK(clk), .RDN(n59412), .Q(
        \pe3/pvq [18]) );
  DRNQHSV4 \pe3/pe5/q_reg[17]  ( .D(pov2[17]), .CK(clk), .RDN(n59444), .Q(
        \pe3/pvq [17]) );
  DRNQHSV4 \pe3/pe5/q_reg[16]  ( .D(n60050), .CK(clk), .RDN(n59453), .Q(
        \pe3/pvq [16]) );
  DRNQHSV4 \pe3/pe5/q_reg[15]  ( .D(pov2[15]), .CK(clk), .RDN(n59457), .Q(
        \pe3/pvq [15]) );
  DRNQHSV4 \pe3/pe5/q_reg[13]  ( .D(n60096), .CK(clk), .RDN(n59444), .Q(
        \pe3/pvq [13]) );
  DRNQHSV4 \pe3/pe5/q_reg[12]  ( .D(n60043), .CK(clk), .RDN(n59925), .Q(
        \pe3/pvq [12]) );
  DRNQHSV4 \pe3/pe5/q_reg[11]  ( .D(n60097), .CK(clk), .RDN(n59445), .Q(
        \pe3/pvq [11]) );
  DRNQHSV4 \pe3/pe5/q_reg[9]  ( .D(n60098), .CK(clk), .RDN(n59411), .Q(
        \pe3/pvq [9]) );
  DRNQHSV4 \pe3/pe5/q_reg[8]  ( .D(n60099), .CK(clk), .RDN(n59445), .Q(
        \pe3/pvq [8]) );
  DRNQHSV4 \pe3/pe5/q_reg[5]  ( .D(n60100), .CK(clk), .RDN(n59402), .Q(
        \pe3/pvq [5]) );
  DRNQHSV4 \pe3/pe5/q_reg[3]  ( .D(n60101), .CK(clk), .RDN(n59408), .Q(
        \pe3/pvq [3]) );
  DRNQHSV4 \pe3/pe6/q_reg[31]  ( .D(poh2[31]), .CK(clk), .RDN(n59492), .Q(
        \pe3/phq [31]) );
  DRNQHSV4 \pe3/pe6/q_reg[30]  ( .D(poh2[30]), .CK(clk), .RDN(n59496), .Q(
        \pe3/phq [30]) );
  DRNQHSV4 \pe3/pe6/q_reg[29]  ( .D(poh2[29]), .CK(clk), .RDN(n59438), .Q(
        \pe3/phq [29]) );
  DRNQHSV4 \pe3/pe6/q_reg[28]  ( .D(poh2[28]), .CK(clk), .RDN(n59653), .Q(
        \pe3/phq [28]) );
  DRNQHSV4 \pe3/pe6/q_reg[27]  ( .D(poh2[27]), .CK(clk), .RDN(n59483), .Q(
        \pe3/phq [27]) );
  DRNQHSV4 \pe3/pe6/q_reg[26]  ( .D(poh2[26]), .CK(clk), .RDN(n59473), .Q(
        \pe3/phq [26]) );
  DRNQHSV4 \pe3/pe6/q_reg[25]  ( .D(poh2[25]), .CK(clk), .RDN(n29730), .Q(
        \pe3/phq [25]) );
  DRNQHSV4 \pe3/pe6/q_reg[24]  ( .D(poh2[24]), .CK(clk), .RDN(n59412), .Q(
        \pe3/phq [24]) );
  DRNQHSV4 \pe3/pe6/q_reg[23]  ( .D(poh2[23]), .CK(clk), .RDN(n59464), .Q(
        \pe3/phq [23]) );
  DRNQHSV4 \pe3/pe6/q_reg[22]  ( .D(poh2[22]), .CK(clk), .RDN(n59437), .Q(
        \pe3/phq [22]) );
  DRNQHSV4 \pe3/pe6/q_reg[21]  ( .D(poh2[21]), .CK(clk), .RDN(n59470), .Q(
        \pe3/phq [21]) );
  DRNQHSV4 \pe3/pe6/q_reg[20]  ( .D(poh2[20]), .CK(clk), .RDN(n59418), .Q(
        \pe3/phq [20]) );
  DRNQHSV4 \pe3/pe6/q_reg[19]  ( .D(poh2[19]), .CK(clk), .RDN(n59432), .Q(
        \pe3/phq [19]) );
  DRNQHSV4 \pe3/pe6/q_reg[18]  ( .D(poh2[18]), .CK(clk), .RDN(n59456), .Q(
        \pe3/phq [18]) );
  DRNQHSV4 \pe3/pe6/q_reg[17]  ( .D(poh2[17]), .CK(clk), .RDN(n59477), .Q(
        \pe3/phq [17]) );
  DRNQHSV4 \pe3/pe6/q_reg[16]  ( .D(poh2[16]), .CK(clk), .RDN(n59416), .Q(
        \pe3/phq [16]) );
  DRNQHSV4 \pe3/pe6/q_reg[15]  ( .D(poh2[15]), .CK(clk), .RDN(n59440), .Q(
        \pe3/phq [15]) );
  DRNQHSV4 \pe3/pe6/q_reg[14]  ( .D(poh2[14]), .CK(clk), .RDN(n59424), .Q(
        \pe3/phq [14]) );
  DRNQHSV4 \pe3/pe6/q_reg[13]  ( .D(poh2[13]), .CK(clk), .RDN(n59923), .Q(
        \pe3/phq [13]) );
  DRNQHSV4 \pe3/pe6/q_reg[12]  ( .D(poh2[12]), .CK(clk), .RDN(n59417), .Q(
        \pe3/phq [12]) );
  DRNQHSV4 \pe3/pe6/q_reg[11]  ( .D(poh2[11]), .CK(clk), .RDN(n59462), .Q(
        \pe3/phq [11]) );
  DRNQHSV4 \pe3/pe6/q_reg[10]  ( .D(poh2[10]), .CK(clk), .RDN(n59450), .Q(
        \pe3/phq [10]) );
  DRNQHSV4 \pe3/pe6/q_reg[9]  ( .D(poh2[9]), .CK(clk), .RDN(n59425), .Q(
        \pe3/phq [9]) );
  DRNQHSV4 \pe3/pe6/q_reg[8]  ( .D(poh2[8]), .CK(clk), .RDN(n59503), .Q(
        \pe3/phq [8]) );
  DRNQHSV4 \pe3/pe6/q_reg[7]  ( .D(poh2[7]), .CK(clk), .RDN(n59407), .Q(
        \pe3/phq [7]) );
  DRNQHSV4 \pe3/pe6/q_reg[6]  ( .D(poh2[6]), .CK(clk), .RDN(n59478), .Q(
        \pe3/phq [6]) );
  DRNQHSV4 \pe3/pe6/q_reg[5]  ( .D(poh2[5]), .CK(clk), .RDN(n59510), .Q(
        \pe3/phq [5]) );
  DRNQHSV4 \pe3/pe6/q_reg[4]  ( .D(poh2[4]), .CK(clk), .RDN(n59922), .Q(
        \pe3/phq [4]) );
  DRNQHSV4 \pe3/pe6/q_reg[3]  ( .D(poh2[3]), .CK(clk), .RDN(n59493), .Q(
        \pe3/phq [3]) );
  DRNQHSV4 \pe3/pe6/q_reg[2]  ( .D(poh2[2]), .CK(clk), .RDN(n29734), .Q(
        \pe3/phq [2]) );
  DRNQHSV4 \pe3/pe7/q_reg  ( .D(n59586), .CK(clk), .RDN(n59479), .Q(\pe3/ctrq ) );
  DRNQHSV4 \pe3/pe8/q_reg  ( .D(n59537), .CK(clk), .RDN(n59467), .Q(ctro3) );
  DRNQHSV4 \pe3/pe12/q_reg[32]  ( .D(n59796), .CK(clk), .RDN(n29734), .Q(
        \pe3/bq[1] ) );
  DRNQHSV4 \pe3/pe12/q_reg[31]  ( .D(n59795), .CK(clk), .RDN(n59416), .Q(
        \pe3/bq[2] ) );
  DRNQHSV4 \pe3/pe12/q_reg[30]  ( .D(\pe3/bqt[3] ), .CK(clk), .RDN(n59414), 
        .Q(\pe3/bq[3] ) );
  DRNQHSV4 \pe3/pe12/q_reg[29]  ( .D(n59561), .CK(clk), .RDN(n59480), .Q(
        \pe3/bq[4] ) );
  DRNQHSV4 \pe3/pe12/q_reg[28]  ( .D(n59793), .CK(clk), .RDN(n59480), .Q(
        \pe3/bq[5] ) );
  DRNQHSV4 \pe3/pe12/q_reg[27]  ( .D(n59791), .CK(clk), .RDN(n59479), .Q(
        \pe3/bq[6] ) );
  DRNQHSV4 \pe3/pe12/q_reg[26]  ( .D(n59560), .CK(clk), .RDN(n59405), .Q(
        \pe3/bq[7] ) );
  DRNQHSV4 \pe3/pe12/q_reg[25]  ( .D(n59785), .CK(clk), .RDN(n59654), .Q(
        \pe3/bq[8] ) );
  DRNQHSV4 \pe3/pe12/q_reg[24]  ( .D(n59786), .CK(clk), .RDN(n59478), .Q(
        \pe3/bq[9] ) );
  DRNQHSV4 \pe3/pe12/q_reg[23]  ( .D(n59784), .CK(clk), .RDN(n59477), .Q(
        \pe3/bq[10] ) );
  DRNQHSV4 \pe3/pe12/q_reg[22]  ( .D(n59781), .CK(clk), .RDN(n59462), .Q(
        \pe3/bq[11] ) );
  DRNQHSV4 \pe3/pe12/q_reg[21]  ( .D(n59782), .CK(clk), .RDN(n59473), .Q(
        \pe3/bq[12] ) );
  DRNQHSV4 \pe3/pe12/q_reg[20]  ( .D(n59788), .CK(clk), .RDN(n59447), .Q(
        \pe3/bq[13] ) );
  DRNQHSV4 \pe3/pe12/q_reg[19]  ( .D(n59787), .CK(clk), .RDN(n59415), .Q(
        \pe3/bq[14] ) );
  DRNQHSV4 \pe3/pe12/q_reg[18]  ( .D(n59779), .CK(clk), .RDN(n59407), .Q(
        \pe3/bq[15] ) );
  DRNQHSV4 \pe3/pe12/q_reg[17]  ( .D(n59780), .CK(clk), .RDN(n59406), .Q(
        \pe3/bq[16] ) );
  DRNQHSV4 \pe3/pe12/q_reg[16]  ( .D(n59776), .CK(clk), .RDN(n59484), .Q(
        \pe3/bq[17] ) );
  DRNQHSV4 \pe3/pe12/q_reg[15]  ( .D(n59559), .CK(clk), .RDN(n59483), .Q(
        \pe3/bq[18] ) );
  DRNQHSV4 \pe3/pe12/q_reg[14]  ( .D(n59770), .CK(clk), .RDN(n59409), .Q(
        \pe3/bq[19] ) );
  DRNQHSV4 \pe3/pe12/q_reg[13]  ( .D(n59771), .CK(clk), .RDN(n59448), .Q(
        \pe3/bq[20] ) );
  DRNQHSV4 \pe3/pe12/q_reg[12]  ( .D(n59772), .CK(clk), .RDN(n59410), .Q(
        \pe3/bq[21] ) );
  DRNQHSV4 \pe3/pe12/q_reg[11]  ( .D(n59762), .CK(clk), .RDN(n59492), .Q(
        \pe3/bq[22] ) );
  DRNQHSV4 \pe3/pe12/q_reg[10]  ( .D(n59558), .CK(clk), .RDN(n59657), .Q(
        \pe3/bq[23] ) );
  DRNQHSV4 \pe3/pe12/q_reg[9]  ( .D(n59557), .CK(clk), .RDN(n59923), .Q(
        \pe3/bq[24] ) );
  DRNQHSV4 \pe3/pe12/q_reg[8]  ( .D(n59556), .CK(clk), .RDN(n59447), .Q(
        \pe3/bq[25] ) );
  DRNQHSV4 \pe3/pe12/q_reg[7]  ( .D(n59555), .CK(clk), .RDN(n59403), .Q(
        \pe3/bq[26] ) );
  DRNQHSV4 \pe3/pe12/q_reg[6]  ( .D(n59765), .CK(clk), .RDN(n59418), .Q(
        \pe3/bq[27] ) );
  DRNQHSV4 \pe3/pe12/q_reg[5]  ( .D(n59764), .CK(clk), .RDN(n59448), .Q(
        \pe3/bq[28] ) );
  DRNQHSV4 \pe3/pe12/q_reg[4]  ( .D(n59763), .CK(clk), .RDN(n59503), .Q(
        \pe3/bq[29] ) );
  DRNQHSV4 \pe3/pe12/q_reg[3]  ( .D(n59760), .CK(clk), .RDN(n59474), .Q(
        \pe3/bq[30] ) );
  DRNQHSV4 \pe3/pe12/q_reg[2]  ( .D(n59554), .CK(clk), .RDN(n29733), .Q(
        \pe3/bq[31] ) );
  DRNQHSV4 \pe3/pe12/q_reg[1]  ( .D(n59688), .CK(clk), .RDN(n29734), .Q(
        \pe3/bq[32] ) );
  DRNQHSV4 \pe3/pe14/q_reg[1]  ( .D(n59648), .CK(clk), .RDN(n59481), .Q(
        \pe3/ti_7t [1]) );
  DRNQHSV4 \pe3/pe14/q_reg[2]  ( .D(n59797), .CK(clk), .RDN(n59405), .Q(
        \pe3/ti_7t [2]) );
  DRNQHSV4 \pe3/pe14/q_reg[3]  ( .D(n59671), .CK(clk), .RDN(n59480), .Q(
        \pe3/ti_7t [3]) );
  DRNQHSV4 \pe4/pe1/q_reg[32]  ( .D(ao3[1]), .CK(clk), .RDN(n59656), .Q(
        \pe4/aot [1]) );
  DRNQHSV4 \pe4/pe1/q_reg[31]  ( .D(ao3[2]), .CK(clk), .RDN(n59503), .Q(
        \pe4/aot [2]) );
  DRNQHSV4 \pe4/pe1/q_reg[30]  ( .D(ao3[3]), .CK(clk), .RDN(n59466), .Q(
        \pe4/aot [3]) );
  DRNQHSV4 \pe4/pe1/q_reg[29]  ( .D(ao3[4]), .CK(clk), .RDN(n59924), .Q(
        \pe4/aot [4]) );
  DRNQHSV4 \pe4/pe1/q_reg[28]  ( .D(ao3[5]), .CK(clk), .RDN(n59654), .Q(
        \pe4/aot [5]) );
  DRNQHSV4 \pe4/pe1/q_reg[27]  ( .D(ao3[6]), .CK(clk), .RDN(n59490), .Q(
        \pe4/aot [6]) );
  DRNQHSV4 \pe4/pe1/q_reg[26]  ( .D(ao3[7]), .CK(clk), .RDN(n59450), .Q(
        \pe4/aot [7]) );
  DRNQHSV4 \pe4/pe1/q_reg[25]  ( .D(ao3[8]), .CK(clk), .RDN(n29731), .Q(
        \pe4/aot [8]) );
  DRNQHSV4 \pe4/pe1/q_reg[24]  ( .D(ao3[9]), .CK(clk), .RDN(n59481), .Q(
        \pe4/aot [9]) );
  DRNQHSV4 \pe4/pe1/q_reg[23]  ( .D(ao3[10]), .CK(clk), .RDN(n59444), .Q(
        \pe4/aot [10]) );
  DRNQHSV4 \pe4/pe1/q_reg[22]  ( .D(ao3[11]), .CK(clk), .RDN(n59412), .Q(
        \pe4/aot [11]) );
  DRNQHSV4 \pe4/pe1/q_reg[21]  ( .D(ao3[12]), .CK(clk), .RDN(n59510), .Q(
        \pe4/aot [12]) );
  DRNQHSV4 \pe4/pe1/q_reg[20]  ( .D(ao3[13]), .CK(clk), .RDN(n59410), .Q(
        \pe4/aot [13]) );
  DRNQHSV4 \pe4/pe1/q_reg[19]  ( .D(ao3[14]), .CK(clk), .RDN(n59446), .Q(
        \pe4/aot [14]) );
  DRNQHSV4 \pe4/pe1/q_reg[18]  ( .D(ao3[15]), .CK(clk), .RDN(n59414), .Q(
        \pe4/aot [15]) );
  DRNQHSV4 \pe4/pe1/q_reg[17]  ( .D(ao3[16]), .CK(clk), .RDN(n59479), .Q(
        \pe4/aot [16]) );
  DRNQHSV4 \pe4/pe1/q_reg[16]  ( .D(ao3[17]), .CK(clk), .RDN(n59464), .Q(
        \pe4/aot [17]) );
  DRNQHSV4 \pe4/pe1/q_reg[15]  ( .D(ao3[18]), .CK(clk), .RDN(n59461), .Q(
        \pe4/aot [18]) );
  DRNQHSV4 \pe4/pe1/q_reg[14]  ( .D(ao3[19]), .CK(clk), .RDN(n59659), .Q(
        \pe4/aot [19]) );
  DRNQHSV4 \pe4/pe1/q_reg[13]  ( .D(ao3[20]), .CK(clk), .RDN(n59659), .Q(
        \pe4/aot [20]) );
  DRNQHSV4 \pe4/pe1/q_reg[12]  ( .D(ao3[21]), .CK(clk), .RDN(n59658), .Q(
        \pe4/aot [21]) );
  DRNQHSV4 \pe4/pe1/q_reg[11]  ( .D(ao3[22]), .CK(clk), .RDN(n59406), .Q(
        \pe4/aot [22]) );
  DRNQHSV4 \pe4/pe1/q_reg[10]  ( .D(ao3[23]), .CK(clk), .RDN(n59657), .Q(
        \pe4/aot [23]) );
  DRNQHSV4 \pe4/pe1/q_reg[9]  ( .D(ao3[24]), .CK(clk), .RDN(n59478), .Q(
        \pe4/aot [24]) );
  DRNQHSV4 \pe4/pe1/q_reg[8]  ( .D(ao3[25]), .CK(clk), .RDN(n59411), .Q(
        \pe4/aot [25]) );
  DRNQHSV4 \pe4/pe1/q_reg[7]  ( .D(ao3[26]), .CK(clk), .RDN(n59921), .Q(
        \pe4/aot [26]) );
  DRNQHSV4 \pe4/pe1/q_reg[6]  ( .D(ao3[27]), .CK(clk), .RDN(n59925), .Q(
        \pe4/aot [27]) );
  DRNQHSV4 \pe4/pe1/q_reg[5]  ( .D(ao3[28]), .CK(clk), .RDN(n59424), .Q(
        \pe4/aot [28]) );
  DRNQHSV4 \pe4/pe1/q_reg[4]  ( .D(ao3[29]), .CK(clk), .RDN(n59455), .Q(
        \pe4/aot [29]) );
  DRNQHSV4 \pe4/pe1/q_reg[3]  ( .D(ao3[30]), .CK(clk), .RDN(n59446), .Q(
        \pe4/aot [30]) );
  DRNQHSV4 \pe4/pe1/q_reg[2]  ( .D(ao3[31]), .CK(clk), .RDN(n29729), .Q(
        \pe4/aot [31]) );
  DRNQHSV4 \pe4/pe1/q_reg[1]  ( .D(ao3[32]), .CK(clk), .RDN(n59407), .Q(
        \pe4/aot [32]) );
  DRNQHSV4 \pe4/pe2/q_reg[32]  ( .D(go3[1]), .CK(clk), .RDN(n59474), .Q(
        \pe4/got [1]) );
  DRNQHSV4 \pe4/pe2/q_reg[31]  ( .D(go3[2]), .CK(clk), .RDN(n59655), .Q(
        \pe4/got [2]) );
  DRNQHSV4 \pe4/pe2/q_reg[30]  ( .D(go3[3]), .CK(clk), .RDN(n59493), .Q(
        \pe4/got [3]) );
  DRNQHSV4 \pe4/pe2/q_reg[29]  ( .D(go3[4]), .CK(clk), .RDN(n59442), .Q(
        \pe4/got [4]) );
  DRNQHSV4 \pe4/pe2/q_reg[28]  ( .D(go3[5]), .CK(clk), .RDN(n59921), .Q(
        \pe4/got [5]) );
  DRNQHSV4 \pe4/pe2/q_reg[27]  ( .D(go3[6]), .CK(clk), .RDN(n59436), .Q(
        \pe4/got [6]) );
  DRNQHSV4 \pe4/pe2/q_reg[26]  ( .D(go3[7]), .CK(clk), .RDN(n59657), .Q(
        \pe4/got [7]) );
  DRNQHSV4 \pe4/pe2/q_reg[25]  ( .D(go3[8]), .CK(clk), .RDN(n59434), .Q(
        \pe4/got [8]) );
  DRNQHSV4 \pe4/pe2/q_reg[24]  ( .D(go3[9]), .CK(clk), .RDN(n59483), .Q(
        \pe4/got [9]) );
  DRNQHSV4 \pe4/pe2/q_reg[23]  ( .D(go3[10]), .CK(clk), .RDN(n59459), .Q(
        \pe4/got [10]) );
  DRNQHSV4 \pe4/pe2/q_reg[22]  ( .D(go3[11]), .CK(clk), .RDN(n59400), .Q(
        \pe4/got [11]) );
  DRNQHSV4 \pe4/pe2/q_reg[21]  ( .D(go3[12]), .CK(clk), .RDN(n59922), .Q(
        \pe4/got [12]) );
  DRNQHSV4 \pe4/pe2/q_reg[20]  ( .D(go3[13]), .CK(clk), .RDN(n59401), .Q(
        \pe4/got [13]) );
  DRNQHSV4 \pe4/pe2/q_reg[19]  ( .D(go3[14]), .CK(clk), .RDN(n59431), .Q(
        \pe4/got [14]) );
  DRNQHSV4 \pe4/pe2/q_reg[18]  ( .D(go3[15]), .CK(clk), .RDN(n59444), .Q(
        \pe4/got [15]) );
  DRNQHSV4 \pe4/pe2/q_reg[17]  ( .D(go3[16]), .CK(clk), .RDN(n59490), .Q(
        \pe4/got [16]) );
  DRNQHSV4 \pe4/pe2/q_reg[16]  ( .D(go3[17]), .CK(clk), .RDN(n59414), .Q(
        \pe4/got [17]) );
  DRNQHSV4 \pe4/pe2/q_reg[15]  ( .D(go3[18]), .CK(clk), .RDN(n59400), .Q(
        \pe4/got [18]) );
  DRNQHSV4 \pe4/pe2/q_reg[14]  ( .D(go3[19]), .CK(clk), .RDN(n59924), .Q(
        \pe4/got [19]) );
  DRNQHSV4 \pe4/pe2/q_reg[13]  ( .D(go3[20]), .CK(clk), .RDN(n59432), .Q(
        \pe4/got [20]) );
  DRNQHSV4 \pe4/pe2/q_reg[12]  ( .D(go3[21]), .CK(clk), .RDN(n59658), .Q(
        \pe4/got [21]) );
  DRNQHSV4 \pe4/pe2/q_reg[11]  ( .D(go3[22]), .CK(clk), .RDN(n59658), .Q(
        \pe4/got [22]) );
  DRNQHSV4 \pe4/pe2/q_reg[10]  ( .D(go3[23]), .CK(clk), .RDN(n59925), .Q(
        \pe4/got [23]) );
  DRNQHSV4 \pe4/pe2/q_reg[9]  ( .D(go3[24]), .CK(clk), .RDN(n59925), .Q(
        \pe4/got [24]) );
  DRNQHSV4 \pe4/pe2/q_reg[8]  ( .D(go3[25]), .CK(clk), .RDN(n59657), .Q(
        \pe4/got [25]) );
  DRNQHSV4 \pe4/pe2/q_reg[7]  ( .D(go3[26]), .CK(clk), .RDN(n59657), .Q(
        \pe4/got [26]) );
  DRNQHSV4 \pe4/pe2/q_reg[6]  ( .D(go3[27]), .CK(clk), .RDN(n59476), .Q(
        \pe4/got [27]) );
  DRNQHSV4 \pe4/pe2/q_reg[5]  ( .D(go3[28]), .CK(clk), .RDN(n59483), .Q(
        \pe4/got [28]) );
  DRNQHSV4 \pe4/pe2/q_reg[4]  ( .D(go3[29]), .CK(clk), .RDN(n59399), .Q(
        \pe4/got [29]) );
  DRNQHSV4 \pe4/pe2/q_reg[3]  ( .D(go3[30]), .CK(clk), .RDN(n59444), .Q(
        \pe4/got [30]) );
  DRNQHSV4 \pe4/pe2/q_reg[2]  ( .D(go3[31]), .CK(clk), .RDN(n59401), .Q(
        \pe4/got [31]) );
  DRNQHSV4 \pe4/pe2/q_reg[1]  ( .D(go3[32]), .CK(clk), .RDN(n59471), .Q(
        \pe4/got [32]) );
  DRNQHSV4 \pe4/pe5/q_reg[22]  ( .D(pov3[22]), .CK(clk), .RDN(n59484), .Q(
        \pe4/pvq [22]) );
  DRNQHSV4 \pe4/pe5/q_reg[19]  ( .D(n60056), .CK(clk), .RDN(n59484), .Q(
        \pe4/pvq [19]) );
  DRNQHSV4 \pe4/pe5/q_reg[17]  ( .D(pov3[17]), .CK(clk), .RDN(n59429), .Q(
        \pe4/pvq [17]) );
  DRNQHSV4 \pe4/pe5/q_reg[15]  ( .D(n60087), .CK(clk), .RDN(n59445), .Q(
        \pe4/pvq [15]) );
  DRNQHSV4 \pe4/pe5/q_reg[13]  ( .D(n60059), .CK(clk), .RDN(n59415), .Q(
        \pe4/pvq [13]) );
  DRNQHSV4 \pe4/pe5/q_reg[11]  ( .D(n60089), .CK(clk), .RDN(n59460), .Q(
        \pe4/pvq [11]) );
  DRNQHSV4 \pe4/pe5/q_reg[10]  ( .D(n60090), .CK(clk), .RDN(n59400), .Q(
        \pe4/pvq [10]) );
  DRNQHSV4 \pe4/pe5/q_reg[9]  ( .D(pov3[9]), .CK(clk), .RDN(n59484), .Q(
        \pe4/pvq [9]) );
  DRNQHSV4 \pe4/pe5/q_reg[8]  ( .D(n60048), .CK(clk), .RDN(n59430), .Q(
        \pe4/pvq [8]) );
  DRNQHSV4 \pe4/pe5/q_reg[5]  ( .D(n60091), .CK(clk), .RDN(n59474), .Q(
        \pe4/pvq [5]) );
  DRNQHSV4 \pe4/pe5/q_reg[3]  ( .D(n60029), .CK(clk), .RDN(n59451), .Q(
        \pe4/pvq [3]) );
  DRNQHSV4 \pe4/pe6/q_reg[31]  ( .D(poh3[31]), .CK(clk), .RDN(n59408), .Q(
        \pe4/phq [31]) );
  DRNQHSV4 \pe4/pe6/q_reg[30]  ( .D(poh3[30]), .CK(clk), .RDN(n59476), .Q(
        \pe4/phq [30]) );
  DRNQHSV4 \pe4/pe6/q_reg[29]  ( .D(poh3[29]), .CK(clk), .RDN(n29729), .Q(
        \pe4/phq [29]) );
  DRNQHSV4 \pe4/pe6/q_reg[28]  ( .D(poh3[28]), .CK(clk), .RDN(n59449), .Q(
        \pe4/phq [28]) );
  DRNQHSV4 \pe4/pe6/q_reg[27]  ( .D(poh3[27]), .CK(clk), .RDN(n59454), .Q(
        \pe4/phq [27]) );
  DRNQHSV4 \pe4/pe6/q_reg[26]  ( .D(poh3[26]), .CK(clk), .RDN(n59408), .Q(
        \pe4/phq [26]) );
  DRNQHSV4 \pe4/pe6/q_reg[25]  ( .D(poh3[25]), .CK(clk), .RDN(n59445), .Q(
        \pe4/phq [25]) );
  DRNQHSV4 \pe4/pe6/q_reg[24]  ( .D(poh3[24]), .CK(clk), .RDN(n29729), .Q(
        \pe4/phq [24]) );
  DRNQHSV4 \pe4/pe6/q_reg[23]  ( .D(poh3[23]), .CK(clk), .RDN(n59453), .Q(
        \pe4/phq [23]) );
  DRNQHSV4 \pe4/pe6/q_reg[22]  ( .D(poh3[22]), .CK(clk), .RDN(n59479), .Q(
        \pe4/phq [22]) );
  DRNQHSV4 \pe4/pe6/q_reg[21]  ( .D(poh3[21]), .CK(clk), .RDN(n59483), .Q(
        \pe4/phq [21]) );
  DRNQHSV4 \pe4/pe6/q_reg[20]  ( .D(poh3[20]), .CK(clk), .RDN(n59478), .Q(
        \pe4/phq [20]) );
  DRNQHSV4 \pe4/pe6/q_reg[19]  ( .D(poh3[19]), .CK(clk), .RDN(n59481), .Q(
        \pe4/phq [19]) );
  DRNQHSV4 \pe4/pe6/q_reg[18]  ( .D(poh3[18]), .CK(clk), .RDN(n59449), .Q(
        \pe4/phq [18]) );
  DRNQHSV4 \pe4/pe6/q_reg[17]  ( .D(poh3[17]), .CK(clk), .RDN(n59429), .Q(
        \pe4/phq [17]) );
  DRNQHSV4 \pe4/pe6/q_reg[16]  ( .D(poh3[16]), .CK(clk), .RDN(n59414), .Q(
        \pe4/phq [16]) );
  DRNQHSV4 \pe4/pe6/q_reg[15]  ( .D(poh3[15]), .CK(clk), .RDN(n59461), .Q(
        \pe4/phq [15]) );
  DRNQHSV4 \pe4/pe6/q_reg[14]  ( .D(poh3[14]), .CK(clk), .RDN(n59925), .Q(
        \pe4/phq [14]) );
  DRNQHSV4 \pe4/pe6/q_reg[13]  ( .D(poh3[13]), .CK(clk), .RDN(n59404), .Q(
        \pe4/phq [13]) );
  DRNQHSV4 \pe4/pe6/q_reg[12]  ( .D(poh3[12]), .CK(clk), .RDN(n59425), .Q(
        \pe4/phq [12]) );
  DRNQHSV4 \pe4/pe6/q_reg[11]  ( .D(poh3[11]), .CK(clk), .RDN(n29731), .Q(
        \pe4/phq [11]) );
  DRNQHSV4 \pe4/pe6/q_reg[10]  ( .D(poh3[10]), .CK(clk), .RDN(n59493), .Q(
        \pe4/phq [10]) );
  DRNQHSV4 \pe4/pe6/q_reg[9]  ( .D(poh3[9]), .CK(clk), .RDN(n59925), .Q(
        \pe4/phq [9]) );
  DRNQHSV4 \pe4/pe6/q_reg[8]  ( .D(poh3[8]), .CK(clk), .RDN(n29734), .Q(
        \pe4/phq [8]) );
  DRNQHSV4 \pe4/pe6/q_reg[7]  ( .D(poh3[7]), .CK(clk), .RDN(n59438), .Q(
        \pe4/phq [7]) );
  DRNQHSV4 \pe4/pe6/q_reg[6]  ( .D(poh3[6]), .CK(clk), .RDN(n59462), .Q(
        \pe4/phq [6]) );
  DRNQHSV4 \pe4/pe6/q_reg[5]  ( .D(poh3[5]), .CK(clk), .RDN(n59402), .Q(
        \pe4/phq [5]) );
  DRNQHSV4 \pe4/pe6/q_reg[4]  ( .D(poh3[4]), .CK(clk), .RDN(n59433), .Q(
        \pe4/phq [4]) );
  DRNQHSV4 \pe4/pe6/q_reg[3]  ( .D(poh3[3]), .CK(clk), .RDN(n59442), .Q(
        \pe4/phq [3]) );
  DRNQHSV4 \pe4/pe6/q_reg[2]  ( .D(poh3[2]), .CK(clk), .RDN(n29734), .Q(
        \pe4/phq [2]) );
  DRNQHSV4 \pe4/pe6/q_reg[1]  ( .D(poh3[1]), .CK(clk), .RDN(n59459), .Q(
        \pe4/phq [1]) );
  DRNQHSV4 \pe4/pe7/q_reg  ( .D(n59998), .CK(clk), .RDN(n59403), .Q(\pe4/ctrq ) );
  DRNQHSV4 \pe4/pe12/q_reg[32]  ( .D(n59829), .CK(clk), .RDN(n59925), .Q(
        \pe4/bq[1] ) );
  DRNQHSV4 \pe4/pe12/q_reg[31]  ( .D(n59553), .CK(clk), .RDN(n59458), .Q(
        \pe4/bq[2] ) );
  DRNQHSV4 \pe4/pe12/q_reg[30]  ( .D(n59828), .CK(clk), .RDN(n59409), .Q(
        \pe4/bq[3] ) );
  DRNQHSV4 \pe4/pe12/q_reg[29]  ( .D(n59552), .CK(clk), .RDN(n59417), .Q(
        \pe4/bq[4] ) );
  DRNQHSV4 \pe4/pe12/q_reg[28]  ( .D(n59825), .CK(clk), .RDN(n59494), .Q(
        \pe4/bq[5] ) );
  DRNQHSV4 \pe4/pe12/q_reg[27]  ( .D(n59827), .CK(clk), .RDN(n59408), .Q(
        \pe4/bq[6] ) );
  DRNQHSV4 \pe4/pe12/q_reg[26]  ( .D(n59826), .CK(clk), .RDN(n59409), .Q(
        \pe4/bq[7] ) );
  DRNQHSV4 \pe4/pe12/q_reg[25]  ( .D(n59824), .CK(clk), .RDN(n59503), .Q(
        \pe4/bq[8] ) );
  DRNQHSV4 \pe4/pe12/q_reg[24]  ( .D(n59551), .CK(clk), .RDN(n59396), .Q(
        \pe4/bq[9] ) );
  DRNQHSV4 \pe4/pe12/q_reg[23]  ( .D(n59550), .CK(clk), .RDN(n59470), .Q(
        \pe4/bq[10] ) );
  DRNQHSV4 \pe4/pe12/q_reg[22]  ( .D(n59549), .CK(clk), .RDN(n59440), .Q(
        \pe4/bq[11] ) );
  DRNQHSV4 \pe4/pe12/q_reg[21]  ( .D(n59822), .CK(clk), .RDN(n59472), .Q(
        \pe4/bq[12] ) );
  DRNQHSV4 \pe4/pe12/q_reg[20]  ( .D(n59548), .CK(clk), .RDN(n59451), .Q(
        \pe4/bq[13] ) );
  DRNQHSV4 \pe4/pe12/q_reg[19]  ( .D(n59547), .CK(clk), .RDN(n59456), .Q(
        \pe4/bq[14] ) );
  DRNQHSV4 \pe4/pe12/q_reg[18]  ( .D(n59820), .CK(clk), .RDN(n59496), .Q(
        \pe4/bq[15] ) );
  DRNQHSV4 \pe4/pe12/q_reg[17]  ( .D(n59819), .CK(clk), .RDN(n59449), .Q(
        \pe4/bq[16] ) );
  DRNQHSV4 \pe4/pe12/q_reg[16]  ( .D(n59546), .CK(clk), .RDN(n59439), .Q(
        \pe4/bq[17] ) );
  DRNQHSV4 \pe4/pe12/q_reg[15]  ( .D(n59818), .CK(clk), .RDN(n59442), .Q(
        \pe4/bq[18] ) );
  DRNQHSV4 \pe4/pe12/q_reg[14]  ( .D(n59817), .CK(clk), .RDN(n59467), .Q(
        \pe4/bq[19] ) );
  DRNQHSV4 \pe4/pe12/q_reg[13]  ( .D(n59815), .CK(clk), .RDN(n59443), .Q(
        \pe4/bq[20] ) );
  DRNQHSV4 \pe4/pe12/q_reg[12]  ( .D(n59545), .CK(clk), .RDN(n59409), .Q(
        \pe4/bq[21] ) );
  DRNQHSV4 \pe4/pe12/q_reg[11]  ( .D(n59813), .CK(clk), .RDN(n59443), .Q(
        \pe4/bq[22] ) );
  DRNQHSV4 \pe4/pe12/q_reg[10]  ( .D(n59812), .CK(clk), .RDN(n59450), .Q(
        \pe4/bq[23] ) );
  DRNQHSV4 \pe4/pe12/q_reg[9]  ( .D(n59814), .CK(clk), .RDN(n59414), .Q(
        \pe4/bq[24] ) );
  DRNQHSV4 \pe4/pe12/q_reg[8]  ( .D(n59801), .CK(clk), .RDN(n59430), .Q(
        \pe4/bq[25] ) );
  DRNQHSV4 \pe4/pe12/q_reg[7]  ( .D(n59803), .CK(clk), .RDN(n59460), .Q(
        \pe4/bq[26] ) );
  DRNQHSV4 \pe4/pe12/q_reg[6]  ( .D(n59802), .CK(clk), .RDN(n59430), .Q(
        \pe4/bq[27] ) );
  DRNQHSV4 \pe4/pe12/q_reg[5]  ( .D(n59806), .CK(clk), .RDN(n59493), .Q(
        \pe4/bq[28] ) );
  DRNQHSV4 \pe4/pe12/q_reg[4]  ( .D(n59805), .CK(clk), .RDN(n59650), .Q(
        \pe4/bq[29] ) );
  DRNQHSV4 \pe4/pe12/q_reg[3]  ( .D(n59804), .CK(clk), .RDN(n59452), .Q(
        \pe4/bq[30] ) );
  DRNQHSV4 \pe4/pe12/q_reg[2]  ( .D(n59800), .CK(clk), .RDN(n59401), .Q(
        \pe4/bq[31] ) );
  DRNQHSV4 \pe4/pe12/q_reg[1]  ( .D(n59798), .CK(clk), .RDN(n59496), .Q(
        \pe4/bq[32] ) );
  DRNQHSV4 \pe4/pe13/q_reg  ( .D(\pe4/ti_1t ), .CK(clk), .RDN(n59457), .Q(
        \pe4/ti_1 ) );
  DRNQHSV4 \pe4/pe14/q_reg[2]  ( .D(n59382), .CK(clk), .RDN(n59655), .Q(
        \pe4/ti_7t [2]) );
  DRNQHSV4 \pe4/pe14/q_reg[4]  ( .D(n59524), .CK(clk), .RDN(n59434), .Q(
        \pe4/ti_7t [4]) );
  DRNQHSV4 \pe5/pe1/q_reg[32]  ( .D(ao4[1]), .CK(clk), .RDN(n59433), .Q(
        \pe5/aot [1]) );
  DRNQHSV4 \pe5/pe1/q_reg[31]  ( .D(ao4[2]), .CK(clk), .RDN(n59470), .Q(
        \pe5/aot [2]) );
  DRNQHSV4 \pe5/pe1/q_reg[30]  ( .D(ao4[3]), .CK(clk), .RDN(n59399), .Q(
        \pe5/aot [3]) );
  DRNQHSV4 \pe5/pe1/q_reg[29]  ( .D(ao4[4]), .CK(clk), .RDN(n59401), .Q(
        \pe5/aot [4]) );
  DRNQHSV4 \pe5/pe1/q_reg[28]  ( .D(ao4[5]), .CK(clk), .RDN(n59925), .Q(
        \pe5/aot [5]) );
  DRNQHSV4 \pe5/pe1/q_reg[27]  ( .D(ao4[6]), .CK(clk), .RDN(n59471), .Q(
        \pe5/aot [6]) );
  DRNQHSV4 \pe5/pe1/q_reg[26]  ( .D(ao4[7]), .CK(clk), .RDN(n59471), .Q(
        \pe5/aot [7]) );
  DRNQHSV4 \pe5/pe1/q_reg[25]  ( .D(ao4[8]), .CK(clk), .RDN(n59396), .Q(
        \pe5/aot [8]) );
  DRNQHSV4 \pe5/pe1/q_reg[24]  ( .D(ao4[9]), .CK(clk), .RDN(n59410), .Q(
        \pe5/aot [9]) );
  DRNQHSV4 \pe5/pe1/q_reg[23]  ( .D(ao4[10]), .CK(clk), .RDN(n59472), .Q(
        \pe5/aot [10]) );
  DRNQHSV4 \pe5/pe1/q_reg[22]  ( .D(ao4[11]), .CK(clk), .RDN(n59472), .Q(
        \pe5/aot [11]) );
  DRNQHSV4 \pe5/pe1/q_reg[21]  ( .D(ao4[12]), .CK(clk), .RDN(n59472), .Q(
        \pe5/aot [12]) );
  DRNQHSV4 \pe5/pe1/q_reg[20]  ( .D(ao4[13]), .CK(clk), .RDN(n59471), .Q(
        \pe5/aot [13]) );
  DRNQHSV4 \pe5/pe1/q_reg[19]  ( .D(ao4[14]), .CK(clk), .RDN(n59397), .Q(
        \pe5/aot [14]) );
  DRNQHSV4 \pe5/pe1/q_reg[18]  ( .D(ao4[15]), .CK(clk), .RDN(n59471), .Q(
        \pe5/aot [15]) );
  DRNQHSV4 \pe5/pe1/q_reg[17]  ( .D(ao4[16]), .CK(clk), .RDN(n59410), .Q(
        \pe5/aot [16]) );
  DRNQHSV4 \pe5/pe1/q_reg[16]  ( .D(ao4[17]), .CK(clk), .RDN(n59397), .Q(
        \pe5/aot [17]) );
  DRNQHSV4 \pe5/pe1/q_reg[15]  ( .D(ao4[18]), .CK(clk), .RDN(n59396), .Q(
        \pe5/aot [18]) );
  DRNQHSV4 \pe5/pe1/q_reg[14]  ( .D(ao4[19]), .CK(clk), .RDN(n59470), .Q(
        \pe5/aot [19]) );
  DRNQHSV4 \pe5/pe1/q_reg[13]  ( .D(ao4[20]), .CK(clk), .RDN(n59471), .Q(
        \pe5/aot [20]) );
  DRNQHSV4 \pe5/pe1/q_reg[12]  ( .D(ao4[21]), .CK(clk), .RDN(n59654), .Q(
        \pe5/aot [21]) );
  DRNQHSV4 \pe5/pe1/q_reg[11]  ( .D(ao4[22]), .CK(clk), .RDN(n59654), .Q(
        \pe5/aot [22]) );
  DRNQHSV4 \pe5/pe1/q_reg[10]  ( .D(ao4[23]), .CK(clk), .RDN(n59655), .Q(
        \pe5/aot [23]) );
  DRNQHSV4 \pe5/pe1/q_reg[9]  ( .D(ao4[24]), .CK(clk), .RDN(n59434), .Q(
        \pe5/aot [24]) );
  DRNQHSV4 \pe5/pe1/q_reg[8]  ( .D(ao4[25]), .CK(clk), .RDN(n59653), .Q(
        \pe5/aot [25]) );
  DRNQHSV4 \pe5/pe1/q_reg[7]  ( .D(ao4[26]), .CK(clk), .RDN(n59653), .Q(
        \pe5/aot [26]) );
  DRNQHSV4 \pe5/pe1/q_reg[6]  ( .D(ao4[27]), .CK(clk), .RDN(n59480), .Q(
        \pe5/aot [27]) );
  DRNQHSV4 \pe5/pe1/q_reg[5]  ( .D(ao4[28]), .CK(clk), .RDN(n29733), .Q(
        \pe5/aot [28]) );
  DRNQHSV4 \pe5/pe1/q_reg[4]  ( .D(ao4[29]), .CK(clk), .RDN(n59405), .Q(
        \pe5/aot [29]) );
  DRNQHSV4 \pe5/pe1/q_reg[3]  ( .D(ao4[30]), .CK(clk), .RDN(n59396), .Q(
        \pe5/aot [30]) );
  DRNQHSV4 \pe5/pe1/q_reg[2]  ( .D(ao4[31]), .CK(clk), .RDN(n59461), .Q(
        \pe5/aot [31]) );
  DRNQHSV4 \pe5/pe1/q_reg[1]  ( .D(ao4[32]), .CK(clk), .RDN(n59473), .Q(
        \pe5/aot [32]) );
  DRNQHSV4 \pe5/pe2/q_reg[32]  ( .D(go4[1]), .CK(clk), .RDN(n59466), .Q(
        \pe5/got [1]) );
  DRNQHSV4 \pe5/pe2/q_reg[31]  ( .D(go4[2]), .CK(clk), .RDN(n59444), .Q(
        \pe5/got [2]) );
  DRNQHSV4 \pe5/pe2/q_reg[30]  ( .D(go4[3]), .CK(clk), .RDN(n59437), .Q(
        \pe5/got [3]) );
  DRNQHSV4 \pe5/pe2/q_reg[29]  ( .D(go4[4]), .CK(clk), .RDN(n59654), .Q(
        \pe5/got [4]) );
  DRNQHSV4 \pe5/pe2/q_reg[28]  ( .D(go4[5]), .CK(clk), .RDN(n59655), .Q(
        \pe5/got [5]) );
  DRNQHSV4 \pe5/pe2/q_reg[27]  ( .D(go4[6]), .CK(clk), .RDN(n59654), .Q(
        \pe5/got [6]) );
  DRNQHSV4 \pe5/pe2/q_reg[26]  ( .D(go4[7]), .CK(clk), .RDN(n59477), .Q(
        \pe5/got [7]) );
  DRNQHSV4 \pe5/pe2/q_reg[25]  ( .D(go4[8]), .CK(clk), .RDN(n59452), .Q(
        \pe5/got [8]) );
  DRNQHSV4 \pe5/pe2/q_reg[24]  ( .D(go4[9]), .CK(clk), .RDN(n59465), .Q(
        \pe5/got [9]) );
  DRNQHSV4 \pe5/pe2/q_reg[23]  ( .D(go4[10]), .CK(clk), .RDN(n59490), .Q(
        \pe5/got [10]) );
  DRNQHSV4 \pe5/pe2/q_reg[22]  ( .D(go4[11]), .CK(clk), .RDN(n59652), .Q(
        \pe5/got [11]) );
  DRNQHSV4 \pe5/pe2/q_reg[21]  ( .D(go4[12]), .CK(clk), .RDN(n59652), .Q(
        \pe5/got [12]) );
  DRNQHSV4 \pe5/pe2/q_reg[20]  ( .D(go4[13]), .CK(clk), .RDN(n59925), .Q(
        \pe5/got [13]) );
  DRNQHSV4 \pe5/pe2/q_reg[19]  ( .D(go4[14]), .CK(clk), .RDN(n59432), .Q(
        \pe5/got [14]) );
  DRNQHSV4 \pe5/pe2/q_reg[18]  ( .D(go4[15]), .CK(clk), .RDN(n59408), .Q(
        \pe5/got [15]) );
  DRNQHSV4 \pe5/pe2/q_reg[17]  ( .D(go4[16]), .CK(clk), .RDN(n59923), .Q(
        \pe5/got [16]) );
  DRNQHSV4 \pe5/pe2/q_reg[16]  ( .D(go4[17]), .CK(clk), .RDN(n59401), .Q(
        \pe5/got [17]) );
  DRNQHSV4 \pe5/pe2/q_reg[15]  ( .D(go4[18]), .CK(clk), .RDN(n59437), .Q(
        \pe5/got [18]) );
  DRNQHSV4 \pe5/pe2/q_reg[14]  ( .D(go4[19]), .CK(clk), .RDN(n59463), .Q(
        \pe5/got [19]) );
  DRNQHSV4 \pe5/pe2/q_reg[13]  ( .D(go4[20]), .CK(clk), .RDN(n59477), .Q(
        \pe5/got [20]) );
  DRNQHSV4 \pe5/pe2/q_reg[12]  ( .D(go4[21]), .CK(clk), .RDN(n59436), .Q(
        \pe5/got [21]) );
  DRNQHSV4 \pe5/pe2/q_reg[11]  ( .D(go4[22]), .CK(clk), .RDN(n59651), .Q(
        \pe5/got [22]) );
  DRNQHSV4 \pe5/pe2/q_reg[10]  ( .D(go4[23]), .CK(clk), .RDN(n59651), .Q(
        \pe5/got [23]) );
  DRNQHSV4 \pe5/pe2/q_reg[9]  ( .D(go4[24]), .CK(clk), .RDN(n59651), .Q(
        \pe5/got [24]) );
  DRNQHSV4 \pe5/pe2/q_reg[8]  ( .D(go4[25]), .CK(clk), .RDN(n59444), .Q(
        \pe5/got [25]) );
  DRNQHSV4 \pe5/pe2/q_reg[7]  ( .D(go4[26]), .CK(clk), .RDN(n59490), .Q(
        \pe5/got [26]) );
  DRNQHSV4 \pe5/pe2/q_reg[6]  ( .D(go4[27]), .CK(clk), .RDN(n59451), .Q(
        \pe5/got [27]) );
  DRNQHSV4 \pe5/pe2/q_reg[5]  ( .D(go4[28]), .CK(clk), .RDN(n59464), .Q(
        \pe5/got [28]) );
  DRNQHSV4 \pe5/pe2/q_reg[4]  ( .D(go4[29]), .CK(clk), .RDN(n59430), .Q(
        \pe5/got [29]) );
  DRNQHSV4 \pe5/pe2/q_reg[3]  ( .D(go4[30]), .CK(clk), .RDN(n59488), .Q(
        \pe5/got [30]) );
  DRNQHSV4 \pe5/pe2/q_reg[2]  ( .D(go4[31]), .CK(clk), .RDN(n59413), .Q(
        \pe5/got [31]) );
  DRNQHSV4 \pe5/pe2/q_reg[1]  ( .D(go4[32]), .CK(clk), .RDN(n29734), .Q(
        \pe5/got [32]) );
  DRNQHSV4 \pe5/pe5/q_reg[24]  ( .D(n60057), .CK(clk), .RDN(n59510), .Q(
        \pe5/pvq [24]) );
  DRNQHSV4 \pe5/pe5/q_reg[23]  ( .D(pov4[23]), .CK(clk), .RDN(n59467), .Q(
        \pe5/pvq [23]) );
  DRNQHSV4 \pe5/pe5/q_reg[21]  ( .D(n60061), .CK(clk), .RDN(n59435), .Q(
        \pe5/pvq [21]) );
  DRNQHSV4 \pe5/pe5/q_reg[20]  ( .D(pov4[20]), .CK(clk), .RDN(n59488), .Q(
        \pe5/pvq [20]) );
  DRNQHSV4 \pe5/pe5/q_reg[19]  ( .D(n60066), .CK(clk), .RDN(n59425), .Q(
        \pe5/pvq [19]) );
  DRNQHSV4 \pe5/pe5/q_reg[18]  ( .D(n60064), .CK(clk), .RDN(n29732), .Q(
        \pe5/pvq [18]) );
  DRNQHSV4 \pe5/pe5/q_reg[17]  ( .D(n60011), .CK(clk), .RDN(n59424), .Q(
        \pe5/pvq [17]) );
  DRNQHSV4 \pe5/pe5/q_reg[15]  ( .D(pov4[15]), .CK(clk), .RDN(n59409), .Q(
        \pe5/pvq [15]) );
  DRNQHSV4 \pe5/pe5/q_reg[13]  ( .D(n60023), .CK(clk), .RDN(n59451), .Q(
        \pe5/pvq [13]) );
  DRNQHSV4 \pe5/pe5/q_reg[12]  ( .D(n60027), .CK(clk), .RDN(n59437), .Q(
        \pe5/pvq [12]) );
  DRNQHSV4 \pe5/pe5/q_reg[10]  ( .D(n60049), .CK(clk), .RDN(n59433), .Q(
        \pe5/pvq [10]) );
  DRNQHSV4 \pe5/pe5/q_reg[8]  ( .D(n60079), .CK(clk), .RDN(n59447), .Q(
        \pe5/pvq [8]) );
  DRNQHSV4 \pe5/pe5/q_reg[7]  ( .D(n60080), .CK(clk), .RDN(n59656), .Q(
        \pe5/pvq [7]) );
  DRNQHSV4 \pe5/pe5/q_reg[6]  ( .D(n60081), .CK(clk), .RDN(n59440), .Q(
        \pe5/pvq [6]) );
  DRNQHSV4 \pe5/pe5/q_reg[3]  ( .D(n60034), .CK(clk), .RDN(n59458), .Q(
        \pe5/pvq [3]) );
  DRNQHSV4 \pe5/pe5/q_reg[2]  ( .D(n60083), .CK(clk), .RDN(n59479), .Q(
        \pe5/pvq [2]) );
  DRNQHSV4 \pe5/pe6/q_reg[31]  ( .D(poh4[31]), .CK(clk), .RDN(n59457), .Q(
        \pe5/phq [31]) );
  DRNQHSV4 \pe5/pe6/q_reg[29]  ( .D(poh4[29]), .CK(clk), .RDN(n59459), .Q(
        \pe5/phq [29]) );
  DRNQHSV4 \pe5/pe6/q_reg[28]  ( .D(poh4[28]), .CK(clk), .RDN(n59400), .Q(
        \pe5/phq [28]) );
  DRNQHSV4 \pe5/pe6/q_reg[27]  ( .D(poh4[27]), .CK(clk), .RDN(n59459), .Q(
        \pe5/phq [27]) );
  DRNQHSV4 \pe5/pe6/q_reg[26]  ( .D(poh4[26]), .CK(clk), .RDN(n59466), .Q(
        \pe5/phq [26]) );
  DRNQHSV4 \pe5/pe6/q_reg[25]  ( .D(poh4[25]), .CK(clk), .RDN(n59655), .Q(
        \pe5/phq [25]) );
  DRNQHSV4 \pe5/pe6/q_reg[24]  ( .D(poh4[24]), .CK(clk), .RDN(n59449), .Q(
        \pe5/phq [24]) );
  DRNQHSV4 \pe5/pe6/q_reg[23]  ( .D(poh4[23]), .CK(clk), .RDN(n59459), .Q(
        \pe5/phq [23]) );
  DRNQHSV4 \pe5/pe6/q_reg[22]  ( .D(poh4[22]), .CK(clk), .RDN(n59477), .Q(
        \pe5/phq [22]) );
  DRNQHSV4 \pe5/pe6/q_reg[21]  ( .D(poh4[21]), .CK(clk), .RDN(n59401), .Q(
        \pe5/phq [21]) );
  DRNQHSV4 \pe5/pe6/q_reg[20]  ( .D(poh4[20]), .CK(clk), .RDN(n59466), .Q(
        \pe5/phq [20]) );
  DRNQHSV4 \pe5/pe6/q_reg[19]  ( .D(poh4[19]), .CK(clk), .RDN(n59438), .Q(
        \pe5/phq [19]) );
  DRNQHSV4 \pe5/pe6/q_reg[18]  ( .D(poh4[18]), .CK(clk), .RDN(n59447), .Q(
        \pe5/phq [18]) );
  DRNQHSV4 \pe5/pe6/q_reg[17]  ( .D(poh4[17]), .CK(clk), .RDN(n59401), .Q(
        \pe5/phq [17]) );
  DRNQHSV4 \pe5/pe6/q_reg[16]  ( .D(poh4[16]), .CK(clk), .RDN(n59436), .Q(
        \pe5/phq [16]) );
  DRNQHSV4 \pe5/pe6/q_reg[15]  ( .D(poh4[15]), .CK(clk), .RDN(n59400), .Q(
        \pe5/phq [15]) );
  DRNQHSV4 \pe5/pe6/q_reg[14]  ( .D(poh4[14]), .CK(clk), .RDN(n59436), .Q(
        \pe5/phq [14]) );
  DRNQHSV4 \pe5/pe6/q_reg[13]  ( .D(poh4[13]), .CK(clk), .RDN(n59466), .Q(
        \pe5/phq [13]) );
  DRNQHSV4 \pe5/pe6/q_reg[12]  ( .D(poh4[12]), .CK(clk), .RDN(n59409), .Q(
        \pe5/phq [12]) );
  DRNQHSV4 \pe5/pe6/q_reg[11]  ( .D(poh4[11]), .CK(clk), .RDN(n59491), .Q(
        \pe5/phq [11]) );
  DRNQHSV4 \pe5/pe6/q_reg[10]  ( .D(poh4[10]), .CK(clk), .RDN(n59408), .Q(
        \pe5/phq [10]) );
  DRNQHSV4 \pe5/pe6/q_reg[9]  ( .D(poh4[9]), .CK(clk), .RDN(n59658), .Q(
        \pe5/phq [9]) );
  DRNQHSV4 \pe5/pe6/q_reg[8]  ( .D(poh4[8]), .CK(clk), .RDN(n59448), .Q(
        \pe5/phq [8]) );
  DRNQHSV4 \pe5/pe6/q_reg[7]  ( .D(poh4[7]), .CK(clk), .RDN(n59472), .Q(
        \pe5/phq [7]) );
  DRNQHSV4 \pe5/pe6/q_reg[6]  ( .D(poh4[6]), .CK(clk), .RDN(n59445), .Q(
        \pe5/phq [6]) );
  DRNQHSV4 \pe5/pe6/q_reg[5]  ( .D(poh4[5]), .CK(clk), .RDN(n29731), .Q(
        \pe5/phq [5]) );
  DRNQHSV4 \pe5/pe6/q_reg[4]  ( .D(poh4[4]), .CK(clk), .RDN(n59438), .Q(
        \pe5/phq [4]) );
  DRNQHSV4 \pe5/pe6/q_reg[3]  ( .D(poh4[3]), .CK(clk), .RDN(n59406), .Q(
        \pe5/phq [3]) );
  DRNQHSV4 \pe5/pe6/q_reg[2]  ( .D(poh4[2]), .CK(clk), .RDN(n59656), .Q(
        \pe5/phq [2]) );
  DRNQHSV4 \pe5/pe6/q_reg[1]  ( .D(poh4[1]), .CK(clk), .RDN(n59460), .Q(
        \pe5/phq [1]) );
  DRNQHSV4 \pe5/pe12/q_reg[32]  ( .D(n59865), .CK(clk), .RDN(n59412), .Q(
        \pe5/bq[1] ) );
  DRNQHSV4 \pe5/pe12/q_reg[31]  ( .D(n59544), .CK(clk), .RDN(n59456), .Q(
        \pe5/bq[2] ) );
  DRNQHSV4 \pe5/pe12/q_reg[29]  ( .D(n59543), .CK(clk), .RDN(n59445), .Q(
        \pe5/bq[4] ) );
  DRNQHSV4 \pe5/pe12/q_reg[28]  ( .D(n59862), .CK(clk), .RDN(n59448), .Q(
        \pe5/bq[5] ) );
  DRNQHSV4 \pe5/pe12/q_reg[27]  ( .D(n59863), .CK(clk), .RDN(n29732), .Q(
        \pe5/bq[6] ) );
  DRNQHSV4 \pe5/pe12/q_reg[26]  ( .D(n59861), .CK(clk), .RDN(n59921), .Q(
        \pe5/bq[7] ) );
  DRNQHSV4 \pe5/pe12/q_reg[25]  ( .D(n59859), .CK(clk), .RDN(n59470), .Q(
        \pe5/bq[8] ) );
  DRNQHSV4 \pe5/pe12/q_reg[24]  ( .D(n59858), .CK(clk), .RDN(n59502), .Q(
        \pe5/bq[9] ) );
  DRNQHSV4 \pe5/pe12/q_reg[23]  ( .D(n59542), .CK(clk), .RDN(n59491), .Q(
        \pe5/bq[10] ) );
  DRNQHSV4 \pe5/pe12/q_reg[22]  ( .D(n59541), .CK(clk), .RDN(n59502), .Q(
        \pe5/bq[11] ) );
  DRNQHSV4 \pe5/pe12/q_reg[21]  ( .D(n59860), .CK(clk), .RDN(n59415), .Q(
        \pe5/bq[12] ) );
  DRNQHSV4 \pe5/pe12/q_reg[20]  ( .D(n59854), .CK(clk), .RDN(n29733), .Q(
        \pe5/bq[13] ) );
  DRNQHSV4 \pe5/pe12/q_reg[19]  ( .D(n59852), .CK(clk), .RDN(n59477), .Q(
        \pe5/bq[14] ) );
  DRNQHSV4 \pe5/pe12/q_reg[18]  ( .D(n59856), .CK(clk), .RDN(n59655), .Q(
        \pe5/bq[15] ) );
  DRNQHSV4 \pe5/pe12/q_reg[17]  ( .D(n59851), .CK(clk), .RDN(n29732), .Q(
        \pe5/bq[16] ) );
  DRNQHSV4 \pe5/pe12/q_reg[16]  ( .D(n59853), .CK(clk), .RDN(n59465), .Q(
        \pe5/bq[17] ) );
  DRNQHSV4 \pe5/pe12/q_reg[15]  ( .D(n59855), .CK(clk), .RDN(n59658), .Q(
        \pe5/bq[18] ) );
  DRNQHSV4 \pe5/pe12/q_reg[14]  ( .D(n59850), .CK(clk), .RDN(n59417), .Q(
        \pe5/bq[19] ) );
  DRNQHSV4 \pe5/pe12/q_reg[13]  ( .D(n59848), .CK(clk), .RDN(n59444), .Q(
        \pe5/bq[20] ) );
  DRNQHSV4 \pe5/pe12/q_reg[12]  ( .D(n59847), .CK(clk), .RDN(n59448), .Q(
        \pe5/bq[21] ) );
  DRNQHSV4 \pe5/pe12/q_reg[11]  ( .D(n59849), .CK(clk), .RDN(n59478), .Q(
        \pe5/bq[22] ) );
  DRNQHSV4 \pe5/pe12/q_reg[10]  ( .D(n59846), .CK(clk), .RDN(n59461), .Q(
        \pe5/bq[23] ) );
  DRNQHSV4 \pe5/pe12/q_reg[9]  ( .D(n59842), .CK(clk), .RDN(n59429), .Q(
        \pe5/bq[24] ) );
  DRNQHSV4 \pe5/pe12/q_reg[8]  ( .D(n59843), .CK(clk), .RDN(n59467), .Q(
        \pe5/bq[25] ) );
  DRNQHSV4 \pe5/pe12/q_reg[7]  ( .D(n59844), .CK(clk), .RDN(n59453), .Q(
        \pe5/bq[26] ) );
  DRNQHSV4 \pe5/pe12/q_reg[6]  ( .D(n59841), .CK(clk), .RDN(n29733), .Q(
        \pe5/bq[27] ) );
  DRNQHSV4 \pe5/pe12/q_reg[5]  ( .D(n59840), .CK(clk), .RDN(n59418), .Q(
        \pe5/bq[28] ) );
  DRNQHSV4 \pe5/pe12/q_reg[4]  ( .D(n59836), .CK(clk), .RDN(n59921), .Q(
        \pe5/bq[29] ) );
  DRNQHSV4 \pe5/pe12/q_reg[3]  ( .D(n59568), .CK(clk), .RDN(n59458), .Q(
        \pe5/bq[30] ) );
  DRNQHSV4 \pe5/pe12/q_reg[2]  ( .D(n59540), .CK(clk), .RDN(n59409), .Q(
        \pe5/bq[31] ) );
  DRNQHSV4 \pe5/pe12/q_reg[1]  ( .D(n59830), .CK(clk), .RDN(n59432), .Q(
        \pe5/bq[32] ) );
  DRNQHSV4 \pe5/pe13/q_reg  ( .D(\pe5/ti_1t ), .CK(clk), .RDN(n59492), .Q(
        \pe5/ti_1 ) );
  DRNQHSV4 \pe5/pe14/q_reg[6]  ( .D(n37723), .CK(clk), .RDN(n59419), .Q(
        \pe5/ti_7t [6]) );
  DRNQHSV4 \pe5/pe14/q_reg[7]  ( .D(n47338), .CK(clk), .RDN(n59454), .Q(
        \pe5/ti_7t [7]) );
  DRNQHSV4 \pe6/pe1/q_reg[32]  ( .D(ao5[1]), .CK(clk), .RDN(n59409), .Q(
        \pe6/aot [1]) );
  DRNQHSV4 \pe6/pe1/q_reg[31]  ( .D(ao5[2]), .CK(clk), .RDN(n59443), .Q(
        \pe6/aot [2]) );
  DRNQHSV4 \pe6/pe1/q_reg[30]  ( .D(ao5[3]), .CK(clk), .RDN(n59403), .Q(
        \pe6/aot [3]) );
  DRNQHSV4 \pe6/pe1/q_reg[29]  ( .D(ao5[4]), .CK(clk), .RDN(n59467), .Q(
        \pe6/aot [4]) );
  DRNQHSV4 \pe6/pe1/q_reg[28]  ( .D(ao5[5]), .CK(clk), .RDN(n59407), .Q(
        \pe6/aot [5]) );
  DRNQHSV4 \pe6/pe1/q_reg[27]  ( .D(ao5[6]), .CK(clk), .RDN(n59462), .Q(
        \pe6/aot [6]) );
  DRNQHSV4 \pe6/pe1/q_reg[26]  ( .D(ao5[7]), .CK(clk), .RDN(n59467), .Q(
        \pe6/aot [7]) );
  DRNQHSV4 \pe6/pe1/q_reg[25]  ( .D(ao5[8]), .CK(clk), .RDN(n59455), .Q(
        \pe6/aot [8]) );
  DRNQHSV4 \pe6/pe1/q_reg[24]  ( .D(ao5[9]), .CK(clk), .RDN(n59481), .Q(
        \pe6/aot [9]) );
  DRNQHSV4 \pe6/pe1/q_reg[23]  ( .D(ao5[10]), .CK(clk), .RDN(n59404), .Q(
        \pe6/aot [10]) );
  DRNQHSV4 \pe6/pe1/q_reg[22]  ( .D(ao5[11]), .CK(clk), .RDN(n59653), .Q(
        \pe6/aot [11]) );
  DRNQHSV4 \pe6/pe1/q_reg[21]  ( .D(ao5[12]), .CK(clk), .RDN(n59415), .Q(
        \pe6/aot [12]) );
  DRNQHSV4 \pe6/pe1/q_reg[20]  ( .D(ao5[13]), .CK(clk), .RDN(n59418), .Q(
        \pe6/aot [13]) );
  DRNQHSV4 \pe6/pe1/q_reg[19]  ( .D(ao5[14]), .CK(clk), .RDN(n59659), .Q(
        \pe6/aot [14]) );
  DRNQHSV4 \pe6/pe1/q_reg[18]  ( .D(ao5[15]), .CK(clk), .RDN(n59440), .Q(
        \pe6/aot [15]) );
  DRNQHSV4 \pe6/pe1/q_reg[17]  ( .D(ao5[16]), .CK(clk), .RDN(n59406), .Q(
        \pe6/aot [16]) );
  DRNQHSV4 \pe6/pe1/q_reg[16]  ( .D(ao5[17]), .CK(clk), .RDN(n59429), .Q(
        \pe6/aot [17]) );
  DRNQHSV4 \pe6/pe1/q_reg[15]  ( .D(ao5[18]), .CK(clk), .RDN(n59479), .Q(
        \pe6/aot [18]) );
  DRNQHSV4 \pe6/pe1/q_reg[14]  ( .D(ao5[19]), .CK(clk), .RDN(n59925), .Q(
        \pe6/aot [19]) );
  DRNQHSV4 \pe6/pe1/q_reg[13]  ( .D(ao5[20]), .CK(clk), .RDN(n29729), .Q(
        \pe6/aot [20]) );
  DRNQHSV4 \pe6/pe1/q_reg[12]  ( .D(ao5[21]), .CK(clk), .RDN(n59493), .Q(
        \pe6/aot [21]) );
  DRNQHSV4 \pe6/pe1/q_reg[11]  ( .D(ao5[22]), .CK(clk), .RDN(n59448), .Q(
        \pe6/aot [22]) );
  DRNQHSV4 \pe6/pe1/q_reg[10]  ( .D(ao5[23]), .CK(clk), .RDN(n59455), .Q(
        \pe6/aot [23]) );
  DRNQHSV4 \pe6/pe1/q_reg[9]  ( .D(ao5[24]), .CK(clk), .RDN(n59482), .Q(
        \pe6/aot [24]) );
  DRNQHSV4 \pe6/pe1/q_reg[8]  ( .D(ao5[25]), .CK(clk), .RDN(n59481), .Q(
        \pe6/aot [25]) );
  DRNQHSV4 \pe6/pe1/q_reg[7]  ( .D(ao5[26]), .CK(clk), .RDN(n59463), .Q(
        \pe6/aot [26]) );
  DRNQHSV4 \pe6/pe1/q_reg[6]  ( .D(ao5[27]), .CK(clk), .RDN(n59411), .Q(
        \pe6/aot [27]) );
  DRNQHSV4 \pe6/pe1/q_reg[5]  ( .D(ao5[28]), .CK(clk), .RDN(n59652), .Q(
        \pe6/aot [28]) );
  DRNQHSV4 \pe6/pe1/q_reg[4]  ( .D(ao5[29]), .CK(clk), .RDN(n59649), .Q(
        \pe6/aot [29]) );
  DRNQHSV4 \pe6/pe1/q_reg[3]  ( .D(ao5[30]), .CK(clk), .RDN(n59481), .Q(
        \pe6/aot [30]) );
  DRNQHSV4 \pe6/pe1/q_reg[2]  ( .D(ao5[31]), .CK(clk), .RDN(n59416), .Q(
        \pe6/aot [31]) );
  DRNQHSV4 \pe6/pe1/q_reg[1]  ( .D(ao5[32]), .CK(clk), .RDN(n59482), .Q(
        \pe6/aot [32]) );
  DRNQHSV4 \pe6/pe2/q_reg[32]  ( .D(go5[1]), .CK(clk), .RDN(n59482), .Q(
        \pe6/got [1]) );
  DRNQHSV4 \pe6/pe2/q_reg[31]  ( .D(go5[2]), .CK(clk), .RDN(n29734), .Q(
        \pe6/got [2]) );
  DRNQHSV4 \pe6/pe2/q_reg[30]  ( .D(go5[3]), .CK(clk), .RDN(n59416), .Q(
        \pe6/got [3]) );
  DRNQHSV4 \pe6/pe2/q_reg[29]  ( .D(go5[4]), .CK(clk), .RDN(n59494), .Q(
        \pe6/got [4]) );
  DRNQHSV4 \pe6/pe2/q_reg[28]  ( .D(go5[5]), .CK(clk), .RDN(n59463), .Q(
        \pe6/got [5]) );
  DRNQHSV4 \pe6/pe2/q_reg[27]  ( .D(go5[6]), .CK(clk), .RDN(n59419), .Q(
        \pe6/got [6]) );
  DRNQHSV4 \pe6/pe2/q_reg[26]  ( .D(go5[7]), .CK(clk), .RDN(n59463), .Q(
        \pe6/got [7]) );
  DRNQHSV4 \pe6/pe2/q_reg[25]  ( .D(go5[8]), .CK(clk), .RDN(n59440), .Q(
        \pe6/got [8]) );
  DRNQHSV4 \pe6/pe2/q_reg[24]  ( .D(go5[9]), .CK(clk), .RDN(n59502), .Q(
        \pe6/got [9]) );
  DRNQHSV4 \pe6/pe2/q_reg[23]  ( .D(go5[10]), .CK(clk), .RDN(n59922), .Q(
        \pe6/got [10]) );
  DRNQHSV4 \pe6/pe2/q_reg[22]  ( .D(go5[11]), .CK(clk), .RDN(n59403), .Q(
        \pe6/got [11]) );
  DRNQHSV4 \pe6/pe2/q_reg[21]  ( .D(go5[12]), .CK(clk), .RDN(n59409), .Q(
        \pe6/got [12]) );
  DRNQHSV4 \pe6/pe2/q_reg[20]  ( .D(go5[13]), .CK(clk), .RDN(n59650), .Q(
        \pe6/got [13]) );
  DRNQHSV4 \pe6/pe2/q_reg[19]  ( .D(go5[14]), .CK(clk), .RDN(n59433), .Q(
        \pe6/got [14]) );
  DRNQHSV4 \pe6/pe2/q_reg[18]  ( .D(go5[15]), .CK(clk), .RDN(n59404), .Q(
        \pe6/got [15]) );
  DRNQHSV4 \pe6/pe2/q_reg[17]  ( .D(go5[16]), .CK(clk), .RDN(n59429), .Q(
        \pe6/got [16]) );
  DRNQHSV4 \pe6/pe2/q_reg[16]  ( .D(go5[17]), .CK(clk), .RDN(n59454), .Q(
        \pe6/got [17]) );
  DRNQHSV4 \pe6/pe2/q_reg[15]  ( .D(go5[18]), .CK(clk), .RDN(n29731), .Q(
        \pe6/got [18]) );
  DRNQHSV4 \pe6/pe2/q_reg[14]  ( .D(go5[19]), .CK(clk), .RDN(n59402), .Q(
        \pe6/got [19]) );
  DRNQHSV4 \pe6/pe2/q_reg[13]  ( .D(go5[20]), .CK(clk), .RDN(n59453), .Q(
        \pe6/got [20]) );
  DRNQHSV4 \pe6/pe2/q_reg[12]  ( .D(go5[21]), .CK(clk), .RDN(n59451), .Q(
        \pe6/got [21]) );
  DRNQHSV4 \pe6/pe2/q_reg[11]  ( .D(go5[22]), .CK(clk), .RDN(n59925), .Q(
        \pe6/got [22]) );
  DRNQHSV4 \pe6/pe2/q_reg[10]  ( .D(go5[23]), .CK(clk), .RDN(n59404), .Q(
        \pe6/got [23]) );
  DRNQHSV4 \pe6/pe2/q_reg[9]  ( .D(go5[24]), .CK(clk), .RDN(n59408), .Q(
        \pe6/got [24]) );
  DRNQHSV4 \pe6/pe2/q_reg[8]  ( .D(go5[25]), .CK(clk), .RDN(n59396), .Q(
        \pe6/got [25]) );
  DRNQHSV4 \pe6/pe2/q_reg[7]  ( .D(go5[26]), .CK(clk), .RDN(n59467), .Q(
        \pe6/got [26]) );
  DRNQHSV4 \pe6/pe2/q_reg[6]  ( .D(go5[27]), .CK(clk), .RDN(n59404), .Q(
        \pe6/got [27]) );
  DRNQHSV4 \pe6/pe2/q_reg[5]  ( .D(go5[28]), .CK(clk), .RDN(n59481), .Q(
        \pe6/got [28]) );
  DRNQHSV4 \pe6/pe2/q_reg[4]  ( .D(go5[29]), .CK(clk), .RDN(n59454), .Q(
        \pe6/got [29]) );
  DRNQHSV4 \pe6/pe2/q_reg[3]  ( .D(go5[30]), .CK(clk), .RDN(n59512), .Q(
        \pe6/got [30]) );
  DRNQHSV4 \pe6/pe2/q_reg[2]  ( .D(go5[31]), .CK(clk), .RDN(n59481), .Q(
        \pe6/got [31]) );
  DRNQHSV4 \pe6/pe2/q_reg[1]  ( .D(go5[32]), .CK(clk), .RDN(n29734), .Q(
        \pe6/got [32]) );
  DRNQHSV4 \pe6/pe5/q_reg[19]  ( .D(n60032), .CK(clk), .RDN(n59463), .Q(
        \pe6/pvq [19]) );
  DRNQHSV4 \pe6/pe5/q_reg[17]  ( .D(n60069), .CK(clk), .RDN(n59649), .Q(
        \pe6/pvq [17]) );
  DRNQHSV4 \pe6/pe5/q_reg[16]  ( .D(n60070), .CK(clk), .RDN(n59650), .Q(
        \pe6/pvq [16]) );
  DRNQHSV4 \pe6/pe5/q_reg[14]  ( .D(n60033), .CK(clk), .RDN(n59650), .Q(
        \pe6/pvq [14]) );
  DRNQHSV4 \pe6/pe5/q_reg[12]  ( .D(pov5[12]), .CK(clk), .RDN(n59445), .Q(
        \pe6/pvq [12]) );
  DRNQHSV4 \pe6/pe5/q_reg[10]  ( .D(n60058), .CK(clk), .RDN(n59424), .Q(
        \pe6/pvq [10]) );
  DRNQHSV4 \pe6/pe5/q_reg[9]  ( .D(n60071), .CK(clk), .RDN(n59457), .Q(
        \pe6/pvq [9]) );
  DRNQHSV4 \pe6/pe5/q_reg[8]  ( .D(n60072), .CK(clk), .RDN(n59456), .Q(
        \pe6/pvq [8]) );
  DRNQHSV4 \pe6/pe5/q_reg[7]  ( .D(n60073), .CK(clk), .RDN(n59414), .Q(
        \pe6/pvq [7]) );
  DRNQHSV4 \pe6/pe5/q_reg[3]  ( .D(n60075), .CK(clk), .RDN(n59649), .Q(
        \pe6/pvq [3]) );
  DRNQHSV4 \pe6/pe5/q_reg[2]  ( .D(n60076), .CK(clk), .RDN(n59477), .Q(
        \pe6/pvq [2]) );
  DRNQHSV4 \pe6/pe6/q_reg[31]  ( .D(poh5[31]), .CK(clk), .RDN(n59452), .Q(
        \pe6/phq [31]) );
  DRNQHSV4 \pe6/pe6/q_reg[30]  ( .D(poh5[30]), .CK(clk), .RDN(n59430), .Q(
        \pe6/phq [30]) );
  DRNQHSV4 \pe6/pe6/q_reg[29]  ( .D(poh5[29]), .CK(clk), .RDN(n59436), .Q(
        \pe6/phq [29]) );
  DRNQHSV4 \pe6/pe6/q_reg[28]  ( .D(poh5[28]), .CK(clk), .RDN(n59510), .Q(
        \pe6/phq [28]) );
  DRNQHSV4 \pe6/pe6/q_reg[27]  ( .D(poh5[27]), .CK(clk), .RDN(n59435), .Q(
        \pe6/phq [27]) );
  DRNQHSV4 \pe6/pe6/q_reg[26]  ( .D(poh5[26]), .CK(clk), .RDN(n59442), .Q(
        \pe6/phq [26]) );
  DRNQHSV4 \pe6/pe6/q_reg[25]  ( .D(poh5[25]), .CK(clk), .RDN(n59405), .Q(
        \pe6/phq [25]) );
  DRNQHSV4 \pe6/pe6/q_reg[24]  ( .D(poh5[24]), .CK(clk), .RDN(n59439), .Q(
        \pe6/phq [24]) );
  DRNQHSV4 \pe6/pe6/q_reg[23]  ( .D(poh5[23]), .CK(clk), .RDN(n59924), .Q(
        \pe6/phq [23]) );
  DRNQHSV4 \pe6/pe6/q_reg[22]  ( .D(poh5[22]), .CK(clk), .RDN(n59443), .Q(
        \pe6/phq [22]) );
  DRNQHSV4 \pe6/pe6/q_reg[21]  ( .D(poh5[21]), .CK(clk), .RDN(n59410), .Q(
        \pe6/phq [21]) );
  DRNQHSV4 \pe6/pe6/q_reg[20]  ( .D(poh5[20]), .CK(clk), .RDN(n29729), .Q(
        \pe6/phq [20]) );
  DRNQHSV4 \pe6/pe6/q_reg[19]  ( .D(poh5[19]), .CK(clk), .RDN(n59493), .Q(
        \pe6/phq [19]) );
  DRNQHSV4 \pe6/pe6/q_reg[18]  ( .D(poh5[18]), .CK(clk), .RDN(n59468), .Q(
        \pe6/phq [18]) );
  DRNQHSV4 \pe6/pe6/q_reg[17]  ( .D(poh5[17]), .CK(clk), .RDN(n59494), .Q(
        \pe6/phq [17]) );
  DRNQHSV4 \pe6/pe6/q_reg[16]  ( .D(poh5[16]), .CK(clk), .RDN(n59414), .Q(
        \pe6/phq [16]) );
  DRNQHSV4 \pe6/pe6/q_reg[15]  ( .D(poh5[15]), .CK(clk), .RDN(n59432), .Q(
        \pe6/phq [15]) );
  DRNQHSV4 \pe6/pe6/q_reg[14]  ( .D(poh5[14]), .CK(clk), .RDN(n59456), .Q(
        \pe6/phq [14]) );
  DRNQHSV4 \pe6/pe6/q_reg[13]  ( .D(poh5[13]), .CK(clk), .RDN(n59454), .Q(
        \pe6/phq [13]) );
  DRNQHSV4 \pe6/pe6/q_reg[12]  ( .D(poh5[12]), .CK(clk), .RDN(n59457), .Q(
        \pe6/phq [12]) );
  DRNQHSV4 \pe6/pe6/q_reg[11]  ( .D(poh5[11]), .CK(clk), .RDN(n59456), .Q(
        \pe6/phq [11]) );
  DRNQHSV4 \pe6/pe6/q_reg[10]  ( .D(poh5[10]), .CK(clk), .RDN(n59440), .Q(
        \pe6/phq [10]) );
  DRNQHSV4 \pe6/pe6/q_reg[9]  ( .D(poh5[9]), .CK(clk), .RDN(n59472), .Q(
        \pe6/phq [9]) );
  DRNQHSV4 \pe6/pe6/q_reg[8]  ( .D(poh5[8]), .CK(clk), .RDN(n59460), .Q(
        \pe6/phq [8]) );
  DRNQHSV4 \pe6/pe6/q_reg[7]  ( .D(poh5[7]), .CK(clk), .RDN(n59512), .Q(
        \pe6/phq [7]) );
  DRNQHSV4 \pe6/pe6/q_reg[6]  ( .D(poh5[6]), .CK(clk), .RDN(n59655), .Q(
        \pe6/phq [6]) );
  DRNQHSV4 \pe6/pe6/q_reg[5]  ( .D(poh5[5]), .CK(clk), .RDN(n59924), .Q(
        \pe6/phq [5]) );
  DRNQHSV4 \pe6/pe6/q_reg[4]  ( .D(poh5[4]), .CK(clk), .RDN(n59446), .Q(
        \pe6/phq [4]) );
  DRNQHSV4 \pe6/pe6/q_reg[3]  ( .D(poh5[3]), .CK(clk), .RDN(n59435), .Q(
        \pe6/phq [3]) );
  DRNQHSV4 \pe6/pe6/q_reg[2]  ( .D(poh5[2]), .CK(clk), .RDN(n59435), .Q(
        \pe6/phq [2]) );
  DRNQHSV4 \pe6/pe6/q_reg[1]  ( .D(poh5[1]), .CK(clk), .RDN(n59431), .Q(
        \pe6/phq [1]) );
  DRNQHSV4 \pe6/pe7/q_reg  ( .D(n39730), .CK(clk), .RDN(n59397), .Q(\pe6/ctrq ) );
  DRNQHSV4 \pe6/pe12/q_reg[32]  ( .D(n59687), .CK(clk), .RDN(n59925), .Q(
        \pe6/bq[1] ) );
  DRNQHSV4 \pe6/pe12/q_reg[31]  ( .D(n59539), .CK(clk), .RDN(n59502), .Q(
        \pe6/bq[2] ) );
  DRNQHSV4 \pe6/pe12/q_reg[30]  ( .D(n59913), .CK(clk), .RDN(n59466), .Q(
        \pe6/bq[3] ) );
  DRNQHSV4 \pe6/pe12/q_reg[29]  ( .D(n59912), .CK(clk), .RDN(n29732), .Q(
        \pe6/bq[4] ) );
  DRNQHSV4 \pe6/pe12/q_reg[28]  ( .D(n59911), .CK(clk), .RDN(n59655), .Q(
        \pe6/bq[5] ) );
  DRNQHSV4 \pe6/pe12/q_reg[27]  ( .D(n59910), .CK(clk), .RDN(n59424), .Q(
        \pe6/bq[6] ) );
  DRNQHSV4 \pe6/pe12/q_reg[26]  ( .D(n59909), .CK(clk), .RDN(n29730), .Q(
        \pe6/bq[7] ) );
  DRNQHSV4 \pe6/pe12/q_reg[25]  ( .D(n59907), .CK(clk), .RDN(n59433), .Q(
        \pe6/bq[8] ) );
  DRNQHSV4 \pe6/pe12/q_reg[24]  ( .D(n59908), .CK(clk), .RDN(n29733), .Q(
        \pe6/bq[9] ) );
  DRNQHSV4 \pe6/pe12/q_reg[23]  ( .D(n59906), .CK(clk), .RDN(n59405), .Q(
        \pe6/bq[10] ) );
  DRNQHSV4 \pe6/pe12/q_reg[22]  ( .D(n59904), .CK(clk), .RDN(n59925), .Q(
        \pe6/bq[11] ) );
  DRNQHSV4 \pe6/pe12/q_reg[21]  ( .D(n59899), .CK(clk), .RDN(n59431), .Q(
        \pe6/bq[12] ) );
  DRNQHSV4 \pe6/pe12/q_reg[20]  ( .D(n59901), .CK(clk), .RDN(n59401), .Q(
        \pe6/bq[13] ) );
  DRNQHSV4 \pe6/pe12/q_reg[19]  ( .D(n59538), .CK(clk), .RDN(n29732), .Q(
        \pe6/bq[14] ) );
  DRNQHSV4 \pe6/pe12/q_reg[18]  ( .D(n59900), .CK(clk), .RDN(n59446), .Q(
        \pe6/bq[15] ) );
  DRNQHSV4 \pe6/pe12/q_reg[17]  ( .D(n59898), .CK(clk), .RDN(n29731), .Q(
        \pe6/bq[16] ) );
  DRNQHSV4 \pe6/pe12/q_reg[16]  ( .D(n59890), .CK(clk), .RDN(n59653), .Q(
        \pe6/bq[17] ) );
  DRNQHSV4 \pe6/pe12/q_reg[15]  ( .D(n59885), .CK(clk), .RDN(n59399), .Q(
        \pe6/bq[18] ) );
  DRNQHSV4 \pe6/pe12/q_reg[14]  ( .D(n59889), .CK(clk), .RDN(n59473), .Q(
        \pe6/bq[19] ) );
  DRNQHSV4 \pe6/pe12/q_reg[13]  ( .D(n59888), .CK(clk), .RDN(n59399), .Q(
        \pe6/bq[20] ) );
  DRNQHSV4 \pe6/pe12/q_reg[12]  ( .D(n59886), .CK(clk), .RDN(n59481), .Q(
        \pe6/bq[21] ) );
  DRNQHSV4 \pe6/pe12/q_reg[11]  ( .D(n59884), .CK(clk), .RDN(n59484), .Q(
        \pe6/bq[22] ) );
  DRNQHSV4 \pe6/pe12/q_reg[10]  ( .D(n59887), .CK(clk), .RDN(n59409), .Q(
        \pe6/bq[23] ) );
  DRNQHSV4 \pe6/pe12/q_reg[9]  ( .D(n59874), .CK(clk), .RDN(n59922), .Q(
        \pe6/bq[24] ) );
  DRNQHSV4 \pe6/pe12/q_reg[8]  ( .D(n59877), .CK(clk), .RDN(n59467), .Q(
        \pe6/bq[25] ) );
  DRNQHSV4 \pe6/pe12/q_reg[7]  ( .D(n59875), .CK(clk), .RDN(n59656), .Q(
        \pe6/bq[26] ) );
  DRNQHSV4 \pe6/pe12/q_reg[6]  ( .D(n59876), .CK(clk), .RDN(n59460), .Q(
        \pe6/bq[27] ) );
  DRNQHSV4 \pe6/pe12/q_reg[5]  ( .D(n59873), .CK(clk), .RDN(n59430), .Q(
        \pe6/bq[28] ) );
  DRNQHSV4 \pe6/pe12/q_reg[4]  ( .D(n59872), .CK(clk), .RDN(n59452), .Q(
        \pe6/bq[29] ) );
  DRNQHSV4 \pe6/pe12/q_reg[3]  ( .D(n59870), .CK(clk), .RDN(n59484), .Q(
        \pe6/bq[30] ) );
  DRNQHSV4 \pe6/pe12/q_reg[2]  ( .D(n59868), .CK(clk), .RDN(n59447), .Q(
        \pe6/bq[31] ) );
  DRNQHSV4 \pe6/pe12/q_reg[1]  ( .D(n59867), .CK(clk), .RDN(n59924), .Q(
        \pe6/bq[32] ) );
  DRNQHSV4 \pe6/pe13/q_reg  ( .D(\pe6/ti_1t ), .CK(clk), .RDN(n59448), .Q(
        \pe6/ti_1 ) );
  DRNQHSV4 \pe6/pe14/q_reg[2]  ( .D(n59038), .CK(clk), .RDN(n59465), .Q(
        \pe6/ti_7t [2]) );
  DRNQHSV4 \pe6/pe14/q_reg[4]  ( .D(n59670), .CK(clk), .RDN(n59649), .Q(
        \pe6/ti_7t [4]) );
  DRNQHSV1 \pe5/pe5/q_reg[4]  ( .D(n59578), .CK(clk), .RDN(n59401), .Q(
        \pe5/pvq [4]) );
  DRNQHSV1 \pe4/pe14/q_reg[31]  ( .D(n57900), .CK(clk), .RDN(n59925), .Q(
        \pe4/ti_7t [31]) );
  DRNQHSV1 \pe5/pe14/q_reg[29]  ( .D(n29777), .CK(clk), .RDN(n59460), .Q(
        \pe5/ti_7t [29]) );
  DRNQHSV2 \pe6/pe3/q_reg[31]  ( .D(bo5[2]), .CK(clk), .RDN(n59414), .Q(bo6[2]) );
  DRNQHSV2 \pe6/pe3/q_reg[19]  ( .D(bo5[14]), .CK(clk), .RDN(n29729), .Q(
        bo6[14]) );
  DRNQHSV2 \pe1/pe14/q_reg[29]  ( .D(n26467), .CK(clk), .RDN(n59925), .Q(
        \pe1/ti_7t [29]) );
  DRNQHSV1 \pe1/pe15/q_reg[30]  ( .D(n59389), .CK(clk), .RDN(n59442), .Q(
        ao1[3]) );
  DRNQHSV1 \pe1/pe15/q_reg[28]  ( .D(n59993), .CK(clk), .RDN(n59430), .Q(
        ao1[5]) );
  DRNQHSV1 \pe1/pe15/q_reg[27]  ( .D(n59992), .CK(clk), .RDN(n59424), .Q(
        ao1[6]) );
  DRNQHSV1 \pe1/pe15/q_reg[26]  ( .D(n54578), .CK(clk), .RDN(n59494), .Q(
        ao1[7]) );
  DRNQHSV1 \pe1/pe15/q_reg[25]  ( .D(n54904), .CK(clk), .RDN(n59512), .Q(
        ao1[8]) );
  DRNQHSV1 \pe1/pe15/q_reg[24]  ( .D(n59495), .CK(clk), .RDN(n59463), .Q(
        ao1[9]) );
  DRNQHSV1 \pe1/pe15/q_reg[23]  ( .D(n59991), .CK(clk), .RDN(n59654), .Q(
        ao1[10]) );
  DRNQHSV1 \pe1/pe15/q_reg[22]  ( .D(n59593), .CK(clk), .RDN(n59430), .Q(
        ao1[11]) );
  DRNQHSV1 \pe1/pe15/q_reg[20]  ( .D(n59990), .CK(clk), .RDN(n59462), .Q(
        ao1[13]) );
  DRNQHSV2 \pe1/pe15/q_reg[19]  ( .D(\pe1/aot [14]), .CK(clk), .RDN(n59494), 
        .Q(ao1[14]) );
  DRNQHSV1 \pe1/pe15/q_reg[18]  ( .D(n42132), .CK(clk), .RDN(rst), .Q(ao1[15])
         );
  DRNQHSV1 \pe1/pe15/q_reg[17]  ( .D(n59989), .CK(clk), .RDN(n59651), .Q(
        ao1[16]) );
  DRNQHSV1 \pe1/pe15/q_reg[16]  ( .D(n59988), .CK(clk), .RDN(n59459), .Q(
        ao1[17]) );
  DRNQHSV1 \pe1/pe15/q_reg[15]  ( .D(n59733), .CK(clk), .RDN(n59432), .Q(
        ao1[18]) );
  DRNQHSV1 \pe1/pe15/q_reg[13]  ( .D(n54669), .CK(clk), .RDN(n59449), .Q(
        ao1[20]) );
  DRNQHSV1 \pe1/pe15/q_reg[11]  ( .D(n54078), .CK(clk), .RDN(n59493), .Q(
        ao1[22]) );
  DRNQHSV1 \pe1/pe15/q_reg[10]  ( .D(n42255), .CK(clk), .RDN(n59491), .Q(
        ao1[23]) );
  DRNQHSV1 \pe1/pe15/q_reg[9]  ( .D(\pe1/aot [24]), .CK(clk), .RDN(n59483), 
        .Q(ao1[24]) );
  DRNQHSV1 \pe1/pe15/q_reg[8]  ( .D(n59589), .CK(clk), .RDN(n59429), .Q(
        ao1[25]) );
  DRNQHSV2 \pe1/pe15/q_reg[7]  ( .D(n41153), .CK(clk), .RDN(n59397), .Q(
        ao1[26]) );
  DRNQHSV1 \pe1/pe15/q_reg[6]  ( .D(n59986), .CK(clk), .RDN(n59439), .Q(
        ao1[27]) );
  DRNQHSV1 \pe1/pe15/q_reg[5]  ( .D(n40683), .CK(clk), .RDN(n59400), .Q(
        ao1[28]) );
  DRNQHSV1 \pe1/pe15/q_reg[4]  ( .D(n59385), .CK(clk), .RDN(n59479), .Q(
        ao1[29]) );
  DRNQHSV1 \pe1/pe15/q_reg[3]  ( .D(n59985), .CK(clk), .RDN(n59469), .Q(
        ao1[30]) );
  DRNQHSV1 \pe1/pe15/q_reg[2]  ( .D(n59376), .CK(clk), .RDN(n59439), .Q(
        ao1[31]) );
  DRNQHSV1 \pe1/pe16/q_reg[31]  ( .D(n59756), .CK(clk), .RDN(n59404), .Q(
        go1[2]) );
  DRNQHSV1 \pe1/pe16/q_reg[30]  ( .D(n55319), .CK(clk), .RDN(n59400), .Q(
        go1[3]) );
  DRNQHSV1 \pe1/pe16/q_reg[29]  ( .D(n55410), .CK(clk), .RDN(n59449), .Q(
        go1[4]) );
  DRNQHSV1 \pe1/pe16/q_reg[28]  ( .D(n55475), .CK(clk), .RDN(n59482), .Q(
        go1[5]) );
  DRNQHSV1 \pe1/pe16/q_reg[27]  ( .D(n55448), .CK(clk), .RDN(n59447), .Q(
        go1[6]) );
  DRNQHSV1 \pe1/pe16/q_reg[26]  ( .D(n59750), .CK(clk), .RDN(n59491), .Q(
        go1[7]) );
  DRNQHSV1 \pe1/pe16/q_reg[25]  ( .D(n55339), .CK(clk), .RDN(n59461), .Q(
        go1[8]) );
  DRNQHSV1 \pe1/pe16/q_reg[23]  ( .D(n55088), .CK(clk), .RDN(n59496), .Q(
        go1[10]) );
  DRNQHSV1 \pe1/pe16/q_reg[19]  ( .D(n54969), .CK(clk), .RDN(rst), .Q(go1[14])
         );
  DRNQHSV1 \pe1/pe16/q_reg[18]  ( .D(n48339), .CK(clk), .RDN(n59649), .Q(
        go1[15]) );
  DRNQHSV1 \pe1/pe16/q_reg[17]  ( .D(n42162), .CK(clk), .RDN(n59921), .Q(
        go1[16]) );
  DRNQHSV1 \pe1/pe16/q_reg[15]  ( .D(n42359), .CK(clk), .RDN(n59651), .Q(
        go1[18]) );
  DRNQHSV1 \pe1/pe16/q_reg[14]  ( .D(n59995), .CK(clk), .RDN(n59924), .Q(
        go1[19]) );
  DRNQHSV1 \pe1/pe16/q_reg[13]  ( .D(n41676), .CK(clk), .RDN(n59466), .Q(
        go1[20]) );
  DRNQHSV1 \pe1/pe16/q_reg[12]  ( .D(n54724), .CK(clk), .RDN(n59406), .Q(
        go1[21]) );
  DRNQHSV1 \pe1/pe16/q_reg[11]  ( .D(n54452), .CK(clk), .RDN(n59492), .Q(
        go1[22]) );
  DRNQHSV1 \pe1/pe16/q_reg[9]  ( .D(n53520), .CK(clk), .RDN(n59446), .Q(
        go1[24]) );
  DRNQHSV1 \pe1/pe16/q_reg[8]  ( .D(\pe1/got [25]), .CK(clk), .RDN(n59453), 
        .Q(go1[25]) );
  DRNQHSV1 \pe1/pe16/q_reg[7]  ( .D(n41689), .CK(clk), .RDN(n59399), .Q(
        go1[26]) );
  DRNQHSV1 \pe1/pe16/q_reg[6]  ( .D(n59374), .CK(clk), .RDN(n59413), .Q(
        go1[27]) );
  DRNQHSV1 \pe1/pe16/q_reg[5]  ( .D(n40873), .CK(clk), .RDN(n59402), .Q(
        go1[28]) );
  DRNQHSV1 \pe1/pe16/q_reg[4]  ( .D(n59994), .CK(clk), .RDN(n59436), .Q(
        go1[29]) );
  DRNQHSV1 \pe1/pe16/q_reg[3]  ( .D(n59394), .CK(clk), .RDN(n59433), .Q(
        go1[30]) );
  DRNQHSV1 \pe1/pe16/q_reg[1]  ( .D(n52831), .CK(clk), .RDN(n59484), .Q(
        go1[32]) );
  DRNQHSV2 \pe1/pe17/q_reg[29]  ( .D(\pe1/poht [29]), .CK(clk), .RDN(n29731), 
        .Q(poh1[29]) );
  DRNQHSV2 \pe1/pe17/q_reg[22]  ( .D(\pe1/poht [22]), .CK(clk), .RDN(n59397), 
        .Q(poh1[22]) );
  DRNQHSV2 \pe1/pe17/q_reg[6]  ( .D(\pe1/poht [6]), .CK(clk), .RDN(n59921), 
        .Q(poh1[6]) );
  DRNQHSV2 \pe1/pe17/q_reg[3]  ( .D(\pe1/poht [3]), .CK(clk), .RDN(n59490), 
        .Q(poh1[3]) );
  DRNQHSV2 \pe1/pe17/q_reg[1]  ( .D(\pe1/poht [1]), .CK(clk), .RDN(n59478), 
        .Q(poh1[1]) );
  DRNQHSV1 \pe2/pe15/q_reg[32]  ( .D(n59783), .CK(clk), .RDN(n59403), .Q(
        ao2[1]) );
  DRNQHSV1 \pe2/pe15/q_reg[31]  ( .D(\pe2/aot [2]), .CK(clk), .RDN(n59401), 
        .Q(ao2[2]) );
  DRNQHSV1 \pe2/pe15/q_reg[30]  ( .D(n59792), .CK(clk), .RDN(n59413), .Q(
        ao2[3]) );
  DRNQHSV1 \pe2/pe15/q_reg[29]  ( .D(n59978), .CK(clk), .RDN(n59653), .Q(
        ao2[4]) );
  DRNQHSV1 \pe2/pe15/q_reg[28]  ( .D(n59499), .CK(clk), .RDN(n59484), .Q(
        ao2[5]) );
  DRNQHSV1 \pe2/pe15/q_reg[27]  ( .D(n52456), .CK(clk), .RDN(n59468), .Q(
        ao2[6]) );
  DRNQHSV1 \pe2/pe15/q_reg[26]  ( .D(n59633), .CK(clk), .RDN(n59413), .Q(
        ao2[7]) );
  DRNQHSV1 \pe2/pe15/q_reg[25]  ( .D(n52951), .CK(clk), .RDN(n59439), .Q(
        ao2[8]) );
  DRNQHSV1 \pe2/pe15/q_reg[24]  ( .D(n59768), .CK(clk), .RDN(n59471), .Q(
        ao2[9]) );
  DRNQHSV1 \pe2/pe15/q_reg[23]  ( .D(n59977), .CK(clk), .RDN(n59924), .Q(
        ao2[10]) );
  DRNQHSV1 \pe2/pe15/q_reg[22]  ( .D(n59976), .CK(clk), .RDN(n59925), .Q(
        ao2[11]) );
  DRNQHSV1 \pe2/pe15/q_reg[21]  ( .D(\pe2/aot [12]), .CK(clk), .RDN(n59461), 
        .Q(ao2[12]) );
  DRNQHSV1 \pe2/pe15/q_reg[20]  ( .D(n59975), .CK(clk), .RDN(n59468), .Q(
        ao2[13]) );
  DRNQHSV1 \pe2/pe15/q_reg[19]  ( .D(n59636), .CK(clk), .RDN(n59468), .Q(
        ao2[14]) );
  DRNQHSV1 \pe2/pe15/q_reg[18]  ( .D(n59974), .CK(clk), .RDN(n59405), .Q(
        ao2[15]) );
  DRNQHSV1 \pe2/pe15/q_reg[17]  ( .D(n59973), .CK(clk), .RDN(n59403), .Q(
        ao2[16]) );
  DRNQHSV1 \pe2/pe15/q_reg[16]  ( .D(\pe2/aot [17]), .CK(clk), .RDN(n59413), 
        .Q(ao2[17]) );
  DRNQHSV1 \pe2/pe15/q_reg[15]  ( .D(n59358), .CK(clk), .RDN(n59477), .Q(
        ao2[18]) );
  DRNQHSV1 \pe2/pe15/q_reg[14]  ( .D(\pe2/aot [19]), .CK(clk), .RDN(n59448), 
        .Q(ao2[19]) );
  DRNQHSV1 \pe2/pe15/q_reg[13]  ( .D(n59587), .CK(clk), .RDN(n59447), .Q(
        ao2[20]) );
  DRNQHSV1 \pe2/pe15/q_reg[12]  ( .D(n59758), .CK(clk), .RDN(n59465), .Q(
        ao2[21]) );
  DRNQHSV1 \pe2/pe15/q_reg[11]  ( .D(\pe2/aot [22]), .CK(clk), .RDN(n59490), 
        .Q(ao2[22]) );
  DRNQHSV1 \pe2/pe15/q_reg[9]  ( .D(n59972), .CK(clk), .RDN(n59465), .Q(
        ao2[24]) );
  DRNQHSV1 \pe2/pe15/q_reg[8]  ( .D(n59971), .CK(clk), .RDN(n59658), .Q(
        ao2[25]) );
  DRNQHSV1 \pe2/pe15/q_reg[7]  ( .D(n59970), .CK(clk), .RDN(n59465), .Q(
        ao2[26]) );
  DRNQHSV1 \pe2/pe15/q_reg[5]  ( .D(n59759), .CK(clk), .RDN(n29730), .Q(
        ao2[28]) );
  DRNQHSV1 \pe2/pe15/q_reg[4]  ( .D(n59588), .CK(clk), .RDN(n59429), .Q(
        ao2[29]) );
  DRNQHSV1 \pe2/pe15/q_reg[3]  ( .D(n59969), .CK(clk), .RDN(n59924), .Q(
        ao2[30]) );
  DRNQHSV1 \pe2/pe15/q_reg[2]  ( .D(n59968), .CK(clk), .RDN(n59465), .Q(
        ao2[31]) );
  DRNQHSV1 \pe2/pe15/q_reg[1]  ( .D(n59582), .CK(clk), .RDN(n59465), .Q(
        ao2[32]) );
  DRNQHSV1 \pe2/pe16/q_reg[32]  ( .D(n59767), .CK(clk), .RDN(n59442), .Q(
        go2[1]) );
  DRNQHSV1 \pe2/pe16/q_reg[31]  ( .D(n51932), .CK(clk), .RDN(n59445), .Q(
        go2[2]) );
  DRNQHSV1 \pe2/pe16/q_reg[29]  ( .D(n59984), .CK(clk), .RDN(n59442), .Q(
        go2[4]) );
  DRNQHSV1 \pe2/pe16/q_reg[28]  ( .D(n59778), .CK(clk), .RDN(n59469), .Q(
        go2[5]) );
  DRNQHSV1 \pe2/pe16/q_reg[27]  ( .D(n59777), .CK(clk), .RDN(n59416), .Q(
        go2[6]) );
  DRNQHSV1 \pe2/pe16/q_reg[26]  ( .D(n59757), .CK(clk), .RDN(n59457), .Q(
        go2[7]) );
  DRNQHSV1 \pe2/pe16/q_reg[25]  ( .D(n59371), .CK(clk), .RDN(n59470), .Q(
        go2[8]) );
  DRNQHSV1 \pe2/pe16/q_reg[24]  ( .D(n52052), .CK(clk), .RDN(n59459), .Q(
        go2[9]) );
  DRNQHSV1 \pe2/pe16/q_reg[23]  ( .D(\pe2/got [10]), .CK(clk), .RDN(n59478), 
        .Q(go2[10]) );
  DRNQHSV1 \pe2/pe16/q_reg[22]  ( .D(n51892), .CK(clk), .RDN(n59431), .Q(
        go2[11]) );
  DRNQHSV1 \pe2/pe16/q_reg[21]  ( .D(n52172), .CK(clk), .RDN(n59481), .Q(
        go2[12]) );
  DRNQHSV1 \pe2/pe16/q_reg[20]  ( .D(n59375), .CK(clk), .RDN(n59451), .Q(
        go2[13]) );
  DRNQHSV1 \pe2/pe16/q_reg[19]  ( .D(n59354), .CK(clk), .RDN(n59430), .Q(
        go2[14]) );
  DRNQHSV1 \pe2/pe16/q_reg[18]  ( .D(n52051), .CK(clk), .RDN(n59469), .Q(
        go2[15]) );
  DRNQHSV1 \pe2/pe16/q_reg[17]  ( .D(n51796), .CK(clk), .RDN(n59407), .Q(
        go2[16]) );
  DRNQHSV1 \pe2/pe16/q_reg[16]  ( .D(n59983), .CK(clk), .RDN(n59473), .Q(
        go2[17]) );
  DRNQHSV1 \pe2/pe16/q_reg[15]  ( .D(n44712), .CK(clk), .RDN(n59469), .Q(
        go2[18]) );
  DRNQHSV1 \pe2/pe16/q_reg[14]  ( .D(n59982), .CK(clk), .RDN(n59430), .Q(
        go2[19]) );
  DRNQHSV1 \pe2/pe16/q_reg[13]  ( .D(n59685), .CK(clk), .RDN(n59473), .Q(
        go2[20]) );
  DRNQHSV1 \pe2/pe16/q_reg[12]  ( .D(n52167), .CK(clk), .RDN(n59448), .Q(
        go2[21]) );
  DRNQHSV1 \pe2/pe16/q_reg[11]  ( .D(n43925), .CK(clk), .RDN(n59447), .Q(
        go2[22]) );
  DRNQHSV1 \pe2/pe16/q_reg[9]  ( .D(n59584), .CK(clk), .RDN(n59478), .Q(
        go2[24]) );
  DRNQHSV1 \pe2/pe16/q_reg[8]  ( .D(n44711), .CK(clk), .RDN(n59400), .Q(
        go2[25]) );
  DRNQHSV1 \pe2/pe16/q_reg[7]  ( .D(n38778), .CK(clk), .RDN(n59479), .Q(
        go2[26]) );
  DRNQHSV1 \pe2/pe16/q_reg[6]  ( .D(n59981), .CK(clk), .RDN(n59453), .Q(
        go2[27]) );
  DRNQHSV2 \pe2/pe16/q_reg[5]  ( .D(n38327), .CK(clk), .RDN(n59502), .Q(
        go2[28]) );
  DRNQHSV1 \pe2/pe16/q_reg[4]  ( .D(n59635), .CK(clk), .RDN(n59418), .Q(
        go2[29]) );
  DRNQHSV1 \pe2/pe16/q_reg[3]  ( .D(n59980), .CK(clk), .RDN(n59491), .Q(
        go2[30]) );
  DRNQHSV1 \pe2/pe16/q_reg[2]  ( .D(n59979), .CK(clk), .RDN(n59477), .Q(
        go2[31]) );
  DRNQHSV1 \pe2/pe16/q_reg[1]  ( .D(n47997), .CK(clk), .RDN(n59424), .Q(
        go2[32]) );
  DRNQHSV2 \pe2/pe17/q_reg[31]  ( .D(\pe2/poht [31]), .CK(clk), .RDN(n59473), 
        .Q(poh2[31]) );
  DRNQHSV2 \pe2/pe17/q_reg[29]  ( .D(\pe2/poht [29]), .CK(clk), .RDN(n59408), 
        .Q(poh2[29]) );
  DRNQHSV1 \pe2/pe17/q_reg[28]  ( .D(\pe2/poht [28]), .CK(clk), .RDN(n59478), 
        .Q(poh2[28]) );
  DRNQHSV2 \pe2/pe17/q_reg[27]  ( .D(\pe2/poht [27]), .CK(clk), .RDN(n59470), 
        .Q(poh2[27]) );
  DRNQHSV1 \pe2/pe17/q_reg[26]  ( .D(\pe2/poht [26]), .CK(clk), .RDN(n59924), 
        .Q(poh2[26]) );
  DRNQHSV2 \pe2/pe17/q_reg[25]  ( .D(\pe2/poht [25]), .CK(clk), .RDN(n59480), 
        .Q(poh2[25]) );
  DRNQHSV2 \pe2/pe17/q_reg[14]  ( .D(\pe2/poht [14]), .CK(clk), .RDN(n59449), 
        .Q(poh2[14]) );
  DRNQHSV2 \pe2/pe17/q_reg[7]  ( .D(\pe2/poht [7]), .CK(clk), .RDN(n59657), 
        .Q(poh2[7]) );
  DRNQHSV2 \pe2/pe17/q_reg[4]  ( .D(\pe2/poht [4]), .CK(clk), .RDN(n59446), 
        .Q(poh2[4]) );
  DRNQHSV2 \pe2/pe17/q_reg[3]  ( .D(\pe2/poht [3]), .CK(clk), .RDN(n59460), 
        .Q(poh2[3]) );
  DRNQHSV1 \pe3/pe15/q_reg[32]  ( .D(n59511), .CK(clk), .RDN(n59471), .Q(
        ao3[1]) );
  DRNQHSV1 \pe3/pe15/q_reg[31]  ( .D(n59961), .CK(clk), .RDN(n59458), .Q(
        ao3[2]) );
  DRNQHSV1 \pe3/pe15/q_reg[30]  ( .D(n56434), .CK(clk), .RDN(n59419), .Q(
        ao3[3]) );
  DRNQHSV1 \pe3/pe15/q_reg[29]  ( .D(n59646), .CK(clk), .RDN(n59408), .Q(
        ao3[4]) );
  DRNQHSV1 \pe3/pe15/q_reg[28]  ( .D(n59816), .CK(clk), .RDN(n59437), .Q(
        ao3[5]) );
  DRNQHSV1 \pe3/pe15/q_reg[27]  ( .D(\pe3/aot [6]), .CK(clk), .RDN(n59453), 
        .Q(ao3[6]) );
  DRNQHSV1 \pe3/pe15/q_reg[26]  ( .D(n59627), .CK(clk), .RDN(n59407), .Q(
        ao3[7]) );
  DRNQHSV1 \pe3/pe15/q_reg[25]  ( .D(\pe3/aot [8]), .CK(clk), .RDN(n59433), 
        .Q(ao3[8]) );
  DRNQHSV1 \pe3/pe15/q_reg[24]  ( .D(n59808), .CK(clk), .RDN(n59400), .Q(
        ao3[9]) );
  DRNQHSV1 \pe3/pe15/q_reg[23]  ( .D(n59960), .CK(clk), .RDN(n59442), .Q(
        ao3[10]) );
  DRNQHSV1 \pe3/pe15/q_reg[22]  ( .D(n59623), .CK(clk), .RDN(n59417), .Q(
        ao3[11]) );
  DRNQHSV1 \pe3/pe15/q_reg[21]  ( .D(n59959), .CK(clk), .RDN(n59458), .Q(
        ao3[12]) );
  DRNQHSV1 \pe3/pe15/q_reg[20]  ( .D(\pe3/aot [13]), .CK(clk), .RDN(n59412), 
        .Q(ao3[13]) );
  DRNQHSV1 \pe3/pe15/q_reg[19]  ( .D(\pe3/aot [14]), .CK(clk), .RDN(n29730), 
        .Q(ao3[14]) );
  DRNQHSV1 \pe3/pe15/q_reg[18]  ( .D(\pe3/aot [15]), .CK(clk), .RDN(n59449), 
        .Q(ao3[15]) );
  DRNQHSV1 \pe3/pe15/q_reg[17]  ( .D(n45645), .CK(clk), .RDN(n59492), .Q(
        ao3[16]) );
  DRNQHSV1 \pe3/pe15/q_reg[16]  ( .D(n59344), .CK(clk), .RDN(n59476), .Q(
        ao3[17]) );
  DRNQHSV1 \pe3/pe15/q_reg[15]  ( .D(n42950), .CK(clk), .RDN(n59451), .Q(
        ao3[18]) );
  DRNQHSV1 \pe3/pe15/q_reg[14]  ( .D(n56464), .CK(clk), .RDN(n59432), .Q(
        ao3[19]) );
  DRNQHSV1 \pe3/pe15/q_reg[13]  ( .D(n56204), .CK(clk), .RDN(n59411), .Q(
        ao3[20]) );
  DRNQHSV1 \pe3/pe15/q_reg[12]  ( .D(\pe3/aot [21]), .CK(clk), .RDN(n59649), 
        .Q(ao3[21]) );
  DRNQHSV1 \pe3/pe15/q_reg[11]  ( .D(n59618), .CK(clk), .RDN(n59922), .Q(
        ao3[22]) );
  DRNQHSV1 \pe3/pe15/q_reg[10]  ( .D(n59612), .CK(clk), .RDN(n59451), .Q(
        ao3[23]) );
  DRNQHSV1 \pe3/pe15/q_reg[9]  ( .D(\pe3/aot [24]), .CK(clk), .RDN(n59502), 
        .Q(ao3[24]) );
  DRNQHSV1 \pe3/pe15/q_reg[8]  ( .D(n59368), .CK(clk), .RDN(n59476), .Q(
        ao3[25]) );
  DRNQHSV1 \pe3/pe15/q_reg[7]  ( .D(n59610), .CK(clk), .RDN(n59413), .Q(
        ao3[26]) );
  DRNQHSV1 \pe3/pe15/q_reg[6]  ( .D(n59622), .CK(clk), .RDN(n59457), .Q(
        ao3[27]) );
  DRNQHSV1 \pe3/pe15/q_reg[5]  ( .D(n59809), .CK(clk), .RDN(n59415), .Q(
        ao3[28]) );
  DRNQHSV1 \pe3/pe15/q_reg[4]  ( .D(n48500), .CK(clk), .RDN(n59429), .Q(
        ao3[29]) );
  DRNQHSV1 \pe3/pe15/q_reg[3]  ( .D(n59609), .CK(clk), .RDN(n59439), .Q(
        ao3[30]) );
  DRNQHSV1 \pe3/pe15/q_reg[2]  ( .D(n59608), .CK(clk), .RDN(n59453), .Q(
        ao3[31]) );
  DRNQHSV1 \pe3/pe15/q_reg[1]  ( .D(n59614), .CK(clk), .RDN(n59437), .Q(
        ao3[32]) );
  DRNQHSV1 \pe3/pe16/q_reg[32]  ( .D(\pe3/got [1]), .CK(clk), .RDN(n59453), 
        .Q(go3[1]) );
  DRNQHSV1 \pe3/pe16/q_reg[31]  ( .D(n59807), .CK(clk), .RDN(n59476), .Q(
        go3[2]) );
  DRNQHSV1 \pe3/pe16/q_reg[30]  ( .D(n59356), .CK(clk), .RDN(n59494), .Q(
        go3[3]) );
  DRNQHSV1 \pe3/pe16/q_reg[29]  ( .D(n56684), .CK(clk), .RDN(n59659), .Q(
        go3[4]) );
  DRNQHSV1 \pe3/pe16/q_reg[28]  ( .D(n59799), .CK(clk), .RDN(n59416), .Q(
        go3[5]) );
  DRNQHSV1 \pe3/pe16/q_reg[27]  ( .D(n56779), .CK(clk), .RDN(n59453), .Q(
        go3[6]) );
  DRNQHSV1 \pe3/pe16/q_reg[26]  ( .D(n59647), .CK(clk), .RDN(n59491), .Q(
        go3[7]) );
  DRNQHSV1 \pe3/pe16/q_reg[25]  ( .D(n56855), .CK(clk), .RDN(n59476), .Q(
        go3[8]) );
  DRNQHSV1 \pe3/pe16/q_reg[24]  ( .D(n59645), .CK(clk), .RDN(n59510), .Q(
        go3[9]) );
  DRNQHSV1 \pe3/pe16/q_reg[23]  ( .D(n59644), .CK(clk), .RDN(n59476), .Q(
        go3[10]) );
  DRNQHSV1 \pe3/pe16/q_reg[22]  ( .D(n59967), .CK(clk), .RDN(n59650), .Q(
        go3[11]) );
  DRNQHSV1 \pe3/pe16/q_reg[21]  ( .D(n59966), .CK(clk), .RDN(n59457), .Q(
        go3[12]) );
  DRNQHSV1 \pe3/pe16/q_reg[20]  ( .D(n56421), .CK(clk), .RDN(n29730), .Q(
        go3[13]) );
  DRNQHSV1 \pe3/pe16/q_reg[19]  ( .D(n56493), .CK(clk), .RDN(n29729), .Q(
        go3[14]) );
  DRNQHSV1 \pe3/pe16/q_reg[18]  ( .D(n59624), .CK(clk), .RDN(n29730), .Q(
        go3[15]) );
  DRNQHSV1 \pe3/pe16/q_reg[17]  ( .D(n49252), .CK(clk), .RDN(n59451), .Q(
        go3[16]) );
  DRNQHSV1 \pe3/pe16/q_reg[16]  ( .D(n56064), .CK(clk), .RDN(n59453), .Q(
        go3[17]) );
  DRNQHSV1 \pe3/pe16/q_reg[15]  ( .D(n43374), .CK(clk), .RDN(n29729), .Q(
        go3[18]) );
  DRNQHSV1 \pe3/pe16/q_reg[14]  ( .D(n59965), .CK(clk), .RDN(n59476), .Q(
        go3[19]) );
  DRNQHSV1 \pe3/pe16/q_reg[13]  ( .D(n45581), .CK(clk), .RDN(n59402), .Q(
        go3[20]) );
  DRNQHSV1 \pe3/pe16/q_reg[12]  ( .D(n43262), .CK(clk), .RDN(n59451), .Q(
        go3[21]) );
  DRNQHSV1 \pe3/pe16/q_reg[11]  ( .D(n55821), .CK(clk), .RDN(n29733), .Q(
        go3[22]) );
  DRNQHSV1 \pe3/pe16/q_reg[10]  ( .D(n42673), .CK(clk), .RDN(n59442), .Q(
        go3[23]) );
  DRNQHSV1 \pe3/pe16/q_reg[9]  ( .D(n59617), .CK(clk), .RDN(n59411), .Q(
        go3[24]) );
  DRNQHSV1 \pe3/pe16/q_reg[8]  ( .D(n59384), .CK(clk), .RDN(n59434), .Q(
        go3[25]) );
  DRNQHSV1 \pe3/pe16/q_reg[7]  ( .D(n59616), .CK(clk), .RDN(n59491), .Q(
        go3[26]) );
  DRNQHSV1 \pe3/pe16/q_reg[6]  ( .D(n37516), .CK(clk), .RDN(n59405), .Q(
        go3[27]) );
  DRNQHSV1 \pe3/pe16/q_reg[3]  ( .D(n59347), .CK(clk), .RDN(n59510), .Q(
        go3[30]) );
  DRNQHSV1 \pe3/pe16/q_reg[2]  ( .D(n45755), .CK(clk), .RDN(n59424), .Q(
        go3[31]) );
  DRNQHSV1 \pe3/pe16/q_reg[1]  ( .D(n59962), .CK(clk), .RDN(n59458), .Q(
        go3[32]) );
  DRNQHSV1 \pe3/pe17/q_reg[27]  ( .D(\pe3/poht [27]), .CK(clk), .RDN(n59425), 
        .Q(poh3[27]) );
  DRNQHSV1 \pe3/pe17/q_reg[14]  ( .D(\pe3/poht [14]), .CK(clk), .RDN(n59436), 
        .Q(poh3[14]) );
  DRNQHSV2 \pe3/pe17/q_reg[12]  ( .D(\pe3/poht [12]), .CK(clk), .RDN(n59437), 
        .Q(poh3[12]) );
  DRNQHSV2 \pe3/pe17/q_reg[11]  ( .D(\pe3/poht [11]), .CK(clk), .RDN(n59438), 
        .Q(poh3[11]) );
  DRNQHSV1 \pe3/pe17/q_reg[10]  ( .D(\pe3/poht [10]), .CK(clk), .RDN(n59925), 
        .Q(poh3[10]) );
  DRNQHSV1 \pe3/pe17/q_reg[9]  ( .D(\pe3/poht [9]), .CK(clk), .RDN(n59418), 
        .Q(poh3[9]) );
  DRNQHSV1 \pe3/pe17/q_reg[2]  ( .D(\pe3/poht [2]), .CK(clk), .RDN(n59454), 
        .Q(poh3[2]) );
  DRNQHSV1 \pe4/pe15/q_reg[32]  ( .D(\pe4/aot [1]), .CK(clk), .RDN(n59443), 
        .Q(ao4[1]) );
  DRNQHSV1 \pe4/pe15/q_reg[31]  ( .D(\pe4/aot [2]), .CK(clk), .RDN(n29730), 
        .Q(ao4[2]) );
  DRNQHSV1 \pe4/pe15/q_reg[30]  ( .D(n59954), .CK(clk), .RDN(n59925), .Q(
        ao4[3]) );
  DRNQHSV1 \pe4/pe15/q_reg[28]  ( .D(n59831), .CK(clk), .RDN(n59482), .Q(
        ao4[5]) );
  DRNQHSV1 \pe4/pe15/q_reg[27]  ( .D(n59352), .CK(clk), .RDN(n59472), .Q(
        ao4[6]) );
  DRNQHSV1 \pe4/pe15/q_reg[26]  ( .D(n59632), .CK(clk), .RDN(n59417), .Q(
        ao4[7]) );
  DRNQHSV1 \pe4/pe15/q_reg[25]  ( .D(n59668), .CK(clk), .RDN(n59921), .Q(
        ao4[8]) );
  DRNQHSV1 \pe4/pe15/q_reg[24]  ( .D(\pe4/aot [9]), .CK(clk), .RDN(n59410), 
        .Q(ao4[9]) );
  DRNQHSV1 \pe4/pe15/q_reg[23]  ( .D(n47718), .CK(clk), .RDN(n59452), .Q(
        ao4[10]) );
  DRNQHSV1 \pe4/pe15/q_reg[22]  ( .D(n59683), .CK(clk), .RDN(n59491), .Q(
        ao4[11]) );
  DRNQHSV2 \pe4/pe15/q_reg[21]  ( .D(n59343), .CK(clk), .RDN(n59473), .Q(
        ao4[12]) );
  DRNQHSV1 \pe4/pe15/q_reg[20]  ( .D(n59857), .CK(clk), .RDN(n59456), .Q(
        ao4[13]) );
  DRNQHSV1 \pe4/pe15/q_reg[19]  ( .D(\pe4/aot [14]), .CK(clk), .RDN(n59418), 
        .Q(ao4[14]) );
  DRNQHSV1 \pe4/pe15/q_reg[18]  ( .D(n59953), .CK(clk), .RDN(n59440), .Q(
        ao4[15]) );
  DRNQHSV1 \pe4/pe15/q_reg[17]  ( .D(n59952), .CK(clk), .RDN(n59462), .Q(
        ao4[16]) );
  DRNQHSV1 \pe4/pe15/q_reg[16]  ( .D(\pe4/aot [17]), .CK(clk), .RDN(n59492), 
        .Q(ao4[17]) );
  DRNQHSV1 \pe4/pe15/q_reg[15]  ( .D(n59605), .CK(clk), .RDN(n59656), .Q(
        ao4[18]) );
  DRNQHSV1 \pe4/pe15/q_reg[12]  ( .D(n59951), .CK(clk), .RDN(n59406), .Q(
        ao4[21]) );
  DRNQHSV1 \pe4/pe15/q_reg[11]  ( .D(\pe4/aot [22]), .CK(clk), .RDN(n59465), 
        .Q(ao4[22]) );
  DRNQHSV1 \pe4/pe15/q_reg[10]  ( .D(n34022), .CK(clk), .RDN(n59433), .Q(
        ao4[23]) );
  DRNQHSV1 \pe4/pe15/q_reg[9]  ( .D(n59388), .CK(clk), .RDN(n59494), .Q(
        ao4[24]) );
  DRNQHSV1 \pe4/pe15/q_reg[8]  ( .D(n59838), .CK(clk), .RDN(n59503), .Q(
        ao4[25]) );
  DRNQHSV1 \pe4/pe15/q_reg[6]  ( .D(n59598), .CK(clk), .RDN(n59502), .Q(
        ao4[27]) );
  DRNQHSV1 \pe4/pe15/q_reg[5]  ( .D(n59390), .CK(clk), .RDN(n59407), .Q(
        ao4[28]) );
  DRNQHSV1 \pe4/pe15/q_reg[4]  ( .D(n59834), .CK(clk), .RDN(n59429), .Q(
        ao4[29]) );
  DRNQHSV1 \pe4/pe15/q_reg[3]  ( .D(n59383), .CK(clk), .RDN(n59429), .Q(
        ao4[30]) );
  DRNQHSV1 \pe4/pe15/q_reg[2]  ( .D(n59523), .CK(clk), .RDN(n59411), .Q(
        ao4[31]) );
  DRNQHSV1 \pe4/pe15/q_reg[1]  ( .D(n59485), .CK(clk), .RDN(n59429), .Q(
        ao4[32]) );
  DRNQHSV1 \pe4/pe16/q_reg[32]  ( .D(n59958), .CK(clk), .RDN(n59432), .Q(
        go4[1]) );
  DRNQHSV1 \pe4/pe16/q_reg[31]  ( .D(n59346), .CK(clk), .RDN(n59921), .Q(
        go4[2]) );
  DRNQHSV1 \pe4/pe16/q_reg[30]  ( .D(n58298), .CK(clk), .RDN(n59476), .Q(
        go4[3]) );
  DRNQHSV1 \pe4/pe16/q_reg[29]  ( .D(n59832), .CK(clk), .RDN(n59496), .Q(
        go4[4]) );
  DRNQHSV1 \pe4/pe16/q_reg[28]  ( .D(n57951), .CK(clk), .RDN(n59412), .Q(
        go4[5]) );
  DRNQHSV1 \pe4/pe16/q_reg[27]  ( .D(n58184), .CK(clk), .RDN(n59481), .Q(
        go4[6]) );
  DRNQHSV1 \pe4/pe16/q_reg[26]  ( .D(n59957), .CK(clk), .RDN(n59924), .Q(
        go4[7]) );
  DRNQHSV1 \pe4/pe16/q_reg[25]  ( .D(n58111), .CK(clk), .RDN(n59407), .Q(
        go4[8]) );
  DRNQHSV1 \pe4/pe16/q_reg[23]  ( .D(n59663), .CK(clk), .RDN(n29732), .Q(
        go4[10]) );
  DRNQHSV1 \pe4/pe16/q_reg[22]  ( .D(n58153), .CK(clk), .RDN(n59490), .Q(
        go4[11]) );
  DRNQHSV1 \pe4/pe16/q_reg[21]  ( .D(n59631), .CK(clk), .RDN(n59480), .Q(
        go4[12]) );
  DRNQHSV1 \pe4/pe16/q_reg[20]  ( .D(n59629), .CK(clk), .RDN(n59921), .Q(
        go4[13]) );
  DRNQHSV1 \pe4/pe16/q_reg[19]  ( .D(n59630), .CK(clk), .RDN(n59416), .Q(
        go4[14]) );
  DRNQHSV1 \pe4/pe16/q_reg[18]  ( .D(n59664), .CK(clk), .RDN(n59450), .Q(
        go4[15]) );
  DRNQHSV1 \pe4/pe16/q_reg[17]  ( .D(n59604), .CK(clk), .RDN(n29730), .Q(
        go4[16]) );
  DRNQHSV1 \pe4/pe16/q_reg[16]  ( .D(n59353), .CK(clk), .RDN(n59923), .Q(
        go4[17]) );
  DRNQHSV1 \pe4/pe16/q_reg[15]  ( .D(n59372), .CK(clk), .RDN(n59447), .Q(
        go4[18]) );
  DRNQHSV1 \pe4/pe16/q_reg[14]  ( .D(n59602), .CK(clk), .RDN(n59458), .Q(
        go4[19]) );
  DRNQHSV1 \pe4/pe16/q_reg[13]  ( .D(n59386), .CK(clk), .RDN(n59409), .Q(
        go4[20]) );
  DRNQHSV1 \pe4/pe16/q_reg[12]  ( .D(n59370), .CK(clk), .RDN(n59482), .Q(
        go4[21]) );
  DRNQHSV1 \pe4/pe16/q_reg[11]  ( .D(n59601), .CK(clk), .RDN(n59510), .Q(
        go4[22]) );
  DRNQHSV1 \pe4/pe16/q_reg[10]  ( .D(n59369), .CK(clk), .RDN(n59465), .Q(
        go4[23]) );
  DRNQHSV1 \pe4/pe16/q_reg[9]  ( .D(n59603), .CK(clk), .RDN(n59407), .Q(
        go4[24]) );
  DRNQHSV1 \pe4/pe16/q_reg[8]  ( .D(n59600), .CK(clk), .RDN(n59405), .Q(
        go4[25]) );
  DRNQHSV1 \pe4/pe16/q_reg[7]  ( .D(n59599), .CK(clk), .RDN(n59650), .Q(
        go4[26]) );
  DRNQHSV1 \pe4/pe16/q_reg[6]  ( .D(n59350), .CK(clk), .RDN(n59466), .Q(
        go4[27]) );
  DRNQHSV1 \pe4/pe16/q_reg[5]  ( .D(n57195), .CK(clk), .RDN(n59476), .Q(
        go4[28]) );
  DRNQHSV1 \pe4/pe16/q_reg[4]  ( .D(n59956), .CK(clk), .RDN(n59419), .Q(
        go4[29]) );
  DRNQHSV1 \pe4/pe16/q_reg[3]  ( .D(n59955), .CK(clk), .RDN(n59402), .Q(
        go4[30]) );
  DRNQHSV1 \pe4/pe16/q_reg[2]  ( .D(n59345), .CK(clk), .RDN(n59922), .Q(
        go4[31]) );
  DRNQHSV1 \pe4/pe16/q_reg[1]  ( .D(n47772), .CK(clk), .RDN(n59649), .Q(
        go4[32]) );
  DRNQHSV2 \pe4/pe17/q_reg[3]  ( .D(\pe4/poht [3]), .CK(clk), .RDN(n59418), 
        .Q(poh4[3]) );
  DRNQHSV2 \pe4/pe17/q_reg[1]  ( .D(\pe4/poht [1]), .CK(clk), .RDN(n59493), 
        .Q(poh4[1]) );
  DRNQHSV1 \pe5/pe15/q_reg[32]  ( .D(n59895), .CK(clk), .RDN(n59401), .Q(
        ao5[1]) );
  DRNQHSV1 \pe5/pe15/q_reg[31]  ( .D(n59866), .CK(clk), .RDN(n59415), .Q(
        ao5[2]) );
  DRNQHSV1 \pe5/pe15/q_reg[29]  ( .D(\pe5/aot [4]), .CK(clk), .RDN(n59419), 
        .Q(ao5[4]) );
  DRNQHSV1 \pe5/pe15/q_reg[28]  ( .D(n59945), .CK(clk), .RDN(n59432), .Q(
        ao5[5]) );
  DRNQHSV1 \pe5/pe15/q_reg[27]  ( .D(n53295), .CK(clk), .RDN(n59469), .Q(
        ao5[6]) );
  DRNQHSV1 \pe5/pe15/q_reg[26]  ( .D(n59944), .CK(clk), .RDN(n59492), .Q(
        ao5[7]) );
  DRNQHSV1 \pe5/pe15/q_reg[25]  ( .D(n59880), .CK(clk), .RDN(n59433), .Q(
        ao5[8]) );
  DRNQHSV1 \pe5/pe15/q_reg[24]  ( .D(n39887), .CK(clk), .RDN(n59447), .Q(
        ao5[9]) );
  DRNQHSV1 \pe5/pe15/q_reg[23]  ( .D(n59642), .CK(clk), .RDN(n59397), .Q(
        ao5[10]) );
  DRNQHSV1 \pe5/pe15/q_reg[21]  ( .D(n59896), .CK(clk), .RDN(n59457), .Q(
        ao5[12]) );
  DRNQHSV1 \pe5/pe15/q_reg[20]  ( .D(\pe5/aot [13]), .CK(clk), .RDN(n59494), 
        .Q(ao5[13]) );
  DRNQHSV1 \pe5/pe15/q_reg[18]  ( .D(n59943), .CK(clk), .RDN(n59488), .Q(
        ao5[15]) );
  DRNQHSV1 \pe5/pe15/q_reg[17]  ( .D(n59640), .CK(clk), .RDN(n59488), .Q(
        ao5[16]) );
  DRNQHSV1 \pe5/pe15/q_reg[16]  ( .D(n59881), .CK(clk), .RDN(n59396), .Q(
        ao5[17]) );
  DRNQHSV1 \pe5/pe15/q_reg[15]  ( .D(\pe5/aot [18]), .CK(clk), .RDN(n59474), 
        .Q(ao5[18]) );
  DRNQHSV1 \pe5/pe15/q_reg[14]  ( .D(n59942), .CK(clk), .RDN(n59464), .Q(
        ao5[19]) );
  DRNQHSV1 \pe5/pe15/q_reg[13]  ( .D(n52591), .CK(clk), .RDN(n59650), .Q(
        ao5[20]) );
  DRNQHSV1 \pe5/pe15/q_reg[12]  ( .D(n59638), .CK(clk), .RDN(n59488), .Q(
        ao5[21]) );
  DRNQHSV1 \pe5/pe15/q_reg[11]  ( .D(n59941), .CK(clk), .RDN(n59437), .Q(
        ao5[22]) );
  DRNQHSV1 \pe5/pe15/q_reg[10]  ( .D(\pe5/aot [23]), .CK(clk), .RDN(n59399), 
        .Q(ao5[23]) );
  DRNQHSV1 \pe5/pe15/q_reg[9]  ( .D(n59940), .CK(clk), .RDN(n59925), .Q(
        ao5[24]) );
  DRNQHSV1 \pe5/pe15/q_reg[8]  ( .D(n59387), .CK(clk), .RDN(n59653), .Q(
        ao5[25]) );
  DRNQHSV1 \pe5/pe15/q_reg[7]  ( .D(n59879), .CK(clk), .RDN(n59412), .Q(
        ao5[26]) );
  DRNQHSV1 \pe5/pe15/q_reg[6]  ( .D(n59939), .CK(clk), .RDN(n59435), .Q(
        ao5[27]) );
  DRNQHSV1 \pe5/pe15/q_reg[5]  ( .D(n39266), .CK(clk), .RDN(n59464), .Q(
        ao5[28]) );
  DRNQHSV1 \pe5/pe15/q_reg[4]  ( .D(n59938), .CK(clk), .RDN(n59464), .Q(
        ao5[29]) );
  DRNQHSV1 \pe5/pe15/q_reg[3]  ( .D(n59427), .CK(clk), .RDN(n59502), .Q(
        ao5[30]) );
  DRNQHSV1 \pe5/pe15/q_reg[2]  ( .D(n59937), .CK(clk), .RDN(n59456), .Q(
        ao5[31]) );
  DRNQHSV1 \pe5/pe16/q_reg[32]  ( .D(\pe5/got [1]), .CK(clk), .RDN(n59433), 
        .Q(go5[1]) );
  DRNQHSV1 \pe5/pe16/q_reg[31]  ( .D(n59357), .CK(clk), .RDN(n59400), .Q(
        go5[2]) );
  DRNQHSV1 \pe5/pe16/q_reg[30]  ( .D(n59355), .CK(clk), .RDN(n59461), .Q(
        go5[3]) );
  DRNQHSV1 \pe5/pe16/q_reg[29]  ( .D(n52577), .CK(clk), .RDN(n59396), .Q(
        go5[4]) );
  DRNQHSV1 \pe5/pe16/q_reg[28]  ( .D(n51334), .CK(clk), .RDN(n59415), .Q(
        go5[5]) );
  DRNQHSV1 \pe5/pe16/q_reg[27]  ( .D(n51200), .CK(clk), .RDN(n59656), .Q(
        go5[6]) );
  DRNQHSV1 \pe5/pe16/q_reg[26]  ( .D(n59905), .CK(clk), .RDN(n59413), .Q(
        go5[7]) );
  DRNQHSV1 \pe5/pe16/q_reg[25]  ( .D(n50698), .CK(clk), .RDN(n59471), .Q(
        go5[8]) );
  DRNQHSV1 \pe5/pe16/q_reg[24]  ( .D(n59891), .CK(clk), .RDN(n59474), .Q(
        go5[9]) );
  DRNQHSV1 \pe5/pe16/q_reg[23]  ( .D(\pe5/got [10]), .CK(clk), .RDN(n59477), 
        .Q(go5[10]) );
  DRNQHSV1 \pe5/pe16/q_reg[22]  ( .D(n59643), .CK(clk), .RDN(n29731), .Q(
        go5[11]) );
  DRNQHSV1 \pe5/pe16/q_reg[21]  ( .D(n48167), .CK(clk), .RDN(n59467), .Q(
        go5[12]) );
  DRNQHSV1 \pe5/pe16/q_reg[20]  ( .D(n59367), .CK(clk), .RDN(n59654), .Q(
        go5[13]) );
  DRNQHSV1 \pe5/pe16/q_reg[19]  ( .D(n40186), .CK(clk), .RDN(n59478), .Q(
        go5[14]) );
  DRNQHSV1 \pe5/pe16/q_reg[18]  ( .D(n50643), .CK(clk), .RDN(n59652), .Q(
        go5[15]) );
  DRNQHSV1 \pe5/pe16/q_reg[17]  ( .D(n39881), .CK(clk), .RDN(n59400), .Q(
        go5[16]) );
  DRNQHSV1 \pe5/pe16/q_reg[16]  ( .D(n59949), .CK(clk), .RDN(n29731), .Q(
        go5[17]) );
  DRNQHSV1 \pe5/pe16/q_reg[15]  ( .D(n39433), .CK(clk), .RDN(n59653), .Q(
        go5[18]) );
  DRNQHSV1 \pe5/pe16/q_reg[14]  ( .D(n47056), .CK(clk), .RDN(n59657), .Q(
        go5[19]) );
  DRNQHSV1 \pe5/pe16/q_reg[13]  ( .D(n45816), .CK(clk), .RDN(n29733), .Q(
        go5[20]) );
  DRNQHSV1 \pe5/pe16/q_reg[12]  ( .D(n40170), .CK(clk), .RDN(n59491), .Q(
        go5[21]) );
  DRNQHSV1 \pe5/pe16/q_reg[11]  ( .D(n47267), .CK(clk), .RDN(n59409), .Q(
        go5[22]) );
  DRNQHSV1 \pe5/pe16/q_reg[10]  ( .D(n59948), .CK(clk), .RDN(n59657), .Q(
        go5[23]) );
  DRNQHSV1 \pe5/pe16/q_reg[9]  ( .D(n59637), .CK(clk), .RDN(n59450), .Q(
        go5[24]) );
  DRNQHSV1 \pe5/pe16/q_reg[8]  ( .D(n37630), .CK(clk), .RDN(n59401), .Q(
        go5[25]) );
  DRNQHSV1 \pe5/pe16/q_reg[7]  ( .D(n48742), .CK(clk), .RDN(n59451), .Q(
        go5[26]) );
  DRNQHSV1 \pe5/pe16/q_reg[6]  ( .D(\pe5/got [27]), .CK(clk), .RDN(n59407), 
        .Q(go5[27]) );
  DRNQHSV1 \pe5/pe16/q_reg[5]  ( .D(n59947), .CK(clk), .RDN(n59434), .Q(
        go5[28]) );
  DRNQHSV1 \pe5/pe16/q_reg[4]  ( .D(n30046), .CK(clk), .RDN(n29734), .Q(
        go5[29]) );
  DRNQHSV1 \pe5/pe16/q_reg[3]  ( .D(n59395), .CK(clk), .RDN(n59433), .Q(
        go5[30]) );
  DRNQHSV1 \pe5/pe16/q_reg[2]  ( .D(n59946), .CK(clk), .RDN(n59419), .Q(
        go5[31]) );
  DRNQHSV1 \pe5/pe16/q_reg[1]  ( .D(n59507), .CK(clk), .RDN(n59494), .Q(
        go5[32]) );
  DRNQHSV2 \pe5/pe17/q_reg[31]  ( .D(\pe5/poht [31]), .CK(clk), .RDN(n59491), 
        .Q(poh5[31]) );
  DRNQHSV2 \pe5/pe17/q_reg[30]  ( .D(\pe5/poht [30]), .CK(clk), .RDN(n59459), 
        .Q(poh5[30]) );
  DRNQHSV2 \pe5/pe17/q_reg[28]  ( .D(\pe5/poht [28]), .CK(clk), .RDN(n59445), 
        .Q(poh5[28]) );
  DRNQHSV2 \pe5/pe17/q_reg[27]  ( .D(\pe5/poht [27]), .CK(clk), .RDN(n59459), 
        .Q(poh5[27]) );
  DRNQHSV2 \pe5/pe17/q_reg[26]  ( .D(\pe5/poht [26]), .CK(clk), .RDN(n59468), 
        .Q(poh5[26]) );
  DRNQHSV2 \pe5/pe17/q_reg[25]  ( .D(\pe5/poht [25]), .CK(clk), .RDN(n59440), 
        .Q(poh5[25]) );
  DRNQHSV2 \pe5/pe17/q_reg[24]  ( .D(\pe5/poht [24]), .CK(clk), .RDN(n59464), 
        .Q(poh5[24]) );
  DRNQHSV2 \pe5/pe17/q_reg[23]  ( .D(\pe5/poht [23]), .CK(clk), .RDN(n59464), 
        .Q(poh5[23]) );
  DRNQHSV2 \pe5/pe17/q_reg[22]  ( .D(\pe5/poht [22]), .CK(clk), .RDN(n59435), 
        .Q(poh5[22]) );
  DRNQHSV2 \pe5/pe17/q_reg[21]  ( .D(\pe5/poht [21]), .CK(clk), .RDN(n59488), 
        .Q(poh5[21]) );
  DRNQHSV2 \pe5/pe17/q_reg[20]  ( .D(\pe5/poht [20]), .CK(clk), .RDN(n59437), 
        .Q(poh5[20]) );
  DRNQHSV2 \pe5/pe17/q_reg[19]  ( .D(\pe5/poht [19]), .CK(clk), .RDN(n59413), 
        .Q(poh5[19]) );
  DRNQHSV2 \pe5/pe17/q_reg[17]  ( .D(\pe5/poht [17]), .CK(clk), .RDN(n59464), 
        .Q(poh5[17]) );
  DRNQHSV1 \pe5/pe17/q_reg[16]  ( .D(\pe5/poht [16]), .CK(clk), .RDN(n59474), 
        .Q(poh5[16]) );
  DRNQHSV2 \pe5/pe17/q_reg[15]  ( .D(\pe5/poht [15]), .CK(clk), .RDN(n59464), 
        .Q(poh5[15]) );
  DRNQHSV2 \pe5/pe17/q_reg[14]  ( .D(\pe5/poht [14]), .CK(clk), .RDN(n59483), 
        .Q(poh5[14]) );
  DRNQHSV2 \pe5/pe17/q_reg[13]  ( .D(\pe5/poht [13]), .CK(clk), .RDN(n59650), 
        .Q(poh5[13]) );
  DRNQHSV2 \pe5/pe17/q_reg[12]  ( .D(\pe5/poht [12]), .CK(clk), .RDN(n59656), 
        .Q(poh5[12]) );
  DRNQHSV2 \pe5/pe17/q_reg[11]  ( .D(\pe5/poht [11]), .CK(clk), .RDN(n59455), 
        .Q(poh5[11]) );
  DRNQHSV2 \pe5/pe17/q_reg[9]  ( .D(\pe5/poht [9]), .CK(clk), .RDN(n59452), 
        .Q(poh5[9]) );
  DRNQHSV2 \pe5/pe17/q_reg[7]  ( .D(\pe5/poht [7]), .CK(clk), .RDN(n59397), 
        .Q(poh5[7]) );
  DRNQHSV2 \pe5/pe17/q_reg[6]  ( .D(\pe5/poht [6]), .CK(clk), .RDN(n59512), 
        .Q(poh5[6]) );
  DRNQHSV2 \pe5/pe17/q_reg[2]  ( .D(\pe5/poht [2]), .CK(clk), .RDN(n59445), 
        .Q(poh5[2]) );
  DRNQHSV1 \pe4/pe14/q_reg[30]  ( .D(n59579), .CK(clk), .RDN(n59925), .Q(
        \pe4/ti_7t [30]) );
  DRNQHSV1 \pe2/pe14/q_reg[31]  ( .D(n59794), .CK(clk), .RDN(n59488), .Q(
        \pe2/ti_7t [31]) );
  DRNQHSV2 \pe6/pe3/q_reg[32]  ( .D(bo5[1]), .CK(clk), .RDN(n59656), .Q(bo6[1]) );
  DRNQHSV2 \pe6/pe3/q_reg[30]  ( .D(bo5[3]), .CK(clk), .RDN(n59458), .Q(bo6[3]) );
  DRNQHSV2 \pe6/pe3/q_reg[29]  ( .D(bo5[4]), .CK(clk), .RDN(n29729), .Q(bo6[4]) );
  DRNQHSV2 \pe6/pe3/q_reg[28]  ( .D(bo5[5]), .CK(clk), .RDN(n59402), .Q(bo6[5]) );
  DRNQHSV2 \pe6/pe3/q_reg[27]  ( .D(bo5[6]), .CK(clk), .RDN(n59473), .Q(bo6[6]) );
  DRNQHSV2 \pe6/pe3/q_reg[26]  ( .D(bo5[7]), .CK(clk), .RDN(n59411), .Q(bo6[7]) );
  DRNQHSV2 \pe6/pe3/q_reg[25]  ( .D(bo5[8]), .CK(clk), .RDN(n59474), .Q(bo6[8]) );
  DRNQHSV2 \pe6/pe3/q_reg[24]  ( .D(bo5[9]), .CK(clk), .RDN(n59655), .Q(bo6[9]) );
  DRNQHSV2 \pe6/pe3/q_reg[22]  ( .D(bo5[11]), .CK(clk), .RDN(n59503), .Q(
        bo6[11]) );
  DRNQHSV2 \pe6/pe3/q_reg[21]  ( .D(bo5[12]), .CK(clk), .RDN(n59652), .Q(
        bo6[12]) );
  DRNQHSV2 \pe6/pe3/q_reg[20]  ( .D(bo5[13]), .CK(clk), .RDN(n59461), .Q(
        bo6[13]) );
  DRNQHSV2 \pe6/pe3/q_reg[18]  ( .D(bo5[15]), .CK(clk), .RDN(n59460), .Q(
        bo6[15]) );
  DRNQHSV2 \pe6/pe3/q_reg[17]  ( .D(bo5[16]), .CK(clk), .RDN(n59482), .Q(
        bo6[16]) );
  DRNQHSV2 \pe6/pe3/q_reg[16]  ( .D(bo5[17]), .CK(clk), .RDN(n59407), .Q(
        bo6[17]) );
  DRNQHSV2 \pe6/pe3/q_reg[15]  ( .D(bo5[18]), .CK(clk), .RDN(n59925), .Q(
        bo6[18]) );
  DRNQHSV2 \pe6/pe3/q_reg[14]  ( .D(bo5[19]), .CK(clk), .RDN(n29729), .Q(
        bo6[19]) );
  DRNQHSV2 \pe6/pe3/q_reg[13]  ( .D(bo5[20]), .CK(clk), .RDN(n59466), .Q(
        bo6[20]) );
  DRNQHSV2 \pe6/pe3/q_reg[12]  ( .D(bo5[21]), .CK(clk), .RDN(n59482), .Q(
        bo6[21]) );
  DRNQHSV2 \pe6/pe3/q_reg[11]  ( .D(bo5[22]), .CK(clk), .RDN(n59442), .Q(
        bo6[22]) );
  DRNQHSV2 \pe6/pe3/q_reg[10]  ( .D(bo5[23]), .CK(clk), .RDN(n59483), .Q(
        bo6[23]) );
  DRNQHSV2 \pe6/pe3/q_reg[9]  ( .D(bo5[24]), .CK(clk), .RDN(n59653), .Q(
        bo6[24]) );
  DRNQHSV2 \pe6/pe3/q_reg[8]  ( .D(bo5[25]), .CK(clk), .RDN(n59512), .Q(
        bo6[25]) );
  DRNQHSV2 \pe6/pe3/q_reg[7]  ( .D(bo5[26]), .CK(clk), .RDN(n59469), .Q(
        bo6[26]) );
  DRNQHSV2 \pe6/pe3/q_reg[6]  ( .D(bo5[27]), .CK(clk), .RDN(n29729), .Q(
        bo6[27]) );
  DRNQHSV2 \pe6/pe3/q_reg[5]  ( .D(bo5[28]), .CK(clk), .RDN(n59464), .Q(
        bo6[28]) );
  DRNQHSV2 \pe6/pe3/q_reg[4]  ( .D(bo5[29]), .CK(clk), .RDN(n59450), .Q(
        bo6[29]) );
  DRNQHSV2 \pe6/pe3/q_reg[3]  ( .D(bo5[30]), .CK(clk), .RDN(n59419), .Q(
        bo6[30]) );
  DRNQHSV2 \pe6/pe3/q_reg[2]  ( .D(bo5[31]), .CK(clk), .RDN(n59922), .Q(
        bo6[31]) );
  DRNQHSV2 \pe6/pe3/q_reg[1]  ( .D(bo5[32]), .CK(clk), .RDN(n59410), .Q(
        bo6[32]) );
  DRNQHSV2 \pe6/pe17/q_reg[31]  ( .D(\pe6/poht [31]), .CK(clk), .RDN(n59443), 
        .Q(poh6[31]) );
  DRNQHSV2 \pe6/pe17/q_reg[12]  ( .D(\pe6/poht [12]), .CK(clk), .RDN(n59450), 
        .Q(poh6[12]) );
  DRNQHSV2 \pe6/pe17/q_reg[11]  ( .D(\pe6/poht [11]), .CK(clk), .RDN(n29732), 
        .Q(poh6[11]) );
  DRNQHSV1 \pe1/pe14/q_reg[30]  ( .D(n59428), .CK(clk), .RDN(n59464), .Q(
        \pe1/ti_7t [30]) );
  DRNQHSV1 \pe3/pe14/q_reg[31]  ( .D(n56676), .CK(clk), .RDN(n59445), .Q(
        \pe3/ti_7t [31]) );
  DRNQHSV1 \pe4/pe14/q_reg[29]  ( .D(n26417), .CK(clk), .RDN(n59456), .Q(
        \pe4/ti_7t [29]) );
  DRNQHSV1 \pe5/pe14/q_reg[31]  ( .D(n59421), .CK(clk), .RDN(n59472), .Q(
        \pe5/ti_7t [31]) );
  DRNQHSV1 \pe6/pe14/q_reg[29]  ( .D(n58712), .CK(clk), .RDN(n59452), .Q(
        \pe6/ti_7t [29]) );
  DRNQHSV1 \pe6/pe14/q_reg[30]  ( .D(n59167), .CK(clk), .RDN(n59484), .Q(
        \pe6/ti_7t [30]) );
  DRNQHSV1 \pe6/pe14/q_reg[31]  ( .D(n59023), .CK(clk), .RDN(n59480), .Q(
        \pe6/ti_7t [31]) );
  DRNQHSV1 \pe6/pe17/q_reg[24]  ( .D(\pe6/poht [24]), .CK(clk), .RDN(n59923), 
        .Q(poh6[24]) );
  DRNQHSV2 \pe6/pe17/q_reg[10]  ( .D(\pe6/poht [10]), .CK(clk), .RDN(n59461), 
        .Q(poh6[10]) );
  DRNQHSV2 \pe2/pe3/q_reg[31]  ( .D(bo1[2]), .CK(clk), .RDN(n59461), .Q(bo2[2]) );
  DRNQHSV2 \pe2/pe3/q_reg[28]  ( .D(bo1[5]), .CK(clk), .RDN(n59408), .Q(bo2[5]) );
  DRNQHSV2 \pe2/pe3/q_reg[25]  ( .D(bo1[8]), .CK(clk), .RDN(n59470), .Q(bo2[8]) );
  DRNQHSV2 \pe2/pe3/q_reg[21]  ( .D(bo1[12]), .CK(clk), .RDN(n59473), .Q(
        bo2[12]) );
  DRNQHSV2 \pe2/pe3/q_reg[14]  ( .D(bo1[19]), .CK(clk), .RDN(n29732), .Q(
        bo2[19]) );
  DRNQHSV2 \pe2/pe3/q_reg[10]  ( .D(bo1[23]), .CK(clk), .RDN(n59418), .Q(
        bo2[23]) );
  DRNQHSV2 \pe3/pe3/q_reg[29]  ( .D(bo2[4]), .CK(clk), .RDN(n59462), .Q(bo3[4]) );
  DRNQHSV2 \pe3/pe3/q_reg[26]  ( .D(bo2[7]), .CK(clk), .RDN(n59459), .Q(bo3[7]) );
  DRNQHSV2 \pe3/pe3/q_reg[15]  ( .D(bo2[18]), .CK(clk), .RDN(n59417), .Q(
        bo3[18]) );
  DRNQHSV2 \pe3/pe3/q_reg[10]  ( .D(bo2[23]), .CK(clk), .RDN(n59657), .Q(
        bo3[23]) );
  DRNQHSV2 \pe3/pe3/q_reg[9]  ( .D(bo2[24]), .CK(clk), .RDN(n59432), .Q(
        bo3[24]) );
  DRNQHSV2 \pe3/pe3/q_reg[8]  ( .D(bo2[25]), .CK(clk), .RDN(n59457), .Q(
        bo3[25]) );
  DRNQHSV2 \pe3/pe3/q_reg[7]  ( .D(bo2[26]), .CK(clk), .RDN(n59413), .Q(
        bo3[26]) );
  DRNQHSV2 \pe3/pe3/q_reg[2]  ( .D(bo2[31]), .CK(clk), .RDN(n59490), .Q(
        bo3[31]) );
  DRNQHSV2 \pe4/pe3/q_reg[31]  ( .D(bo3[2]), .CK(clk), .RDN(n59655), .Q(bo4[2]) );
  DRNQHSV2 \pe4/pe3/q_reg[29]  ( .D(bo3[4]), .CK(clk), .RDN(n59658), .Q(bo4[4]) );
  DRNQHSV2 \pe4/pe3/q_reg[24]  ( .D(bo3[9]), .CK(clk), .RDN(n59659), .Q(bo4[9]) );
  DRNQHSV2 \pe4/pe3/q_reg[23]  ( .D(bo3[10]), .CK(clk), .RDN(n59468), .Q(
        bo4[10]) );
  DRNQHSV2 \pe4/pe3/q_reg[22]  ( .D(bo3[11]), .CK(clk), .RDN(n59658), .Q(
        bo4[11]) );
  DRNQHSV2 \pe4/pe3/q_reg[20]  ( .D(bo3[13]), .CK(clk), .RDN(n59924), .Q(
        bo4[13]) );
  DRNQHSV2 \pe4/pe3/q_reg[19]  ( .D(bo3[14]), .CK(clk), .RDN(n59923), .Q(
        bo4[14]) );
  DRNQHSV2 \pe4/pe3/q_reg[16]  ( .D(bo3[17]), .CK(clk), .RDN(n59921), .Q(
        bo4[17]) );
  DRNQHSV2 \pe4/pe3/q_reg[12]  ( .D(bo3[21]), .CK(clk), .RDN(n59922), .Q(
        bo4[21]) );
  DRNQHSV2 \pe5/pe3/q_reg[31]  ( .D(bo4[2]), .CK(clk), .RDN(n59925), .Q(bo5[2]) );
  DRNQHSV2 \pe5/pe3/q_reg[29]  ( .D(bo4[4]), .CK(clk), .RDN(n59655), .Q(bo5[4]) );
  DRNQHSV2 \pe5/pe3/q_reg[23]  ( .D(bo4[10]), .CK(clk), .RDN(n59449), .Q(
        bo5[10]) );
  DRNQHSV2 \pe5/pe3/q_reg[22]  ( .D(bo4[11]), .CK(clk), .RDN(n59439), .Q(
        bo5[11]) );
  DRNQHSV2 \pe5/pe3/q_reg[3]  ( .D(bo4[30]), .CK(clk), .RDN(n59410), .Q(
        bo5[30]) );
  DRNQHSV2 \pe5/pe3/q_reg[2]  ( .D(bo4[31]), .CK(clk), .RDN(n59482), .Q(
        bo5[31]) );
  DRNQHSV2 \pe1/pe3/q_reg[32]  ( .D(bi[1]), .CK(clk), .RDN(n59654), .Q(bo1[1])
         );
  DRNQHSV2 \pe1/pe3/q_reg[31]  ( .D(bi[2]), .CK(clk), .RDN(rst), .Q(bo1[2]) );
  DRNQHSV2 \pe1/pe3/q_reg[30]  ( .D(bi[3]), .CK(clk), .RDN(rst), .Q(bo1[3]) );
  DRNQHSV2 \pe1/pe3/q_reg[26]  ( .D(bi[7]), .CK(clk), .RDN(n59410), .Q(bo1[7])
         );
  DRNQHSV2 \pe1/pe3/q_reg[25]  ( .D(bi[8]), .CK(clk), .RDN(n59410), .Q(bo1[8])
         );
  DRNQHSV2 \pe1/pe3/q_reg[24]  ( .D(bi[9]), .CK(clk), .RDN(rst), .Q(bo1[9]) );
  DRNQHSV2 \pe1/pe3/q_reg[23]  ( .D(bi[10]), .CK(clk), .RDN(n59469), .Q(
        bo1[10]) );
  DRNQHSV2 \pe1/pe3/q_reg[21]  ( .D(bi[12]), .CK(clk), .RDN(n59488), .Q(
        bo1[12]) );
  DRNQHSV2 \pe1/pe3/q_reg[20]  ( .D(bi[13]), .CK(clk), .RDN(n59455), .Q(
        bo1[13]) );
  DRNQHSV2 \pe1/pe3/q_reg[17]  ( .D(bi[16]), .CK(clk), .RDN(n59488), .Q(
        bo1[16]) );
  DRNQHSV2 \pe1/pe3/q_reg[16]  ( .D(bi[17]), .CK(clk), .RDN(n59400), .Q(
        bo1[17]) );
  DRNQHSV2 \pe1/pe3/q_reg[15]  ( .D(bi[18]), .CK(clk), .RDN(n59494), .Q(
        bo1[18]) );
  DRNQHSV2 \pe1/pe3/q_reg[14]  ( .D(bi[19]), .CK(clk), .RDN(n59488), .Q(
        bo1[19]) );
  DRNQHSV2 \pe1/pe3/q_reg[13]  ( .D(bi[20]), .CK(clk), .RDN(n59469), .Q(
        bo1[20]) );
  DRNQHSV2 \pe1/pe3/q_reg[7]  ( .D(bi[26]), .CK(clk), .RDN(rst), .Q(bo1[26])
         );
  DRNQHSV2 \pe1/pe3/q_reg[6]  ( .D(bi[27]), .CK(clk), .RDN(rst), .Q(bo1[27])
         );
  DRNQHSV2 \pe1/pe3/q_reg[4]  ( .D(bi[29]), .CK(clk), .RDN(n59925), .Q(bo1[29]) );
  DRNQHSV2 \pe1/pe3/q_reg[3]  ( .D(bi[30]), .CK(clk), .RDN(rst), .Q(bo1[30])
         );
  DRNQHSV2 \pe2/pe3/q_reg[32]  ( .D(bo1[1]), .CK(clk), .RDN(n59436), .Q(bo2[1]) );
  DRNQHSV2 \pe2/pe3/q_reg[30]  ( .D(bo1[3]), .CK(clk), .RDN(n59494), .Q(bo2[3]) );
  DRNQHSV2 \pe2/pe3/q_reg[29]  ( .D(bo1[4]), .CK(clk), .RDN(n59438), .Q(bo2[4]) );
  DRNQHSV2 \pe2/pe3/q_reg[27]  ( .D(bo1[6]), .CK(clk), .RDN(n59453), .Q(bo2[6]) );
  DRNQHSV2 \pe2/pe3/q_reg[26]  ( .D(bo1[7]), .CK(clk), .RDN(n59452), .Q(bo2[7]) );
  DRNQHSV2 \pe2/pe3/q_reg[24]  ( .D(bo1[9]), .CK(clk), .RDN(n59430), .Q(bo2[9]) );
  DRNQHSV2 \pe2/pe3/q_reg[23]  ( .D(bo1[10]), .CK(clk), .RDN(n59401), .Q(
        bo2[10]) );
  DRNQHSV2 \pe2/pe3/q_reg[22]  ( .D(bo1[11]), .CK(clk), .RDN(n59440), .Q(
        bo2[11]) );
  DRNQHSV2 \pe2/pe3/q_reg[20]  ( .D(bo1[13]), .CK(clk), .RDN(n59658), .Q(
        bo2[13]) );
  DRNQHSV2 \pe2/pe3/q_reg[17]  ( .D(bo1[16]), .CK(clk), .RDN(n59429), .Q(
        bo2[16]) );
  DRNQHSV2 \pe2/pe3/q_reg[16]  ( .D(bo1[17]), .CK(clk), .RDN(n59454), .Q(
        bo2[17]) );
  DRNQHSV2 \pe2/pe3/q_reg[15]  ( .D(bo1[18]), .CK(clk), .RDN(n59472), .Q(
        bo2[18]) );
  DRNQHSV2 \pe2/pe3/q_reg[13]  ( .D(bo1[20]), .CK(clk), .RDN(n59448), .Q(
        bo2[20]) );
  DRNQHSV2 \pe2/pe3/q_reg[12]  ( .D(bo1[21]), .CK(clk), .RDN(n59655), .Q(
        bo2[21]) );
  DRNQHSV2 \pe2/pe3/q_reg[11]  ( .D(bo1[22]), .CK(clk), .RDN(n59653), .Q(
        bo2[22]) );
  DRNQHSV2 \pe2/pe3/q_reg[9]  ( .D(bo1[24]), .CK(clk), .RDN(n29733), .Q(
        bo2[24]) );
  DRNQHSV2 \pe2/pe3/q_reg[8]  ( .D(bo1[25]), .CK(clk), .RDN(n59477), .Q(
        bo2[25]) );
  DRNQHSV2 \pe2/pe3/q_reg[7]  ( .D(bo1[26]), .CK(clk), .RDN(n59657), .Q(
        bo2[26]) );
  DRNQHSV2 \pe2/pe3/q_reg[6]  ( .D(bo1[27]), .CK(clk), .RDN(n59406), .Q(
        bo2[27]) );
  DRNQHSV2 \pe2/pe3/q_reg[5]  ( .D(bo1[28]), .CK(clk), .RDN(n59496), .Q(
        bo2[28]) );
  DRNQHSV2 \pe2/pe3/q_reg[4]  ( .D(bo1[29]), .CK(clk), .RDN(n59477), .Q(
        bo2[29]) );
  DRNQHSV2 \pe2/pe3/q_reg[3]  ( .D(bo1[30]), .CK(clk), .RDN(n59484), .Q(
        bo2[30]) );
  DRNQHSV2 \pe2/pe3/q_reg[2]  ( .D(bo1[31]), .CK(clk), .RDN(n59473), .Q(
        bo2[31]) );
  DRNQHSV2 \pe2/pe3/q_reg[1]  ( .D(bo1[32]), .CK(clk), .RDN(n59492), .Q(
        bo2[32]) );
  DRNQHSV2 \pe3/pe3/q_reg[32]  ( .D(bo2[1]), .CK(clk), .RDN(n59450), .Q(bo3[1]) );
  DRNQHSV1 \pe3/pe3/q_reg[31]  ( .D(bo2[2]), .CK(clk), .RDN(n59491), .Q(bo3[2]) );
  DRNQHSV2 \pe3/pe3/q_reg[30]  ( .D(bo2[3]), .CK(clk), .RDN(n59417), .Q(bo3[3]) );
  DRNQHSV2 \pe3/pe3/q_reg[28]  ( .D(bo2[5]), .CK(clk), .RDN(n59465), .Q(bo3[5]) );
  DRNQHSV2 \pe3/pe3/q_reg[27]  ( .D(bo2[6]), .CK(clk), .RDN(n59476), .Q(bo3[6]) );
  DRNQHSV2 \pe3/pe3/q_reg[25]  ( .D(bo2[8]), .CK(clk), .RDN(n59651), .Q(bo3[8]) );
  DRNQHSV2 \pe3/pe3/q_reg[24]  ( .D(bo2[9]), .CK(clk), .RDN(n59462), .Q(bo3[9]) );
  DRNQHSV2 \pe3/pe3/q_reg[23]  ( .D(bo2[10]), .CK(clk), .RDN(n59438), .Q(
        bo3[10]) );
  DRNQHSV2 \pe3/pe3/q_reg[22]  ( .D(bo2[11]), .CK(clk), .RDN(n59462), .Q(
        bo3[11]) );
  DRNQHSV2 \pe3/pe3/q_reg[21]  ( .D(bo2[12]), .CK(clk), .RDN(n59656), .Q(
        bo3[12]) );
  DRNQHSV2 \pe3/pe3/q_reg[20]  ( .D(bo2[13]), .CK(clk), .RDN(n59410), .Q(
        bo3[13]) );
  DRNQHSV2 \pe3/pe3/q_reg[19]  ( .D(bo2[14]), .CK(clk), .RDN(n59436), .Q(
        bo3[14]) );
  DRNQHSV2 \pe3/pe3/q_reg[18]  ( .D(bo2[15]), .CK(clk), .RDN(n59462), .Q(
        bo3[15]) );
  DRNQHSV2 \pe3/pe3/q_reg[17]  ( .D(bo2[16]), .CK(clk), .RDN(n59921), .Q(
        bo3[16]) );
  DRNQHSV2 \pe3/pe3/q_reg[16]  ( .D(bo2[17]), .CK(clk), .RDN(n59488), .Q(
        bo3[17]) );
  DRNQHSV2 \pe3/pe3/q_reg[14]  ( .D(bo2[19]), .CK(clk), .RDN(n59438), .Q(
        bo3[19]) );
  DRNQHSV2 \pe3/pe3/q_reg[13]  ( .D(bo2[20]), .CK(clk), .RDN(n59462), .Q(
        bo3[20]) );
  DRNQHSV2 \pe3/pe3/q_reg[6]  ( .D(bo2[27]), .CK(clk), .RDN(n59443), .Q(
        bo3[27]) );
  DRNQHSV2 \pe3/pe3/q_reg[4]  ( .D(bo2[29]), .CK(clk), .RDN(n59406), .Q(
        bo3[29]) );
  DRNQHSV2 \pe4/pe3/q_reg[32]  ( .D(bo3[1]), .CK(clk), .RDN(n59412), .Q(bo4[1]) );
  DRNQHSV2 \pe4/pe3/q_reg[30]  ( .D(bo3[3]), .CK(clk), .RDN(n59656), .Q(bo4[3]) );
  DRNQHSV2 \pe4/pe3/q_reg[28]  ( .D(bo3[5]), .CK(clk), .RDN(n59655), .Q(bo4[5]) );
  DRNQHSV2 \pe4/pe3/q_reg[27]  ( .D(bo3[6]), .CK(clk), .RDN(n59658), .Q(bo4[6]) );
  DRNQHSV2 \pe4/pe3/q_reg[26]  ( .D(bo3[7]), .CK(clk), .RDN(n59649), .Q(bo4[7]) );
  DRNQHSV2 \pe4/pe3/q_reg[25]  ( .D(bo3[8]), .CK(clk), .RDN(n59654), .Q(bo4[8]) );
  DRNQHSV2 \pe4/pe3/q_reg[21]  ( .D(bo3[12]), .CK(clk), .RDN(n59490), .Q(
        bo4[12]) );
  DRNQHSV2 \pe4/pe3/q_reg[18]  ( .D(bo3[15]), .CK(clk), .RDN(n59922), .Q(
        bo4[15]) );
  DRNQHSV2 \pe4/pe3/q_reg[17]  ( .D(bo3[16]), .CK(clk), .RDN(n59653), .Q(
        bo4[16]) );
  DRNQHSV2 \pe4/pe3/q_reg[15]  ( .D(bo3[18]), .CK(clk), .RDN(n59444), .Q(
        bo4[18]) );
  DRNQHSV2 \pe4/pe3/q_reg[14]  ( .D(bo3[19]), .CK(clk), .RDN(n59479), .Q(
        bo4[19]) );
  DRNQHSV2 \pe4/pe3/q_reg[13]  ( .D(bo3[20]), .CK(clk), .RDN(n59412), .Q(
        bo4[20]) );
  DRNQHSV2 \pe4/pe3/q_reg[11]  ( .D(bo3[22]), .CK(clk), .RDN(n59923), .Q(
        bo4[22]) );
  DRNQHSV2 \pe4/pe3/q_reg[10]  ( .D(bo3[23]), .CK(clk), .RDN(n59456), .Q(
        bo4[23]) );
  DRNQHSV2 \pe4/pe3/q_reg[9]  ( .D(bo3[24]), .CK(clk), .RDN(n59431), .Q(
        bo4[24]) );
  DRNQHSV2 \pe4/pe3/q_reg[8]  ( .D(bo3[25]), .CK(clk), .RDN(n59417), .Q(
        bo4[25]) );
  DRNQHSV2 \pe4/pe3/q_reg[7]  ( .D(bo3[26]), .CK(clk), .RDN(n59503), .Q(
        bo4[26]) );
  DRNQHSV2 \pe4/pe3/q_reg[6]  ( .D(bo3[27]), .CK(clk), .RDN(n59455), .Q(
        bo4[27]) );
  DRNQHSV2 \pe4/pe3/q_reg[5]  ( .D(bo3[28]), .CK(clk), .RDN(n59471), .Q(
        bo4[28]) );
  DRNQHSV2 \pe4/pe3/q_reg[4]  ( .D(bo3[29]), .CK(clk), .RDN(n59482), .Q(
        bo4[29]) );
  DRNQHSV2 \pe4/pe3/q_reg[3]  ( .D(bo3[30]), .CK(clk), .RDN(n59460), .Q(
        bo4[30]) );
  DRNQHSV1 \pe4/pe3/q_reg[2]  ( .D(bo3[31]), .CK(clk), .RDN(n59417), .Q(
        bo4[31]) );
  DRNQHSV2 \pe4/pe3/q_reg[1]  ( .D(bo3[32]), .CK(clk), .RDN(n59649), .Q(
        bo4[32]) );
  DRNQHSV2 \pe5/pe3/q_reg[32]  ( .D(bo4[1]), .CK(clk), .RDN(n59470), .Q(bo5[1]) );
  DRNQHSV2 \pe5/pe3/q_reg[30]  ( .D(bo4[3]), .CK(clk), .RDN(n59459), .Q(bo5[3]) );
  DRNQHSV2 \pe5/pe3/q_reg[28]  ( .D(bo4[5]), .CK(clk), .RDN(n59490), .Q(bo5[5]) );
  DRNQHSV2 \pe5/pe3/q_reg[27]  ( .D(bo4[6]), .CK(clk), .RDN(n59462), .Q(bo5[6]) );
  DRNQHSV2 \pe5/pe3/q_reg[26]  ( .D(bo4[7]), .CK(clk), .RDN(n59425), .Q(bo5[7]) );
  DRNQHSV2 \pe5/pe3/q_reg[25]  ( .D(bo4[8]), .CK(clk), .RDN(n59416), .Q(bo5[8]) );
  DRNQHSV1 \pe5/pe3/q_reg[24]  ( .D(bo4[9]), .CK(clk), .RDN(n59432), .Q(bo5[9]) );
  DRNQHSV2 \pe5/pe3/q_reg[21]  ( .D(bo4[12]), .CK(clk), .RDN(n59651), .Q(
        bo5[12]) );
  DRNQHSV1 \pe5/pe3/q_reg[20]  ( .D(bo4[13]), .CK(clk), .RDN(n29734), .Q(
        bo5[13]) );
  DRNQHSV1 \pe5/pe3/q_reg[19]  ( .D(bo4[14]), .CK(clk), .RDN(n59413), .Q(
        bo5[14]) );
  DRNQHSV2 \pe5/pe3/q_reg[18]  ( .D(bo4[15]), .CK(clk), .RDN(n59480), .Q(
        bo5[15]) );
  DRNQHSV2 \pe5/pe3/q_reg[17]  ( .D(bo4[16]), .CK(clk), .RDN(n59433), .Q(
        bo5[16]) );
  DRNQHSV1 \pe5/pe3/q_reg[16]  ( .D(bo4[17]), .CK(clk), .RDN(n29729), .Q(
        bo5[17]) );
  DRNQHSV2 \pe5/pe3/q_reg[15]  ( .D(bo4[18]), .CK(clk), .RDN(n59496), .Q(
        bo5[18]) );
  DRNQHSV2 \pe5/pe3/q_reg[13]  ( .D(bo4[20]), .CK(clk), .RDN(n59411), .Q(
        bo5[20]) );
  DRNQHSV1 \pe5/pe3/q_reg[12]  ( .D(bo4[21]), .CK(clk), .RDN(n59454), .Q(
        bo5[21]) );
  DRNQHSV2 \pe5/pe3/q_reg[10]  ( .D(bo4[23]), .CK(clk), .RDN(n59496), .Q(
        bo5[23]) );
  DRNQHSV2 \pe5/pe3/q_reg[9]  ( .D(bo4[24]), .CK(clk), .RDN(n59438), .Q(
        bo5[24]) );
  DRNQHSV2 \pe5/pe3/q_reg[8]  ( .D(bo4[25]), .CK(clk), .RDN(n59452), .Q(
        bo5[25]) );
  DRNQHSV2 \pe5/pe3/q_reg[7]  ( .D(bo4[26]), .CK(clk), .RDN(n59651), .Q(
        bo5[26]) );
  DRNQHSV2 \pe5/pe3/q_reg[6]  ( .D(bo4[27]), .CK(clk), .RDN(n59468), .Q(
        bo5[27]) );
  DRNQHSV2 \pe5/pe3/q_reg[5]  ( .D(bo4[28]), .CK(clk), .RDN(n59463), .Q(
        bo5[28]) );
  DRNQHSV2 \pe5/pe3/q_reg[4]  ( .D(bo4[29]), .CK(clk), .RDN(n59470), .Q(
        bo5[29]) );
  DRNQHSV2 \pe5/pe3/q_reg[1]  ( .D(bo4[32]), .CK(clk), .RDN(n59445), .Q(
        bo5[32]) );
  DRNQHSV1 \pe1/pe14/q_reg[31]  ( .D(n25848), .CK(clk), .RDN(n59925), .Q(
        \pe1/ti_7t [31]) );
  DRNQHSV1 \pe5/pe14/q_reg[30]  ( .D(n52668), .CK(clk), .RDN(n59396), .Q(
        \pe5/ti_7t [30]) );
  DRNQHSV1 \pe2/pe14/q_reg[29]  ( .D(n52414), .CK(clk), .RDN(n59474), .Q(
        \pe2/ti_7t [29]) );
  DRNQHSV1 \pe5/pe14/q_reg[24]  ( .D(n59516), .CK(clk), .RDN(n59655), .Q(
        \pe5/ti_7t [24]) );
  DRNQHSV1 \pe2/pe14/q_reg[26]  ( .D(n59929), .CK(clk), .RDN(n59434), .Q(
        \pe2/ti_7t [26]) );
  DRNQHSV1 \pe5/pe14/q_reg[26]  ( .D(n59535), .CK(clk), .RDN(n59455), .Q(
        \pe5/ti_7t [26]) );
  DRNQHSV1 \pe6/pe14/q_reg[24]  ( .D(n59487), .CK(clk), .RDN(n59659), .Q(
        \pe6/ti_7t [24]) );
  DRNQHSV1 \pe6/pe14/q_reg[26]  ( .D(n59528), .CK(clk), .RDN(n59424), .Q(
        \pe6/ti_7t [26]) );
  DRNQHSV1 \pe3/pe14/q_reg[26]  ( .D(n56173), .CK(clk), .RDN(n59458), .Q(
        \pe3/ti_7t [26]) );
  DRNQHSV1 \pe1/pe14/q_reg[24]  ( .D(n59751), .CK(clk), .RDN(n59404), .Q(
        \pe1/ti_7t [24]) );
  DRNQHSV1 \pe1/pe14/q_reg[25]  ( .D(n59736), .CK(clk), .RDN(n59492), .Q(
        \pe1/ti_7t [25]) );
  DRNQHSV1 \pe3/pe14/q_reg[28]  ( .D(n56953), .CK(clk), .RDN(n29730), .Q(
        \pe3/ti_7t [28]) );
  DRNQHSV1 \pe4/pe14/q_reg[25]  ( .D(n59837), .CK(clk), .RDN(n59437), .Q(
        \pe4/ti_7t [25]) );
  DRNQHSV1 \pe4/pe14/q_reg[28]  ( .D(n26596), .CK(clk), .RDN(n59436), .Q(
        \pe4/ti_7t [28]) );
  DRNQHSV1 \pe6/pe14/q_reg[28]  ( .D(n59514), .CK(clk), .RDN(n59419), .Q(
        \pe6/ti_7t [28]) );
  DRNQHSV1 \pe2/pe14/q_reg[27]  ( .D(n52168), .CK(clk), .RDN(n59424), .Q(
        \pe2/ti_7t [27]) );
  DRNQHSV1 \pe3/pe14/q_reg[29]  ( .D(n56172), .CK(clk), .RDN(n59416), .Q(
        \pe3/ti_7t [29]) );
  DRNQHSV1 \pe4/pe14/q_reg[26]  ( .D(n58141), .CK(clk), .RDN(n59436), .Q(
        \pe4/ti_7t [26]) );
  DRNQHSV1 \pe5/pe14/q_reg[27]  ( .D(n52564), .CK(clk), .RDN(n59443), .Q(
        \pe5/ti_7t [27]) );
  DRNQHSV1 \pe6/pe14/q_reg[27]  ( .D(n58809), .CK(clk), .RDN(n59924), .Q(
        \pe6/ti_7t [27]) );
  DRNQHSV2 \pe1/pe14/q_reg[26]  ( .D(n54146), .CK(clk), .RDN(n59496), .Q(
        \pe1/ti_7t [26]) );
  DRNQHSV1 \pe2/pe14/q_reg[28]  ( .D(n59475), .CK(clk), .RDN(n59445), .Q(
        \pe2/ti_7t [28]) );
  DRNQHSV1 \pe4/pe14/q_reg[27]  ( .D(n59348), .CK(clk), .RDN(n59451), .Q(
        \pe4/ti_7t [27]) );
  DRNQHSV1 \pe2/pe14/q_reg[25]  ( .D(n59927), .CK(clk), .RDN(n59414), .Q(
        \pe2/ti_7t [25]) );
  DRNQHSV1 \pe5/pe14/q_reg[25]  ( .D(n59892), .CK(clk), .RDN(n59512), .Q(
        \pe5/ti_7t [25]) );
  DRNQHSV1 \pe5/pe14/q_reg[28]  ( .D(n59933), .CK(clk), .RDN(n59396), .Q(
        \pe5/ti_7t [28]) );
  DRNQHSV1 \pe4/pe14/q_reg[24]  ( .D(n35033), .CK(clk), .RDN(n59406), .Q(
        \pe4/ti_7t [24]) );
  DRNQHSV1 \pe6/pe14/q_reg[25]  ( .D(n58716), .CK(clk), .RDN(n59512), .Q(
        \pe6/ti_7t [25]) );
  DRNQHSV1 \pe2/pe14/q_reg[22]  ( .D(n59774), .CK(clk), .RDN(n59436), .Q(
        \pe2/ti_7t [22]) );
  DRNQHSV1 \pe2/pe14/q_reg[23]  ( .D(n59522), .CK(clk), .RDN(n29731), .Q(
        \pe2/ti_7t [23]) );
  DRNQHSV1 \pe3/pe14/q_reg[20]  ( .D(n59500), .CK(clk), .RDN(n59400), .Q(
        \pe3/ti_7t [20]) );
  DRNQHSV1 \pe3/pe14/q_reg[21]  ( .D(n59920), .CK(clk), .RDN(n59457), .Q(
        \pe3/ti_7t [21]) );
  DRNQHSV1 \pe4/pe14/q_reg[22]  ( .D(n47841), .CK(clk), .RDN(n59477), .Q(
        \pe4/ti_7t [22]) );
  DRNQHSV1 \pe5/pe14/q_reg[19]  ( .D(n52653), .CK(clk), .RDN(n59435), .Q(
        \pe5/ti_7t [19]) );
  DRNQHSV1 \pe2/pe14/q_reg[24]  ( .D(n59790), .CK(clk), .RDN(n59403), .Q(
        \pe2/ti_7t [24]) );
  DRNQHSV1 \pe4/pe14/q_reg[23]  ( .D(n25427), .CK(clk), .RDN(n59476), .Q(
        \pe4/ti_7t [23]) );
  DRNQHSV1 \pe2/pe14/q_reg[21]  ( .D(n60002), .CK(clk), .RDN(n59510), .Q(
        \pe2/ti_7t [21]) );
  DRNQHSV1 \pe3/pe14/q_reg[23]  ( .D(n59930), .CK(clk), .RDN(n59458), .Q(
        \pe3/ti_7t [23]) );
  DRNQHSV1 \pe4/pe14/q_reg[20]  ( .D(n50065), .CK(clk), .RDN(n59442), .Q(
        \pe4/ti_7t [20]) );
  DRNQHSV1 \pe6/pe14/q_reg[22]  ( .D(n59918), .CK(clk), .RDN(n59452), .Q(
        \pe6/ti_7t [22]) );
  DRNQHSV1 \pe6/pe14/q_reg[23]  ( .D(n59677), .CK(clk), .RDN(n59460), .Q(
        \pe6/ti_7t [23]) );
  DRNQHSV1 \pe3/pe14/q_reg[22]  ( .D(n49253), .CK(clk), .RDN(n59451), .Q(
        \pe3/ti_7t [22]) );
  DRNQHSV1 \pe5/pe14/q_reg[21]  ( .D(n59903), .CK(clk), .RDN(n59412), .Q(
        \pe5/ti_7t [21]) );
  DRNQHSV1 \pe1/pe14/q_reg[20]  ( .D(n59391), .CK(clk), .RDN(n59459), .Q(
        \pe1/ti_7t [20]) );
  DRNQHSV1 \pe1/pe14/q_reg[23]  ( .D(n59521), .CK(clk), .RDN(n59439), .Q(
        \pe1/ti_7t [23]) );
  DRNQHSV1 \pe4/pe14/q_reg[21]  ( .D(n59672), .CK(clk), .RDN(n59443), .Q(
        \pe4/ti_7t [21]) );
  DRNQHSV1 \pe3/pe14/q_reg[24]  ( .D(n59359), .CK(clk), .RDN(n59476), .Q(
        \pe3/ti_7t [24]) );
  DRNQHSV1 \pe5/pe14/q_reg[23]  ( .D(n59893), .CK(clk), .RDN(n59431), .Q(
        \pe5/ti_7t [23]) );
  DRNQHSV1 \pe5/pe14/q_reg[22]  ( .D(n59926), .CK(clk), .RDN(n59416), .Q(
        \pe5/ti_7t [22]) );
  DRNQHSV1 \pe2/pe14/q_reg[15]  ( .D(n59773), .CK(clk), .RDN(n59468), .Q(
        \pe2/ti_7t [15]) );
  DRNQHSV1 \pe2/pe14/q_reg[18]  ( .D(n59769), .CK(clk), .RDN(n59474), .Q(
        \pe2/ti_7t [18]) );
  DRNQHSV1 \pe3/pe14/q_reg[17]  ( .D(n55824), .CK(clk), .RDN(n59925), .Q(
        \pe3/ti_7t [17]) );
  DRNQHSV1 \pe6/pe14/q_reg[16]  ( .D(n59676), .CK(clk), .RDN(n59494), .Q(
        \pe6/ti_7t [16]) );
  DRNQHSV1 \pe6/pe14/q_reg[17]  ( .D(n53113), .CK(clk), .RDN(n59458), .Q(
        \pe6/ti_7t [17]) );
  DRNQHSV1 \pe6/pe14/q_reg[18]  ( .D(n59916), .CK(clk), .RDN(n59437), .Q(
        \pe6/ti_7t [18]) );
  DRNQHSV1 \pe1/pe14/q_reg[15]  ( .D(n54521), .CK(clk), .RDN(n59471), .Q(
        \pe1/ti_7t [15]) );
  DRNQHSV1 \pe2/pe14/q_reg[17]  ( .D(n59506), .CK(clk), .RDN(n59469), .Q(
        \pe2/ti_7t [17]) );
  DRNQHSV1 \pe3/pe14/q_reg[15]  ( .D(n59810), .CK(clk), .RDN(n59470), .Q(
        \pe3/ti_7t [15]) );
  DRNQHSV1 \pe4/pe14/q_reg[17]  ( .D(n49951), .CK(clk), .RDN(n59651), .Q(
        \pe4/ti_7t [17]) );
  DRNQHSV1 \pe5/pe14/q_reg[17]  ( .D(n59882), .CK(clk), .RDN(n59482), .Q(
        \pe5/ti_7t [17]) );
  DRNQHSV1 \pe1/pe14/q_reg[18]  ( .D(n55230), .CK(clk), .RDN(n29732), .Q(
        \pe1/ti_7t [18]) );
  DRNQHSV1 \pe5/pe14/q_reg[16]  ( .D(n59517), .CK(clk), .RDN(n59431), .Q(
        \pe5/ti_7t [16]) );
  DRNQHSV1 \pe6/pe14/q_reg[19]  ( .D(n53111), .CK(clk), .RDN(n59465), .Q(
        \pe6/ti_7t [19]) );
  DRNQHSV1 \pe2/pe14/q_reg[16]  ( .D(n59505), .CK(clk), .RDN(n59406), .Q(
        \pe2/ti_7t [16]) );
  DRNQHSV1 \pe2/pe14/q_reg[20]  ( .D(n59775), .CK(clk), .RDN(n59464), .Q(
        \pe2/ti_7t [20]) );
  DRNQHSV1 \pe3/pe14/q_reg[16]  ( .D(n59811), .CK(clk), .RDN(n59479), .Q(
        \pe3/ti_7t [16]) );
  DRNQHSV1 \pe6/pe14/q_reg[20]  ( .D(n59915), .CK(clk), .RDN(n59402), .Q(
        \pe6/ti_7t [20]) );
  DRNQHSV1 \pe4/pe14/q_reg[16]  ( .D(n59526), .CK(clk), .RDN(n59415), .Q(
        \pe4/ti_7t [16]) );
  DRNQHSV1 \pe5/pe14/q_reg[15]  ( .D(n59525), .CK(clk), .RDN(n59450), .Q(
        \pe5/ti_7t [15]) );
  DRNQHSV1 \pe4/pe14/q_reg[18]  ( .D(n59935), .CK(clk), .RDN(n59407), .Q(
        \pe4/ti_7t [18]) );
  DRNQHSV1 \pe5/pe14/q_reg[18]  ( .D(n59894), .CK(clk), .RDN(n59431), .Q(
        \pe5/ti_7t [18]) );
  DRNQHSV1 \pe5/pe14/q_reg[13]  ( .D(n59878), .CK(clk), .RDN(n59455), .Q(
        \pe5/ti_7t [13]) );
  DRNQHSV1 \pe1/pe14/q_reg[16]  ( .D(n53657), .CK(clk), .RDN(n59471), .Q(
        \pe1/ti_7t [16]) );
  DRNQHSV1 \pe3/pe14/q_reg[18]  ( .D(n43754), .CK(clk), .RDN(n59483), .Q(
        \pe3/ti_7t [18]) );
  DRNQHSV1 \pe1/pe14/q_reg[17]  ( .D(n59592), .CK(clk), .RDN(n59406), .Q(
        \pe1/ti_7t [17]) );
  DRNQHSV1 \pe1/pe14/q_reg[11]  ( .D(n59934), .CK(clk), .RDN(n59468), .Q(
        \pe1/ti_7t [11]) );
  DRNQHSV1 \pe1/pe14/q_reg[12]  ( .D(n59534), .CK(clk), .RDN(n59493), .Q(
        \pe1/ti_7t [12]) );
  DRNQHSV1 \pe2/pe14/q_reg[13]  ( .D(n44713), .CK(clk), .RDN(n59399), .Q(
        \pe2/ti_7t [13]) );
  DRNQHSV1 \pe3/pe14/q_reg[11]  ( .D(n59620), .CK(clk), .RDN(n59480), .Q(
        \pe3/ti_7t [11]) );
  DRNQHSV1 \pe4/pe14/q_reg[13]  ( .D(n34949), .CK(clk), .RDN(n59488), .Q(
        \pe4/ti_7t [13]) );
  DRNQHSV1 \pe4/pe14/q_reg[14]  ( .D(n59378), .CK(clk), .RDN(n59468), .Q(
        \pe4/ti_7t [14]) );
  DRNQHSV1 \pe5/pe14/q_reg[12]  ( .D(n59392), .CK(clk), .RDN(n59447), .Q(
        \pe5/ti_7t [12]) );
  DRNQHSV2 \pe2/pe6/q_reg[31]  ( .D(poh1[31]), .CK(clk), .RDN(n59414), .Q(
        \pe2/phq [31]) );
  DRNQHSV2 \pe5/pe6/q_reg[30]  ( .D(poh4[30]), .CK(clk), .RDN(n59415), .Q(
        \pe5/phq [30]) );
  DRNQHSV2 \pe2/pe5/q_reg[31]  ( .D(n60044), .CK(clk), .RDN(n59921), .Q(
        \pe2/pvq [31]) );
  DRNQHSV1 \pe2/pe5/q_reg[30]  ( .D(n60036), .CK(clk), .RDN(n59409), .Q(
        \pe2/pvq [30]) );
  DRNQHSV2 \pe4/pe5/q_reg[31]  ( .D(n60022), .CK(clk), .RDN(n59921), .Q(
        \pe4/pvq [31]) );
  DRNQHSV2 \pe4/pe5/q_reg[26]  ( .D(n60085), .CK(clk), .RDN(n59396), .Q(
        \pe4/pvq [26]) );
  DRNQHSV1 \pe4/pe14/q_reg[10]  ( .D(n59928), .CK(clk), .RDN(n59435), .Q(
        \pe4/ti_7t [10]) );
  DRNQHSV1 \pe4/pe14/q_reg[15]  ( .D(n57547), .CK(clk), .RDN(n59452), .Q(
        \pe4/ti_7t [15]) );
  DRNQHSV1 \pe5/pe5/q_reg[31]  ( .D(pov4[31]), .CK(clk), .RDN(n59467), .Q(
        \pe5/pvq [31]) );
  DRNQHSV1 \pe5/pe5/q_reg[30]  ( .D(n60077), .CK(clk), .RDN(n59440), .Q(
        \pe5/pvq [30]) );
  DRNQHSV1 \pe5/pe14/q_reg[9]  ( .D(n51162), .CK(clk), .RDN(n59429), .Q(
        \pe5/ti_7t [9]) );
  DRNQHSV1 \pe5/pe14/q_reg[11]  ( .D(n59871), .CK(clk), .RDN(n59448), .Q(
        \pe5/ti_7t [11]) );
  DRNQHSV1 \pe6/pe5/q_reg[22]  ( .D(n60007), .CK(clk), .RDN(n59413), .Q(
        \pe6/pvq [22]) );
  DRNQHSV1 \pe6/pe14/q_reg[10]  ( .D(n59596), .CK(clk), .RDN(n59461), .Q(
        \pe6/ti_7t [10]) );
  DRNQHSV1 \pe6/pe14/q_reg[15]  ( .D(n35898), .CK(clk), .RDN(n59430), .Q(
        \pe6/ti_7t [15]) );
  DRNQHSV1 \pe1/pe14/q_reg[10]  ( .D(n44532), .CK(clk), .RDN(n59473), .Q(
        \pe1/ti_7t [10]) );
  DRNQHSV1 \pe1/pe14/q_reg[14]  ( .D(n59518), .CK(clk), .RDN(n59480), .Q(
        \pe1/ti_7t [14]) );
  DRNQHSV1 \pe3/pe14/q_reg[10]  ( .D(n59625), .CK(clk), .RDN(n59469), .Q(
        \pe3/ti_7t [10]) );
  DRNQHSV1 \pe5/pe14/q_reg[10]  ( .D(n29770), .CK(clk), .RDN(n59436), .Q(
        \pe5/ti_7t [10]) );
  DRNQHSV1 \pe3/pe14/q_reg[14]  ( .D(n59362), .CK(clk), .RDN(n59410), .Q(
        \pe3/ti_7t [14]) );
  DRNQHSV2 \pe2/pe4/q_reg  ( .D(po1), .CK(clk), .RDN(n59925), .Q(\pe2/pq ) );
  DRNQHSV1 \pe2/pe14/q_reg[14]  ( .D(n59634), .CK(clk), .RDN(n59921), .Q(
        \pe2/ti_7t [14]) );
  DRNQHSV1 \pe3/pe4/q_reg  ( .D(po2), .CK(clk), .RDN(n59471), .Q(\pe3/pq ) );
  DRNQHSV1 \pe6/pe14/q_reg[12]  ( .D(n59420), .CK(clk), .RDN(n59470), .Q(
        \pe6/ti_7t [12]) );
  DRNQHSV2 \pe6/pe4/q_reg  ( .D(po5), .CK(clk), .RDN(n59464), .Q(\pe6/pq ) );
  DRNQHSV1 \pe2/pe14/q_reg[12]  ( .D(n59761), .CK(clk), .RDN(n29729), .Q(
        \pe2/ti_7t [12]) );
  DRNQHSV1 \pe4/pe14/q_reg[11]  ( .D(n59833), .CK(clk), .RDN(n59925), .Q(
        \pe4/ti_7t [11]) );
  DRNQHSV1 \pe4/pe14/q_reg[12]  ( .D(n59835), .CK(clk), .RDN(n59419), .Q(
        \pe4/ti_7t [12]) );
  DRNQHSV1 \pe3/pe14/q_reg[12]  ( .D(n59380), .CK(clk), .RDN(n59470), .Q(
        \pe3/ti_7t [12]) );
  DRNQHSV1 \pe2/pe14/q_reg[10]  ( .D(n52287), .CK(clk), .RDN(n59502), .Q(
        \pe2/ti_7t [10]) );
  DRNQHSV1 \pe6/pe14/q_reg[13]  ( .D(n59379), .CK(clk), .RDN(n59435), .Q(
        \pe6/ti_7t [13]) );
  DRNQHSV1 \pe6/pe14/q_reg[8]  ( .D(n59917), .CK(clk), .RDN(n29729), .Q(
        \pe6/ti_7t [8]) );
  DRNQHSV1 \pe1/pe14/q_reg[8]  ( .D(n41332), .CK(clk), .RDN(n59403), .Q(
        \pe1/ti_7t [8]) );
  DRNQHSV1 \pe1/pe14/q_reg[9]  ( .D(n29773), .CK(clk), .RDN(n59399), .Q(
        \pe1/ti_7t [9]) );
  DRNQHSV1 \pe3/pe14/q_reg[7]  ( .D(n59364), .CK(clk), .RDN(n59415), .Q(
        \pe3/ti_7t [7]) );
  DRNQHSV1 \pe3/pe14/q_reg[9]  ( .D(n59519), .CK(clk), .RDN(n59469), .Q(
        \pe3/ti_7t [9]) );
  DRNQHSV1 \pe6/pe14/q_reg[5]  ( .D(n59595), .CK(clk), .RDN(n59457), .Q(
        \pe6/ti_7t [5]) );
  DRNQHSV1 \pe2/pe14/q_reg[8]  ( .D(n59766), .CK(clk), .RDN(n59439), .Q(
        \pe2/ti_7t [8]) );
  DRNQHSV2 \pe2/pe5/q_reg[29]  ( .D(n60103), .CK(clk), .RDN(n59397), .Q(
        \pe2/pvq [29]) );
  DRNQHSV1 \pe2/pe5/q_reg[28]  ( .D(n60015), .CK(clk), .RDN(n59496), .Q(
        \pe2/pvq [28]) );
  DRNQHSV2 \pe2/pe5/q_reg[27]  ( .D(n60063), .CK(clk), .RDN(n59404), .Q(
        \pe2/pvq [27]) );
  DRNQHSV1 \pe2/pe5/q_reg[26]  ( .D(n60018), .CK(clk), .RDN(n59491), .Q(
        \pe2/pvq [26]) );
  DRNQHSV1 \pe2/pe5/q_reg[25]  ( .D(pov1[25]), .CK(clk), .RDN(n59503), .Q(
        \pe2/pvq [25]) );
  DRNQHSV1 \pe2/pe5/q_reg[24]  ( .D(n29760), .CK(clk), .RDN(n59465), .Q(
        \pe2/pvq [24]) );
  DRNQHSV1 \pe2/pe5/q_reg[23]  ( .D(pov1[23]), .CK(clk), .RDN(n59415), .Q(
        \pe2/pvq [23]) );
  DRNQHSV1 \pe2/pe5/q_reg[22]  ( .D(pov1[22]), .CK(clk), .RDN(n59494), .Q(
        \pe2/pvq [22]) );
  DRNQHSV1 \pe2/pe5/q_reg[19]  ( .D(pov1[19]), .CK(clk), .RDN(n59468), .Q(
        \pe2/pvq [19]) );
  DRNQHSV1 \pe2/pe5/q_reg[18]  ( .D(n60106), .CK(clk), .RDN(n29733), .Q(
        \pe2/pvq [18]) );
  DRNQHSV1 \pe2/pe5/q_reg[17]  ( .D(n60107), .CK(clk), .RDN(n59456), .Q(
        \pe2/pvq [17]) );
  DRNQHSV1 \pe2/pe5/q_reg[16]  ( .D(n60026), .CK(clk), .RDN(n59403), .Q(
        \pe2/pvq [16]) );
  DRNQHSV2 \pe3/pe5/q_reg[31]  ( .D(n60014), .CK(clk), .RDN(n59659), .Q(
        \pe3/pvq [31]) );
  DRNQHSV1 \pe3/pe5/q_reg[30]  ( .D(n60013), .CK(clk), .RDN(n59407), .Q(
        \pe3/pvq [30]) );
  DRNQHSV1 \pe3/pe5/q_reg[29]  ( .D(n60012), .CK(clk), .RDN(n59401), .Q(
        \pe3/pvq [29]) );
  DRNQHSV1 \pe3/pe5/q_reg[28]  ( .D(pov2[28]), .CK(clk), .RDN(n59657), .Q(
        \pe3/pvq [28]) );
  DRNQHSV2 \pe3/pe5/q_reg[27]  ( .D(n60092), .CK(clk), .RDN(n59922), .Q(
        \pe3/pvq [27]) );
  DRNQHSV1 \pe3/pe5/q_reg[26]  ( .D(n29764), .CK(clk), .RDN(n59415), .Q(
        \pe3/pvq [26]) );
  DRNQHSV1 \pe3/pe5/q_reg[22]  ( .D(n60095), .CK(clk), .RDN(n59469), .Q(
        \pe3/pvq [22]) );
  DRNQHSV1 \pe3/pe5/q_reg[20]  ( .D(n60021), .CK(clk), .RDN(n59654), .Q(
        \pe3/pvq [20]) );
  DRNQHSV1 \pe4/pe5/q_reg[30]  ( .D(n60001), .CK(clk), .RDN(n59466), .Q(
        \pe4/pvq [30]) );
  DRNQHSV2 \pe4/pe5/q_reg[29]  ( .D(pov3[29]), .CK(clk), .RDN(n59924), .Q(
        \pe4/pvq [29]) );
  DRNQHSV1 \pe4/pe5/q_reg[28]  ( .D(n60060), .CK(clk), .RDN(n59405), .Q(
        \pe4/pvq [28]) );
  DRNQHSV2 \pe4/pe5/q_reg[27]  ( .D(n60084), .CK(clk), .RDN(n59404), .Q(
        \pe4/pvq [27]) );
  DRNQHSV1 \pe4/pe5/q_reg[24]  ( .D(pov3[24]), .CK(clk), .RDN(n59403), .Q(
        \pe4/pvq [24]) );
  DRNQHSV1 \pe4/pe5/q_reg[23]  ( .D(n59575), .CK(clk), .RDN(n59453), .Q(
        \pe4/pvq [23]) );
  DRNQHSV1 \pe4/pe5/q_reg[20]  ( .D(n43137), .CK(clk), .RDN(n59925), .Q(
        \pe4/pvq [20]) );
  DRNQHSV1 \pe4/pe5/q_reg[18]  ( .D(n60086), .CK(clk), .RDN(n59465), .Q(
        \pe4/pvq [18]) );
  DRNQHSV1 \pe4/pe5/q_reg[16]  ( .D(pov3[16]), .CK(clk), .RDN(n59454), .Q(
        \pe4/pvq [16]) );
  DRNQHSV1 \pe4/pe14/q_reg[8]  ( .D(n33608), .CK(clk), .RDN(n59483), .Q(
        \pe4/ti_7t [8]) );
  DRNQHSV1 \pe5/pe5/q_reg[29]  ( .D(pov4[29]), .CK(clk), .RDN(n59923), .Q(
        \pe5/pvq [29]) );
  DRNQHSV2 \pe5/pe5/q_reg[28]  ( .D(n60055), .CK(clk), .RDN(n59413), .Q(
        \pe5/pvq [28]) );
  DRNQHSV2 \pe5/pe5/q_reg[27]  ( .D(n60053), .CK(clk), .RDN(n59657), .Q(
        \pe5/pvq [27]) );
  DRNQHSV2 \pe5/pe5/q_reg[26]  ( .D(n60078), .CK(clk), .RDN(n59443), .Q(
        \pe5/pvq [26]) );
  DRNQHSV1 \pe5/pe5/q_reg[22]  ( .D(n60045), .CK(clk), .RDN(n59467), .Q(
        \pe5/pvq [22]) );
  DRNQHSV1 \pe5/pe5/q_reg[16]  ( .D(pov4[16]), .CK(clk), .RDN(n59401), .Q(
        \pe5/pvq [16]) );
  DRNQHSV1 \pe5/pe5/q_reg[14]  ( .D(n60042), .CK(clk), .RDN(n59455), .Q(
        \pe5/pvq [14]) );
  DRNQHSV1 \pe5/pe14/q_reg[8]  ( .D(n59381), .CK(clk), .RDN(n59479), .Q(
        \pe5/ti_7t [8]) );
  DRNQHSV2 \pe6/pe5/q_reg[29]  ( .D(n60006), .CK(clk), .RDN(n59425), .Q(
        \pe6/pvq [29]) );
  DRNQHSV1 \pe6/pe5/q_reg[28]  ( .D(n60000), .CK(clk), .RDN(n59430), .Q(
        \pe6/pvq [28]) );
  DRNQHSV2 \pe6/pe5/q_reg[27]  ( .D(pov5[27]), .CK(clk), .RDN(n59659), .Q(
        \pe6/pvq [27]) );
  DRNQHSV1 \pe6/pe5/q_reg[26]  ( .D(n59423), .CK(clk), .RDN(n59417), .Q(
        \pe6/pvq [26]) );
  DRNQHSV1 \pe6/pe5/q_reg[25]  ( .D(n60068), .CK(clk), .RDN(n59649), .Q(
        \pe6/pvq [25]) );
  DRNQHSV1 \pe6/pe5/q_reg[21]  ( .D(n60025), .CK(clk), .RDN(n59465), .Q(
        \pe6/pvq [21]) );
  DRNQHSV1 \pe6/pe5/q_reg[20]  ( .D(pov5[20]), .CK(clk), .RDN(n59658), .Q(
        \pe6/pvq [20]) );
  DRNQHSV1 \pe3/pe14/q_reg[5]  ( .D(n55951), .CK(clk), .RDN(n59470), .Q(
        \pe3/ti_7t [5]) );
  DRNQHSV1 \pe4/pe14/q_reg[7]  ( .D(n59681), .CK(clk), .RDN(n59453), .Q(
        \pe4/ti_7t [7]) );
  DRNQHSV1 \pe3/pe14/q_reg[8]  ( .D(n59581), .CK(clk), .RDN(n59472), .Q(
        \pe3/ti_7t [8]) );
  DRNQHSV1 \pe6/pe14/q_reg[6]  ( .D(n59597), .CK(clk), .RDN(n59451), .Q(
        \pe6/ti_7t [6]) );
  DRNQHSV2 \pe6/pe14/q_reg[7]  ( .D(n59678), .CK(clk), .RDN(n59396), .Q(
        \pe6/ti_7t [7]) );
  DRNQHSV1 \pe5/pe14/q_reg[5]  ( .D(n59936), .CK(clk), .RDN(n59400), .Q(
        \pe5/ti_7t [5]) );
  DRNQHSV1 \pe2/pe14/q_reg[6]  ( .D(n45150), .CK(clk), .RDN(n59442), .Q(
        \pe2/ti_7t [6]) );
  DRNQHSV1 \pe4/pe14/q_reg[9]  ( .D(n59682), .CK(clk), .RDN(n59410), .Q(
        \pe4/ti_7t [9]) );
  DRNQHSV1 \pe4/pe14/q_reg[6]  ( .D(n59667), .CK(clk), .RDN(n59416), .Q(
        \pe4/ti_7t [6]) );
  DRNQHSV1 \pe6/pe14/q_reg[9]  ( .D(n26109), .CK(clk), .RDN(n59417), .Q(
        \pe6/ti_7t [9]) );
  DRNQHSV1 \pe1/pe14/q_reg[2]  ( .D(n59590), .CK(clk), .RDN(n59448), .Q(
        \pe1/ti_7t [2]) );
  DRNQHSV1 \pe5/pe14/q_reg[4]  ( .D(n59639), .CK(clk), .RDN(n59651), .Q(
        \pe5/ti_7t [4]) );
  DRNQHSV1 \pe6/pe14/q_reg[3]  ( .D(n59594), .CK(clk), .RDN(n59460), .Q(
        \pe6/ti_7t [3]) );
  DRNQHSV1 \pe2/pe5/q_reg[13]  ( .D(n59576), .CK(clk), .RDN(n59411), .Q(
        \pe2/pvq [13]) );
  DRNQHSV1 \pe2/pe5/q_reg[10]  ( .D(n60008), .CK(clk), .RDN(n59437), .Q(
        \pe2/pvq [10]) );
  DRNQHSV1 \pe2/pe5/q_reg[8]  ( .D(n59504), .CK(clk), .RDN(n59925), .Q(
        \pe2/pvq [8]) );
  DRNQHSV1 \pe2/pe5/q_reg[5]  ( .D(n59498), .CK(clk), .RDN(n59425), .Q(
        \pe2/pvq [5]) );
  DRNQHSV1 \pe2/pe5/q_reg[4]  ( .D(n60108), .CK(clk), .RDN(n59450), .Q(
        \pe2/pvq [4]) );
  DRNQHSV1 \pe2/pe5/q_reg[3]  ( .D(n60009), .CK(clk), .RDN(n59449), .Q(
        \pe2/pvq [3]) );
  DRNQHSV1 \pe3/pe5/q_reg[14]  ( .D(n60020), .CK(clk), .RDN(n59417), .Q(
        \pe3/pvq [14]) );
  DRNQHSV1 \pe3/pe5/q_reg[10]  ( .D(n60019), .CK(clk), .RDN(n59402), .Q(
        \pe3/pvq [10]) );
  DRNQHSV1 \pe3/pe5/q_reg[7]  ( .D(n60005), .CK(clk), .RDN(n59459), .Q(
        \pe3/pvq [7]) );
  DRNQHSV1 \pe3/pe5/q_reg[6]  ( .D(n60004), .CK(clk), .RDN(n59655), .Q(
        \pe3/pvq [6]) );
  DRNQHSV1 \pe3/pe5/q_reg[2]  ( .D(n60003), .CK(clk), .RDN(n59649), .Q(
        \pe3/pvq [2]) );
  DRNQHSV1 \pe3/pe14/q_reg[4]  ( .D(n59621), .CK(clk), .RDN(n59480), .Q(
        \pe3/ti_7t [4]) );
  DRNQHSV1 \pe4/pe5/q_reg[14]  ( .D(n60088), .CK(clk), .RDN(n59492), .Q(
        \pe4/pvq [14]) );
  DRNQHSV1 \pe4/pe5/q_reg[12]  ( .D(n60046), .CK(clk), .RDN(n59512), .Q(
        \pe4/pvq [12]) );
  DRNQHSV1 \pe4/pe5/q_reg[6]  ( .D(n60024), .CK(clk), .RDN(n59430), .Q(
        \pe4/pvq [6]) );
  DRNQHSV1 \pe5/pe5/q_reg[11]  ( .D(n60031), .CK(clk), .RDN(n59405), .Q(
        \pe5/pvq [11]) );
  DRNQHSV1 \pe5/pe5/q_reg[9]  ( .D(n60038), .CK(clk), .RDN(n59442), .Q(
        \pe5/pvq [9]) );
  DRNQHSV1 \pe5/pe5/q_reg[5]  ( .D(n60082), .CK(clk), .RDN(n59478), .Q(
        \pe5/pvq [5]) );
  DRNQHSV1 \pe6/pe5/q_reg[15]  ( .D(n60035), .CK(clk), .RDN(n59433), .Q(
        \pe6/pvq [15]) );
  DRNQHSV1 \pe6/pe5/q_reg[13]  ( .D(n60041), .CK(clk), .RDN(n59482), .Q(
        \pe6/pvq [13]) );
  DRNQHSV1 \pe6/pe5/q_reg[11]  ( .D(n59426), .CK(clk), .RDN(n59463), .Q(
        \pe6/pvq [11]) );
  DRNQHSV1 \pe6/pe5/q_reg[6]  ( .D(n60074), .CK(clk), .RDN(n59463), .Q(
        \pe6/pvq [6]) );
  DRNQHSV1 \pe6/pe5/q_reg[5]  ( .D(n60040), .CK(clk), .RDN(n59494), .Q(
        \pe6/pvq [5]) );
  DRNQHSV1 \pe6/pe5/q_reg[4]  ( .D(n60037), .CK(clk), .RDN(n59412), .Q(
        \pe6/pvq [4]) );
  DRNQHSV1 \pe1/pe14/q_reg[3]  ( .D(n59529), .CK(clk), .RDN(n59439), .Q(
        \pe1/ti_7t [3]) );
  DRNQHSV1 \pe2/pe14/q_reg[1]  ( .D(n39061), .CK(clk), .RDN(n59414), .Q(
        \pe2/ti_7t [1]) );
  DRNQHSV1 \pe5/pe14/q_reg[1]  ( .D(n59393), .CK(clk), .RDN(n59413), .Q(
        \pe5/ti_7t [1]) );
  DRNQHSV1 \pe6/pe14/q_reg[1]  ( .D(n31325), .CK(clk), .RDN(n59473), .Q(
        \pe6/ti_7t [1]) );
  DRNQHSV1 \pe5/pe14/q_reg[3]  ( .D(n40187), .CK(clk), .RDN(n59460), .Q(
        \pe5/ti_7t [3]) );
  DRNQHSV1 \pe4/pe17/q_reg[18]  ( .D(\pe4/poht [18]), .CK(clk), .RDN(n59405), 
        .Q(poh4[18]) );
  DRNQHSV4 \pe5/pe5/q_reg[25]  ( .D(n29768), .CK(clk), .RDN(n59925), .Q(
        \pe5/pvq [25]) );
  DRNQHSV1 \pe2/pe17/q_reg[10]  ( .D(\pe2/poht [10]), .CK(clk), .RDN(n59418), 
        .Q(poh2[10]) );
  DRNQHSV2 \pe2/pe14/q_reg[30]  ( .D(n25709), .CK(clk), .RDN(n59412), .Q(
        \pe2/ti_7t [30]) );
  DRNQHSV1 \pe3/pe17/q_reg[4]  ( .D(\pe3/poht [4]), .CK(clk), .RDN(n59469), 
        .Q(poh3[4]) );
  DRNQHSV2 \pe6/pe14/q_reg[14]  ( .D(n49667), .CK(clk), .RDN(n59451), .Q(
        \pe6/ti_7t [14]) );
  DRNQHSV4 \pe4/pe14/q_reg[19]  ( .D(n59665), .CK(clk), .RDN(n59654), .Q(
        \pe4/ti_7t [19]) );
  DRNQHSV2 \pe6/pe5/q_reg[31]  ( .D(pov5[31]), .CK(clk), .RDN(n59650), .Q(
        \pe6/pvq [31]) );
  DRNQHSV1 \pe4/pe17/q_reg[31]  ( .D(\pe4/poht [31]), .CK(clk), .RDN(n59657), 
        .Q(poh4[31]) );
  DRNQHSV1 \pe1/pe17/q_reg[31]  ( .D(\pe1/poht [31]), .CK(clk), .RDN(n59659), 
        .Q(poh1[31]) );
  DRNQHSV4 \pe4/pe8/q_reg  ( .D(n59486), .CK(clk), .RDN(n59923), .Q(ctro4) );
  DRNQHSV2 \pe6/pe17/q_reg[16]  ( .D(\pe6/poht [16]), .CK(clk), .RDN(n59459), 
        .Q(poh6[16]) );
  DRNQHSV1 \pe4/pe4/q_reg  ( .D(po3), .CK(clk), .RDN(n59478), .Q(\pe4/pq ) );
  DRNQHSV4 \pe6/pe8/q_reg  ( .D(n59902), .CK(clk), .RDN(n59925), .Q(ctro6) );
  DRNQHSV1 \pe4/pe17/q_reg[26]  ( .D(\pe4/poht [26]), .CK(clk), .RDN(n59657), 
        .Q(poh4[26]) );
  DRNQHSV1 \pe4/pe17/q_reg[14]  ( .D(\pe4/poht [14]), .CK(clk), .RDN(n59438), 
        .Q(poh4[14]) );
  DRNQHSV1 \pe4/pe17/q_reg[30]  ( .D(\pe4/poht [30]), .CK(clk), .RDN(n59512), 
        .Q(poh4[30]) );
  DRNQHSV1 \pe4/pe17/q_reg[21]  ( .D(\pe4/poht [21]), .CK(clk), .RDN(n59435), 
        .Q(poh4[21]) );
  DRNQHSV1 \pe4/pe17/q_reg[23]  ( .D(\pe4/poht [23]), .CK(clk), .RDN(n59397), 
        .Q(poh4[23]) );
  DRNQHSV1 \pe4/pe17/q_reg[22]  ( .D(\pe4/poht [22]), .CK(clk), .RDN(n59494), 
        .Q(poh4[22]) );
  DRNQHSV1 \pe4/pe17/q_reg[17]  ( .D(\pe4/poht [17]), .CK(clk), .RDN(n59442), 
        .Q(poh4[17]) );
  DRNQHSV1 \pe3/pe17/q_reg[21]  ( .D(\pe3/poht [21]), .CK(clk), .RDN(n59449), 
        .Q(poh3[21]) );
  DRNQHSV1 \pe3/pe17/q_reg[18]  ( .D(\pe3/poht [18]), .CK(clk), .RDN(n59438), 
        .Q(poh3[18]) );
  DRNQHSV1 \pe3/pe17/q_reg[23]  ( .D(\pe3/poht [23]), .CK(clk), .RDN(n59437), 
        .Q(poh3[23]) );
  DRNQHSV1 \pe3/pe17/q_reg[15]  ( .D(\pe3/poht [15]), .CK(clk), .RDN(n59413), 
        .Q(poh3[15]) );
  DRNQHSV1 \pe3/pe17/q_reg[20]  ( .D(\pe3/poht [20]), .CK(clk), .RDN(n59488), 
        .Q(poh3[20]) );
  DRNQHSV1 \pe3/pe17/q_reg[25]  ( .D(\pe3/poht [25]), .CK(clk), .RDN(n59425), 
        .Q(poh3[25]) );
  DRNQHSV1 \pe3/pe17/q_reg[29]  ( .D(\pe3/poht [29]), .CK(clk), .RDN(n59652), 
        .Q(poh3[29]) );
  DRNQHSV1 \pe3/pe17/q_reg[13]  ( .D(\pe3/poht [13]), .CK(clk), .RDN(n59412), 
        .Q(poh3[13]) );
  DRNQHSV1 \pe3/pe17/q_reg[3]  ( .D(\pe3/poht [3]), .CK(clk), .RDN(n59923), 
        .Q(poh3[3]) );
  DRNQHSV4 \pe2/pe17/q_reg[11]  ( .D(\pe2/poht [11]), .CK(clk), .RDN(n59467), 
        .Q(poh2[11]) );
  DRNQHSV4 \pe2/pe17/q_reg[5]  ( .D(\pe2/poht [5]), .CK(clk), .RDN(n59416), 
        .Q(poh2[5]) );
  DRNQHSV4 \pe2/pe17/q_reg[12]  ( .D(\pe2/poht [12]), .CK(clk), .RDN(n59465), 
        .Q(poh2[12]) );
  DRNQHSV1 \pe1/pe17/q_reg[30]  ( .D(\pe1/poht [30]), .CK(clk), .RDN(n59476), 
        .Q(poh1[30]) );
  DRNQHSV4 \pe2/pe17/q_reg[16]  ( .D(\pe2/poht [16]), .CK(clk), .RDN(n59651), 
        .Q(poh2[16]) );
  DRNQHSV1 \pe6/pe17/q_reg[1]  ( .D(\pe6/poht [1]), .CK(clk), .RDN(n59443), 
        .Q(poh6[1]) );
  DRNQHSV1 \pe6/pe17/q_reg[3]  ( .D(\pe6/poht [3]), .CK(clk), .RDN(n59446), 
        .Q(poh6[3]) );
  DRNQHSV1 \pe6/pe17/q_reg[27]  ( .D(\pe6/poht [27]), .CK(clk), .RDN(n59455), 
        .Q(poh6[27]) );
  DRNQHSV1 \pe6/pe17/q_reg[21]  ( .D(\pe6/poht [21]), .CK(clk), .RDN(n59480), 
        .Q(poh6[21]) );
  DRNQHSV1 \pe6/pe17/q_reg[17]  ( .D(\pe6/poht [17]), .CK(clk), .RDN(n59922), 
        .Q(poh6[17]) );
  DRNQHSV1 \pe6/pe17/q_reg[8]  ( .D(\pe6/poht [8]), .CK(clk), .RDN(n59435), 
        .Q(poh6[8]) );
  DRNQHSV1 \pe6/pe17/q_reg[26]  ( .D(\pe6/poht [26]), .CK(clk), .RDN(n59460), 
        .Q(poh6[26]) );
  DRNQHSV1 \pe6/pe17/q_reg[28]  ( .D(\pe6/poht [28]), .CK(clk), .RDN(n59650), 
        .Q(poh6[28]) );
  DRNQHSV2 \pe6/pe17/q_reg[14]  ( .D(\pe6/poht [14]), .CK(clk), .RDN(n59439), 
        .Q(poh6[14]) );
  DRNQHSV2 \pe6/pe17/q_reg[13]  ( .D(\pe6/poht [13]), .CK(clk), .RDN(n59419), 
        .Q(poh6[13]) );
  DRNQHSV2 \pe6/pe17/q_reg[9]  ( .D(\pe6/poht [9]), .CK(clk), .RDN(n59461), 
        .Q(poh6[9]) );
  DRNQHSV1 \pe6/pe17/q_reg[30]  ( .D(\pe6/poht [30]), .CK(clk), .RDN(n59450), 
        .Q(poh6[30]) );
  DRNQHSV1 \pe6/pe17/q_reg[25]  ( .D(\pe6/poht [25]), .CK(clk), .RDN(n59493), 
        .Q(poh6[25]) );
  DRNQHSV1 \pe6/pe17/q_reg[29]  ( .D(\pe6/poht [29]), .CK(clk), .RDN(n59482), 
        .Q(poh6[29]) );
  DRNQHSV1 \pe6/pe17/q_reg[20]  ( .D(\pe6/poht [20]), .CK(clk), .RDN(n59446), 
        .Q(poh6[20]) );
  DRNQHSV4 \pe3/pe14/q_reg[27]  ( .D(n25989), .CK(clk), .RDN(n59476), .Q(
        \pe3/ti_7t [27]) );
  DSNHSV4 \pe4/pe5/q_reg[2]  ( .D(n59533), .CK(clk), .SDN(n59652), .QN(
        \pe4/pvq [2]) );
  DSNHSV4 \pe4/pe5/q_reg[7]  ( .D(n59569), .CK(clk), .SDN(n59652), .QN(
        \pe4/pvq [7]) );
  DSNHSV4 \pe3/pe13/q_reg  ( .D(\pe3/ti_1t ), .CK(clk), .SDN(rst), .Q(n59607), 
        .QN(\pe3/ti_1 ) );
  DSNHSV4 \pe3/pe2/q_reg[2]  ( .D(n59532), .CK(clk), .SDN(n59429), .Q(n59615), 
        .QN(\pe3/got [31]) );
  DSNHSV4 \pe3/pe1/q_reg[1]  ( .D(n59531), .CK(clk), .SDN(n59415), .Q(n59606), 
        .QN(\pe3/aot [32]) );
  DSNHSV4 \pe4/pe5/q_reg[1]  ( .D(n59530), .CK(clk), .SDN(n59492), .QN(
        \pe4/pvq [1]) );
  DRNQHSV1 \pe3/pe17/q_reg[1]  ( .D(\pe3/poht [1]), .CK(clk), .RDN(n59406), 
        .Q(poh3[1]) );
  DRNQHSV2 \pe5/pe15/q_reg[22]  ( .D(n59897), .CK(clk), .RDN(n59436), .Q(
        ao5[11]) );
  DRNQHSV2 \pe2/pe17/q_reg[20]  ( .D(\pe2/poht [20]), .CK(clk), .RDN(n59409), 
        .Q(poh2[20]) );
  DRNQHSV4 \pe1/pe3/q_reg[5]  ( .D(bi[28]), .CK(clk), .RDN(n59432), .Q(bo1[28]) );
  DRNQHSV4 \pe1/pe3/q_reg[2]  ( .D(bi[31]), .CK(clk), .RDN(rst), .Q(bo1[31])
         );
  DRNQHSV2 \pe1/pe14/q_reg[22]  ( .D(n59422), .CK(clk), .RDN(n59403), .Q(
        \pe1/ti_7t [22]) );
  DRNQHSV2 \pe2/pe17/q_reg[22]  ( .D(\pe2/poht [22]), .CK(clk), .RDN(n59477), 
        .Q(poh2[22]) );
  DRNQHSV1 \pe1/pe17/q_reg[8]  ( .D(\pe1/poht [8]), .CK(clk), .RDN(n59456), 
        .Q(poh1[8]) );
  DRNQHSV1 \pe1/pe17/q_reg[9]  ( .D(\pe1/poht [9]), .CK(clk), .RDN(n59418), 
        .Q(poh1[9]) );
  DRNQHSV1 \pe1/pe17/q_reg[24]  ( .D(\pe1/poht [24]), .CK(clk), .RDN(n59425), 
        .Q(poh1[24]) );
  DRNQHSV4 \pe3/pe14/q_reg[6]  ( .D(n59626), .CK(clk), .RDN(n59406), .Q(
        \pe3/ti_7t [6]) );
  DRNQHSV1 \pe1/pe17/q_reg[21]  ( .D(\pe1/poht [21]), .CK(clk), .RDN(n59474), 
        .Q(poh1[21]) );
  DRNQHSV1 \pe1/pe17/q_reg[18]  ( .D(\pe1/poht [18]), .CK(clk), .RDN(n59399), 
        .Q(poh1[18]) );
  DRNQHSV1 \pe1/pe17/q_reg[20]  ( .D(\pe1/poht [20]), .CK(clk), .RDN(n59472), 
        .Q(poh1[20]) );
  DRNQHSV1 \pe1/pe17/q_reg[27]  ( .D(\pe1/poht [27]), .CK(clk), .RDN(n59418), 
        .Q(poh1[27]) );
  DRNQHSV1 \pe1/pe17/q_reg[17]  ( .D(\pe1/poht [17]), .CK(clk), .RDN(n59923), 
        .Q(poh1[17]) );
  DRNQHSV1 \pe1/pe17/q_reg[12]  ( .D(\pe1/poht [12]), .CK(clk), .RDN(n59406), 
        .Q(poh1[12]) );
  DRNQHSV4 \pe5/pe3/q_reg[14]  ( .D(bo4[19]), .CK(clk), .RDN(n59434), .Q(
        bo5[19]) );
  DRNQHSV4 \pe5/pe3/q_reg[11]  ( .D(bo4[22]), .CK(clk), .RDN(n59473), .Q(
        bo5[22]) );
  DRNQHSV4 \pe6/pe14/q_reg[11]  ( .D(n59363), .CK(clk), .RDN(n59462), .Q(
        \pe6/ti_7t [11]) );
  DRNQHSV2 \pe1/pe16/q_reg[24]  ( .D(n55331), .CK(clk), .RDN(n59653), .Q(
        go1[9]) );
  DRNQHSV2 \pe1/pe15/q_reg[32]  ( .D(n59373), .CK(clk), .RDN(n59455), .Q(
        ao1[1]) );
  DRNQHSV4 \pe1/pe7/q_reg  ( .D(ctr), .CK(clk), .RDN(n59502), .Q(\pe1/ctrq )
         );
  DRNQHSV2 \pe1/pe16/q_reg[32]  ( .D(n59755), .CK(clk), .RDN(n59925), .Q(
        go1[1]) );
  DRNQHSV2 \pe1/pe15/q_reg[12]  ( .D(n59987), .CK(clk), .RDN(n59925), .Q(
        ao1[21]) );
  DRNQHSV4 \pe1/pe3/q_reg[9]  ( .D(bi[24]), .CK(clk), .RDN(rst), .Q(bo1[24])
         );
  DRNQHSV4 \pe1/pe3/q_reg[10]  ( .D(bi[23]), .CK(clk), .RDN(rst), .Q(bo1[23])
         );
  DRNQHSV4 \pe3/pe5/q_reg[4]  ( .D(n59509), .CK(clk), .RDN(n59450), .Q(
        \pe3/pvq [4]) );
  DRNQHSV2 \pe1/pe15/q_reg[14]  ( .D(n59737), .CK(clk), .RDN(n59479), .Q(
        ao1[19]) );
  DRNQHSV2 \pe1/pe16/q_reg[21]  ( .D(n55087), .CK(clk), .RDN(n59502), .Q(
        go1[12]) );
  DRNQHSV2 \pe1/pe16/q_reg[22]  ( .D(n54970), .CK(clk), .RDN(n59480), .Q(
        go1[11]) );
  DRNQHSV2 \pe1/pe15/q_reg[21]  ( .D(n44533), .CK(clk), .RDN(n59431), .Q(
        ao1[12]) );
  DRNQHSV4 \pe1/pe3/q_reg[1]  ( .D(bi[32]), .CK(clk), .RDN(n29734), .Q(bo1[32]) );
  DRNQHSV4 \pe1/pe3/q_reg[27]  ( .D(bi[6]), .CK(clk), .RDN(n29733), .Q(bo1[6])
         );
  DRNQHSV4 \pe1/pe3/q_reg[28]  ( .D(bi[5]), .CK(clk), .RDN(n59452), .Q(bo1[5])
         );
  DRNQHSV2 \pe1/pe15/q_reg[29]  ( .D(n59619), .CK(clk), .RDN(n59439), .Q(
        ao1[4]) );
  DRNQHSV4 \pe1/pe3/q_reg[11]  ( .D(bi[22]), .CK(clk), .RDN(n59440), .Q(
        bo1[22]) );
  DRNQHSV4 \pe1/pe3/q_reg[12]  ( .D(bi[21]), .CK(clk), .RDN(n59411), .Q(
        bo1[21]) );
  DRNQHSV2 \pe1/pe14/q_reg[5]  ( .D(n40552), .CK(clk), .RDN(n59446), .Q(
        \pe1/ti_7t [5]) );
  DRNQHSV4 \pe1/pe3/q_reg[22]  ( .D(bi[11]), .CK(clk), .RDN(rst), .Q(bo1[11])
         );
  DRNQHSV1 \pe1/pe14/q_reg[6]  ( .D(n59686), .CK(clk), .RDN(n59444), .Q(
        \pe1/ti_7t [6]) );
  DRNQHSV4 \pe4/pe14/q_reg[3]  ( .D(n59501), .CK(clk), .RDN(n59657), .Q(
        \pe4/ti_7t [3]) );
  DRNQHSV1 \pe1/pe14/q_reg[27]  ( .D(n59931), .CK(clk), .RDN(n59403), .Q(
        \pe1/ti_7t [27]) );
  DRNQHSV1 \pe4/pe17/q_reg[29]  ( .D(\pe4/poht [29]), .CK(clk), .RDN(n59484), 
        .Q(poh4[29]) );
  DRNQHSV2 \pe3/pe14/q_reg[25]  ( .D(n59527), .CK(clk), .RDN(n59403), .Q(
        \pe3/ti_7t [25]) );
  DRNQHSV4 \pe1/pe14/q_reg[13]  ( .D(n59725), .CK(clk), .RDN(n59439), .Q(
        \pe1/ti_7t [13]) );
  DRNQHSV4 \pe1/pe3/q_reg[19]  ( .D(bi[14]), .CK(clk), .RDN(n29732), .Q(
        bo1[14]) );
  DRNQHSV4 \pe1/pe3/q_reg[18]  ( .D(bi[15]), .CK(clk), .RDN(rst), .Q(bo1[15])
         );
  DRNQHSV4 \pe1/pe3/q_reg[8]  ( .D(bi[25]), .CK(clk), .RDN(n59925), .Q(bo1[25]) );
  DRNQHSV4 \pe1/pe3/q_reg[29]  ( .D(bi[4]), .CK(clk), .RDN(n59407), .Q(bo1[4])
         );
  DRNQHSV4 \pe3/pe3/q_reg[1]  ( .D(bo2[32]), .CK(clk), .RDN(n59493), .Q(
        bo3[32]) );
  DRNQHSV2 \pe3/pe16/q_reg[5]  ( .D(n59964), .CK(clk), .RDN(n59503), .Q(
        go3[28]) );
  DRNQHSV2 \pe2/pe14/q_reg[11]  ( .D(n51966), .CK(clk), .RDN(n59410), .Q(
        \pe2/ti_7t [11]) );
  DRNQHSV4 \pe1/pe1/q_reg[31]  ( .D(ai[2]), .CK(clk), .RDN(rst), .Q(
        \pe1/aot [2]) );
  DRNQHSV4 \pe2/pe3/q_reg[18]  ( .D(bo1[15]), .CK(clk), .RDN(n59462), .Q(
        bo2[15]) );
  DRNQHSV4 \pe2/pe3/q_reg[19]  ( .D(bo1[14]), .CK(clk), .RDN(n59650), .Q(
        bo2[14]) );
  DRNQHSV4 \pe3/pe3/q_reg[11]  ( .D(bo2[22]), .CK(clk), .RDN(n59408), .Q(
        bo3[22]) );
  DRNQHSV4 \pe3/pe3/q_reg[12]  ( .D(bo2[21]), .CK(clk), .RDN(n59411), .Q(
        bo3[21]) );
  DRNQHSV4 \pe3/pe3/q_reg[5]  ( .D(bo2[28]), .CK(clk), .RDN(n29730), .Q(
        bo3[28]) );
  DRNQHSV2 \pe4/pe15/q_reg[7]  ( .D(n59661), .CK(clk), .RDN(n59425), .Q(
        ao4[26]) );
  DRNQHSV1 \pe1/pe17/q_reg[2]  ( .D(\pe1/poht [2]), .CK(clk), .RDN(n59439), 
        .Q(poh1[2]) );
  DRNQHSV1 \pe1/pe17/q_reg[5]  ( .D(\pe1/poht [5]), .CK(clk), .RDN(n59412), 
        .Q(poh1[5]) );
  DRNQHSV2 \pe3/pe16/q_reg[4]  ( .D(n59963), .CK(clk), .RDN(n59451), .Q(
        go3[29]) );
  DRNQHSV1 \pe3/pe17/q_reg[31]  ( .D(\pe3/poht [31]), .CK(clk), .RDN(n59407), 
        .Q(poh3[31]) );
  DRNQHSV1 \pe2/pe17/q_reg[15]  ( .D(\pe2/poht [15]), .CK(clk), .RDN(n59473), 
        .Q(poh2[15]) );
  DRNQHSV1 \pe3/pe5/q_reg[25]  ( .D(n60051), .CK(clk), .RDN(n59399), .Q(
        \pe3/pvq [25]) );
  DRNQHSV1 \pe1/pe17/q_reg[10]  ( .D(\pe1/poht [10]), .CK(clk), .RDN(n59399), 
        .Q(poh1[10]) );
  DRNQHSV1 \pe6/pe5/q_reg[23]  ( .D(n59573), .CK(clk), .RDN(n59415), .Q(
        \pe6/pvq [23]) );
  DRNQHSV1 \pe4/pe17/q_reg[24]  ( .D(\pe4/poht [24]), .CK(clk), .RDN(n59490), 
        .Q(poh4[24]) );
  DRNQHSV1 \pe1/pe14/q_reg[19]  ( .D(n59360), .CK(clk), .RDN(n59492), .Q(
        \pe1/ti_7t [19]) );
  DRNQHSV1 \pe1/pe14/q_reg[4]  ( .D(n59674), .CK(clk), .RDN(n59924), .Q(
        \pe1/ti_7t [4]) );
  DRNQHSV1 \pe4/pe17/q_reg[28]  ( .D(\pe4/poht [28]), .CK(clk), .RDN(n59404), 
        .Q(poh4[28]) );
  DRNQHSV4 \pe1/pe12/q_reg[15]  ( .D(n59704), .CK(clk), .RDN(n59494), .Q(
        \pe1/bq[18] ) );
  DRNQHSV1 \pe3/pe17/q_reg[16]  ( .D(\pe3/poht [16]), .CK(clk), .RDN(n59925), 
        .Q(poh3[16]) );
  DRNQHSV1 \pe1/pe14/q_reg[21]  ( .D(n59377), .CK(clk), .RDN(n59503), .Q(
        \pe1/ti_7t [21]) );
  DRNQHSV2 \pe4/pe15/q_reg[13]  ( .D(n59839), .CK(clk), .RDN(n59435), .Q(
        ao4[20]) );
  DRNQHSV1 \pe4/pe17/q_reg[5]  ( .D(\pe4/poht [5]), .CK(clk), .RDN(n59438), 
        .Q(poh4[5]) );
  DRNQHSV1 \pe4/pe17/q_reg[4]  ( .D(\pe4/poht [4]), .CK(clk), .RDN(n29732), 
        .Q(poh4[4]) );
  DRNQHSV1 \pe4/pe17/q_reg[8]  ( .D(\pe4/poht [8]), .CK(clk), .RDN(n59479), 
        .Q(poh4[8]) );
  DRNQHSV1 \pe5/pe17/q_reg[4]  ( .D(\pe5/poht [4]), .CK(clk), .RDN(n59425), 
        .Q(poh5[4]) );
  DRNQHSV1 \pe5/pe17/q_reg[8]  ( .D(\pe5/poht [8]), .CK(clk), .RDN(n59413), 
        .Q(poh5[8]) );
  DRNQHSV2 \pe2/pe15/q_reg[10]  ( .D(n59585), .CK(clk), .RDN(n59652), .Q(
        ao2[23]) );
  DRNQHSV2 \pe2/pe16/q_reg[30]  ( .D(n59351), .CK(clk), .RDN(n59396), .Q(
        go2[3]) );
  DRNQHSV2 \pe1/pe16/q_reg[2]  ( .D(n59365), .CK(clk), .RDN(n59405), .Q(
        go1[31]) );
  DRNQHSV1 \pe4/pe5/q_reg[4]  ( .D(n36775), .CK(clk), .RDN(n59470), .Q(
        \pe4/pvq [4]) );
  DRNQHSV1 \pe6/pe17/q_reg[5]  ( .D(\pe6/poht [5]), .CK(clk), .RDN(n59478), 
        .Q(poh6[5]) );
  DRNQHSV4 \pe6/pe5/q_reg[24]  ( .D(n60010), .CK(clk), .RDN(n59649), .Q(
        \pe6/pvq [24]) );
  DRNQHSV1 \pe6/pe5/q_reg[18]  ( .D(n60054), .CK(clk), .RDN(n59649), .Q(
        \pe6/pvq [18]) );
  DRNQHSV1 \pe1/pe17/q_reg[26]  ( .D(\pe1/poht [26]), .CK(clk), .RDN(n59396), 
        .Q(poh1[26]) );
  DRNQHSV1 \pe5/pe17/q_reg[1]  ( .D(\pe5/poht [1]), .CK(clk), .RDN(n29734), 
        .Q(poh5[1]) );
  DRNQHSV1 \pe1/pe17/q_reg[15]  ( .D(\pe1/poht [15]), .CK(clk), .RDN(n59454), 
        .Q(poh1[15]) );
  DRNQHSV1 \pe1/pe17/q_reg[4]  ( .D(\pe1/poht [4]), .CK(clk), .RDN(n59438), 
        .Q(poh1[4]) );
  DRNQHSV1 \pe1/pe15/q_reg[1]  ( .D(n59591), .CK(clk), .RDN(n59492), .Q(
        ao1[32]) );
  DSNHSV1 \pe5/pe15/q_reg[30]  ( .D(n59869), .CK(clk), .SDN(rst), .QN(ao5[3])
         );
  DSNHSV1 \pe4/pe15/q_reg[14]  ( .D(n57605), .CK(clk), .SDN(n59432), .QN(
        ao4[19]) );
  DSNHSV1 \pe4/pe15/q_reg[29]  ( .D(n57011), .CK(clk), .SDN(n59443), .QN(
        ao4[4]) );
  DSNHSV1 \pe4/pe16/q_reg[24]  ( .D(n59628), .CK(clk), .SDN(rst), .QN(go4[9])
         );
  DSNHSV1 \pe5/pe15/q_reg[19]  ( .D(n59641), .CK(clk), .SDN(n59471), .QN(
        ao5[14]) );
  DSNHSV1 \pe3/pe14/q_reg[13]  ( .D(n46519), .CK(clk), .SDN(n59479), .QN(
        \pe3/ti_7t [13]) );
  DRSNHSV4 \pe3/pe6/q_reg[1]  ( .D(poh2[1]), .CK(clk), .SDN(1'b1), .RDN(rst), 
        .QN(n59572) );
  DSNHSV4 \pe3/pe2/q_reg[1]  ( .D(n59341), .CK(clk), .SDN(rst), .Q(n59611), 
        .QN(\pe3/got [32]) );
  DRNQHSV2 \pe2/pe17/q_reg[19]  ( .D(\pe2/poht [19]), .CK(clk), .RDN(n59408), 
        .Q(poh2[19]) );
  DRNQHSV1 \pe1/pe16/q_reg[10]  ( .D(\pe1/got [23]), .CK(clk), .RDN(n29734), 
        .Q(go1[23]) );
  DRNQHSV4 \pe5/pe12/q_reg[30]  ( .D(n59864), .CK(clk), .RDN(n59470), .Q(
        \pe5/bq[3] ) );
  DRNQHSV1 \pe1/pe17/q_reg[28]  ( .D(\pe1/poht [28]), .CK(clk), .RDN(n59406), 
        .Q(poh1[28]) );
  DRNQHSV1 \pe1/pe17/q_reg[11]  ( .D(\pe1/poht [11]), .CK(clk), .RDN(n59432), 
        .Q(poh1[11]) );
  DRNQHSV2 \pe2/pe14/q_reg[4]  ( .D(n59669), .CK(clk), .RDN(n59481), .Q(
        \pe2/ti_7t [4]) );
  DRNQHSV2 \pe2/pe16/q_reg[10]  ( .D(n45249), .CK(clk), .RDN(n59483), .Q(
        go2[23]) );
  DRNQHSV2 \pe2/pe17/q_reg[23]  ( .D(n60016), .CK(clk), .RDN(n59483), .Q(
        poh2[23]) );
  DRNQHSV2 \pe2/pe17/q_reg[9]  ( .D(\pe2/poht [9]), .CK(clk), .RDN(n59483), 
        .Q(poh2[9]) );
  DRNQHSV1 \pe2/pe15/q_reg[6]  ( .D(n49530), .CK(clk), .RDN(n59650), .Q(
        ao2[27]) );
  DRNQHSV1 \pe1/pe17/q_reg[13]  ( .D(\pe1/poht [13]), .CK(clk), .RDN(n59463), 
        .Q(poh1[13]) );
  DRNQHSV1 \pe5/pe15/q_reg[1]  ( .D(n59366), .CK(clk), .RDN(n59473), .Q(
        ao5[32]) );
  DRNQHSV4 \pe6/pe3/q_reg[23]  ( .D(bo5[10]), .CK(clk), .RDN(n59472), .Q(
        bo6[10]) );
  DRNQHSV1 \pe2/pe14/q_reg[2]  ( .D(n59349), .CK(clk), .RDN(n59921), .Q(
        \pe2/ti_7t [2]) );
  DRNQHSV1 \pe2/pe17/q_reg[21]  ( .D(\pe2/poht [21]), .CK(clk), .RDN(n59503), 
        .Q(poh2[21]) );
  DRNQHSV2 \pe2/pe17/q_reg[1]  ( .D(\pe2/poht [1]), .CK(clk), .RDN(n59415), 
        .Q(poh2[1]) );
  DRNQHSV2 \pe2/pe17/q_reg[6]  ( .D(\pe2/poht [6]), .CK(clk), .RDN(n59415), 
        .Q(poh2[6]) );
  DRNQHSV1 \pe6/pe5/q_reg[1]  ( .D(n59398), .CK(clk), .RDN(n59434), .Q(
        \pe6/pvq [1]) );
  DRNQHSV1 \pe1/pe16/q_reg[16]  ( .D(n59996), .CK(clk), .RDN(n59463), .Q(
        go1[17]) );
  DRNQHSV2 \pe1/pe14/q_reg[28]  ( .D(n59489), .CK(clk), .RDN(n59474), .Q(
        \pe1/ti_7t [28]) );
  DRNQHSV2 \pe1/pe14/q_reg[7]  ( .D(n59919), .CK(clk), .RDN(n59453), .Q(
        \pe1/ti_7t [7]) );
  DRNQHSV2 \pe3/pe3/q_reg[3]  ( .D(bo2[30]), .CK(clk), .RDN(n59923), .Q(
        bo3[30]) );
  DSNHSV2 \pe4/pe5/q_reg[21]  ( .D(n59571), .CK(clk), .SDN(n59483), .QN(
        \pe4/pvq [21]) );
  DRNQHSV1 \pe1/pe15/q_reg[31]  ( .D(n59730), .CK(clk), .RDN(n59503), .Q(
        ao1[2]) );
  DRNQHSV1 \pe1/pe16/q_reg[20]  ( .D(n54812), .CK(clk), .RDN(n59503), .Q(
        go1[13]) );
  DRNQHSV1 \pe2/pe14/q_reg[19]  ( .D(n59361), .CK(clk), .RDN(n59418), .Q(
        \pe2/ti_7t [19]) );
  DRNQHSV1 \pe1/pe17/q_reg[25]  ( .D(\pe1/poht [25]), .CK(clk), .RDN(n59924), 
        .Q(poh1[25]) );
  DRNQHSV1 \pe5/pe14/q_reg[20]  ( .D(n59883), .CK(clk), .RDN(n59481), .Q(
        \pe5/ti_7t [20]) );
  DRNQHSV4 \pe2/pe12/q_reg[32]  ( .D(n59753), .CK(clk), .RDN(n59469), .Q(
        \pe2/bq[1] ) );
  DRNQHSV4 \pe2/pe1/q_reg[31]  ( .D(ao1[2]), .CK(clk), .RDN(n59431), .Q(
        \pe2/aot [2]) );
  DRNQHSV4 \pe1/pe12/q_reg[24]  ( .D(n59710), .CK(clk), .RDN(n59468), .Q(
        \pe1/bq[9] ) );
  DRNQHSV2 \pe2/pe5/q_reg[1]  ( .D(n60110), .CK(clk), .RDN(n59419), .Q(
        \pe2/pvq [1]) );
  DRNQHSV4 \pe1/pe12/q_reg[22]  ( .D(n59712), .CK(clk), .RDN(n59434), .Q(
        \pe1/bq[11] ) );
  DRNQHSV4 \pe1/pe12/q_reg[3]  ( .D(n59691), .CK(clk), .RDN(n59432), .Q(
        \pe1/bq[30] ) );
  DRNQHSV4 \pe5/pe7/q_reg  ( .D(n59997), .CK(clk), .RDN(n59419), .Q(\pe5/ctrq ) );
  DRNQHSV4 \pe1/pe12/q_reg[12]  ( .D(n59699), .CK(clk), .RDN(n59490), .Q(
        \pe1/bq[21] ) );
  DRNQHSV2 \pe2/pe14/q_reg[9]  ( .D(n45218), .CK(clk), .RDN(n59419), .Q(
        \pe2/ti_7t [9]) );
  DRNQHSV1 \pe4/pe14/q_reg[1]  ( .D(n33976), .CK(clk), .RDN(n59457), .Q(
        \pe4/ti_7t [1]) );
  DRNQHSV2 \pe5/pe14/q_reg[2]  ( .D(n37608), .CK(clk), .RDN(n59466), .Q(
        \pe5/ti_7t [2]) );
  DRNQHSV2 \pe4/pe14/q_reg[5]  ( .D(n59662), .CK(clk), .RDN(n59404), .Q(
        \pe4/ti_7t [5]) );
  DRNQHSV2 \pe5/pe17/q_reg[18]  ( .D(\pe5/poht [18]), .CK(clk), .RDN(n59464), 
        .Q(poh5[18]) );
  DRNQHSV2 \pe3/pe17/q_reg[6]  ( .D(\pe3/poht [6]), .CK(clk), .RDN(n59447), 
        .Q(poh3[6]) );
  DRNQHSV2 \pe6/pe14/q_reg[21]  ( .D(n59680), .CK(clk), .RDN(n59466), .Q(
        \pe6/ti_7t [21]) );
  DRNQHSV1 \pe5/pe8/q_reg  ( .D(n44335), .CK(clk), .RDN(n59496), .Q(ctro5) );
  DRNQHSV1 \pe4/pe5/q_reg[25]  ( .D(n59515), .CK(clk), .RDN(n59435), .Q(
        \pe4/pvq [25]) );
  DRNQHSV2 \pe3/pe5/q_reg[1]  ( .D(n60102), .CK(clk), .RDN(n59481), .Q(
        \pe3/pvq [1]) );
  DRNQHSV2 \pe5/pe17/q_reg[3]  ( .D(\pe5/poht [3]), .CK(clk), .RDN(n59477), 
        .Q(poh5[3]) );
  DRNQHSV2 \pe6/pe17/q_reg[22]  ( .D(\pe6/poht [22]), .CK(clk), .RDN(n59502), 
        .Q(poh6[22]) );
  DRNQHSV2 \pe2/pe5/q_reg[20]  ( .D(n60105), .CK(clk), .RDN(n59502), .Q(
        \pe2/pvq [20]) );
  DRNQHSV1 \pe5/pe14/q_reg[14]  ( .D(n44694), .CK(clk), .RDN(n59459), .Q(
        \pe5/ti_7t [14]) );
  DRNQHSV1 \pe4/pe17/q_reg[2]  ( .D(\pe4/poht [2]), .CK(clk), .RDN(n59462), 
        .Q(poh4[2]) );
  DRNQHSV2 \pe1/pe17/q_reg[23]  ( .D(\pe1/poht [23]), .CK(clk), .RDN(n59451), 
        .Q(poh1[23]) );
  DRNQHSV2 \pe1/pe17/q_reg[19]  ( .D(\pe1/poht [19]), .CK(clk), .RDN(n59924), 
        .Q(poh1[19]) );
  DRNQHSV2 \pe3/pe14/q_reg[30]  ( .D(n59823), .CK(clk), .RDN(n59402), .Q(
        \pe3/ti_7t [30]) );
  DRNQHSV2 \pe6/pe5/q_reg[30]  ( .D(n29761), .CK(clk), .RDN(n59650), .Q(
        \pe6/pvq [30]) );
  DRNQHSV1 \pe4/pe17/q_reg[19]  ( .D(\pe4/poht [19]), .CK(clk), .RDN(n59424), 
        .Q(poh4[19]) );
  DRNQHSV2 \pe6/pe17/q_reg[23]  ( .D(\pe6/poht [23]), .CK(clk), .RDN(n59447), 
        .Q(poh6[23]) );
  DRNQHSV2 \pe3/pe17/q_reg[5]  ( .D(\pe3/poht [5]), .CK(clk), .RDN(n59512), 
        .Q(poh3[5]) );
  DRNQHSV2 \pe3/pe17/q_reg[24]  ( .D(\pe3/poht [24]), .CK(clk), .RDN(n29729), 
        .Q(poh3[24]) );
  DRNQHSV2 \pe3/pe17/q_reg[8]  ( .D(\pe3/poht [8]), .CK(clk), .RDN(n29734), 
        .Q(poh3[8]) );
  DRNQHSV1 \pe3/pe17/q_reg[30]  ( .D(\pe3/poht [30]), .CK(clk), .RDN(n59456), 
        .Q(poh3[30]) );
  DRNQHSV2 \pe3/pe17/q_reg[28]  ( .D(\pe3/poht [28]), .CK(clk), .RDN(n59481), 
        .Q(poh3[28]) );
  DRNQHSV2 \pe3/pe17/q_reg[22]  ( .D(\pe3/poht [22]), .CK(clk), .RDN(n29734), 
        .Q(poh3[22]) );
  DRNQHSV2 \pe3/pe17/q_reg[17]  ( .D(\pe3/poht [17]), .CK(clk), .RDN(n59444), 
        .Q(poh3[17]) );
  DRNQHSV2 \pe6/pe17/q_reg[18]  ( .D(\pe6/poht [18]), .CK(clk), .RDN(n59923), 
        .Q(poh6[18]) );
  DRNQHSV2 \pe6/pe17/q_reg[19]  ( .D(\pe6/poht [19]), .CK(clk), .RDN(n59453), 
        .Q(poh6[19]) );
  DRNQHSV1 \pe4/pe17/q_reg[27]  ( .D(\pe4/poht [27]), .CK(clk), .RDN(n59654), 
        .Q(poh4[27]) );
  DRNQHSV1 \pe4/pe17/q_reg[25]  ( .D(\pe4/poht [25]), .CK(clk), .RDN(n59468), 
        .Q(poh4[25]) );
  DRNQHSV1 \pe4/pe17/q_reg[11]  ( .D(\pe4/poht [11]), .CK(clk), .RDN(n59467), 
        .Q(poh4[11]) );
  DRNQHSV1 \pe4/pe17/q_reg[20]  ( .D(\pe4/poht [20]), .CK(clk), .RDN(n59449), 
        .Q(poh4[20]) );
  DRNQHSV1 \pe4/pe17/q_reg[10]  ( .D(\pe4/poht [10]), .CK(clk), .RDN(n59405), 
        .Q(poh4[10]) );
  DRNQHSV1 \pe4/pe17/q_reg[6]  ( .D(\pe4/poht [6]), .CK(clk), .RDN(n59512), 
        .Q(poh4[6]) );
  DRNQHSV1 \pe5/pe4/q_reg  ( .D(po4), .CK(clk), .RDN(n59400), .Q(\pe5/pq ) );
  DRNQHSV1 \pe4/pe17/q_reg[9]  ( .D(\pe4/poht [9]), .CK(clk), .RDN(n59502), 
        .Q(poh4[9]) );
  DRNQHSV1 \pe4/pe17/q_reg[13]  ( .D(\pe4/poht [13]), .CK(clk), .RDN(n59659), 
        .Q(poh4[13]) );
  DRNQHSV1 \pe4/pe17/q_reg[15]  ( .D(\pe4/poht [15]), .CK(clk), .RDN(n59399), 
        .Q(poh4[15]) );
  DRNQHSV1 \pe4/pe17/q_reg[16]  ( .D(\pe4/poht [16]), .CK(clk), .RDN(n59649), 
        .Q(poh4[16]) );
  DRNQHSV1 \pe5/pe17/q_reg[29]  ( .D(\pe5/poht [29]), .CK(clk), .RDN(n59503), 
        .Q(poh5[29]) );
  DRNQHSV2 \pe6/pe17/q_reg[2]  ( .D(\pe6/poht [2]), .CK(clk), .RDN(n59656), 
        .Q(poh6[2]) );
  DRNQHSV2 \pe22/q_reg  ( .D(po6), .CK(clk), .RDN(n59443), .Q(po[1]) );
  DRNQHSV2 \pe1/pe17/q_reg[7]  ( .D(\pe1/poht [7]), .CK(clk), .RDN(n59439), 
        .Q(poh1[7]) );
  DRNQHSV2 \pe1/pe17/q_reg[16]  ( .D(\pe1/poht [16]), .CK(clk), .RDN(n59405), 
        .Q(poh1[16]) );
  DRNQHSV2 \pe2/pe17/q_reg[8]  ( .D(\pe2/poht [8]), .CK(clk), .RDN(n59924), 
        .Q(poh2[8]) );
  DRNQHSV2 \pe2/pe17/q_reg[30]  ( .D(\pe2/poht [30]), .CK(clk), .RDN(n59469), 
        .Q(poh2[30]) );
  DRNQHSV4 \pe5/pe5/q_reg[1]  ( .D(n59577), .CK(clk), .RDN(n59435), .Q(
        \pe5/pvq [1]) );
  DRNQHSV1 \pe4/pe17/q_reg[7]  ( .D(\pe4/poht [7]), .CK(clk), .RDN(n59925), 
        .Q(poh4[7]) );
  DRNQHSV1 \pe4/pe17/q_reg[12]  ( .D(\pe4/poht [12]), .CK(clk), .RDN(n59460), 
        .Q(poh4[12]) );
  DRNQHSV2 \pe1/pe17/q_reg[14]  ( .D(\pe1/poht [14]), .CK(clk), .RDN(n59457), 
        .Q(poh1[14]) );
  DRNQHSV2 \pe5/pe17/q_reg[10]  ( .D(\pe5/poht [10]), .CK(clk), .RDN(n59429), 
        .Q(poh5[10]) );
  DRNQHSV2 \pe5/pe17/q_reg[5]  ( .D(\pe5/poht [5]), .CK(clk), .RDN(n59658), 
        .Q(poh5[5]) );
  DRNQHSV2 \pe2/pe17/q_reg[24]  ( .D(\pe2/poht [24]), .CK(clk), .RDN(n59456), 
        .Q(poh2[24]) );
  DRNQHSV4 \pe6/pe17/q_reg[6]  ( .D(\pe6/poht [6]), .CK(clk), .RDN(n59406), 
        .Q(poh6[6]) );
  DRNQHSV2 \pe3/pe17/q_reg[7]  ( .D(\pe3/poht [7]), .CK(clk), .RDN(n59443), 
        .Q(poh3[7]) );
  DRNQHSV2 \pe2/pe17/q_reg[18]  ( .D(\pe2/poht [18]), .CK(clk), .RDN(n59435), 
        .Q(poh2[18]) );
  DRNQHSV1 \pe2/pe17/q_reg[17]  ( .D(\pe2/poht [17]), .CK(clk), .RDN(n59477), 
        .Q(poh2[17]) );
  DRNQHSV2 \pe6/pe17/q_reg[4]  ( .D(\pe6/poht [4]), .CK(clk), .RDN(n59483), 
        .Q(poh6[4]) );
  DRNQHSV4 \pe2/pe17/q_reg[2]  ( .D(\pe2/poht [2]), .CK(clk), .RDN(n59416), 
        .Q(poh2[2]) );
  DRNQHSV1 \pe3/pe17/q_reg[19]  ( .D(\pe3/poht [19]), .CK(clk), .RDN(n59417), 
        .Q(poh3[19]) );
  DRNQHSV2 \pe3/pe14/q_reg[19]  ( .D(n43463), .CK(clk), .RDN(n29732), .Q(
        \pe3/ti_7t [19]) );
  DRNQHSV1 \pe6/pe17/q_reg[15]  ( .D(\pe6/poht [15]), .CK(clk), .RDN(n59654), 
        .Q(poh6[15]) );
  DRNQHSV2 \pe6/pe17/q_reg[7]  ( .D(\pe6/poht [7]), .CK(clk), .RDN(n59425), 
        .Q(poh6[7]) );
  DRNQHSV4 \pe3/pe17/q_reg[26]  ( .D(\pe3/poht [26]), .CK(clk), .RDN(n59446), 
        .Q(poh3[26]) );
  DRNQHSV2 \pe2/pe17/q_reg[13]  ( .D(\pe2/poht [13]), .CK(clk), .RDN(n59456), 
        .Q(poh2[13]) );
  CLKNHSV4 U25899 ( .I(n42916), .ZN(n42925) );
  XNOR2HSV4 U25900 ( .A1(n26581), .A2(n26580), .ZN(n42916) );
  NOR2HSV4 U25901 ( .A1(n25137), .A2(n45621), .ZN(n42933) );
  XNOR2HSV4 U25902 ( .A1(n42915), .A2(n42925), .ZN(n25137) );
  CLKNAND2HSV2 U25903 ( .A1(n42784), .A2(n42785), .ZN(n42915) );
  CLKNAND2HSV2 U25904 ( .A1(n25138), .A2(n43128), .ZN(n43129) );
  CLKNAND2HSV2 U25905 ( .A1(n25151), .A2(n25138), .ZN(n25693) );
  INHSV2 U25906 ( .I(n43344), .ZN(n25138) );
  MOAI22HSV4 U25907 ( .A1(n25591), .A2(n26027), .B1(n31869), .B2(n32422), .ZN(
        n26026) );
  INHSV4 U25908 ( .I(n33602), .ZN(n59928) );
  NAND2HSV4 U25909 ( .A1(n26103), .A2(n31759), .ZN(n26102) );
  INHSV4 U25910 ( .I(n34457), .ZN(n34409) );
  CLKNAND2HSV2 U25911 ( .A1(n34409), .A2(n59350), .ZN(n34412) );
  MUX2NHSV2 U25912 ( .I0(n41216), .I1(n41215), .S(n41214), .ZN(n41224) );
  NAND2HSV4 U25913 ( .A1(n26481), .A2(n26482), .ZN(n42605) );
  NAND2HSV4 U25914 ( .A1(n25693), .A2(n25692), .ZN(n59536) );
  NAND2HSV4 U25915 ( .A1(n43895), .A2(n43894), .ZN(n43909) );
  CLKNAND2HSV2 U25916 ( .A1(n44678), .A2(n44677), .ZN(n44686) );
  NOR2HSV2 U25917 ( .A1(n45503), .A2(n43893), .ZN(n43894) );
  NAND2HSV4 U25918 ( .A1(n43908), .A2(n59515), .ZN(n45506) );
  INHSV6 U25919 ( .I(n43749), .ZN(n44683) );
  CLKNAND2HSV8 U25920 ( .A1(n45618), .A2(\pe3/ti_7t [25]), .ZN(n45596) );
  XNOR2HSV4 U25921 ( .A1(n43861), .A2(n43860), .ZN(n43863) );
  CLKNAND2HSV2 U25922 ( .A1(n43133), .A2(n42815), .ZN(n42816) );
  NAND2HSV4 U25923 ( .A1(n33153), .A2(n26182), .ZN(n26181) );
  NAND3HSV4 U25924 ( .A1(n26839), .A2(n41409), .A3(n40957), .ZN(n41595) );
  INHSV4 U25925 ( .I(n41595), .ZN(n41596) );
  XNOR2HSV4 U25926 ( .A1(n41818), .A2(n41817), .ZN(n41819) );
  INHSV2 U25927 ( .I(n25139), .ZN(n25768) );
  CLKNAND2HSV2 U25928 ( .A1(n43493), .A2(n43464), .ZN(n25139) );
  NAND2HSV4 U25929 ( .A1(n45102), .A2(n45101), .ZN(n44181) );
  XNOR2HSV4 U25930 ( .A1(n25957), .A2(n25956), .ZN(n45094) );
  CLKNAND2HSV4 U25931 ( .A1(n39378), .A2(n25140), .ZN(n51115) );
  NAND3HSV3 U25932 ( .A1(n39377), .A2(n39375), .A3(n39376), .ZN(n25140) );
  INHSV2 U25933 ( .I(n25763), .ZN(n43364) );
  NAND2HSV2 U25934 ( .A1(n25207), .A2(n25255), .ZN(n25763) );
  INAND2HSV4 U25935 ( .A1(n45396), .B1(n45394), .ZN(n45398) );
  NOR2HSV4 U25936 ( .A1(n45270), .A2(n25141), .ZN(n45396) );
  NOR2HSV4 U25937 ( .A1(n25143), .A2(n25142), .ZN(n25141) );
  CLKNHSV2 U25938 ( .I(n45271), .ZN(n25142) );
  CLKNHSV2 U25939 ( .I(n45272), .ZN(n25143) );
  INHSV6 U25940 ( .I(n26070), .ZN(n43887) );
  CLKNAND2HSV4 U25941 ( .A1(n39739), .A2(n40017), .ZN(n29744) );
  INHSV2 U25942 ( .I(n29744), .ZN(n25458) );
  NAND2HSV4 U25943 ( .A1(n47932), .A2(n44350), .ZN(n44351) );
  INHSV2 U25944 ( .I(n44351), .ZN(n44368) );
  NAND2HSV2 U25945 ( .A1(n34319), .A2(n25144), .ZN(n34350) );
  CLKNHSV2 U25946 ( .I(n25145), .ZN(n25144) );
  CLKNAND2HSV2 U25947 ( .A1(n34320), .A2(n34318), .ZN(n25145) );
  NAND2HSV2 U25948 ( .A1(n46122), .A2(n25146), .ZN(n38609) );
  NOR2HSV2 U25949 ( .A1(n25350), .A2(n46120), .ZN(n25146) );
  CLKNAND2HSV2 U25950 ( .A1(n25172), .A2(n37264), .ZN(n25152) );
  NAND2HSV2 U25951 ( .A1(n29753), .A2(n49741), .ZN(n49160) );
  XOR3HSV4 U25952 ( .A1(n49162), .A2(n49161), .A3(n49160), .Z(n49163) );
  CLKNAND2HSV3 U25953 ( .A1(n43020), .A2(n43019), .ZN(n43236) );
  CLKNAND2HSV4 U25954 ( .A1(n26001), .A2(n29698), .ZN(n43884) );
  INHSV8 U25955 ( .I(n56059), .ZN(n56490) );
  CLKNAND2HSV3 U25956 ( .A1(n25770), .A2(n43465), .ZN(n43471) );
  CLKNAND2HSV3 U25957 ( .A1(n45584), .A2(n43753), .ZN(n25165) );
  INHSV6 U25958 ( .I(n50757), .ZN(n48484) );
  AOI21HSV2 U25959 ( .A1(n45596), .A2(n36967), .B(n43744), .ZN(n43745) );
  OAI21HSV1 U25960 ( .A1(n29443), .A2(n29444), .B(n29445), .ZN(\pe3/poht [12])
         );
  NAND2HSV4 U25961 ( .A1(n25709), .A2(n51958), .ZN(n51959) );
  NOR2HSV4 U25962 ( .A1(n46561), .A2(n46115), .ZN(n26072) );
  CLKNAND2HSV2 U25963 ( .A1(n25148), .A2(n25147), .ZN(n29899) );
  CLKNAND2HSV2 U25964 ( .A1(n29895), .A2(n29896), .ZN(n25147) );
  CLKNHSV2 U25965 ( .I(n29897), .ZN(n25148) );
  NAND2HSV2 U25966 ( .A1(n25709), .A2(n52418), .ZN(n26714) );
  CLKNHSV2 U25967 ( .I(n30975), .ZN(n30761) );
  XNOR2HSV4 U25968 ( .A1(n26043), .A2(n30995), .ZN(n30975) );
  OAI21HSV2 U25969 ( .A1(n25149), .A2(n30508), .B(n30510), .ZN(n30511) );
  CLKNAND2HSV2 U25970 ( .A1(n30649), .A2(n29699), .ZN(n25149) );
  NOR3HSV2 U25971 ( .A1(n30433), .A2(n30435), .A3(n29950), .ZN(n30410) );
  NOR2HSV2 U25972 ( .A1(n30399), .A2(n30400), .ZN(n30433) );
  INHSV4 U25973 ( .I(n44952), .ZN(n25595) );
  NAND2HSV4 U25974 ( .A1(n25595), .A2(n25596), .ZN(n25594) );
  CLKNHSV6 U25975 ( .I(n53095), .ZN(n52840) );
  NAND2HSV4 U25976 ( .A1(n41136), .A2(n41137), .ZN(n41220) );
  NAND2HSV2 U25977 ( .A1(n36035), .A2(n36033), .ZN(n36031) );
  XOR2HSV2 U25978 ( .A1(n25150), .A2(n48163), .Z(\pe2/poht [10]) );
  XNOR2HSV4 U25979 ( .A1(n25710), .A2(n25711), .ZN(n25150) );
  INHSV4 U25980 ( .I(n42817), .ZN(n55701) );
  INHSV2 U25981 ( .I(n25152), .ZN(n25151) );
  CLKNAND2HSV4 U25982 ( .A1(n41321), .A2(n41320), .ZN(n41327) );
  CLKNAND2HSV8 U25983 ( .A1(n41327), .A2(n41326), .ZN(n41699) );
  BUFHSV6 U25984 ( .I(n26734), .Z(n48049) );
  BUFHSV6 U25985 ( .I(n26734), .Z(n48029) );
  INHSV2 U25986 ( .I(n37928), .ZN(n25153) );
  CLKNAND2HSV2 U25987 ( .A1(n25153), .A2(n26836), .ZN(n26898) );
  INHSV2 U25988 ( .I(n45408), .ZN(n25154) );
  IOA21HSV4 U25989 ( .A1(n25154), .A2(n45145), .B(n45407), .ZN(n26137) );
  NAND2HSV4 U25990 ( .A1(n43614), .A2(n37272), .ZN(n26341) );
  NAND2HSV4 U25991 ( .A1(n39120), .A2(n30779), .ZN(n30853) );
  INHSV4 U25992 ( .I(n45147), .ZN(n25832) );
  CLKNHSV6 U25993 ( .I(n25832), .ZN(n25833) );
  CLKNAND2HSV3 U25994 ( .A1(n43879), .A2(n43878), .ZN(n45599) );
  INHSV4 U25995 ( .I(n43884), .ZN(n43885) );
  NAND3HSV4 U25996 ( .A1(n44708), .A2(n44707), .A3(n44706), .ZN(n45389) );
  INOR2HSV1 U25997 ( .A1(\pe6/ti_7t [17]), .B1(n35797), .ZN(n32533) );
  CLKNAND2HSV3 U25998 ( .A1(n30586), .A2(n30585), .ZN(n30753) );
  NAND2HSV8 U25999 ( .A1(n35806), .A2(\pe6/ti_7t [19]), .ZN(n32551) );
  CLKNAND2HSV2 U26000 ( .A1(n43730), .A2(n43729), .ZN(n43725) );
  NAND2HSV4 U26001 ( .A1(n47988), .A2(n26162), .ZN(n26158) );
  INHSV2 U26002 ( .I(n53227), .ZN(n56175) );
  INHSV6 U26003 ( .I(n45931), .ZN(n44669) );
  CLKNAND2HSV3 U26004 ( .A1(n44670), .A2(n44669), .ZN(n44671) );
  CLKNHSV6 U26005 ( .I(n55705), .ZN(n53227) );
  CLKNAND2HSV2 U26006 ( .A1(n29765), .A2(n58372), .ZN(n59340) );
  NAND2HSV4 U26007 ( .A1(n25695), .A2(n25694), .ZN(n43352) );
  NAND2HSV2 U26008 ( .A1(n38730), .A2(n38731), .ZN(n38746) );
  NAND3HSV3 U26009 ( .A1(n29671), .A2(n30436), .A3(n52799), .ZN(n30408) );
  NOR2HSV8 U26010 ( .A1(n43885), .A2(n43469), .ZN(n43888) );
  XNOR2HSV4 U26011 ( .A1(n44285), .A2(n44284), .ZN(n44286) );
  INHSV4 U26012 ( .I(n26258), .ZN(n26259) );
  INHSV8 U26013 ( .I(n42051), .ZN(n42069) );
  INHSV3 U26014 ( .I(n43365), .ZN(n43366) );
  NAND2HSV8 U26015 ( .A1(n43610), .A2(n29747), .ZN(n25960) );
  CLKNAND2HSV4 U26016 ( .A1(n41908), .A2(n42200), .ZN(n41822) );
  CLKNAND2HSV4 U26017 ( .A1(n30200), .A2(n30199), .ZN(n30397) );
  CLKAND2HSV4 U26018 ( .A1(n30403), .A2(n39403), .Z(n29671) );
  INHSV2 U26019 ( .I(n26721), .ZN(n26720) );
  INHSV2 U26020 ( .I(n25155), .ZN(n38364) );
  CLKNAND2HSV2 U26021 ( .A1(n38363), .A2(n38108), .ZN(n25155) );
  CLKNAND2HSV4 U26022 ( .A1(n41908), .A2(n42084), .ZN(n41909) );
  CLKXOR2HSV4 U26023 ( .A1(n41910), .A2(n41909), .Z(n25827) );
  CLKNHSV3 U26024 ( .I(n45509), .ZN(n43750) );
  CLKNHSV8 U26025 ( .I(n45618), .ZN(n44664) );
  INHSV2 U26026 ( .I(n42321), .ZN(n25156) );
  NAND3HSV4 U26027 ( .A1(n25156), .A2(n44650), .A3(n44523), .ZN(n42489) );
  INHSV2 U26028 ( .I(n43127), .ZN(n43135) );
  XNOR2HSV4 U26029 ( .A1(n25158), .A2(n25157), .ZN(\pe1/poht [12]) );
  CLKNAND2HSV2 U26030 ( .A1(n55423), .A2(\pe1/got [20]), .ZN(n25157) );
  XNOR2HSV4 U26031 ( .A1(n54633), .A2(n54634), .ZN(n25158) );
  CLKNAND2HSV4 U26032 ( .A1(n36572), .A2(n36571), .ZN(n36655) );
  INHSV4 U26033 ( .I(n39698), .ZN(n39721) );
  INHSV6 U26034 ( .I(n25961), .ZN(n43899) );
  NAND2HSV4 U26035 ( .A1(n43356), .A2(n26134), .ZN(n43353) );
  CLKNAND2HSV4 U26036 ( .A1(n43348), .A2(n43347), .ZN(n43357) );
  NAND2HSV4 U26037 ( .A1(n43255), .A2(n43254), .ZN(n25959) );
  NAND2HSV2 U26038 ( .A1(n36651), .A2(n36650), .ZN(n36653) );
  INHSV4 U26039 ( .I(n43123), .ZN(n43124) );
  CLKNAND2HSV4 U26040 ( .A1(n43134), .A2(n25256), .ZN(n43125) );
  CLKNAND2HSV8 U26041 ( .A1(n43125), .A2(n43124), .ZN(n43143) );
  AOI22HSV4 U26042 ( .A1(n35316), .A2(n35472), .B1(n35471), .B2(n35470), .ZN(
        n35473) );
  CLKNAND2HSV4 U26043 ( .A1(n36471), .A2(n36470), .ZN(n36557) );
  XNOR2HSV4 U26044 ( .A1(n33525), .A2(n25159), .ZN(n33607) );
  CLKNAND2HSV2 U26045 ( .A1(n45801), .A2(n33805), .ZN(n25159) );
  NAND2HSV4 U26046 ( .A1(n34867), .A2(n33707), .ZN(n33756) );
  INHSV2 U26047 ( .I(n41232), .ZN(n29057) );
  AOI21HSV2 U26048 ( .A1(n35008), .A2(n35007), .B(n35482), .ZN(n35009) );
  CLKNAND2HSV2 U26049 ( .A1(n25160), .A2(n38622), .ZN(n38875) );
  CLKNAND2HSV2 U26050 ( .A1(n38624), .A2(n38635), .ZN(n25160) );
  INHSV4 U26051 ( .I(n52778), .ZN(n38377) );
  CLKNAND2HSV2 U26052 ( .A1(n38602), .A2(n38601), .ZN(n38610) );
  NAND2HSV2 U26053 ( .A1(n26098), .A2(n38778), .ZN(n38722) );
  BUFHSV6 U26054 ( .I(n49253), .Z(n56622) );
  BUFHSV8 U26055 ( .I(n49253), .Z(n56561) );
  AND2HSV4 U26056 ( .A1(n48620), .A2(n36972), .Z(n37103) );
  CLKNAND2HSV0 U26057 ( .A1(n52163), .A2(n38782), .ZN(n47568) );
  INOR2HSV2 U26058 ( .A1(n41322), .B1(n41324), .ZN(n41320) );
  OAI21HSV4 U26059 ( .A1(n59573), .A2(n39688), .B(n39242), .ZN(n39574) );
  OAI21HSV2 U26060 ( .A1(n41134), .A2(\pe1/ti_7t [17]), .B(n52831), .ZN(n41218) );
  INHSV4 U26061 ( .I(n36652), .ZN(n37837) );
  NOR2HSV4 U26062 ( .A1(n45787), .A2(n32457), .ZN(n44379) );
  CLKNAND2HSV4 U26063 ( .A1(n30338), .A2(n30337), .ZN(n30661) );
  OAI22HSV4 U26064 ( .A1(n34445), .A2(n34560), .B1(n34444), .B2(n33928), .ZN(
        n34556) );
  CLKNHSV6 U26065 ( .I(n50211), .ZN(n58141) );
  NAND2HSV2 U26066 ( .A1(n37550), .A2(n37549), .ZN(n37754) );
  CLKNAND2HSV2 U26067 ( .A1(n52816), .A2(n31242), .ZN(n37549) );
  CLKNAND2HSV4 U26068 ( .A1(n30974), .A2(n30973), .ZN(n31099) );
  CLKAND2HSV4 U26069 ( .A1(n35312), .A2(n35311), .Z(n35314) );
  NAND3HSV4 U26070 ( .A1(n45792), .A2(n25605), .A3(n35314), .ZN(n35461) );
  NAND2HSV4 U26071 ( .A1(n36037), .A2(n36036), .ZN(n36044) );
  NAND2HSV4 U26072 ( .A1(n43357), .A2(n43358), .ZN(n43354) );
  NOR2HSV8 U26073 ( .A1(n43354), .A2(n43353), .ZN(n43479) );
  NAND2HSV4 U26074 ( .A1(n45603), .A2(n45602), .ZN(n45609) );
  NOR2HSV3 U26075 ( .A1(n41140), .A2(n44522), .ZN(n41236) );
  NOR2HSV2 U26076 ( .A1(n46103), .A2(n46071), .ZN(n45927) );
  NOR2HSV4 U26077 ( .A1(n45613), .A2(n45614), .ZN(n46103) );
  CLKNAND2HSV2 U26078 ( .A1(n38882), .A2(n38881), .ZN(n25180) );
  AOI21HSV4 U26079 ( .A1(n38880), .A2(n44309), .B(n38879), .ZN(n38882) );
  INHSV2 U26080 ( .I(n45400), .ZN(n52918) );
  INHSV2 U26081 ( .I(n25161), .ZN(n39426) );
  CLKNAND2HSV2 U26082 ( .A1(n39397), .A2(n39391), .ZN(n25161) );
  INHSV2 U26083 ( .I(n26530), .ZN(n26523) );
  CLKNAND2HSV2 U26084 ( .A1(n53093), .A2(n53092), .ZN(n53096) );
  CLKNAND2HSV4 U26085 ( .A1(n33704), .A2(n33703), .ZN(n33706) );
  NAND2HSV2 U26086 ( .A1(n38387), .A2(\pe2/got [29]), .ZN(n26767) );
  INHSV2 U26087 ( .I(n47784), .ZN(n47780) );
  NAND2HSV4 U26088 ( .A1(n26742), .A2(n47780), .ZN(n26585) );
  INHSV4 U26089 ( .I(n43246), .ZN(n43140) );
  CLKNAND2HSV3 U26090 ( .A1(n43493), .A2(n42694), .ZN(n25760) );
  INAND2HSV4 U26091 ( .A1(n30093), .B1(n30190), .ZN(n52733) );
  AOI21HSV2 U26092 ( .A1(n52733), .A2(n30095), .B(n30094), .ZN(n30096) );
  INHSV2 U26093 ( .I(n43870), .ZN(n59998) );
  CLKNHSV1 U26094 ( .I(n46558), .ZN(n46114) );
  NAND3HSV4 U26095 ( .A1(n26038), .A2(n48313), .A3(n42490), .ZN(n48456) );
  NAND2HSV2 U26096 ( .A1(n48456), .A2(n53512), .ZN(n48457) );
  CLKNAND2HSV4 U26097 ( .A1(n60074), .A2(n30320), .ZN(n30070) );
  CLKNAND2HSV8 U26098 ( .A1(n30070), .A2(n30203), .ZN(n30099) );
  NOR2HSV4 U26099 ( .A1(n43738), .A2(n43485), .ZN(n43486) );
  NAND2HSV4 U26100 ( .A1(n33593), .A2(n33192), .ZN(n33697) );
  CLKNAND2HSV3 U26101 ( .A1(n25237), .A2(n25236), .ZN(n45765) );
  INHSV8 U26102 ( .I(n44678), .ZN(n46310) );
  CLKNAND2HSV3 U26103 ( .A1(n45766), .A2(n45765), .ZN(n45777) );
  NAND2HSV4 U26104 ( .A1(n45626), .A2(n43021), .ZN(n45627) );
  NAND2HSV4 U26105 ( .A1(n43886), .A2(n45596), .ZN(n44328) );
  NAND3HSV3 U26106 ( .A1(n46106), .A2(n46105), .A3(n46104), .ZN(n46110) );
  NOR2HSV4 U26107 ( .A1(n42797), .A2(n26565), .ZN(n25899) );
  NAND2HSV2 U26108 ( .A1(n25899), .A2(n25898), .ZN(n25897) );
  CLKNAND2HSV2 U26109 ( .A1(n45927), .A2(n46104), .ZN(n25211) );
  INHSV4 U26110 ( .I(n25211), .ZN(n45929) );
  CLKNAND2HSV4 U26111 ( .A1(n26264), .A2(n26263), .ZN(n39005) );
  INHSV2 U26112 ( .I(n50717), .ZN(n55946) );
  CLKNAND2HSV4 U26113 ( .A1(n42033), .A2(n41328), .ZN(n26613) );
  NAND2HSV4 U26114 ( .A1(n25164), .A2(n25162), .ZN(n41915) );
  INHSV2 U26115 ( .I(n25163), .ZN(n25162) );
  NAND2HSV2 U26116 ( .A1(n42033), .A2(n41727), .ZN(n25163) );
  NAND2HSV4 U26117 ( .A1(n41729), .A2(n41728), .ZN(n25164) );
  CLKNAND2HSV3 U26118 ( .A1(n43738), .A2(n26169), .ZN(n43879) );
  INHSV4 U26119 ( .I(n38272), .ZN(n44315) );
  BUFHSV8 U26120 ( .I(n41823), .Z(n41828) );
  CLKXOR2HSV4 U26121 ( .A1(n25224), .A2(n26136), .Z(n25442) );
  CLKNAND2HSV4 U26122 ( .A1(n25165), .A2(n43863), .ZN(n26034) );
  XNOR2HSV2 U26123 ( .A1(n51685), .A2(n51684), .ZN(\pe2/poht [12]) );
  NAND2HSV4 U26124 ( .A1(n45508), .A2(n44667), .ZN(n44681) );
  INHSV12 U26125 ( .I(\pe1/got [32]), .ZN(n40329) );
  BUFHSV12 U26126 ( .I(n40329), .Z(n47935) );
  CLKNAND2HSV2 U26127 ( .A1(n38012), .A2(n38109), .ZN(n25851) );
  NOR2HSV4 U26128 ( .A1(n38328), .A2(n45129), .ZN(n38012) );
  NOR2HSV4 U26129 ( .A1(n40361), .A2(n40329), .ZN(n40375) );
  INHSV4 U26130 ( .I(n43601), .ZN(n43610) );
  INHSV6 U26131 ( .I(n40599), .ZN(n40601) );
  NAND2HSV4 U26132 ( .A1(n40601), .A2(n26885), .ZN(n40602) );
  NAND2HSV2 U26133 ( .A1(n38176), .A2(n38179), .ZN(n26721) );
  NOR2HSV4 U26134 ( .A1(n38747), .A2(n52810), .ZN(n38620) );
  NOR2HSV4 U26135 ( .A1(n26148), .A2(n26144), .ZN(n29993) );
  CLKNAND2HSV4 U26136 ( .A1(n30060), .A2(n29984), .ZN(n30143) );
  INHSV4 U26137 ( .I(n30143), .ZN(n29985) );
  MUX2NHSV2 U26138 ( .I0(n45769), .I1(n45767), .S(n45770), .ZN(n45766) );
  XOR2HSV0 U26139 ( .A1(n25167), .A2(n25166), .Z(\pe5/poht [25]) );
  NAND2HSV0 U26140 ( .A1(n53210), .A2(n59905), .ZN(n25166) );
  CLKXOR2HSV2 U26141 ( .A1(n51271), .A2(n51270), .Z(n25167) );
  NAND2HSV4 U26142 ( .A1(n25709), .A2(n51889), .ZN(n51682) );
  CLKNAND2HSV4 U26143 ( .A1(n25197), .A2(n44683), .ZN(n45762) );
  CLKNAND2HSV4 U26144 ( .A1(n45762), .A2(n45763), .ZN(n46092) );
  INHSV2 U26145 ( .I(n41589), .ZN(n41591) );
  INHSV2 U26146 ( .I(n33404), .ZN(n25168) );
  NOR2HSV4 U26147 ( .A1(n25168), .A2(n33405), .ZN(n33400) );
  INHSV4 U26148 ( .I(n26823), .ZN(n26408) );
  NAND2HSV4 U26149 ( .A1(n26839), .A2(n40407), .ZN(n41408) );
  NAND2HSV4 U26150 ( .A1(n41408), .A2(n41407), .ZN(n41593) );
  XNOR2HSV4 U26151 ( .A1(n36021), .A2(n36020), .ZN(n36022) );
  NAND2HSV2 U26152 ( .A1(n46097), .A2(n46096), .ZN(n46098) );
  CLKNAND2HSV2 U26153 ( .A1(n46099), .A2(n46071), .ZN(n45611) );
  OAI21HSV4 U26154 ( .A1(n29922), .A2(n29921), .B(n29920), .ZN(n29924) );
  CLKNHSV0 U26155 ( .I(n42918), .ZN(n59821) );
  CLKNHSV0 U26156 ( .I(n47430), .ZN(n55824) );
  NAND2HSV4 U26157 ( .A1(n36053), .A2(n36083), .ZN(n35912) );
  CLKNHSV6 U26158 ( .I(n40969), .ZN(n40439) );
  CLKNAND2HSV2 U26159 ( .A1(n60031), .A2(n33450), .ZN(n33671) );
  CLKNAND2HSV2 U26160 ( .A1(n33671), .A2(n33670), .ZN(n33673) );
  INHSV4 U26161 ( .I(n52812), .ZN(n38759) );
  NAND2HSV4 U26162 ( .A1(n29946), .A2(n39558), .ZN(n29821) );
  INHSV4 U26163 ( .I(n29821), .ZN(n29822) );
  INHSV4 U26164 ( .I(n43911), .ZN(n43913) );
  CLKNAND2HSV2 U26165 ( .A1(n36071), .A2(n46163), .ZN(n36070) );
  NAND3HSV3 U26166 ( .A1(n35915), .A2(n35802), .A3(n52710), .ZN(n35803) );
  NAND2HSV4 U26167 ( .A1(n26839), .A2(n53514), .ZN(n41586) );
  NOR2HSV8 U26168 ( .A1(n56910), .A2(n43613), .ZN(n45752) );
  CLKNHSV2 U26169 ( .I(n46545), .ZN(n51118) );
  CLKNAND2HSV2 U26170 ( .A1(n43914), .A2(n25169), .ZN(n46545) );
  CLKNAND2HSV2 U26171 ( .A1(n25171), .A2(n25170), .ZN(n25169) );
  CLKNHSV2 U26172 ( .I(n46089), .ZN(n25170) );
  CLKNHSV2 U26173 ( .I(n43915), .ZN(n25171) );
  NAND2HSV4 U26174 ( .A1(n26337), .A2(n26334), .ZN(n26335) );
  CLKNAND2HSV1 U26175 ( .A1(n40432), .A2(n40433), .ZN(n25199) );
  CLKNHSV3 U26176 ( .I(n31519), .ZN(n31513) );
  INAND2HSV4 U26177 ( .A1(n45399), .B1(\pe2/ti_7t [30]), .ZN(n45138) );
  OR2HSV4 U26178 ( .A1(n42335), .A2(n40378), .Z(n40379) );
  CLKNAND2HSV0 U26179 ( .A1(n30884), .A2(n48885), .ZN(n30763) );
  NAND3HSV3 U26180 ( .A1(n34340), .A2(n34333), .A3(n34698), .ZN(n34335) );
  NAND2HSV4 U26181 ( .A1(n47902), .A2(n47901), .ZN(n51151) );
  INHSV2 U26182 ( .I(n43135), .ZN(n43134) );
  CLKNHSV0 U26183 ( .I(n43127), .ZN(n25172) );
  INHSV4 U26184 ( .I(n34994), .ZN(n34999) );
  CLKXOR2HSV4 U26185 ( .A1(n31657), .A2(n31656), .Z(n31660) );
  INHSV6 U26186 ( .I(n32714), .ZN(n32991) );
  CLKNHSV0 U26187 ( .I(n32714), .ZN(n35925) );
  NAND2HSV2 U26188 ( .A1(n36405), .A2(n36404), .ZN(n36407) );
  OAI21HSV2 U26189 ( .A1(n27150), .A2(n27151), .B(n27152), .ZN(\pe6/poht [4])
         );
  BUFHSV8 U26190 ( .I(n34218), .Z(n34865) );
  CLKNAND2HSV4 U26191 ( .A1(n34093), .A2(n34865), .ZN(n34094) );
  NOR2HSV8 U26192 ( .A1(n41913), .A2(n41722), .ZN(n41840) );
  CLKXOR2HSV2 U26193 ( .A1(n29190), .A2(n29203), .Z(n29204) );
  CLKNAND2HSV2 U26194 ( .A1(n59023), .A2(n49665), .ZN(n58931) );
  NOR2HSV4 U26195 ( .A1(n36407), .A2(n36406), .ZN(n36411) );
  NAND2HSV4 U26196 ( .A1(n48454), .A2(n48455), .ZN(n48453) );
  NAND3HSV4 U26197 ( .A1(n29889), .A2(n25562), .A3(n25173), .ZN(n29990) );
  CLKNAND2HSV2 U26198 ( .A1(n25175), .A2(n25174), .ZN(n25173) );
  CLKNHSV2 U26199 ( .I(n29888), .ZN(n25174) );
  CLKNHSV2 U26200 ( .I(n29887), .ZN(n25175) );
  XNOR2HSV4 U26201 ( .A1(n25845), .A2(n42467), .ZN(n42468) );
  NOR2HSV4 U26202 ( .A1(n25507), .A2(n32045), .ZN(n25459) );
  NOR2HSV4 U26203 ( .A1(n29757), .A2(n32158), .ZN(n25507) );
  NAND2HSV2 U26204 ( .A1(n30340), .A2(n30046), .ZN(n30047) );
  INHSV4 U26205 ( .I(n54159), .ZN(n55543) );
  NAND2HSV2 U26206 ( .A1(n55543), .A2(\pe1/got [20]), .ZN(n54446) );
  XNOR2HSV4 U26207 ( .A1(n30393), .A2(n30392), .ZN(n30394) );
  INHSV2 U26208 ( .I(n46101), .ZN(n25216) );
  NAND2HSV4 U26209 ( .A1(n46102), .A2(n25216), .ZN(n46111) );
  NAND3HSV4 U26210 ( .A1(n44691), .A2(n36087), .A3(n36088), .ZN(n44375) );
  NAND3HSV4 U26211 ( .A1(n36063), .A2(n36064), .A3(n36062), .ZN(n36087) );
  CLKNAND2HSV2 U26212 ( .A1(n35154), .A2(n35153), .ZN(n35155) );
  INHSV2 U26213 ( .I(n26279), .ZN(n35156) );
  NOR2HSV2 U26214 ( .A1(n35156), .A2(n35155), .ZN(n35159) );
  CLKNHSV6 U26215 ( .I(n40014), .ZN(n52836) );
  INOR2HSV4 U26216 ( .A1(n39872), .B1(n39874), .ZN(n40138) );
  INHSV2 U26217 ( .I(n37769), .ZN(n25478) );
  OR2HSV4 U26218 ( .A1(n35918), .A2(n59487), .Z(n29649) );
  XOR3HSV2 U26219 ( .A1(n25176), .A2(n55818), .A3(n55819), .Z(\pe3/poht [3])
         );
  XNOR2HSV4 U26220 ( .A1(n55817), .A2(n55816), .ZN(n25176) );
  INHSV2 U26221 ( .I(n25177), .ZN(n35296) );
  NAND3HSV2 U26222 ( .A1(n35161), .A2(n35160), .A3(n47772), .ZN(n25177) );
  XNOR2HSV4 U26223 ( .A1(n35140), .A2(n35139), .ZN(n35142) );
  XNOR2HSV4 U26224 ( .A1(n40887), .A2(n40888), .ZN(n40906) );
  XNOR2HSV4 U26225 ( .A1(n40848), .A2(n40847), .ZN(n40850) );
  INAND2HSV4 U26226 ( .A1(n43743), .B1(n55612), .ZN(n43896) );
  AOI21HSV4 U26227 ( .A1(n45596), .A2(n45932), .B(n43880), .ZN(n43881) );
  NAND3HSV3 U26228 ( .A1(n37423), .A2(n25178), .A3(n37429), .ZN(n37426) );
  INHSV2 U26229 ( .I(n37421), .ZN(n25178) );
  CLKNAND2HSV2 U26230 ( .A1(n42592), .A2(n42591), .ZN(n37431) );
  NAND2HSV4 U26231 ( .A1(n41061), .A2(n40958), .ZN(n40959) );
  INHSV4 U26232 ( .I(n40959), .ZN(n40961) );
  DELHS1 U26233 ( .I(n53526), .Z(n25179) );
  BUFHSV6 U26234 ( .I(n39698), .Z(n26285) );
  NAND2HSV4 U26235 ( .A1(n26285), .A2(n39695), .ZN(n39712) );
  CLKNAND2HSV4 U26236 ( .A1(n34592), .A2(n34017), .ZN(n34106) );
  CLKNAND2HSV3 U26237 ( .A1(n25686), .A2(n44669), .ZN(n44672) );
  INHSV8 U26238 ( .I(n31325), .ZN(n31497) );
  NOR2HSV3 U26239 ( .A1(n25652), .A2(n46076), .ZN(n25322) );
  INHSV6 U26240 ( .I(n50752), .ZN(n56058) );
  INHSV2 U26241 ( .I(n50752), .ZN(n56676) );
  NAND2HSV0 U26242 ( .A1(n56676), .A2(n56560), .ZN(n56932) );
  CLKNAND2HSV4 U26243 ( .A1(n25181), .A2(n25180), .ZN(n44034) );
  NAND2HSV4 U26244 ( .A1(n38883), .A2(n25263), .ZN(n25181) );
  NAND2HSV4 U26245 ( .A1(n52748), .A2(n25182), .ZN(n38112) );
  NOR2HSV8 U26246 ( .A1(n25184), .A2(n25183), .ZN(n25182) );
  INHSV4 U26247 ( .I(n38885), .ZN(n25183) );
  INHSV6 U26248 ( .I(n52747), .ZN(n25184) );
  INHSV4 U26249 ( .I(n45121), .ZN(n45118) );
  XNOR2HSV4 U26250 ( .A1(n52911), .A2(n25185), .ZN(n52913) );
  CLKNAND2HSV2 U26251 ( .A1(n52910), .A2(n52895), .ZN(n25185) );
  CLKNAND2HSV4 U26252 ( .A1(n30754), .A2(n30960), .ZN(n52787) );
  INHSV4 U26253 ( .I(n47853), .ZN(n57835) );
  BUFHSV16 U26254 ( .I(n49661), .Z(n25709) );
  NAND3HSV2 U26255 ( .A1(n25994), .A2(n37245), .A3(n43468), .ZN(n37247) );
  NOR2HSV4 U26256 ( .A1(n37247), .A2(n37246), .ZN(n37256) );
  XOR3HSV2 U26257 ( .A1(n47925), .A2(n47924), .A3(n47923), .Z(\pe4/poht [22])
         );
  XNOR2HSV4 U26258 ( .A1(n35794), .A2(n35795), .ZN(n35801) );
  AOI21HSV2 U26259 ( .A1(n25843), .A2(n47782), .B(n33457), .ZN(n47781) );
  CLKNHSV0 U26260 ( .I(n47781), .ZN(n25555) );
  IOA21HSV4 U26261 ( .A1(n59573), .A2(n39741), .B(n39742), .ZN(n39880) );
  NAND2HSV2 U26262 ( .A1(n48742), .A2(n39880), .ZN(n40275) );
  XNOR2HSV4 U26263 ( .A1(n40703), .A2(n25186), .ZN(n40705) );
  XNOR2HSV4 U26264 ( .A1(n40702), .A2(n40701), .ZN(n25186) );
  NOR2HSV4 U26265 ( .A1(n37223), .A2(n43613), .ZN(n37173) );
  XNOR2HSV4 U26266 ( .A1(n51096), .A2(n51095), .ZN(n51098) );
  XNOR2HSV2 U26267 ( .A1(n51098), .A2(n51097), .ZN(n51099) );
  CLKNAND2HSV1 U26268 ( .A1(n43133), .A2(n45755), .ZN(n25400) );
  NAND2HSV8 U26269 ( .A1(n37432), .A2(n37431), .ZN(n42600) );
  OR2HSV8 U26270 ( .A1(n32968), .A2(n46549), .Z(n32962) );
  CLKNAND2HSV2 U26271 ( .A1(n48309), .A2(n39879), .ZN(n47385) );
  CLKNAND2HSV4 U26272 ( .A1(n37415), .A2(n37269), .ZN(n37270) );
  INHSV1 U26273 ( .I(n40969), .ZN(n41225) );
  AOI21HSV2 U26274 ( .A1(n37088), .A2(n36978), .B(n36985), .ZN(n37034) );
  CLKNAND2HSV2 U26275 ( .A1(n58476), .A2(n32354), .ZN(n50907) );
  CLKNHSV6 U26276 ( .I(n32433), .ZN(n32646) );
  CLKNAND2HSV2 U26277 ( .A1(n59600), .A2(n33498), .ZN(n33653) );
  XNOR2HSV2 U26278 ( .A1(n33654), .A2(n33653), .ZN(n33657) );
  XNOR2HSV4 U26279 ( .A1(n35700), .A2(n35699), .ZN(n35702) );
  INHSV2 U26280 ( .I(n37267), .ZN(n37164) );
  INHSV4 U26281 ( .I(n37164), .ZN(n37167) );
  INHSV2 U26282 ( .I(n37446), .ZN(n37450) );
  INHSV2 U26283 ( .I(n35464), .ZN(n25421) );
  CLKNHSV2 U26284 ( .I(n26546), .ZN(n26511) );
  CLKNAND2HSV2 U26285 ( .A1(n45098), .A2(n45097), .ZN(n26546) );
  NAND2HSV2 U26286 ( .A1(n42616), .A2(n25818), .ZN(n25817) );
  INHSV4 U26287 ( .I(n26416), .ZN(n26690) );
  OAI21HSV2 U26288 ( .A1(n44828), .A2(n44824), .B(n44309), .ZN(n44825) );
  CLKNHSV0 U26289 ( .I(n44825), .ZN(n45274) );
  CLKNAND2HSV4 U26290 ( .A1(n26061), .A2(n37260), .ZN(n37346) );
  NAND2HSV4 U26291 ( .A1(n42499), .A2(n42498), .ZN(n26482) );
  CLKNAND2HSV4 U26292 ( .A1(n44687), .A2(n44686), .ZN(n44685) );
  CLKNAND2HSV4 U26293 ( .A1(n25715), .A2(n26602), .ZN(n46299) );
  NOR2HSV4 U26294 ( .A1(n35704), .A2(n32239), .ZN(n44344) );
  INAND2HSV4 U26295 ( .A1(n32686), .B1(n32685), .ZN(n32687) );
  OAI21HSV4 U26296 ( .A1(n33085), .A2(n35704), .B(n35703), .ZN(n25860) );
  CLKNAND2HSV2 U26297 ( .A1(n59340), .A2(n58384), .ZN(n58373) );
  NOR2HSV2 U26298 ( .A1(n38455), .A2(n25187), .ZN(n38374) );
  INHSV4 U26299 ( .I(n38359), .ZN(n25187) );
  NAND2HSV4 U26300 ( .A1(n38358), .A2(n38362), .ZN(n38359) );
  BUFHSV6 U26301 ( .I(n42596), .Z(n42492) );
  XNOR2HSV4 U26302 ( .A1(n50702), .A2(n50701), .ZN(n50704) );
  XNOR2HSV2 U26303 ( .A1(n50704), .A2(n50703), .ZN(n50705) );
  INHSV6 U26304 ( .I(n36873), .ZN(n36689) );
  CLKXOR2HSV4 U26305 ( .A1(n36750), .A2(n36749), .Z(n26610) );
  NAND3HSV4 U26306 ( .A1(n45775), .A2(n45774), .A3(n45773), .ZN(n45776) );
  OAI21HSV4 U26307 ( .A1(n43360), .A2(\pe3/ti_7t [27]), .B(n59962), .ZN(n44679) );
  NOR2HSV8 U26308 ( .A1(n42592), .A2(n36689), .ZN(n42693) );
  NAND2HSV0 U26309 ( .A1(n58655), .A2(n58711), .ZN(n27624) );
  NAND2HSV0 U26310 ( .A1(n58655), .A2(n58713), .ZN(n27990) );
  INHSV8 U26311 ( .I(n39398), .ZN(n40162) );
  CLKNAND2HSV4 U26312 ( .A1(n40011), .A2(n25830), .ZN(n40159) );
  NAND2HSV4 U26313 ( .A1(n26688), .A2(n42696), .ZN(n26687) );
  INHSV4 U26314 ( .I(\pe5/got [31]), .ZN(n29848) );
  NAND2HSV2 U26315 ( .A1(n40786), .A2(n26554), .ZN(n26553) );
  CLKNAND2HSV4 U26316 ( .A1(n32954), .A2(n32953), .ZN(n32955) );
  NOR2HSV4 U26317 ( .A1(n33994), .A2(n33993), .ZN(n34008) );
  CLKNHSV0 U26318 ( .I(n30441), .ZN(n37659) );
  NAND2HSV4 U26319 ( .A1(n46825), .A2(n32967), .ZN(n32810) );
  XNOR2HSV4 U26320 ( .A1(n43711), .A2(n43710), .ZN(n43713) );
  BUFHSV2 U26321 ( .I(n52789), .Z(n26565) );
  NAND2HSV4 U26322 ( .A1(n25188), .A2(n33986), .ZN(n33788) );
  CLKNHSV2 U26323 ( .I(n48892), .ZN(n25188) );
  INHSV4 U26324 ( .I(n49400), .ZN(n53172) );
  NAND2HSV2 U26325 ( .A1(n53172), .A2(n59166), .ZN(n44515) );
  NAND2HSV4 U26326 ( .A1(n42607), .A2(n26562), .ZN(n26561) );
  INHSV4 U26327 ( .I(n45622), .ZN(n42924) );
  OR2HSV4 U26328 ( .A1(n41225), .A2(n40395), .Z(n40467) );
  NOR2HSV8 U26329 ( .A1(n45268), .A2(n45267), .ZN(n45269) );
  INHSV4 U26330 ( .I(n38613), .ZN(n26889) );
  NAND2HSV4 U26331 ( .A1(n26889), .A2(n26890), .ZN(n26892) );
  INHSV2 U26332 ( .I(n36635), .ZN(n36650) );
  NAND2HSV4 U26333 ( .A1(n47951), .A2(n44344), .ZN(n33071) );
  NAND2HSV2 U26334 ( .A1(n25483), .A2(n32959), .ZN(n47951) );
  CLKNAND2HSV2 U26335 ( .A1(n42192), .A2(n42193), .ZN(n42194) );
  NAND2HSV2 U26336 ( .A1(n25862), .A2(n37554), .ZN(n30405) );
  NAND2HSV2 U26337 ( .A1(n56909), .A2(n56779), .ZN(n50747) );
  CLKNAND2HSV4 U26338 ( .A1(n25685), .A2(n25684), .ZN(n25683) );
  XOR2HSV4 U26339 ( .A1(n44306), .A2(n44305), .Z(n44323) );
  CLKXOR2HSV2 U26340 ( .A1(n26652), .A2(n25469), .Z(\pe2/poht [3]) );
  XNOR2HSV4 U26341 ( .A1(n41237), .A2(n25189), .ZN(n41214) );
  XNOR2HSV4 U26342 ( .A1(n41233), .A2(n41213), .ZN(n25189) );
  NAND3HSV2 U26343 ( .A1(n37104), .A2(n36978), .A3(n37103), .ZN(n36977) );
  NOR2HSV4 U26344 ( .A1(n36984), .A2(n43752), .ZN(n36978) );
  CLKNAND2HSV4 U26345 ( .A1(n39393), .A2(n39392), .ZN(n39395) );
  NAND2HSV2 U26346 ( .A1(n25335), .A2(n27779), .ZN(n27780) );
  OAI21HSV2 U26347 ( .A1(n27780), .A2(n27781), .B(n27782), .ZN(\pe2/poht [19])
         );
  NAND2HSV2 U26348 ( .A1(n25338), .A2(n28795), .ZN(n28796) );
  OAI21HSV2 U26349 ( .A1(n28796), .A2(n28797), .B(n28798), .ZN(\pe2/poht [25])
         );
  NOR2HSV4 U26350 ( .A1(n25191), .A2(n25190), .ZN(n29674) );
  CLKNHSV2 U26351 ( .I(n46603), .ZN(n25190) );
  CLKNHSV2 U26352 ( .I(n33594), .ZN(n25191) );
  XOR2HSV2 U26353 ( .A1(n58349), .A2(n25192), .Z(\pe6/poht [28]) );
  XOR2HSV2 U26354 ( .A1(n58350), .A2(n58351), .Z(n25192) );
  NAND2HSV4 U26355 ( .A1(n42599), .A2(n42600), .ZN(n42701) );
  NOR2HSV4 U26356 ( .A1(n37419), .A2(n37418), .ZN(n42599) );
  CLKNAND2HSV2 U26357 ( .A1(n36451), .A2(n36450), .ZN(n36455) );
  CLKNAND2HSV2 U26358 ( .A1(n25194), .A2(n25193), .ZN(n36302) );
  CLKNAND2HSV2 U26359 ( .A1(n36341), .A2(n36317), .ZN(n25193) );
  AOI21HSV4 U26360 ( .A1(n36315), .A2(n36320), .B(n38272), .ZN(n25194) );
  INHSV2 U26361 ( .I(n55917), .ZN(n45582) );
  INAND2HSV4 U26362 ( .A1(n55917), .B1(n36788), .ZN(n43345) );
  INHSV4 U26363 ( .I(n52763), .ZN(n41114) );
  NAND2HSV4 U26364 ( .A1(n41035), .A2(n41114), .ZN(n41037) );
  CLKNAND2HSV2 U26365 ( .A1(n25527), .A2(n30192), .ZN(n30078) );
  NAND2HSV4 U26366 ( .A1(n25597), .A2(n33089), .ZN(n36207) );
  INHSV3 U26367 ( .I(n26225), .ZN(n26396) );
  CLKNHSV8 U26368 ( .I(n43482), .ZN(n43370) );
  INHSV4 U26369 ( .I(n41124), .ZN(n41127) );
  NAND2HSV2 U26370 ( .A1(n44647), .A2(n44648), .ZN(n25571) );
  NAND2HSV4 U26371 ( .A1(n55490), .A2(n53786), .ZN(n25572) );
  CLKNAND2HSV2 U26372 ( .A1(n25572), .A2(n25571), .ZN(n25573) );
  INHSV4 U26373 ( .I(n25195), .ZN(n43741) );
  CLKNAND2HSV4 U26374 ( .A1(n43739), .A2(n29721), .ZN(n25195) );
  NAND2HSV4 U26375 ( .A1(n43476), .A2(n43612), .ZN(n43739) );
  NAND2HSV4 U26376 ( .A1(n42358), .A2(\pe1/got [26]), .ZN(n41903) );
  XNOR2HSV2 U26377 ( .A1(n41903), .A2(n41902), .ZN(n41904) );
  CLKNHSV6 U26378 ( .I(\pe1/bq[32] ), .ZN(n40558) );
  INHSV2 U26379 ( .I(n47539), .ZN(n29746) );
  BUFHSV6 U26380 ( .I(n45083), .Z(n59774) );
  CLKNAND2HSV4 U26381 ( .A1(n33689), .A2(n35311), .ZN(n33675) );
  NAND2HSV4 U26382 ( .A1(n33675), .A2(n33677), .ZN(n33684) );
  INHSV4 U26383 ( .I(n46299), .ZN(n25671) );
  NAND2HSV4 U26384 ( .A1(n26135), .A2(n56493), .ZN(n56330) );
  NAND3HSV4 U26385 ( .A1(n25323), .A2(n25321), .A3(n25322), .ZN(n46081) );
  XOR2HSV4 U26386 ( .A1(n46167), .A2(n26732), .Z(n46819) );
  CLKNHSV6 U26387 ( .I(n49173), .ZN(n53102) );
  CLKNAND2HSV2 U26388 ( .A1(n56058), .A2(n59384), .ZN(n56169) );
  XOR2HSV4 U26389 ( .A1(n46167), .A2(n26732), .Z(n46302) );
  OAI21HSV2 U26390 ( .A1(n42042), .A2(n41924), .B(n26850), .ZN(n42045) );
  BUFHSV6 U26391 ( .I(n59487), .Z(n58717) );
  NAND2HSV2 U26392 ( .A1(n34098), .A2(n25196), .ZN(n34100) );
  CLKNAND2HSV2 U26393 ( .A1(n34097), .A2(n34210), .ZN(n25196) );
  INHSV4 U26394 ( .I(n43748), .ZN(n25197) );
  NAND2HSV4 U26395 ( .A1(n44681), .A2(n26262), .ZN(n43748) );
  CLKNAND2HSV2 U26396 ( .A1(n48888), .A2(\pe6/got [8]), .ZN(n28758) );
  INHSV2 U26397 ( .I(n41593), .ZN(n41594) );
  NAND2HSV4 U26398 ( .A1(n59639), .A2(n47267), .ZN(n30635) );
  NAND2HSV2 U26399 ( .A1(n44151), .A2(n44152), .ZN(n44153) );
  INHSV6 U26400 ( .I(n45614), .ZN(n51119) );
  NAND2HSV4 U26401 ( .A1(n45610), .A2(n51119), .ZN(n25217) );
  CLKNAND2HSV4 U26402 ( .A1(n25667), .A2(n25666), .ZN(n36218) );
  NAND2HSV4 U26403 ( .A1(n26279), .A2(n35154), .ZN(n25342) );
  CLKNHSV2 U26404 ( .I(n56854), .ZN(n56899) );
  INHSV6 U26405 ( .I(n37351), .ZN(n37271) );
  NAND2HSV4 U26406 ( .A1(n37266), .A2(n42682), .ZN(n37351) );
  OAI21HSV4 U26407 ( .A1(n60004), .A2(n59586), .B(n36633), .ZN(n36634) );
  INHSV4 U26408 ( .I(n36847), .ZN(n36876) );
  INHSV2 U26409 ( .I(n30099), .ZN(n30253) );
  INHSV8 U26410 ( .I(n47992), .ZN(n37332) );
  CLKNAND2HSV4 U26411 ( .A1(n30099), .A2(n30142), .ZN(n30136) );
  CLKNAND2HSV4 U26412 ( .A1(n42332), .A2(n40975), .ZN(n42333) );
  INHSV4 U26413 ( .I(n42333), .ZN(n26283) );
  NAND2HSV2 U26414 ( .A1(n36094), .A2(n36093), .ZN(n36099) );
  CLKNAND2HSV2 U26415 ( .A1(n37453), .A2(n37452), .ZN(n37456) );
  CLKNAND2HSV3 U26416 ( .A1(n37259), .A2(n25670), .ZN(n26061) );
  CLKNAND2HSV3 U26417 ( .A1(n25951), .A2(n37272), .ZN(n37343) );
  CLKNAND2HSV2 U26418 ( .A1(n42917), .A2(n42933), .ZN(n42930) );
  CLKNHSV6 U26419 ( .I(n26418), .ZN(n47902) );
  CLKNAND2HSV4 U26420 ( .A1(n39568), .A2(n26648), .ZN(n39874) );
  NAND2HSV4 U26421 ( .A1(n26015), .A2(n43468), .ZN(n53376) );
  CLKNAND2HSV3 U26422 ( .A1(n25325), .A2(n25324), .ZN(n25323) );
  INHSV6 U26423 ( .I(n33088), .ZN(n35719) );
  NAND2HSV4 U26424 ( .A1(n38841), .A2(n52415), .ZN(n36427) );
  NAND2HSV4 U26425 ( .A1(n41506), .A2(n41505), .ZN(n41420) );
  CLKNHSV2 U26426 ( .I(n60028), .ZN(n44311) );
  XNOR2HSV4 U26427 ( .A1(n26800), .A2(n44181), .ZN(n60028) );
  CLKNAND2HSV2 U26428 ( .A1(n26608), .A2(n44304), .ZN(n44321) );
  CLKNAND2HSV4 U26429 ( .A1(n40511), .A2(n40526), .ZN(n40534) );
  NAND3HSV3 U26430 ( .A1(n46766), .A2(n46817), .A3(n53101), .ZN(n53185) );
  CLKNAND2HSV4 U26431 ( .A1(n26424), .A2(n26426), .ZN(n25982) );
  CLKNAND2HSV4 U26432 ( .A1(n52734), .A2(n30072), .ZN(n26426) );
  XNOR2HSV4 U26433 ( .A1(n34192), .A2(n34191), .ZN(n34227) );
  XNOR2HSV4 U26434 ( .A1(n34188), .A2(n34189), .ZN(n34191) );
  INHSV2 U26435 ( .I(n46302), .ZN(n49177) );
  CLKNAND2HSV2 U26436 ( .A1(n43364), .A2(n43365), .ZN(n43368) );
  CLKNAND2HSV2 U26437 ( .A1(n43600), .A2(n43603), .ZN(n43601) );
  CLKNAND2HSV2 U26438 ( .A1(n25212), .A2(n43890), .ZN(n43895) );
  XNOR2HSV4 U26439 ( .A1(n25198), .A2(n42686), .ZN(n42688) );
  XNOR2HSV4 U26440 ( .A1(n42681), .A2(n42680), .ZN(n25198) );
  NAND2HSV2 U26441 ( .A1(n34578), .A2(n34837), .ZN(n34579) );
  NAND2HSV4 U26442 ( .A1(n40436), .A2(n25199), .ZN(n40479) );
  NAND3HSV4 U26443 ( .A1(n40296), .A2(n40294), .A3(n40295), .ZN(n40317) );
  CLKNAND2HSV2 U26444 ( .A1(n43020), .A2(n43019), .ZN(n43133) );
  AOI22HSV4 U26445 ( .A1(n46559), .A2(\pe3/ti_7t [19]), .B1(n42805), .B2(
        n45799), .ZN(n43020) );
  INHSV8 U26446 ( .I(n25200), .ZN(n46766) );
  NOR2HSV4 U26447 ( .A1(n46307), .A2(n49402), .ZN(n25200) );
  CLKNAND2HSV2 U26448 ( .A1(n43122), .A2(n43121), .ZN(n43123) );
  CLKNAND2HSV2 U26449 ( .A1(n25201), .A2(n33082), .ZN(n33083) );
  CLKNHSV2 U26450 ( .I(n25202), .ZN(n25201) );
  CLKNAND2HSV2 U26451 ( .A1(n33081), .A2(n33080), .ZN(n25202) );
  CLKNHSV2 U26452 ( .I(n25203), .ZN(n33072) );
  CLKNAND2HSV2 U26453 ( .A1(n33084), .A2(n35798), .ZN(n25203) );
  INHSV4 U26454 ( .I(n30017), .ZN(n26141) );
  INHSV8 U26455 ( .I(n25262), .ZN(n34844) );
  OAI21HSV4 U26456 ( .A1(n25204), .A2(n37923), .B(n36250), .ZN(n36666) );
  XNOR2HSV4 U26457 ( .A1(n25205), .A2(n36662), .ZN(n25204) );
  XNOR2HSV4 U26458 ( .A1(n36663), .A2(n36664), .ZN(n25205) );
  INAND2HSV4 U26459 ( .A1(n38002), .B1(n38603), .ZN(n38018) );
  NAND2HSV4 U26460 ( .A1(n44668), .A2(n44666), .ZN(n25647) );
  CLKNHSV2 U26461 ( .I(n51451), .ZN(n25648) );
  XNOR2HSV4 U26462 ( .A1(n33069), .A2(n33068), .ZN(n51451) );
  NAND2HSV4 U26463 ( .A1(n25599), .A2(n35708), .ZN(n35709) );
  XNOR2HSV4 U26464 ( .A1(n44363), .A2(n44362), .ZN(n44364) );
  CLKNAND2HSV4 U26465 ( .A1(n32459), .A2(n36095), .ZN(n32412) );
  CLKAND2HSV2 U26466 ( .A1(n37918), .A2(n38264), .Z(n36660) );
  CLKNAND2HSV4 U26467 ( .A1(n60018), .A2(n53649), .ZN(n29016) );
  XNOR2HSV1 U26468 ( .A1(n26713), .A2(n26712), .ZN(\pe2/poht [18]) );
  NAND2HSV4 U26469 ( .A1(n44650), .A2(n40438), .ZN(n42331) );
  XNOR2HSV4 U26470 ( .A1(n26544), .A2(n25206), .ZN(n40318) );
  CLKNAND2HSV2 U26471 ( .A1(n29744), .A2(n48885), .ZN(n25206) );
  INHSV2 U26472 ( .I(n34320), .ZN(n34325) );
  NOR2HSV4 U26473 ( .A1(n34325), .A2(n34324), .ZN(n34347) );
  CLKNAND2HSV2 U26474 ( .A1(n34575), .A2(n34581), .ZN(n34968) );
  CLKNAND2HSV2 U26475 ( .A1(n34969), .A2(n34968), .ZN(n34973) );
  AOI21HSV4 U26476 ( .A1(n46310), .A2(n26259), .B(n44679), .ZN(n44687) );
  INHSV4 U26477 ( .I(n43870), .ZN(n46559) );
  CLKNAND2HSV2 U26478 ( .A1(n43912), .A2(\pe3/ti_7t [15]), .ZN(n42700) );
  CLKBUFHSV12 U26479 ( .I(n43752), .Z(n46090) );
  BUFHSV2 U26480 ( .I(n31759), .Z(n26586) );
  NAND3HSV4 U26481 ( .A1(n32519), .A2(n32351), .A3(n32352), .ZN(n32459) );
  CLKNAND2HSV4 U26482 ( .A1(n59536), .A2(n43355), .ZN(n43241) );
  INHSV4 U26483 ( .I(n43465), .ZN(n25767) );
  CLKNAND2HSV4 U26484 ( .A1(n25768), .A2(n25767), .ZN(n43472) );
  CLKNAND2HSV2 U26485 ( .A1(n43479), .A2(n43355), .ZN(n25207) );
  CLKNAND2HSV4 U26486 ( .A1(n25208), .A2(n31480), .ZN(n31515) );
  NAND2HSV2 U26487 ( .A1(n31478), .A2(n35914), .ZN(n25208) );
  NAND2HSV4 U26488 ( .A1(n25209), .A2(n38885), .ZN(n38005) );
  NAND2HSV2 U26489 ( .A1(n37864), .A2(n36319), .ZN(n25209) );
  CLKNAND2HSV2 U26490 ( .A1(n38012), .A2(n38109), .ZN(n47979) );
  INHSV2 U26491 ( .I(n25537), .ZN(n25536) );
  MUX2NHSV4 U26492 ( .I0(n25536), .I1(n25534), .S(n26423), .ZN(n25533) );
  INHSV4 U26493 ( .I(n37983), .ZN(n38006) );
  OAI21HSV4 U26494 ( .A1(n46532), .A2(n43891), .B(n43134), .ZN(n25692) );
  CLKNAND2HSV2 U26495 ( .A1(n31949), .A2(n31667), .ZN(n31619) );
  AOI21HSV2 U26496 ( .A1(n33804), .A2(n25725), .B(n33803), .ZN(n33846) );
  CLKNAND2HSV4 U26497 ( .A1(n25920), .A2(n25921), .ZN(n25345) );
  NAND2HSV4 U26498 ( .A1(n25919), .A2(n25345), .ZN(n38894) );
  NAND2HSV4 U26499 ( .A1(n42489), .A2(n42488), .ZN(n26042) );
  INHSV4 U26500 ( .I(n26042), .ZN(n26037) );
  XNOR2HSV4 U26501 ( .A1(n34954), .A2(n34953), .ZN(n34957) );
  INHSV4 U26502 ( .I(n36967), .ZN(n43126) );
  INHSV8 U26503 ( .I(n35704), .ZN(n47934) );
  NAND2HSV4 U26504 ( .A1(n32320), .A2(n32164), .ZN(n32225) );
  INHSV4 U26505 ( .I(n38875), .ZN(n38871) );
  NAND2HSV2 U26506 ( .A1(n26852), .A2(n25210), .ZN(n38641) );
  INHSV4 U26507 ( .I(n38768), .ZN(n25210) );
  NOR2HSV2 U26508 ( .A1(n44043), .A2(n38887), .ZN(n38768) );
  INHSV4 U26509 ( .I(n25628), .ZN(n25629) );
  CLKNHSV6 U26510 ( .I(n31339), .ZN(n31269) );
  NOR2HSV2 U26511 ( .A1(n30140), .A2(n30141), .ZN(n25985) );
  CLKNAND2HSV2 U26512 ( .A1(n26426), .A2(n26425), .ZN(n30141) );
  CLKNAND2HSV4 U26513 ( .A1(n60019), .A2(n44315), .ZN(n38016) );
  CLKNAND2HSV3 U26514 ( .A1(n43883), .A2(n43882), .ZN(n44676) );
  CLKNAND2HSV1 U26515 ( .A1(n45599), .A2(n43484), .ZN(n43889) );
  NAND2HSV2 U26516 ( .A1(n43889), .A2(n43892), .ZN(n25212) );
  INHSV4 U26517 ( .I(n32446), .ZN(n32449) );
  NAND2HSV4 U26518 ( .A1(n32448), .A2(n32449), .ZN(n32450) );
  CLKNAND2HSV2 U26519 ( .A1(n32535), .A2(n32534), .ZN(n32536) );
  NOR2HSV4 U26520 ( .A1(n32814), .A2(n44372), .ZN(n32452) );
  NAND2HSV2 U26521 ( .A1(n32524), .A2(n32523), .ZN(n32525) );
  XNOR2HSV4 U26522 ( .A1(n25213), .A2(n32641), .ZN(n25568) );
  XNOR2HSV4 U26523 ( .A1(n25569), .A2(n32639), .ZN(n25213) );
  CLKAND2HSV4 U26524 ( .A1(n43493), .A2(n36671), .Z(n43488) );
  NAND2HSV4 U26525 ( .A1(n56063), .A2(n43608), .ZN(n45503) );
  CLKNAND2HSV4 U26526 ( .A1(n25214), .A2(n31704), .ZN(n31898) );
  CLKNAND2HSV4 U26527 ( .A1(n31703), .A2(n31702), .ZN(n25214) );
  CLKNAND2HSV4 U26528 ( .A1(n56965), .A2(\pe3/got [20]), .ZN(n26205) );
  CLKNAND2HSV2 U26529 ( .A1(n31591), .A2(n31590), .ZN(n31616) );
  AOI21HSV2 U26530 ( .A1(n31516), .A2(n31517), .B(n31515), .ZN(n31484) );
  NAND2HSV4 U26531 ( .A1(n29870), .A2(n29869), .ZN(n29933) );
  INHSV4 U26532 ( .I(n45930), .ZN(n46116) );
  INHSV4 U26533 ( .I(n31253), .ZN(n59276) );
  CLKNAND2HSV4 U26534 ( .A1(n26834), .A2(n30397), .ZN(n30423) );
  BUFHSV6 U26535 ( .I(n55213), .Z(n55332) );
  NAND3HSV4 U26536 ( .A1(n32525), .A2(n32527), .A3(n32526), .ZN(n32528) );
  NAND2HSV4 U26537 ( .A1(n30023), .A2(n30022), .ZN(n25307) );
  BUFHSV8 U26538 ( .I(n40446), .Z(n40416) );
  CLKNAND2HSV4 U26539 ( .A1(n34583), .A2(n34834), .ZN(n34342) );
  CLKNAND2HSV2 U26540 ( .A1(n34218), .A2(n34436), .ZN(n34097) );
  NOR2HSV4 U26541 ( .A1(n34967), .A2(n34726), .ZN(n34856) );
  INAND2HSV4 U26542 ( .A1(n34856), .B1(n34855), .ZN(n34857) );
  OAI31HSV2 U26543 ( .A1(n50752), .A2(n29521), .A3(n43457), .B(n29522), .ZN(
        n29523) );
  NAND2HSV2 U26544 ( .A1(n29523), .A2(n29524), .ZN(n29525) );
  INHSV2 U26545 ( .I(n45754), .ZN(n25215) );
  NOR2HSV4 U26546 ( .A1(n25215), .A2(n43912), .ZN(n46087) );
  CLKNAND2HSV2 U26547 ( .A1(n25217), .A2(n27521), .ZN(n46101) );
  NAND2HSV4 U26548 ( .A1(n43611), .A2(n43612), .ZN(n43751) );
  CLKNAND2HSV2 U26549 ( .A1(n45599), .A2(n45779), .ZN(n43886) );
  INHSV4 U26550 ( .I(n43912), .ZN(n45779) );
  OAI21HSV4 U26551 ( .A1(n32549), .A2(n32548), .B(n32547), .ZN(n32550) );
  NAND2HSV4 U26552 ( .A1(n31287), .A2(n31286), .ZN(n31353) );
  INHSV4 U26553 ( .I(n31353), .ZN(n31354) );
  NAND2HSV4 U26554 ( .A1(n31259), .A2(n31258), .ZN(n31265) );
  DELHS1 U26555 ( .I(n59011), .Z(n25218) );
  NAND2HSV2 U26556 ( .A1(n40636), .A2(n40700), .ZN(n40469) );
  NOR2HSV2 U26557 ( .A1(n47953), .A2(n32949), .ZN(n29637) );
  MUX2NHSV4 U26558 ( .I0(n25662), .I1(n25219), .S(n25661), .ZN(n25660) );
  INHSV2 U26559 ( .I(n25220), .ZN(n25219) );
  INAND2HSV2 U26560 ( .A1(n32241), .B1(n46824), .ZN(n25220) );
  BUFHSV24 U26561 ( .I(n26413), .Z(n26761) );
  NOR2HSV4 U26562 ( .A1(n26761), .A2(n35319), .ZN(n50061) );
  INHSV6 U26563 ( .I(n46118), .ZN(n55820) );
  INHSV4 U26564 ( .I(n55820), .ZN(n56935) );
  NAND2HSV4 U26565 ( .A1(n40507), .A2(n40508), .ZN(n40526) );
  XNOR2HSV4 U26566 ( .A1(n25221), .A2(n26195), .ZN(n40590) );
  XNOR2HSV4 U26567 ( .A1(n26196), .A2(n26197), .ZN(n25221) );
  CLKNAND2HSV4 U26568 ( .A1(n40360), .A2(n40359), .ZN(n40396) );
  CLKNAND2HSV4 U26569 ( .A1(n40396), .A2(n40467), .ZN(n40410) );
  XNOR2HSV4 U26570 ( .A1(n53209), .A2(n53208), .ZN(n53213) );
  NOR2HSV4 U26571 ( .A1(n26761), .A2(n58253), .ZN(n50124) );
  NAND2HSV4 U26572 ( .A1(n26756), .A2(n25222), .ZN(n26755) );
  INHSV4 U26573 ( .I(n25223), .ZN(n25222) );
  NAND2HSV4 U26574 ( .A1(n35481), .A2(n46566), .ZN(n25223) );
  XNOR2HSV4 U26575 ( .A1(n26138), .A2(n26137), .ZN(n25224) );
  NAND3HSV3 U26576 ( .A1(n25496), .A2(n47953), .A3(n32951), .ZN(n32954) );
  INHSV2 U26577 ( .I(n43494), .ZN(n45583) );
  CLKNHSV0 U26578 ( .I(n43494), .ZN(n56066) );
  XNOR2HSV4 U26579 ( .A1(n40452), .A2(n40451), .ZN(n40463) );
  CLKNAND2HSV2 U26580 ( .A1(n40910), .A2(n40923), .ZN(n40629) );
  INHSV2 U26581 ( .I(n32814), .ZN(n46631) );
  CLKNAND2HSV4 U26582 ( .A1(n46631), .A2(n32815), .ZN(n32825) );
  CLKXOR2HSV4 U26583 ( .A1(n58203), .A2(n58202), .Z(n58205) );
  CLKXOR2HSV4 U26584 ( .A1(n58245), .A2(n58244), .Z(n58248) );
  CLKXOR2HSV4 U26585 ( .A1(n50101), .A2(n50100), .Z(n50103) );
  XOR2HSV4 U26586 ( .A1(n47988), .A2(n30304), .Z(n30200) );
  CLKNAND2HSV4 U26587 ( .A1(n26620), .A2(n26619), .ZN(pov1[22]) );
  CLKNAND2HSV8 U26588 ( .A1(pov1[22]), .A2(n42471), .ZN(n42051) );
  CLKNAND2HSV4 U26589 ( .A1(n29983), .A2(n29982), .ZN(n60040) );
  CLKNAND2HSV4 U26590 ( .A1(n60040), .A2(n31086), .ZN(n30060) );
  NAND2HSV2 U26591 ( .A1(n60028), .A2(n44308), .ZN(n44955) );
  CLKNAND2HSV4 U26592 ( .A1(n36046), .A2(n36045), .ZN(n47940) );
  INHSV4 U26593 ( .I(n47940), .ZN(n36079) );
  NAND2HSV2 U26594 ( .A1(n30099), .A2(n52799), .ZN(n52735) );
  CLKNHSV0 U26595 ( .I(n52735), .ZN(n30071) );
  XNOR2HSV4 U26596 ( .A1(n44811), .A2(n44810), .ZN(n44813) );
  CLKNHSV6 U26597 ( .I(n45617), .ZN(n45610) );
  NAND2HSV2 U26598 ( .A1(n26398), .A2(n26397), .ZN(n45605) );
  NOR2HSV4 U26599 ( .A1(n25281), .A2(n34104), .ZN(n34231) );
  NAND3HSV3 U26600 ( .A1(n53102), .A2(n46766), .A3(n49174), .ZN(n49249) );
  NOR2HSV4 U26601 ( .A1(n30506), .A2(n30419), .ZN(n30420) );
  INHSV4 U26602 ( .I(n49661), .ZN(n53095) );
  OAI31HSV2 U26603 ( .A1(n36799), .A2(n28974), .A3(n28959), .B(n28975), .ZN(
        n28976) );
  NOR2HSV3 U26604 ( .A1(n44668), .A2(n44667), .ZN(n25639) );
  CLKNHSV6 U26605 ( .I(n29890), .ZN(n29815) );
  CLKNAND2HSV8 U26606 ( .A1(n60013), .A2(n44309), .ZN(n26235) );
  CLKNAND2HSV8 U26607 ( .A1(n26235), .A2(n45138), .ZN(n49661) );
  INHSV2 U26608 ( .I(n45584), .ZN(n45586) );
  CLKNAND2HSV2 U26609 ( .A1(n42077), .A2(n42068), .ZN(n42047) );
  NAND2HSV4 U26610 ( .A1(n42048), .A2(n42047), .ZN(n42057) );
  CLKNAND2HSV1 U26611 ( .A1(n59515), .A2(n51011), .ZN(n43890) );
  CLKNHSV2 U26612 ( .I(n25225), .ZN(n46106) );
  CLKNAND2HSV2 U26613 ( .A1(n50716), .A2(n46107), .ZN(n25225) );
  INHSV6 U26614 ( .I(\pe1/bq[30] ), .ZN(n40411) );
  CLKBUFHSV12 U26615 ( .I(n53530), .Z(n25226) );
  NAND3HSV3 U26616 ( .A1(n53102), .A2(n46766), .A3(n46765), .ZN(n46767) );
  CLKNAND2HSV4 U26617 ( .A1(n42075), .A2(n42050), .ZN(n42080) );
  NAND3HSV4 U26618 ( .A1(n42080), .A2(n42055), .A3(n42064), .ZN(n42056) );
  NAND2HSV2 U26619 ( .A1(n25234), .A2(n26224), .ZN(n25233) );
  INOR2HSV4 U26620 ( .A1(n46553), .B1(n46168), .ZN(n46298) );
  CLKNAND2HSV2 U26621 ( .A1(n60086), .A2(n25227), .ZN(n43028) );
  CLKNHSV2 U26622 ( .I(n25801), .ZN(n25227) );
  NAND2HSV4 U26623 ( .A1(n25228), .A2(n38355), .ZN(n38336) );
  INHSV2 U26624 ( .I(n25721), .ZN(n25228) );
  OAI21HSV4 U26625 ( .A1(n29954), .A2(n29953), .B(n29952), .ZN(n29955) );
  NAND2HSV4 U26626 ( .A1(n33673), .A2(n33672), .ZN(n33689) );
  NOR2HSV4 U26627 ( .A1(n38006), .A2(n38007), .ZN(n38008) );
  NAND2HSV4 U26628 ( .A1(n38008), .A2(n38009), .ZN(n38033) );
  AOI22HSV2 U26629 ( .A1(n25229), .A2(n36584), .B1(n36582), .B2(n38340), .ZN(
        n36579) );
  CLKNHSV2 U26630 ( .I(n36576), .ZN(n25229) );
  INHSV4 U26631 ( .I(n43256), .ZN(n59571) );
  INHSV2 U26632 ( .I(n37784), .ZN(n42694) );
  NOR2HSV2 U26633 ( .A1(n43744), .A2(n43891), .ZN(n43141) );
  INHSV2 U26634 ( .I(n43136), .ZN(n43137) );
  AOI21HSV2 U26635 ( .A1(n25230), .A2(n32673), .B(n32552), .ZN(n32553) );
  NOR2HSV4 U26636 ( .A1(n32674), .A2(n32550), .ZN(n25230) );
  INHSV2 U26637 ( .I(n42064), .ZN(n42065) );
  CLKNHSV0 U26638 ( .I(n29826), .ZN(n30918) );
  NAND2HSV4 U26639 ( .A1(n26568), .A2(n38520), .ZN(n38524) );
  NAND2HSV4 U26640 ( .A1(n48049), .A2(\pe5/pvq [4]), .ZN(n29903) );
  XNOR2HSV2 U26641 ( .A1(n50751), .A2(n50750), .ZN(n50755) );
  INHSV8 U26642 ( .I(n55944), .ZN(n56682) );
  NOR2HSV4 U26643 ( .A1(n46100), .A2(n56682), .ZN(n46102) );
  NAND2HSV2 U26644 ( .A1(n26063), .A2(n46092), .ZN(n45758) );
  NOR2HSV2 U26645 ( .A1(n42320), .A2(n42329), .ZN(n42321) );
  XNOR2HSV4 U26646 ( .A1(n42325), .A2(n42324), .ZN(n42320) );
  XNOR2HSV4 U26647 ( .A1(n25232), .A2(n25231), .ZN(n53284) );
  CLKNAND2HSV2 U26648 ( .A1(n53279), .A2(n43829), .ZN(n25231) );
  XNOR2HSV4 U26649 ( .A1(n53281), .A2(n53280), .ZN(n25232) );
  CLKNAND2HSV4 U26650 ( .A1(n35428), .A2(n59956), .ZN(n34562) );
  NAND2HSV4 U26651 ( .A1(n34562), .A2(n34561), .ZN(n34563) );
  CLKNAND2HSV4 U26652 ( .A1(n42057), .A2(n42056), .ZN(n42466) );
  CLKNAND2HSV2 U26653 ( .A1(n42466), .A2(n42200), .ZN(n42201) );
  XNOR2HSV4 U26654 ( .A1(n44275), .A2(n44274), .ZN(n44277) );
  XOR3HSV4 U26655 ( .A1(n44278), .A2(n44277), .A3(n44276), .Z(n44279) );
  NAND2HSV4 U26656 ( .A1(n44677), .A2(n25233), .ZN(n45944) );
  NOR2HSV0 U26657 ( .A1(n25639), .A2(n45607), .ZN(n25234) );
  INHSV4 U26658 ( .I(n56778), .ZN(n56888) );
  CLKNAND2HSV4 U26659 ( .A1(n44514), .A2(n46567), .ZN(n44367) );
  NAND2HSV2 U26660 ( .A1(n44361), .A2(n44360), .ZN(n44514) );
  NAND2HSV4 U26661 ( .A1(n25671), .A2(n46303), .ZN(n46304) );
  INHSV2 U26662 ( .I(n38756), .ZN(n38761) );
  NAND3HSV3 U26663 ( .A1(n38760), .A2(n38761), .A3(n26626), .ZN(n38762) );
  XNOR2HSV4 U26664 ( .A1(n25235), .A2(n25643), .ZN(n29357) );
  CLKNAND2HSV2 U26665 ( .A1(n25644), .A2(n29356), .ZN(n25235) );
  INHSV2 U26666 ( .I(n45771), .ZN(n25236) );
  INHSV2 U26667 ( .I(n45772), .ZN(n25237) );
  NOR2HSV2 U26668 ( .A1(n46089), .A2(n45764), .ZN(n45772) );
  CLKNAND2HSV4 U26669 ( .A1(n48328), .A2(n25238), .ZN(n48335) );
  CLKNHSV2 U26670 ( .I(n48329), .ZN(n25238) );
  NOR2HSV4 U26671 ( .A1(n42476), .A2(n42477), .ZN(n48329) );
  NOR2HSV4 U26672 ( .A1(n58437), .A2(n58435), .ZN(n46301) );
  NOR2HSV4 U26673 ( .A1(n42354), .A2(n42083), .ZN(n26078) );
  NOR2HSV4 U26674 ( .A1(n26079), .A2(n42082), .ZN(n42354) );
  CLKXOR2HSV4 U26675 ( .A1(n56883), .A2(n56882), .Z(n56884) );
  CLKXOR2HSV2 U26676 ( .A1(n56885), .A2(n56884), .Z(n56886) );
  IOA21HSV4 U26677 ( .A1(n26510), .A2(n26512), .B(n26511), .ZN(n26507) );
  XNOR2HSV4 U26678 ( .A1(n44144), .A2(n25239), .ZN(n44147) );
  XNOR2HSV4 U26679 ( .A1(n44141), .A2(n44142), .ZN(n25239) );
  XNOR2HSV4 U26680 ( .A1(n55698), .A2(n25240), .ZN(n55699) );
  XNOR2HSV4 U26681 ( .A1(n55696), .A2(n55697), .ZN(n25240) );
  XNOR2HSV4 U26682 ( .A1(n44365), .A2(n36219), .ZN(n36220) );
  CLKNAND2HSV2 U26683 ( .A1(n28424), .A2(n45593), .ZN(n45594) );
  NAND2HSV4 U26684 ( .A1(n45594), .A2(n25472), .ZN(n45601) );
  NAND2HSV4 U26685 ( .A1(n59576), .A2(n44649), .ZN(n41045) );
  OAI21HSV4 U26686 ( .A1(n37332), .A2(n45622), .B(n37331), .ZN(n37333) );
  INHSV4 U26687 ( .I(n37333), .ZN(n37339) );
  INHSV24 U26688 ( .I(n26097), .ZN(n25241) );
  CLKAND2HSV2 U26689 ( .A1(n60020), .A2(n25241), .Z(n38459) );
  INHSV2 U26690 ( .I(n25242), .ZN(n29677) );
  CLKNAND2HSV2 U26691 ( .A1(n32927), .A2(n32821), .ZN(n25242) );
  CLKAND2HSV4 U26692 ( .A1(n37236), .A2(n43126), .Z(n29691) );
  NAND2HSV4 U26693 ( .A1(n29691), .A2(n37237), .ZN(n37334) );
  NOR2HSV4 U26694 ( .A1(n36975), .A2(n36974), .ZN(n36986) );
  INHSV4 U26695 ( .I(n42683), .ZN(n56057) );
  INHSV4 U26696 ( .I(n56680), .ZN(n56177) );
  INHSV4 U26697 ( .I(n50802), .ZN(n56176) );
  CLKXOR2HSV4 U26698 ( .A1(n43012), .A2(n43011), .Z(n43014) );
  DELHS1 U26699 ( .I(n50384), .Z(n25243) );
  CLKNAND2HSV4 U26700 ( .A1(n45516), .A2(n43141), .ZN(n26551) );
  INHSV4 U26701 ( .I(n56682), .ZN(n26151) );
  INHSV2 U26702 ( .I(n50717), .ZN(n56863) );
  CLKNAND2HSV4 U26703 ( .A1(n37090), .A2(n37513), .ZN(n37098) );
  CLKNAND2HSV4 U26704 ( .A1(n37334), .A2(n37089), .ZN(n37513) );
  NAND2HSV4 U26705 ( .A1(n60015), .A2(n25358), .ZN(n48326) );
  INHSV4 U26706 ( .I(n35560), .ZN(n26795) );
  INHSV4 U26707 ( .I(n32447), .ZN(n32448) );
  OAI21HSV4 U26708 ( .A1(n30163), .A2(n39166), .B(n37664), .ZN(n29896) );
  NAND2HSV2 U26709 ( .A1(n25244), .A2(n42607), .ZN(n25261) );
  NOR2HSV2 U26710 ( .A1(n52789), .A2(n42604), .ZN(n25244) );
  NAND2HSV4 U26711 ( .A1(n36775), .A2(n43905), .ZN(n36774) );
  CLKNAND2HSV2 U26712 ( .A1(n25246), .A2(n25245), .ZN(n52796) );
  CLKNHSV2 U26713 ( .I(n47972), .ZN(n25245) );
  CLKNHSV2 U26714 ( .I(n34002), .ZN(n25246) );
  CLKNAND2HSV2 U26715 ( .A1(n33989), .A2(n25247), .ZN(n34002) );
  CLKNHSV2 U26716 ( .I(n34221), .ZN(n25247) );
  INHSV4 U26717 ( .I(n36537), .ZN(n36547) );
  NAND2HSV4 U26718 ( .A1(n33444), .A2(n33450), .ZN(n33410) );
  INAND2HSV4 U26719 ( .A1(n31044), .B1(n30164), .ZN(n30261) );
  CLKXOR2HSV2 U26720 ( .A1(n29960), .A2(n30261), .Z(n29964) );
  CLKNAND2HSV3 U26721 ( .A1(n36923), .A2(n45612), .ZN(n25941) );
  CLKNHSV3 U26722 ( .I(n46150), .ZN(n46162) );
  INHSV8 U26723 ( .I(n38523), .ZN(n38026) );
  CLKNHSV12 U26724 ( .I(n37931), .ZN(n45265) );
  BUFHSV4 U26725 ( .I(n34446), .Z(n47969) );
  CLKNAND2HSV4 U26726 ( .A1(n46152), .A2(n46151), .ZN(n58369) );
  INHSV4 U26727 ( .I(n40528), .ZN(n40507) );
  NAND2HSV2 U26728 ( .A1(n58812), .A2(n58476), .ZN(n28186) );
  OAI21HSV2 U26729 ( .A1(n28185), .A2(n28186), .B(n28187), .ZN(\pe6/poht [22])
         );
  NAND2HSV4 U26730 ( .A1(n59665), .A2(n34966), .ZN(n34818) );
  INHSV2 U26731 ( .I(\pe1/aot [32]), .ZN(n40493) );
  MUX2NHSV2 U26732 ( .I0(n29949), .I1(n52716), .S(n29948), .ZN(n29953) );
  AOI31HSV2 U26733 ( .A1(n34700), .A2(n59345), .A3(n34701), .B(n25248), .ZN(
        n34703) );
  CLKNAND2HSV2 U26734 ( .A1(n34698), .A2(n25249), .ZN(n25248) );
  CLKNAND2HSV2 U26735 ( .A1(n25251), .A2(n25250), .ZN(n25249) );
  CLKNHSV2 U26736 ( .I(n34699), .ZN(n25250) );
  CLKNHSV2 U26737 ( .I(n34727), .ZN(n25251) );
  CLKNAND2HSV2 U26738 ( .A1(n57308), .A2(n34864), .ZN(n34552) );
  CLKXOR2HSV2 U26739 ( .A1(n34552), .A2(n34551), .Z(n34553) );
  NAND2HSV4 U26740 ( .A1(n32544), .A2(n32545), .ZN(n32462) );
  CLKNAND2HSV4 U26741 ( .A1(n26468), .A2(n25252), .ZN(n32544) );
  NAND2HSV4 U26742 ( .A1(n25254), .A2(n25253), .ZN(n25252) );
  INHSV2 U26743 ( .I(n32458), .ZN(n25253) );
  INHSV2 U26744 ( .I(n26469), .ZN(n25254) );
  INHSV4 U26745 ( .I(n43706), .ZN(n56475) );
  XNOR2HSV2 U26746 ( .A1(n26592), .A2(\pe3/phq [4]), .ZN(n26591) );
  AOI21HSV2 U26747 ( .A1(n29674), .A2(n33697), .B(n33696), .ZN(n33698) );
  CLKNAND2HSV2 U26748 ( .A1(n36861), .A2(n36737), .ZN(n36743) );
  AOI31HSV2 U26749 ( .A1(n43592), .A2(n25800), .A3(n43363), .B(n43362), .ZN(
        n25255) );
  CLKNHSV6 U26750 ( .I(n33594), .ZN(n35560) );
  INHSV4 U26751 ( .I(n35560), .ZN(n33603) );
  INHSV4 U26752 ( .I(n25257), .ZN(n25256) );
  CLKNAND2HSV4 U26753 ( .A1(n43344), .A2(n44664), .ZN(n25257) );
  CLKNAND2HSV2 U26754 ( .A1(n33219), .A2(n33220), .ZN(n33223) );
  NAND3HSV2 U26755 ( .A1(n31129), .A2(n31134), .A3(n31128), .ZN(n31132) );
  XNOR2HSV4 U26756 ( .A1(n25260), .A2(n25258), .ZN(n33580) );
  XNOR2HSV4 U26757 ( .A1(n25259), .A2(n33566), .ZN(n25258) );
  XNOR2HSV4 U26758 ( .A1(n33568), .A2(n33567), .ZN(n25259) );
  NOR2HSV4 U26759 ( .A1(n33529), .A2(n33530), .ZN(n25260) );
  XNOR2HSV4 U26760 ( .A1(n32837), .A2(n32836), .ZN(n32839) );
  MUX2NHSV2 U26761 ( .I0(n32840), .I1(n58901), .S(n32839), .ZN(n32919) );
  OA21HSV4 U26762 ( .A1(n36873), .A2(\pe3/ti_7t [10]), .B(n44669), .Z(n37155)
         );
  BUFHSV4 U26763 ( .I(n43226), .Z(n43453) );
  CLKNAND2HSV3 U26764 ( .A1(n31281), .A2(n31280), .ZN(n31324) );
  NAND2HSV4 U26765 ( .A1(n42797), .A2(n25261), .ZN(n42802) );
  INHSV3 U26766 ( .I(n42611), .ZN(n42615) );
  INHSV6 U26767 ( .I(n34711), .ZN(n25262) );
  INHSV2 U26768 ( .I(n33193), .ZN(n26047) );
  INHSV4 U26769 ( .I(n36780), .ZN(n36928) );
  NAND2HSV2 U26770 ( .A1(n36728), .A2(n36727), .ZN(n36731) );
  INHSV4 U26771 ( .I(n38881), .ZN(n25263) );
  CLKNAND2HSV4 U26772 ( .A1(n25931), .A2(n25264), .ZN(n38881) );
  CLKNAND2HSV4 U26773 ( .A1(n25266), .A2(n25265), .ZN(n25264) );
  INHSV2 U26774 ( .I(n25932), .ZN(n25265) );
  INHSV4 U26775 ( .I(n25934), .ZN(n25266) );
  INHSV2 U26776 ( .I(n43490), .ZN(n25766) );
  OAI21HSV4 U26777 ( .A1(n38172), .A2(n38173), .B(n25267), .ZN(n38182) );
  CLKNAND2HSV2 U26778 ( .A1(n38170), .A2(n25268), .ZN(n25267) );
  CLKNHSV2 U26779 ( .I(n38171), .ZN(n25268) );
  CLKNHSV6 U26780 ( .I(n40443), .ZN(n40324) );
  INHSV6 U26781 ( .I(n40324), .ZN(n40569) );
  NOR2HSV4 U26782 ( .A1(n34684), .A2(n57453), .ZN(n34682) );
  CLKNHSV0 U26783 ( .I(n34682), .ZN(n34680) );
  XNOR2HSV4 U26784 ( .A1(n25269), .A2(n30972), .ZN(n30984) );
  XNOR2HSV4 U26785 ( .A1(n30963), .A2(n30964), .ZN(n25269) );
  NAND2HSV4 U26786 ( .A1(n25270), .A2(n32335), .ZN(n32512) );
  INHSV2 U26787 ( .I(n32333), .ZN(n25270) );
  NAND2HSV2 U26788 ( .A1(n32048), .A2(n32047), .ZN(n32333) );
  INHSV4 U26789 ( .I(n37791), .ZN(n52934) );
  CLKXOR2HSV4 U26790 ( .A1(n32129), .A2(n32128), .Z(n32132) );
  NAND2HSV4 U26791 ( .A1(n60005), .A2(n36509), .ZN(n36510) );
  CLKNAND2HSV2 U26792 ( .A1(n34218), .A2(n35032), .ZN(n34188) );
  XNOR2HSV4 U26793 ( .A1(n25273), .A2(n25271), .ZN(n35266) );
  XOR2HSV2 U26794 ( .A1(n35264), .A2(n25272), .Z(n25271) );
  CLKNHSV2 U26795 ( .I(n35263), .ZN(n25272) );
  CLKNAND2HSV2 U26796 ( .A1(n35577), .A2(n35318), .ZN(n25273) );
  OAI21HSV2 U26797 ( .A1(n45272), .A2(n25274), .B(n45269), .ZN(n45270) );
  CLKNAND2HSV2 U26798 ( .A1(n45266), .A2(n45265), .ZN(n25274) );
  INHSV4 U26799 ( .I(n33219), .ZN(n33222) );
  NAND2HSV4 U26800 ( .A1(n33222), .A2(n33221), .ZN(n25454) );
  XNOR2HSV4 U26801 ( .A1(n45387), .A2(n45386), .ZN(n45391) );
  CLKNAND2HSV4 U26802 ( .A1(n25276), .A2(n25275), .ZN(n32429) );
  CLKNAND2HSV2 U26803 ( .A1(n32309), .A2(n32310), .ZN(n25275) );
  CLKNAND2HSV4 U26804 ( .A1(n32312), .A2(n32311), .ZN(n25276) );
  XNOR2HSV1 U26805 ( .A1(n25279), .A2(n25277), .ZN(n60016) );
  INHSV2 U26806 ( .I(n25278), .ZN(n25277) );
  AOI21HSV2 U26807 ( .A1(n51150), .A2(n51151), .B(n51800), .ZN(n25278) );
  CLKXOR2HSV2 U26808 ( .A1(n25280), .A2(n51153), .Z(n25279) );
  XOR2HSV4 U26809 ( .A1(n51152), .A2(n51154), .Z(n25280) );
  NAND2HSV4 U26810 ( .A1(n40355), .A2(n40354), .ZN(n40360) );
  NAND2HSV4 U26811 ( .A1(n34320), .A2(n34323), .ZN(n25281) );
  CLKNHSV6 U26812 ( .I(n34435), .ZN(n34713) );
  INHSV6 U26813 ( .I(n34713), .ZN(n34440) );
  NAND2HSV2 U26814 ( .A1(n26063), .A2(n46082), .ZN(n46083) );
  NOR2HSV4 U26815 ( .A1(n25283), .A2(n25282), .ZN(n26307) );
  CLKNHSV2 U26816 ( .I(n31540), .ZN(n25282) );
  CLKNHSV2 U26817 ( .I(n31526), .ZN(n25283) );
  NAND2HSV2 U26818 ( .A1(n43492), .A2(n43491), .ZN(n26420) );
  NOR2HSV4 U26819 ( .A1(n52567), .A2(n40020), .ZN(n40121) );
  DELHS1 U26820 ( .I(n34007), .Z(n25284) );
  CLKNAND2HSV4 U26821 ( .A1(n36695), .A2(\pe3/got [29]), .ZN(n26592) );
  CLKNAND2HSV4 U26822 ( .A1(n33388), .A2(n33387), .ZN(n33392) );
  INHSV12 U26823 ( .I(n36940), .ZN(n36816) );
  CLKNAND2HSV8 U26824 ( .A1(n36816), .A2(n36955), .ZN(n25707) );
  BUFHSV6 U26825 ( .I(n59611), .Z(n37265) );
  INHSV2 U26826 ( .I(n39393), .ZN(n39677) );
  INHSV4 U26827 ( .I(n25726), .ZN(n36712) );
  NAND3HSV3 U26828 ( .A1(n25401), .A2(n36896), .A3(n36897), .ZN(n36914) );
  NOR2HSV8 U26829 ( .A1(n25286), .A2(n25285), .ZN(n39392) );
  INHSV4 U26830 ( .I(n37767), .ZN(n25285) );
  INHSV6 U26831 ( .I(n39408), .ZN(n25286) );
  NAND2HSV4 U26832 ( .A1(n39116), .A2(n48741), .ZN(n37759) );
  XNOR2HSV4 U26833 ( .A1(n33197), .A2(n25287), .ZN(n33231) );
  CLKNAND2HSV2 U26834 ( .A1(n29780), .A2(n33507), .ZN(n25287) );
  XNOR2HSV4 U26835 ( .A1(n39666), .A2(n39665), .ZN(n39668) );
  AO21HSV4 U26836 ( .A1(n30017), .A2(n30016), .B(n39240), .Z(n29651) );
  CLKNAND2HSV4 U26837 ( .A1(n45398), .A2(n45397), .ZN(n26066) );
  NAND3HSV3 U26838 ( .A1(n33667), .A2(n33666), .A3(n59955), .ZN(n33668) );
  CLKNAND2HSV2 U26839 ( .A1(n48459), .A2(n48460), .ZN(n48463) );
  CLKAND2HSV4 U26840 ( .A1(n29944), .A2(n30320), .Z(n29940) );
  CLKNAND2HSV4 U26841 ( .A1(n25947), .A2(n25949), .ZN(n48328) );
  CLKBUFHSV12 U26842 ( .I(n32158), .Z(n25288) );
  NAND2HSV2 U26843 ( .A1(n59365), .A2(n42029), .ZN(n26947) );
  MUX2NHSV2 U26844 ( .I0(n37147), .I1(n25972), .S(n25289), .ZN(n25962) );
  CLKNHSV2 U26845 ( .I(n25974), .ZN(n25289) );
  CLKNHSV2 U26846 ( .I(n37146), .ZN(n37147) );
  XNOR2HSV4 U26847 ( .A1(n37144), .A2(n37145), .ZN(n37146) );
  NOR2HSV4 U26848 ( .A1(n25290), .A2(n52829), .ZN(n42346) );
  CLKNAND2HSV2 U26849 ( .A1(n25292), .A2(n25291), .ZN(n25290) );
  CLKNHSV2 U26850 ( .I(n48331), .ZN(n25291) );
  CLKNHSV2 U26851 ( .I(n60104), .ZN(n25292) );
  XNOR2HSV4 U26852 ( .A1(n25294), .A2(n25293), .ZN(n55565) );
  XNOR2HSV4 U26853 ( .A1(n55563), .A2(n55564), .ZN(n25293) );
  CLKNAND2HSV2 U26854 ( .A1(n59931), .A2(n55319), .ZN(n25294) );
  XOR2HSV2 U26855 ( .A1(n54888), .A2(n25295), .Z(n54889) );
  XOR2HSV2 U26856 ( .A1(n54885), .A2(n25296), .Z(n25295) );
  XOR2HSV2 U26857 ( .A1(n54886), .A2(n54887), .Z(n25296) );
  INHSV4 U26858 ( .I(n52789), .ZN(n26560) );
  NAND2HSV4 U26859 ( .A1(n26560), .A2(n42605), .ZN(n26563) );
  CLKNAND2HSV4 U26860 ( .A1(n45136), .A2(n45137), .ZN(n60013) );
  CLKNAND2HSV4 U26861 ( .A1(n36690), .A2(n44333), .ZN(n36783) );
  CLKNAND2HSV4 U26862 ( .A1(n36687), .A2(n36688), .ZN(n44333) );
  INHSV4 U26863 ( .I(n32519), .ZN(n32520) );
  NAND2HSV4 U26864 ( .A1(n32520), .A2(n35808), .ZN(n32527) );
  XNOR2HSV4 U26865 ( .A1(n32342), .A2(n32343), .ZN(n32337) );
  XNOR2HSV4 U26866 ( .A1(n25297), .A2(n32779), .ZN(n32780) );
  XNOR2HSV4 U26867 ( .A1(n32778), .A2(n32777), .ZN(n25297) );
  NAND2HSV4 U26868 ( .A1(n36783), .A2(n36709), .ZN(n36732) );
  INHSV4 U26869 ( .I(n25372), .ZN(n29689) );
  NAND2HSV2 U26870 ( .A1(n25750), .A2(n36705), .ZN(n36708) );
  NAND2HSV4 U26871 ( .A1(n36748), .A2(n25976), .ZN(n36780) );
  NAND2HSV2 U26872 ( .A1(n48075), .A2(\pe3/pvq [4]), .ZN(n26589) );
  XNOR2HSV4 U26873 ( .A1(n25299), .A2(n25298), .ZN(n25996) );
  XOR2HSV2 U26874 ( .A1(n36797), .A2(n36796), .Z(n25298) );
  XNOR2HSV4 U26875 ( .A1(n25998), .A2(n25997), .ZN(n25299) );
  INHSV4 U26876 ( .I(\pe3/aot [31]), .ZN(n36999) );
  INHSV4 U26877 ( .I(n56854), .ZN(n56948) );
  NOR2HSV4 U26878 ( .A1(n48451), .A2(n42196), .ZN(n42198) );
  NOR2HSV4 U26879 ( .A1(n37533), .A2(n37532), .ZN(n37536) );
  NAND2HSV4 U26880 ( .A1(n37536), .A2(n37535), .ZN(n37537) );
  XNOR2HSV4 U26881 ( .A1(n37747), .A2(n37748), .ZN(n37750) );
  NAND3HSV3 U26882 ( .A1(n26523), .A2(n26519), .A3(n26522), .ZN(n26535) );
  MUX2NHSV4 U26883 ( .I0(n29814), .I1(n29813), .S(n25300), .ZN(n29818) );
  NAND2HSV4 U26884 ( .A1(n26736), .A2(n26735), .ZN(n25300) );
  CLKNAND2HSV4 U26885 ( .A1(n34016), .A2(n34015), .ZN(n34218) );
  CLKNAND2HSV4 U26886 ( .A1(n29812), .A2(n29811), .ZN(n29910) );
  CLKNAND2HSV8 U26887 ( .A1(n29910), .A2(n30864), .ZN(n29849) );
  NAND3HSV3 U26888 ( .A1(n29857), .A2(n25302), .A3(n25301), .ZN(n29858) );
  INHSV2 U26889 ( .I(n29854), .ZN(n25301) );
  NAND2HSV4 U26890 ( .A1(n29855), .A2(n39246), .ZN(n25302) );
  XOR2HSV4 U26891 ( .A1(n53096), .A2(n26865), .Z(n25841) );
  XOR2HSV4 U26892 ( .A1(n29640), .A2(n25841), .Z(n53100) );
  INHSV4 U26893 ( .I(n45933), .ZN(n45630) );
  NAND2HSV4 U26894 ( .A1(n45925), .A2(n46108), .ZN(n45933) );
  INHSV4 U26895 ( .I(n30678), .ZN(n30674) );
  NOR2HSV8 U26896 ( .A1(n30674), .A2(n39241), .ZN(n30751) );
  CLKNAND2HSV2 U26897 ( .A1(n31881), .A2(n31880), .ZN(n31878) );
  INHSV2 U26898 ( .I(n31878), .ZN(n31882) );
  XOR3HSV2 U26899 ( .A1(n25303), .A2(n50803), .A3(n50804), .Z(\pe3/poht [19])
         );
  XNOR2HSV4 U26900 ( .A1(n50801), .A2(n50800), .ZN(n25303) );
  XNOR2HSV4 U26901 ( .A1(n56487), .A2(n56488), .ZN(n25320) );
  INHSV2 U26902 ( .I(n31134), .ZN(n25304) );
  CLKNAND2HSV2 U26903 ( .A1(n25304), .A2(n31133), .ZN(n31136) );
  BUFHSV6 U26904 ( .I(n46545), .Z(n48480) );
  CLKNAND2HSV2 U26905 ( .A1(n59573), .A2(n52767), .ZN(n39381) );
  NAND2HSV2 U26906 ( .A1(n56860), .A2(\pe3/got [17]), .ZN(n56488) );
  NAND2HSV2 U26907 ( .A1(n29444), .A2(n29443), .ZN(n29445) );
  INHSV4 U26908 ( .I(\pe4/got [30]), .ZN(n33098) );
  CLKNHSV6 U26909 ( .I(n45943), .ZN(n50716) );
  INHSV4 U26910 ( .I(n33178), .ZN(n26644) );
  CLKAND2HSV2 U26911 ( .A1(n32648), .A2(n32644), .Z(n32535) );
  CLKNHSV0 U26912 ( .I(n30496), .ZN(n39744) );
  CLKNAND2HSV4 U26913 ( .A1(n52818), .A2(n30867), .ZN(n30868) );
  NOR2HSV8 U26914 ( .A1(n30869), .A2(n30868), .ZN(n31100) );
  XNOR2HSV4 U26915 ( .A1(n25305), .A2(n31084), .ZN(n31094) );
  XOR2HSV2 U26916 ( .A1(n31083), .A2(n31082), .Z(n25305) );
  CLKXOR2HSV4 U26917 ( .A1(n56255), .A2(n56254), .Z(n56256) );
  CLKNAND2HSV2 U26918 ( .A1(n57325), .A2(n59599), .ZN(n33497) );
  INHSV4 U26919 ( .I(n33063), .ZN(n48010) );
  XNOR2HSV4 U26920 ( .A1(n48608), .A2(n48609), .ZN(n48610) );
  CLKNAND2HSV3 U26921 ( .A1(n45938), .A2(n45779), .ZN(n45939) );
  CLKNAND2HSV3 U26922 ( .A1(n31406), .A2(n31407), .ZN(n26337) );
  NOR2HSV4 U26923 ( .A1(n39252), .A2(n40130), .ZN(n39253) );
  CLKNAND2HSV1 U26924 ( .A1(n34096), .A2(n34218), .ZN(n34098) );
  INHSV3 U26925 ( .I(n39003), .ZN(n26264) );
  INHSV4 U26926 ( .I(n25306), .ZN(n40579) );
  INHSV4 U26927 ( .I(n40479), .ZN(n25306) );
  NAND2HSV2 U26928 ( .A1(n59609), .A2(n37298), .ZN(n36794) );
  OAI21HSV4 U26929 ( .A1(n36732), .A2(n25995), .B(n36717), .ZN(n36735) );
  CLKNAND2HSV4 U26930 ( .A1(n26621), .A2(n26623), .ZN(n26620) );
  INHSV4 U26931 ( .I(n31425), .ZN(n31368) );
  NAND2HSV4 U26932 ( .A1(n52821), .A2(n47773), .ZN(n34316) );
  INHSV4 U26933 ( .I(n34316), .ZN(n34321) );
  CLKNAND2HSV2 U26934 ( .A1(n25651), .A2(n46558), .ZN(n45934) );
  CLKNAND2HSV2 U26935 ( .A1(n34285), .A2(n59600), .ZN(n33436) );
  NAND2HSV4 U26936 ( .A1(n25307), .A2(n30024), .ZN(n30026) );
  INHSV2 U26937 ( .I(n26821), .ZN(n52698) );
  INHSV2 U26938 ( .I(n52698), .ZN(n33158) );
  INHSV4 U26939 ( .I(\pe1/aot [27]), .ZN(n41442) );
  NAND2HSV4 U26940 ( .A1(n53530), .A2(n53411), .ZN(n40349) );
  NAND2HSV2 U26941 ( .A1(n25418), .A2(n36675), .ZN(n36676) );
  XNOR2HSV4 U26942 ( .A1(n25309), .A2(n25308), .ZN(n25938) );
  CLKNAND2HSV2 U26943 ( .A1(n32469), .A2(n32410), .ZN(n25308) );
  XNOR2HSV4 U26944 ( .A1(n32409), .A2(n32408), .ZN(n25309) );
  CLKNAND2HSV4 U26945 ( .A1(n25843), .A2(n26781), .ZN(n25386) );
  NAND2HSV4 U26946 ( .A1(n25387), .A2(n25386), .ZN(n26779) );
  OAI21HSV4 U26947 ( .A1(n40558), .A2(n40443), .B(n40466), .ZN(n40340) );
  OAI21HSV4 U26948 ( .A1(n45758), .A2(n45759), .B(n45757), .ZN(n45771) );
  INHSV2 U26949 ( .I(n32514), .ZN(n25937) );
  CLKNAND2HSV2 U26950 ( .A1(n25310), .A2(n54161), .ZN(n55159) );
  CLKNHSV2 U26951 ( .I(n55158), .ZN(n25310) );
  NAND2HSV4 U26952 ( .A1(n45609), .A2(n25311), .ZN(n45623) );
  NAND3HSV2 U26953 ( .A1(n45604), .A2(n45606), .A3(n45605), .ZN(n25311) );
  CLKNAND2HSV2 U26954 ( .A1(n25313), .A2(n25312), .ZN(n29949) );
  CLKNHSV2 U26955 ( .I(n29947), .ZN(n25312) );
  CLKNHSV2 U26956 ( .I(n29946), .ZN(n25313) );
  CLKNAND2HSV2 U26957 ( .A1(n29018), .A2(n34212), .ZN(n34206) );
  NAND2HSV4 U26958 ( .A1(n25314), .A2(n38527), .ZN(n38739) );
  NAND2HSV2 U26959 ( .A1(n38526), .A2(n38525), .ZN(n25314) );
  NAND2HSV4 U26960 ( .A1(n25315), .A2(n32322), .ZN(n32160) );
  NAND2HSV2 U26961 ( .A1(n32156), .A2(n25316), .ZN(n25315) );
  NOR2HSV0 U26962 ( .A1(n32325), .A2(n25317), .ZN(n25316) );
  INHSV2 U26963 ( .I(n35908), .ZN(n25317) );
  INHSV2 U26964 ( .I(\pe5/phq [2]), .ZN(n26733) );
  INHSV4 U26965 ( .I(n46310), .ZN(n48481) );
  XNOR2HSV4 U26966 ( .A1(n32428), .A2(n32429), .ZN(n32433) );
  INHSV4 U26967 ( .I(n32310), .ZN(n32311) );
  INHSV4 U26968 ( .I(n29805), .ZN(n29804) );
  XNOR2HSV4 U26969 ( .A1(n56774), .A2(n25318), .ZN(n56777) );
  XOR2HSV2 U26970 ( .A1(n25475), .A2(n56772), .Z(n25318) );
  NAND2HSV4 U26971 ( .A1(n47979), .A2(n38015), .ZN(n38192) );
  XNOR2HSV4 U26972 ( .A1(n25319), .A2(n31745), .ZN(n26655) );
  XOR2HSV2 U26973 ( .A1(n31741), .A2(n31742), .Z(n25319) );
  INHSV4 U26974 ( .I(n31440), .ZN(n31434) );
  INHSV2 U26975 ( .I(n31434), .ZN(n44426) );
  XOR3HSV2 U26976 ( .A1(n25320), .A2(n56491), .A3(n56492), .Z(\pe3/poht [13])
         );
  INHSV4 U26977 ( .I(n39113), .ZN(n26884) );
  NAND3HSV4 U26978 ( .A1(n44148), .A2(n26884), .A3(n36654), .ZN(n39109) );
  OAI21HSV2 U26979 ( .A1(n27448), .A2(n27449), .B(n27450), .ZN(n27451) );
  NAND2HSV2 U26980 ( .A1(n27452), .A2(n27451), .ZN(n27453) );
  CLKNAND2HSV2 U26981 ( .A1(n44668), .A2(n26964), .ZN(n26262) );
  INHSV6 U26982 ( .I(n59883), .ZN(n47057) );
  NOR2HSV4 U26983 ( .A1(n47057), .A2(n30210), .ZN(n39982) );
  CLKNAND2HSV2 U26984 ( .A1(n45943), .A2(n46072), .ZN(n25321) );
  CLKNHSV2 U26985 ( .I(n46075), .ZN(n25324) );
  CLKNAND2HSV2 U26986 ( .A1(n45944), .A2(n45946), .ZN(n46075) );
  CLKNHSV2 U26987 ( .I(n46073), .ZN(n25325) );
  CLKNAND2HSV4 U26988 ( .A1(n45610), .A2(n44685), .ZN(n44689) );
  INHSV4 U26989 ( .I(n29802), .ZN(n26358) );
  NAND2HSV4 U26990 ( .A1(n59508), .A2(n59356), .ZN(n56883) );
  CLKNAND2HSV3 U26991 ( .A1(n36706), .A2(n25733), .ZN(n36707) );
  CLKNAND2HSV3 U26992 ( .A1(n36736), .A2(n36735), .ZN(n25359) );
  BUFHSV2 U26993 ( .I(n33795), .Z(n25326) );
  NAND2HSV4 U26994 ( .A1(n44476), .A2(n49665), .ZN(n31959) );
  NAND2HSV4 U26995 ( .A1(n42084), .A2(n41243), .ZN(n29158) );
  XOR2HSV4 U26996 ( .A1(n30039), .A2(n30038), .Z(n30043) );
  NAND2HSV4 U26997 ( .A1(n26015), .A2(n43898), .ZN(n37525) );
  CLKNAND2HSV4 U26998 ( .A1(n43595), .A2(n43594), .ZN(n43614) );
  NAND2HSV4 U26999 ( .A1(n25328), .A2(n25327), .ZN(n32039) );
  INHSV4 U27000 ( .I(n32038), .ZN(n25327) );
  INHSV4 U27001 ( .I(n32037), .ZN(n25328) );
  INHSV4 U27002 ( .I(n36984), .ZN(n36975) );
  XNOR2HSV4 U27003 ( .A1(n35268), .A2(n35267), .ZN(n35271) );
  NOR2HSV4 U27004 ( .A1(n29774), .A2(n47861), .ZN(n47863) );
  XNOR2HSV4 U27005 ( .A1(n29816), .A2(n25329), .ZN(n29817) );
  NOR2HSV4 U27006 ( .A1(n29959), .A2(n39163), .ZN(n25329) );
  INHSV2 U27007 ( .I(n38623), .ZN(n52810) );
  NAND2HSV2 U27008 ( .A1(n26892), .A2(n26891), .ZN(n38623) );
  CLKNAND2HSV4 U27009 ( .A1(n32328), .A2(n32327), .ZN(n32342) );
  INAND2HSV4 U27010 ( .A1(n32166), .B1(n32833), .ZN(n32142) );
  CLKNAND2HSV2 U27011 ( .A1(n37034), .A2(n37035), .ZN(n37032) );
  NAND2HSV2 U27012 ( .A1(n32650), .A2(n32649), .ZN(n32654) );
  OA21HSV4 U27013 ( .A1(n36899), .A2(\pe3/got [32]), .B(n29713), .Z(n36897) );
  CLKNAND2HSV4 U27014 ( .A1(n25441), .A2(n25440), .ZN(n25980) );
  XNOR2HSV4 U27015 ( .A1(n30002), .A2(\pe5/phq [7]), .ZN(n30003) );
  XOR2HSV4 U27016 ( .A1(n40384), .A2(n40383), .Z(n40390) );
  NAND2HSV4 U27017 ( .A1(n48029), .A2(\pe5/pvq [6]), .ZN(n30039) );
  CLKNAND2HSV2 U27018 ( .A1(n29795), .A2(n29794), .ZN(n29798) );
  XNOR2HSV4 U27019 ( .A1(n37244), .A2(n25330), .ZN(n37258) );
  OAI21HSV4 U27020 ( .A1(n37512), .A2(n37513), .B(n37243), .ZN(n25330) );
  NAND2HSV2 U27021 ( .A1(n41705), .A2(n41704), .ZN(n41846) );
  NAND2HSV2 U27022 ( .A1(n42794), .A2(n25331), .ZN(n42795) );
  CLKNHSV2 U27023 ( .I(n42793), .ZN(n25331) );
  NOR2HSV4 U27024 ( .A1(n42915), .A2(n29705), .ZN(n42793) );
  OAI21HSV4 U27025 ( .A1(n25574), .A2(n25575), .B(n25573), .ZN(n44656) );
  INHSV3 U27026 ( .I(n32522), .ZN(n32235) );
  AOI31HSV2 U27027 ( .A1(n38618), .A2(n38617), .A3(n38611), .B(n52411), .ZN(
        n38466) );
  NAND3HSV4 U27028 ( .A1(n38465), .A2(n38606), .A3(n38519), .ZN(n38617) );
  CLKNAND2HSV2 U27029 ( .A1(n48481), .A2(n42673), .ZN(n55933) );
  BUFHSV8 U27030 ( .I(n59607), .Z(n36940) );
  INHSV2 U27031 ( .I(n59607), .ZN(n25332) );
  NAND3HSV4 U27032 ( .A1(n25332), .A2(n59347), .A3(\pe3/bq[30] ), .ZN(n36677)
         );
  NAND2HSV4 U27033 ( .A1(n40340), .A2(n40341), .ZN(n25431) );
  NAND2HSV4 U27034 ( .A1(n31758), .A2(n26255), .ZN(n26254) );
  NAND2HSV4 U27035 ( .A1(n29999), .A2(n30037), .ZN(n29893) );
  NAND2HSV4 U27036 ( .A1(n31958), .A2(n31902), .ZN(n31813) );
  NOR2HSV4 U27037 ( .A1(n51112), .A2(n41824), .ZN(n40333) );
  CLKNAND2HSV4 U27038 ( .A1(n59376), .A2(n40332), .ZN(n51113) );
  OAI21HSV4 U27039 ( .A1(n51113), .A2(\pe1/got [32]), .B(n40333), .ZN(n40334)
         );
  XNOR2HSV4 U27040 ( .A1(n25334), .A2(n25333), .ZN(n26401) );
  CLKNAND2HSV2 U27041 ( .A1(n39824), .A2(n30254), .ZN(n25333) );
  XNOR2HSV4 U27042 ( .A1(n30296), .A2(n29716), .ZN(n25334) );
  INHSV6 U27043 ( .I(n54155), .ZN(n55608) );
  CLKNAND2HSV2 U27044 ( .A1(n55608), .A2(\pe1/got [23]), .ZN(n54449) );
  INHSV4 U27045 ( .I(n39797), .ZN(n30146) );
  INAND2HSV2 U27046 ( .A1(n53095), .B1(n38603), .ZN(n29640) );
  CLKNAND2HSV4 U27047 ( .A1(n32036), .A2(n44378), .ZN(n32037) );
  CLKNAND2HSV4 U27048 ( .A1(n34831), .A2(n34829), .ZN(n35143) );
  CLKNAND2HSV4 U27049 ( .A1(n35143), .A2(n35011), .ZN(n34827) );
  CLKNAND2HSV2 U27050 ( .A1(n27780), .A2(n27781), .ZN(n27782) );
  CLKNAND2HSV2 U27051 ( .A1(n25337), .A2(n25336), .ZN(n25335) );
  CLKNHSV2 U27052 ( .I(n27777), .ZN(n25336) );
  CLKNHSV2 U27053 ( .I(n27778), .ZN(n25337) );
  CLKNAND2HSV2 U27054 ( .A1(n28796), .A2(n28797), .ZN(n28798) );
  CLKNAND2HSV2 U27055 ( .A1(n25340), .A2(n25339), .ZN(n25338) );
  CLKNHSV2 U27056 ( .I(n28793), .ZN(n25339) );
  CLKNHSV2 U27057 ( .I(n28794), .ZN(n25340) );
  INHSV4 U27058 ( .I(n32309), .ZN(n32312) );
  IOA21HSV4 U27059 ( .A1(\pe5/pvq [2]), .A2(\pe5/ctrq ), .B(\pe5/phq [2]), 
        .ZN(n26735) );
  INHSV4 U27060 ( .I(n32506), .ZN(n59363) );
  INAND2HSV4 U27061 ( .A1(n49315), .B1(n59363), .ZN(n32135) );
  XNOR2HSV4 U27062 ( .A1(n29875), .A2(n25341), .ZN(n29878) );
  OAI22HSV4 U27063 ( .A1(n29873), .A2(n30223), .B1(n29874), .B2(\pe5/phq [3]), 
        .ZN(n25341) );
  CLKAND2HSV2 U27064 ( .A1(n42706), .A2(n42936), .Z(n42687) );
  CLKNAND2HSV4 U27065 ( .A1(n32442), .A2(n32441), .ZN(n32557) );
  CLKNHSV6 U27066 ( .I(n32557), .ZN(n32559) );
  NOR2HSV4 U27067 ( .A1(n29774), .A2(n58294), .ZN(n58296) );
  XNOR2HSV4 U27068 ( .A1(n44947), .A2(n44948), .ZN(n44951) );
  INHSV4 U27069 ( .I(n26734), .ZN(n29800) );
  NOR2HSV4 U27070 ( .A1(n29800), .A2(n29799), .ZN(n29802) );
  CLKNAND2HSV4 U27071 ( .A1(n29999), .A2(n30029), .ZN(n29830) );
  INHSV4 U27072 ( .I(n29830), .ZN(n29832) );
  INHSV4 U27073 ( .I(n56260), .ZN(n56059) );
  CLKNAND2HSV4 U27074 ( .A1(n25698), .A2(n45144), .ZN(n59789) );
  BUFHSV6 U27075 ( .I(n59789), .Z(n52414) );
  NAND2HSV2 U27076 ( .A1(n48481), .A2(n56558), .ZN(n53276) );
  XNOR2HSV2 U27077 ( .A1(n53276), .A2(n53275), .ZN(n53277) );
  NAND3HSV4 U27078 ( .A1(n56418), .A2(n49404), .A3(n56417), .ZN(n29247) );
  OAI21HSV2 U27079 ( .A1(n29246), .A2(n29247), .B(n29248), .ZN(n29249) );
  INHSV4 U27080 ( .I(n26610), .ZN(n25441) );
  OAI21HSV4 U27081 ( .A1(n25342), .A2(n35157), .B(n35306), .ZN(n35019) );
  NOR2HSV4 U27082 ( .A1(n40411), .A2(n40445), .ZN(n40323) );
  XNOR2HSV1 U27083 ( .A1(n40323), .A2(n26170), .ZN(n26172) );
  INHSV2 U27084 ( .I(n25343), .ZN(n35446) );
  CLKNAND2HSV2 U27085 ( .A1(n35284), .A2(n35011), .ZN(n25343) );
  DELHS1 U27086 ( .I(n29848), .Z(n25344) );
  NAND2HSV4 U27087 ( .A1(n36789), .A2(\pe3/aot [29]), .ZN(n36790) );
  INHSV4 U27088 ( .I(n42616), .ZN(n26564) );
  NAND2HSV2 U27089 ( .A1(n50318), .A2(n57646), .ZN(n50107) );
  NAND3HSV3 U27090 ( .A1(n40308), .A2(n40307), .A3(n51411), .ZN(n40313) );
  NAND2HSV4 U27091 ( .A1(n40313), .A2(n40312), .ZN(n40316) );
  CLKNAND2HSV2 U27092 ( .A1(n38749), .A2(n38625), .ZN(n52812) );
  CLKXOR2HSV2 U27093 ( .A1(n47384), .A2(n25887), .Z(n47386) );
  NOR2HSV4 U27094 ( .A1(n58212), .A2(n34851), .ZN(n57322) );
  XNOR2HSV4 U27095 ( .A1(n26864), .A2(n26859), .ZN(\pe5/poht [1]) );
  CLKNAND2HSV4 U27096 ( .A1(n37098), .A2(n37097), .ZN(n37165) );
  INHSV4 U27097 ( .I(\pe1/aot [32]), .ZN(n40443) );
  NAND3HSV4 U27098 ( .A1(n33384), .A2(n33383), .A3(n35604), .ZN(n33388) );
  NAND2HSV4 U27099 ( .A1(n33337), .A2(n33336), .ZN(n33404) );
  CLKNAND2HSV2 U27100 ( .A1(n33404), .A2(n33588), .ZN(n33406) );
  CLKNAND2HSV2 U27101 ( .A1(n52840), .A2(n52052), .ZN(n27963) );
  NAND2HSV2 U27102 ( .A1(n27963), .A2(n27962), .ZN(n27964) );
  NAND2HSV4 U27103 ( .A1(n31625), .A2(n35797), .ZN(n31684) );
  NOR2HSV8 U27104 ( .A1(n40736), .A2(n40556), .ZN(n26174) );
  XNOR2HSV4 U27105 ( .A1(n31955), .A2(n31954), .ZN(n31956) );
  NAND2HSV4 U27106 ( .A1(n32414), .A2(n25346), .ZN(n32558) );
  NAND2HSV2 U27107 ( .A1(n32453), .A2(n32412), .ZN(n25346) );
  INHSV4 U27108 ( .I(n48466), .ZN(n26005) );
  NAND2HSV4 U27109 ( .A1(n25412), .A2(n48463), .ZN(n48466) );
  NAND2HSV4 U27110 ( .A1(n26879), .A2(n26880), .ZN(n26882) );
  XOR2HSV4 U27111 ( .A1(n34315), .A2(n34314), .Z(n34434) );
  CLKNAND2HSV4 U27112 ( .A1(n38601), .A2(n38607), .ZN(n38618) );
  CLKXOR2HSV4 U27113 ( .A1(n41586), .A2(n41587), .Z(n47957) );
  CLKNAND2HSV2 U27114 ( .A1(n33857), .A2(n25347), .ZN(n33780) );
  CLKNHSV2 U27115 ( .I(n25348), .ZN(n25347) );
  CLKNAND2HSV2 U27116 ( .A1(n34949), .A2(n33778), .ZN(n25348) );
  MUX2NHSV2 U27117 ( .I0(n38598), .I1(n38597), .S(n25349), .ZN(n38599) );
  XNOR2HSV4 U27118 ( .A1(n38596), .A2(n38595), .ZN(n25349) );
  NOR2HSV4 U27119 ( .A1(n42617), .A2(n26564), .ZN(n52789) );
  NAND2HSV4 U27120 ( .A1(n25477), .A2(n25816), .ZN(n42784) );
  XNOR2HSV4 U27121 ( .A1(n33563), .A2(n33562), .ZN(n33568) );
  CLKNAND2HSV2 U27122 ( .A1(n38606), .A2(n25351), .ZN(n25350) );
  CLKNHSV2 U27123 ( .I(n38605), .ZN(n25351) );
  CLKNAND2HSV2 U27124 ( .A1(n37642), .A2(n30028), .ZN(n37643) );
  NAND3HSV4 U27125 ( .A1(n31244), .A2(n37540), .A3(n31243), .ZN(n37642) );
  NAND2HSV2 U27126 ( .A1(n34206), .A2(n34205), .ZN(n34214) );
  AOI22HSV4 U27127 ( .A1(n38351), .A2(n38350), .B1(n38352), .B2(n52776), .ZN(
        n38367) );
  CLKNAND2HSV2 U27128 ( .A1(n38267), .A2(n25352), .ZN(n52776) );
  CLKNHSV2 U27129 ( .I(n38452), .ZN(n25352) );
  NAND3HSV3 U27130 ( .A1(n46071), .A2(n46076), .A3(n46072), .ZN(n46080) );
  OAI21HSV4 U27131 ( .A1(n36511), .A2(n60005), .B(n36510), .ZN(n36517) );
  INHSV2 U27132 ( .I(n46089), .ZN(n46095) );
  XOR2HSV2 U27133 ( .A1(n36794), .A2(n25353), .Z(n36798) );
  CLKNAND2HSV2 U27134 ( .A1(n37280), .A2(n25354), .ZN(n25353) );
  CLKNHSV2 U27135 ( .I(n36999), .ZN(n25354) );
  NOR2HSV4 U27136 ( .A1(n32646), .A2(n32530), .ZN(n32534) );
  NAND2HSV2 U27137 ( .A1(n32435), .A2(n32652), .ZN(n32437) );
  NAND3HSV4 U27138 ( .A1(n25826), .A2(n41727), .A3(n41719), .ZN(n41914) );
  CLKXOR2HSV4 U27139 ( .A1(n36818), .A2(n36817), .Z(n36822) );
  XNOR2HSV4 U27140 ( .A1(n36625), .A2(n36624), .ZN(n36628) );
  NAND2HSV4 U27141 ( .A1(n46117), .A2(n25355), .ZN(n46308) );
  CLKNAND2HSV4 U27142 ( .A1(n26072), .A2(n46560), .ZN(n25355) );
  IAO21HSV4 U27143 ( .A1(n32423), .A2(n32421), .B(n32239), .ZN(n29652) );
  CLKNHSV6 U27144 ( .I(n39112), .ZN(n26883) );
  NAND2HSV4 U27145 ( .A1(n32026), .A2(n31899), .ZN(n31966) );
  AOI21HSV4 U27146 ( .A1(n34582), .A2(n29700), .B(n34581), .ZN(n34586) );
  NAND2HSV4 U27147 ( .A1(n34586), .A2(n34585), .ZN(n34969) );
  CLKNAND2HSV2 U27148 ( .A1(n60051), .A2(n53092), .ZN(n44820) );
  CLKNHSV2 U27149 ( .I(n31522), .ZN(n31402) );
  XNOR2HSV4 U27150 ( .A1(n31397), .A2(n31396), .ZN(n31522) );
  CLKNAND2HSV4 U27151 ( .A1(n42042), .A2(n25394), .ZN(n42052) );
  CLKNAND2HSV2 U27152 ( .A1(n59595), .A2(n31667), .ZN(n31668) );
  NAND2HSV0 U27153 ( .A1(n28793), .A2(n28794), .ZN(n28795) );
  NAND2HSV0 U27154 ( .A1(n52910), .A2(n51939), .ZN(n28794) );
  NAND2HSV0 U27155 ( .A1(n27777), .A2(n27778), .ZN(n27779) );
  NAND2HSV0 U27156 ( .A1(n52910), .A2(\pe2/got [12]), .ZN(n27778) );
  INHSV4 U27157 ( .I(n45926), .ZN(n25651) );
  NOR2HSV2 U27158 ( .A1(n31629), .A2(n31681), .ZN(n31630) );
  NAND2HSV4 U27159 ( .A1(n42030), .A2(n42031), .ZN(n42036) );
  CLKNAND2HSV4 U27160 ( .A1(n42036), .A2(n42035), .ZN(n26622) );
  INHSV2 U27161 ( .I(n41908), .ZN(n42206) );
  INHSV4 U27162 ( .I(n42206), .ZN(n42085) );
  NOR2HSV2 U27163 ( .A1(n31497), .A2(n31441), .ZN(n31327) );
  INHSV2 U27164 ( .I(n31327), .ZN(n31328) );
  NAND2HSV4 U27165 ( .A1(n33415), .A2(n33103), .ZN(n33946) );
  XOR2HSV4 U27166 ( .A1(n38440), .A2(n38460), .Z(n26084) );
  NAND2HSV4 U27167 ( .A1(n25356), .A2(n38359), .ZN(n52778) );
  INHSV2 U27168 ( .I(n38371), .ZN(n25356) );
  NAND2HSV2 U27169 ( .A1(\pe4/aot [32]), .A2(\pe4/bq[32] ), .ZN(n26191) );
  XOR3HSV2 U27170 ( .A1(n25357), .A2(n56051), .A3(n56052), .Z(n56053) );
  CLKNHSV2 U27171 ( .I(n56050), .ZN(n25357) );
  CLKNAND2HSV4 U27172 ( .A1(n48464), .A2(n48465), .ZN(n26007) );
  INHSV4 U27173 ( .I(n26007), .ZN(n26006) );
  INHSV2 U27174 ( .I(n37851), .ZN(n37852) );
  CLKNHSV2 U27175 ( .I(n26149), .ZN(n25358) );
  NAND2HSV2 U27176 ( .A1(n44660), .A2(n44527), .ZN(n26530) );
  CLKNAND2HSV4 U27177 ( .A1(n34844), .A2(n34843), .ZN(n34845) );
  NOR2HSV4 U27178 ( .A1(n37863), .A2(n37864), .ZN(n38007) );
  NAND2HSV2 U27179 ( .A1(n36861), .A2(n36840), .ZN(n36842) );
  CLKNAND2HSV2 U27180 ( .A1(n31111), .A2(n39718), .ZN(n31112) );
  INHSV4 U27181 ( .I(n31112), .ZN(n31115) );
  NAND2HSV4 U27182 ( .A1(n31143), .A2(n31142), .ZN(n26493) );
  NAND2HSV2 U27183 ( .A1(n31141), .A2(n31091), .ZN(n31143) );
  CLKNAND2HSV4 U27184 ( .A1(n38373), .A2(n26559), .ZN(n52286) );
  CLKNAND2HSV2 U27185 ( .A1(n52286), .A2(n38777), .ZN(n38262) );
  CLKNAND2HSV4 U27186 ( .A1(n25360), .A2(n25359), .ZN(n25719) );
  NAND2HSV4 U27187 ( .A1(n36726), .A2(n36733), .ZN(n25360) );
  INHSV8 U27188 ( .I(n37020), .ZN(n36748) );
  CLKNAND2HSV8 U27189 ( .A1(n36748), .A2(n45612), .ZN(n25750) );
  INHSV2 U27190 ( .I(n39117), .ZN(n37548) );
  AND2HSV4 U27191 ( .A1(n37642), .A2(n39382), .Z(n29669) );
  NAND2HSV4 U27192 ( .A1(n29669), .A2(n37548), .ZN(n39227) );
  INHSV4 U27193 ( .I(n31277), .ZN(n31273) );
  CLKNAND2HSV2 U27194 ( .A1(n55608), .A2(n59374), .ZN(n54156) );
  NAND2HSV4 U27195 ( .A1(n25361), .A2(n36268), .ZN(n36285) );
  CLKNAND2HSV4 U27196 ( .A1(n36267), .A2(n36266), .ZN(n25361) );
  MUX2NHSV2 U27197 ( .I0(n31342), .I1(n31353), .S(n31352), .ZN(n31347) );
  CLKNAND2HSV2 U27198 ( .A1(n31374), .A2(n31373), .ZN(n31375) );
  NAND2HSV4 U27199 ( .A1(n57510), .A2(n48074), .ZN(n33210) );
  XOR2HSV4 U27200 ( .A1(n33209), .A2(n33210), .Z(n26031) );
  INHSV2 U27201 ( .I(n36787), .ZN(n25362) );
  CLKNAND2HSV2 U27202 ( .A1(n25362), .A2(n43464), .ZN(n25383) );
  NAND2HSV4 U27203 ( .A1(n36433), .A2(\pe2/bq[27] ), .ZN(n36436) );
  CLKNAND2HSV2 U27204 ( .A1(n37109), .A2(n37186), .ZN(n36792) );
  CLKXOR2HSV4 U27205 ( .A1(n36543), .A2(n36542), .Z(n36545) );
  CLKNAND2HSV4 U27206 ( .A1(n36816), .A2(n56057), .ZN(n25997) );
  CLKNAND2HSV4 U27207 ( .A1(n36745), .A2(n36725), .ZN(n37274) );
  INHSV4 U27208 ( .I(n26622), .ZN(n26621) );
  CLKAND2HSV4 U27209 ( .A1(n47947), .A2(n39417), .Z(n39423) );
  CLKNAND2HSV2 U27210 ( .A1(n37235), .A2(n37234), .ZN(n37244) );
  NAND3HSV2 U27211 ( .A1(n40146), .A2(n25364), .A3(n25363), .ZN(n40147) );
  INHSV4 U27212 ( .I(n40144), .ZN(n25363) );
  NAND3HSV2 U27213 ( .A1(n25393), .A2(n40145), .A3(n25392), .ZN(n25364) );
  NAND2HSV4 U27214 ( .A1(n39554), .A2(n39866), .ZN(n39565) );
  NAND2HSV4 U27215 ( .A1(n38041), .A2(n52415), .ZN(n37914) );
  CLKNHSV2 U27216 ( .I(n44644), .ZN(n44645) );
  XNOR2HSV4 U27217 ( .A1(n26058), .A2(n44642), .ZN(n44644) );
  INHSV2 U27218 ( .I(n33437), .ZN(n59501) );
  INHSV4 U27219 ( .I(n26466), .ZN(n43473) );
  MOAI22HSV4 U27220 ( .A1(n36643), .A2(n36561), .B1(n36562), .B2(n36645), .ZN(
        n36524) );
  NAND2HSV2 U27221 ( .A1(n36647), .A2(n36642), .ZN(n36525) );
  NAND2HSV4 U27222 ( .A1(n36525), .A2(n36524), .ZN(n36573) );
  NOR2HSV4 U27223 ( .A1(n31474), .A2(n31473), .ZN(n31301) );
  NAND2HSV4 U27224 ( .A1(n31476), .A2(n31301), .ZN(n31319) );
  CLKNAND2HSV2 U27225 ( .A1(n26683), .A2(n44329), .ZN(n39385) );
  NAND2HSV4 U27226 ( .A1(n39385), .A2(n26650), .ZN(n39869) );
  XNOR2HSV4 U27227 ( .A1(n33293), .A2(n25365), .ZN(n60082) );
  XOR2HSV2 U27228 ( .A1(n29740), .A2(n33292), .Z(n25365) );
  INHSV2 U27229 ( .I(n25366), .ZN(n25829) );
  CLKNAND2HSV2 U27230 ( .A1(n40159), .A2(n40158), .ZN(n25366) );
  XNOR2HSV4 U27231 ( .A1(n40127), .A2(n40126), .ZN(n40129) );
  CLKNAND2HSV2 U27232 ( .A1(n40928), .A2(n25367), .ZN(n47983) );
  CLKNHSV2 U27233 ( .I(n48320), .ZN(n25367) );
  XNOR2HSV4 U27234 ( .A1(n33310), .A2(n33309), .ZN(n25955) );
  NOR2HSV3 U27235 ( .A1(n42914), .A2(n42913), .ZN(n43018) );
  NAND2HSV4 U27236 ( .A1(n31266), .A2(n31267), .ZN(n31271) );
  CLKBUFHSV4 U27237 ( .I(n53188), .Z(n51229) );
  INHSV6 U27238 ( .I(n43021), .ZN(n43912) );
  INHSV8 U27239 ( .I(n36630), .ZN(n36631) );
  INHSV6 U27240 ( .I(n37991), .ZN(n38036) );
  CLKNAND2HSV2 U27241 ( .A1(n41239), .A2(n40972), .ZN(n41049) );
  CLKNAND2HSV2 U27242 ( .A1(n47962), .A2(n34193), .ZN(n34190) );
  OAI21HSV4 U27243 ( .A1(n34231), .A2(n34233), .B(n34345), .ZN(n34193) );
  NAND3HSV3 U27244 ( .A1(n25370), .A2(n31336), .A3(n25368), .ZN(n31337) );
  INAND2HSV4 U27245 ( .A1(n31335), .B1(n25369), .ZN(n25368) );
  CLKNHSV0 U27246 ( .I(\pe6/aot [30]), .ZN(n25369) );
  NAND3HSV4 U27247 ( .A1(n31418), .A2(n31367), .A3(n31335), .ZN(n25370) );
  MUX2NHSV2 U27248 ( .I0(n31434), .I1(n31371), .S(n31372), .ZN(n31376) );
  NOR2HSV4 U27249 ( .A1(n34344), .A2(n34345), .ZN(n34348) );
  XOR3HSV2 U27250 ( .A1(\pe6/phq [7]), .A2(n31415), .A3(n31416), .Z(n31423) );
  CLKNAND2HSV8 U27251 ( .A1(n41847), .A2(n40407), .ZN(n41323) );
  INHSV4 U27252 ( .I(n41323), .ZN(n41321) );
  CLKNAND2HSV4 U27253 ( .A1(n60106), .A2(n41225), .ZN(n41227) );
  CLKNAND2HSV8 U27254 ( .A1(n41227), .A2(n41226), .ZN(n41412) );
  XNOR2HSV4 U27255 ( .A1(n30502), .A2(n25371), .ZN(n30588) );
  CLKNAND2HSV2 U27256 ( .A1(n30884), .A2(n30779), .ZN(n25371) );
  CLKNAND2HSV2 U27257 ( .A1(n55608), .A2(n59996), .ZN(n55037) );
  INHSV4 U27258 ( .I(n31275), .ZN(n31276) );
  CLKNHSV6 U27259 ( .I(n37222), .ZN(n37151) );
  NAND2HSV4 U27260 ( .A1(n51115), .A2(n39382), .ZN(n25372) );
  NAND2HSV4 U27261 ( .A1(n39672), .A2(n25432), .ZN(n45489) );
  NAND2HSV4 U27262 ( .A1(n35370), .A2(n33215), .ZN(n33120) );
  XNOR2HSV4 U27263 ( .A1(n31951), .A2(n31950), .ZN(n31953) );
  XNOR2HSV4 U27264 ( .A1(n31419), .A2(n31420), .ZN(n31421) );
  INHSV2 U27265 ( .I(n31755), .ZN(n26659) );
  NAND2HSV0 U27266 ( .A1(n25373), .A2(n41582), .ZN(n41584) );
  NOR2HSV2 U27267 ( .A1(n41583), .A2(n25374), .ZN(n25373) );
  NAND2HSV4 U27268 ( .A1(n41580), .A2(n41581), .ZN(n25374) );
  NOR2HSV2 U27269 ( .A1(n41847), .A2(n41511), .ZN(n41583) );
  CLKNAND2HSV2 U27270 ( .A1(n40778), .A2(n40776), .ZN(n40775) );
  INHSV4 U27271 ( .I(n44690), .ZN(n50199) );
  BUFHSV6 U27272 ( .I(n50199), .Z(n57970) );
  CLKNAND2HSV4 U27273 ( .A1(n33276), .A2(n33676), .ZN(n33527) );
  NOR2HSV4 U27274 ( .A1(n33527), .A2(n33517), .ZN(n33519) );
  INHSV2 U27275 ( .I(n31365), .ZN(n31363) );
  NAND2HSV4 U27276 ( .A1(n31322), .A2(n31323), .ZN(n31365) );
  NAND3HSV4 U27277 ( .A1(n37758), .A2(n37757), .A3(n39227), .ZN(n39387) );
  XNOR2HSV4 U27278 ( .A1(n25375), .A2(n39117), .ZN(n26789) );
  CLKNAND2HSV2 U27279 ( .A1(n39116), .A2(n52767), .ZN(n25375) );
  INHSV4 U27280 ( .I(n36894), .ZN(n25910) );
  NOR2HSV4 U27281 ( .A1(n25910), .A2(n25908), .ZN(n29713) );
  INHSV4 U27282 ( .I(n32418), .ZN(n32416) );
  CLKNAND2HSV2 U27283 ( .A1(n31289), .A2(n31288), .ZN(n31294) );
  NAND2HSV2 U27284 ( .A1(n26586), .A2(n29644), .ZN(n31892) );
  CLKNAND2HSV2 U27285 ( .A1(n32150), .A2(n32149), .ZN(n32238) );
  INHSV2 U27286 ( .I(n37101), .ZN(n37088) );
  INHSV4 U27287 ( .I(n37088), .ZN(n37237) );
  INHSV24 U27288 ( .I(n39218), .ZN(n25376) );
  NAND3HSV2 U27289 ( .A1(n25376), .A2(n39227), .A3(n37553), .ZN(n29022) );
  INHSV4 U27290 ( .I(n33231), .ZN(n33234) );
  NAND2HSV4 U27291 ( .A1(n33233), .A2(n33234), .ZN(n33235) );
  CLKNAND2HSV4 U27292 ( .A1(n32469), .A2(n32240), .ZN(n32309) );
  NAND3HSV4 U27293 ( .A1(n37339), .A2(n37338), .A3(n37337), .ZN(n37408) );
  CLKNAND2HSV2 U27294 ( .A1(n39880), .A2(n39879), .ZN(n39991) );
  CLKNAND2HSV2 U27295 ( .A1(n39364), .A2(n39363), .ZN(n39372) );
  CLKNHSV2 U27296 ( .I(n25377), .ZN(n31890) );
  CLKNAND2HSV2 U27297 ( .A1(n25912), .A2(n25378), .ZN(n25377) );
  CLKNHSV2 U27298 ( .I(n31885), .ZN(n25378) );
  CLKNAND2HSV4 U27299 ( .A1(n39542), .A2(n39692), .ZN(n31097) );
  CLKNAND2HSV2 U27300 ( .A1(n25379), .A2(n26023), .ZN(n26022) );
  NAND3HSV4 U27301 ( .A1(n25380), .A2(n33172), .A3(n34419), .ZN(n25379) );
  CLKNHSV2 U27302 ( .I(n33108), .ZN(n25380) );
  NAND2HSV2 U27303 ( .A1(n32452), .A2(n32458), .ZN(n32456) );
  INHSV6 U27304 ( .I(n55144), .ZN(n54541) );
  XNOR2HSV4 U27305 ( .A1(n25381), .A2(n33255), .ZN(n33262) );
  XNOR2HSV4 U27306 ( .A1(n25444), .A2(n25445), .ZN(n25381) );
  OAI21HSV4 U27307 ( .A1(n36744), .A2(n36743), .B(n36742), .ZN(n36773) );
  CLKNAND2HSV2 U27308 ( .A1(n30663), .A2(n30662), .ZN(n30664) );
  INHSV4 U27309 ( .I(n37780), .ZN(n37778) );
  CLKNHSV6 U27310 ( .I(n40860), .ZN(n40941) );
  INHSV6 U27311 ( .I(n31255), .ZN(n32881) );
  XNOR2HSV4 U27312 ( .A1(n25382), .A2(n36803), .ZN(n36856) );
  CLKNAND2HSV2 U27313 ( .A1(n36786), .A2(n25383), .ZN(n25382) );
  NAND3HSV3 U27314 ( .A1(n36861), .A2(n36841), .A3(n42806), .ZN(n36777) );
  INHSV2 U27315 ( .I(n36777), .ZN(n36778) );
  XNOR2HSV4 U27316 ( .A1(n25384), .A2(n36764), .ZN(n36766) );
  XNOR2HSV4 U27317 ( .A1(n25385), .A2(n36757), .ZN(n25384) );
  XNOR2HSV4 U27318 ( .A1(n25704), .A2(n25705), .ZN(n25385) );
  OAI22HSV2 U27319 ( .A1(n40866), .A2(n40865), .B1(n40864), .B2(n42478), .ZN(
        n40867) );
  NAND2HSV4 U27320 ( .A1(n40955), .A2(n41727), .ZN(n40868) );
  OAI21HSV4 U27321 ( .A1(n41142), .A2(n40868), .B(n40867), .ZN(n40869) );
  CLKNAND2HSV2 U27322 ( .A1(n26417), .A2(n58052), .ZN(n49961) );
  INHSV4 U27323 ( .I(n38456), .ZN(n38373) );
  NOR2HSV2 U27324 ( .A1(n26504), .A2(n26502), .ZN(n26501) );
  INHSV4 U27325 ( .I(n39872), .ZN(n39569) );
  BUFHSV4 U27326 ( .I(n45794), .Z(n49253) );
  MOAI22HSV4 U27327 ( .A1(n47947), .A2(n26758), .B1(n47387), .B2(
        \pe5/ti_7t [22]), .ZN(n26757) );
  NOR2HSV4 U27328 ( .A1(n26571), .A2(n38518), .ZN(n26570) );
  NAND2HSV4 U27329 ( .A1(n26570), .A2(n38519), .ZN(n26568) );
  CLKNHSV2 U27330 ( .I(n26780), .ZN(n25387) );
  NAND3HSV4 U27331 ( .A1(n35456), .A2(n25389), .A3(n25388), .ZN(n35486) );
  CLKNHSV2 U27332 ( .I(n26693), .ZN(n25388) );
  CLKNAND2HSV2 U27333 ( .A1(n26695), .A2(n26694), .ZN(n25389) );
  NAND2HSV2 U27334 ( .A1(n26536), .A2(n26527), .ZN(n26526) );
  INHSV2 U27335 ( .I(n26213), .ZN(n26212) );
  CLKNHSV6 U27336 ( .I(n32506), .ZN(n49743) );
  NAND2HSV4 U27337 ( .A1(n48484), .A2(n43865), .ZN(n26327) );
  INHSV2 U27338 ( .I(n25390), .ZN(n32027) );
  CLKNAND2HSV2 U27339 ( .A1(n32026), .A2(n29719), .ZN(n25390) );
  XNOR2HSV4 U27340 ( .A1(n48002), .A2(n48003), .ZN(n31709) );
  INHSV8 U27341 ( .I(n43242), .ZN(n42899) );
  NAND2HSV2 U27342 ( .A1(n37652), .A2(n30142), .ZN(n31096) );
  INHSV2 U27343 ( .I(n26083), .ZN(n38602) );
  NAND3HSV4 U27344 ( .A1(n39717), .A2(n39558), .A3(n39722), .ZN(n39568) );
  NAND2HSV2 U27345 ( .A1(n52668), .A2(n51418), .ZN(n51434) );
  CLKNAND2HSV4 U27346 ( .A1(n41417), .A2(n41416), .ZN(pov1[19]) );
  NAND2HSV4 U27347 ( .A1(pov1[19]), .A2(n53787), .ZN(n41588) );
  NOR2HSV4 U27348 ( .A1(n33246), .A2(n26966), .ZN(n33270) );
  NAND3HSV4 U27349 ( .A1(n40299), .A2(n40298), .A3(n40297), .ZN(n40300) );
  CLKNHSV6 U27350 ( .I(n40300), .ZN(n40315) );
  OAI21HSV4 U27351 ( .A1(n37032), .A2(n37033), .B(n37031), .ZN(n37039) );
  NOR2HSV4 U27352 ( .A1(n44042), .A2(n25391), .ZN(n44166) );
  CLKNHSV2 U27353 ( .I(n45105), .ZN(n25391) );
  NAND3HSV4 U27354 ( .A1(n44943), .A2(n44168), .A3(n44177), .ZN(n45105) );
  CLKNAND2HSV2 U27355 ( .A1(n42584), .A2(n42694), .ZN(n42585) );
  INHSV4 U27356 ( .I(n26254), .ZN(n26103) );
  BUFHSV6 U27357 ( .I(n59810), .Z(n45732) );
  INHSV4 U27358 ( .I(n31677), .ZN(n31678) );
  NOR2HSV4 U27359 ( .A1(n31678), .A2(n31685), .ZN(n31679) );
  NAND3HSV2 U27360 ( .A1(n56417), .A2(n56171), .A3(n56418), .ZN(n29098) );
  NAND2HSV2 U27361 ( .A1(n29098), .A2(n29097), .ZN(n29099) );
  INHSV2 U27362 ( .I(n45794), .ZN(n26121) );
  NOR2HSV4 U27363 ( .A1(n26121), .A2(n26120), .ZN(n26126) );
  CLKNAND2HSV2 U27364 ( .A1(n45937), .A2(n45936), .ZN(n45938) );
  INHSV2 U27365 ( .I(n38607), .ZN(n46122) );
  CLKNAND2HSV4 U27366 ( .A1(n40001), .A2(n47199), .ZN(n40296) );
  INHSV4 U27367 ( .I(n32688), .ZN(n32666) );
  XNOR2HSV4 U27368 ( .A1(n50123), .A2(n50122), .ZN(n50126) );
  INHSV2 U27369 ( .I(n53279), .ZN(n28959) );
  CLKNHSV2 U27370 ( .I(n40139), .ZN(n25392) );
  CLKNHSV2 U27371 ( .I(n40140), .ZN(n25393) );
  CLKAND2HSV4 U27372 ( .A1(n32543), .A2(n32542), .Z(n32464) );
  OAI21HSV4 U27373 ( .A1(n32464), .A2(n32686), .B(n32551), .ZN(n32465) );
  INHSV4 U27374 ( .I(n35721), .ZN(n26472) );
  CLKNAND2HSV4 U27375 ( .A1(n37105), .A2(n42899), .ZN(n37156) );
  CLKNAND2HSV4 U27376 ( .A1(n37156), .A2(n37155), .ZN(n37251) );
  INHSV2 U27377 ( .I(n31456), .ZN(n31458) );
  CLKNAND2HSV4 U27378 ( .A1(n31357), .A2(n31356), .ZN(n31456) );
  CLKNHSV2 U27379 ( .I(n29767), .ZN(n25394) );
  XNOR2HSV4 U27380 ( .A1(n41830), .A2(n41829), .ZN(n29767) );
  AOI21HSV4 U27381 ( .A1(n25395), .A2(n30667), .B(n30666), .ZN(n30668) );
  CLKNAND2HSV2 U27382 ( .A1(n30664), .A2(n30665), .ZN(n25395) );
  CLKNAND2HSV2 U27383 ( .A1(n36863), .A2(n36844), .ZN(n36845) );
  CLKNAND2HSV2 U27384 ( .A1(n42512), .A2(n29704), .ZN(n37262) );
  NOR2HSV2 U27385 ( .A1(n44833), .A2(n44969), .ZN(n44288) );
  CLKNAND2HSV2 U27386 ( .A1(n42466), .A2(n59994), .ZN(n42467) );
  INAND2HSV4 U27387 ( .A1(n38455), .B1(n38373), .ZN(n38537) );
  XNOR2HSV4 U27388 ( .A1(n31460), .A2(n25396), .ZN(n31466) );
  CLKNHSV2 U27389 ( .I(n31459), .ZN(n25396) );
  CLKNAND2HSV4 U27390 ( .A1(n49743), .A2(n49665), .ZN(n25486) );
  MUX2NHSV4 U27391 ( .I0(n32307), .I1(n25486), .S(n32308), .ZN(n25485) );
  XNOR2HSV4 U27392 ( .A1(n37746), .A2(n37745), .ZN(n37747) );
  CLKNAND2HSV8 U27393 ( .A1(n53381), .A2(n37786), .ZN(n37918) );
  CLKNAND2HSV2 U27394 ( .A1(n41592), .A2(n42202), .ZN(n41589) );
  INHSV6 U27395 ( .I(n37040), .ZN(n37170) );
  INHSV4 U27396 ( .I(n37040), .ZN(n59364) );
  AOI21HSV4 U27397 ( .A1(n38116), .A2(n38115), .B(n38114), .ZN(n38117) );
  NAND2HSV4 U27398 ( .A1(n26585), .A2(n26584), .ZN(pov4[29]) );
  XNOR2HSV4 U27399 ( .A1(n57664), .A2(n57663), .ZN(n57666) );
  XNOR2HSV2 U27400 ( .A1(n57666), .A2(n57665), .ZN(n57667) );
  XOR2HSV2 U27401 ( .A1(n25397), .A2(n38326), .Z(n38330) );
  XNOR2HSV4 U27402 ( .A1(n26773), .A2(n26771), .ZN(n25397) );
  CLKNAND2HSV4 U27403 ( .A1(n48046), .A2(\pe6/pvq [11]), .ZN(n31565) );
  INHSV4 U27404 ( .I(n26406), .ZN(n26405) );
  CLKAND2HSV4 U27405 ( .A1(n25882), .A2(n42899), .Z(n29641) );
  BUFHSV4 U27406 ( .I(n40657), .Z(n25398) );
  AOI31HSV2 U27407 ( .A1(n48012), .A2(n31524), .A3(n36065), .B(n31405), .ZN(
        n31406) );
  NAND2HSV4 U27408 ( .A1(n46627), .A2(n59087), .ZN(n31604) );
  BUFHSV8 U27409 ( .I(n33218), .Z(n33437) );
  NOR2HSV8 U27410 ( .A1(n33437), .A2(n33928), .ZN(n33267) );
  NAND3HSV4 U27411 ( .A1(n26304), .A2(n26302), .A3(n45145), .ZN(n52917) );
  BUFHSV6 U27412 ( .I(n52917), .Z(n25831) );
  INHSV2 U27413 ( .I(n42338), .ZN(n25399) );
  CLKNAND2HSV2 U27414 ( .A1(n25399), .A2(n42490), .ZN(n42332) );
  INHSV4 U27415 ( .I(\pe6/phq [3]), .ZN(n31335) );
  NAND2HSV4 U27416 ( .A1(n46625), .A2(n32740), .ZN(n31275) );
  CLKNAND2HSV4 U27417 ( .A1(n31593), .A2(\pe6/pvq [6]), .ZN(n26460) );
  INHSV2 U27418 ( .I(n46144), .ZN(n46152) );
  MUX2NHSV4 U27419 ( .I0(n42912), .I1(n25400), .S(n42911), .ZN(n25697) );
  NOR2HSV2 U27420 ( .A1(n43349), .A2(n25891), .ZN(n43245) );
  XNOR2HSV4 U27421 ( .A1(n43241), .A2(n43240), .ZN(n43349) );
  CLKNAND2HSV2 U27422 ( .A1(n36888), .A2(n29695), .ZN(n25401) );
  INHSV8 U27423 ( .I(n33114), .ZN(n57242) );
  NAND2HSV4 U27424 ( .A1(n57242), .A2(n33249), .ZN(n26628) );
  CLKNAND2HSV2 U27425 ( .A1(n42085), .A2(\pe1/got [27]), .ZN(n42184) );
  XNOR2HSV4 U27426 ( .A1(n35714), .A2(n35713), .ZN(n36034) );
  CLKNAND2HSV2 U27427 ( .A1(n36203), .A2(n35808), .ZN(n35713) );
  INHSV4 U27428 ( .I(n34485), .ZN(n33326) );
  INHSV8 U27429 ( .I(n25719), .ZN(n36861) );
  CLKNAND2HSV4 U27430 ( .A1(n47499), .A2(n44709), .ZN(n44957) );
  NOR2HSV4 U27431 ( .A1(n44957), .A2(n44958), .ZN(n44964) );
  XNOR2HSV4 U27432 ( .A1(n25403), .A2(n25402), .ZN(\pe6/poht [21]) );
  CLKNAND2HSV2 U27433 ( .A1(n29772), .A2(n58572), .ZN(n25402) );
  XOR2HSV2 U27434 ( .A1(n58523), .A2(n25404), .Z(n25403) );
  CLKNHSV2 U27435 ( .I(n58524), .ZN(n25404) );
  NOR2HSV4 U27436 ( .A1(n42343), .A2(n42340), .ZN(n42334) );
  XOR2HSV2 U27437 ( .A1(n25405), .A2(n48997), .Z(n26654) );
  NOR2HSV4 U27438 ( .A1(n25833), .A2(n25406), .ZN(n25405) );
  CLKNHSV2 U27439 ( .I(n53086), .ZN(n25406) );
  NOR2HSV4 U27440 ( .A1(n37332), .A2(n37268), .ZN(n37090) );
  INHSV4 U27441 ( .I(n38097), .ZN(n26893) );
  NAND2HSV4 U27442 ( .A1(n50213), .A2(n34441), .ZN(n34443) );
  MUX2NHSV2 U27443 ( .I0(n25407), .I1(n33933), .S(n33932), .ZN(n33981) );
  CLKNAND2HSV2 U27444 ( .A1(n25409), .A2(n25408), .ZN(n25407) );
  CLKNHSV2 U27445 ( .I(n33928), .ZN(n25408) );
  CLKNHSV2 U27446 ( .I(n48892), .ZN(n25409) );
  CLKNHSV6 U27447 ( .I(n26414), .ZN(n45400) );
  INHSV24 U27448 ( .I(n37092), .ZN(n25410) );
  INAND2HSV4 U27449 ( .A1(n37335), .B1(n25410), .ZN(n29707) );
  NAND2HSV4 U27450 ( .A1(n37039), .A2(n37038), .ZN(n37166) );
  XNOR2HSV4 U27451 ( .A1(n37341), .A2(n25411), .ZN(n37342) );
  CLKNAND2HSV2 U27452 ( .A1(n37408), .A2(n37340), .ZN(n25411) );
  CLKNAND2HSV2 U27453 ( .A1(n36072), .A2(n44692), .ZN(n36075) );
  NAND3HSV3 U27454 ( .A1(n46766), .A2(n53102), .A3(n46818), .ZN(n46901) );
  CLKNAND2HSV4 U27455 ( .A1(n48461), .A2(n48462), .ZN(n25412) );
  BUFHSV4 U27456 ( .I(n35479), .Z(n58207) );
  BUFHSV8 U27457 ( .I(n26738), .Z(n26417) );
  CLKAND2HSV8 U27458 ( .A1(n44949), .A2(n45108), .Z(n29696) );
  INHSV8 U27459 ( .I(n41843), .ZN(n41844) );
  CLKNAND2HSV8 U27460 ( .A1(n41845), .A2(n41844), .ZN(n29735) );
  BUFHSV8 U27461 ( .I(n50400), .Z(n58183) );
  XNOR2HSV4 U27462 ( .A1(n42463), .A2(n42462), .ZN(n42464) );
  AOI21HSV4 U27463 ( .A1(n31818), .A2(n32329), .B(n48010), .ZN(n31819) );
  CLKNAND2HSV4 U27464 ( .A1(n25449), .A2(n36735), .ZN(n36726) );
  INHSV4 U27465 ( .I(n52815), .ZN(n26626) );
  AOI21HSV4 U27466 ( .A1(n25415), .A2(n25414), .B(n25413), .ZN(n39362) );
  CLKNHSV2 U27467 ( .I(n39357), .ZN(n25413) );
  CLKNHSV2 U27468 ( .I(n39358), .ZN(n25414) );
  CLKNHSV2 U27469 ( .I(n39359), .ZN(n25415) );
  AOI22HSV4 U27470 ( .A1(n46574), .A2(n32533), .B1(n32532), .B2(n32642), .ZN(
        n32537) );
  NAND2HSV4 U27471 ( .A1(n32537), .A2(n32536), .ZN(n32538) );
  CLKNAND2HSV4 U27472 ( .A1(n39740), .A2(n40131), .ZN(n40285) );
  NAND2HSV2 U27473 ( .A1(n46415), .A2(n42936), .ZN(n42902) );
  OAI21HSV4 U27474 ( .A1(n25416), .A2(n36519), .B(n39007), .ZN(n43916) );
  XNOR2HSV4 U27475 ( .A1(n44034), .A2(n60002), .ZN(n25416) );
  XNOR2HSV4 U27476 ( .A1(n44140), .A2(n44139), .ZN(n44141) );
  XNOR2HSV4 U27477 ( .A1(n39859), .A2(n39858), .ZN(n39862) );
  NAND2HSV2 U27478 ( .A1(n37274), .A2(n46309), .ZN(n36765) );
  NAND2HSV4 U27479 ( .A1(n25417), .A2(n41128), .ZN(n41130) );
  CLKNAND2HSV4 U27480 ( .A1(n41126), .A2(n41127), .ZN(n25417) );
  CLKNAND2HSV2 U27481 ( .A1(n36695), .A2(\pe3/got [30]), .ZN(n25418) );
  CLKNAND2HSV4 U27482 ( .A1(n37774), .A2(n37773), .ZN(n39408) );
  MUX2NHSV4 U27483 ( .I0(n42706), .I1(n53376), .S(n53377), .ZN(n37419) );
  NAND2HSV0 U27484 ( .A1(n25848), .A2(n55514), .ZN(n55602) );
  INAND2HSV4 U27485 ( .A1(n30059), .B1(n25419), .ZN(n30080) );
  CLKNHSV2 U27486 ( .I(n30058), .ZN(n25419) );
  NAND2HSV2 U27487 ( .A1(n55423), .A2(n53390), .ZN(n54725) );
  CLKXOR2HSV4 U27488 ( .A1(n52406), .A2(n52405), .Z(n52407) );
  DELHS1 U27489 ( .I(\pe4/got [32]), .Z(n25420) );
  NAND2HSV4 U27490 ( .A1(n44694), .A2(n30513), .ZN(n30961) );
  CLKNAND2HSV2 U27491 ( .A1(n55423), .A2(\pe1/got [21]), .ZN(n54809) );
  CLKNAND2HSV2 U27492 ( .A1(n25421), .A2(n35454), .ZN(n35020) );
  CLKNAND2HSV2 U27493 ( .A1(n35305), .A2(n35009), .ZN(n35464) );
  NOR2HSV8 U27494 ( .A1(n25425), .A2(n25424), .ZN(n26424) );
  INHSV4 U27495 ( .I(n38023), .ZN(n37853) );
  NAND2HSV4 U27496 ( .A1(n37852), .A2(n37853), .ZN(n25668) );
  NAND2HSV4 U27497 ( .A1(n26080), .A2(n26082), .ZN(n31362) );
  BUFHSV8 U27498 ( .I(n55476), .Z(n59931) );
  NAND2HSV2 U27499 ( .A1(n59931), .A2(n54965), .ZN(n54802) );
  CLKNHSV6 U27500 ( .I(n36916), .ZN(n59569) );
  NAND2HSV4 U27501 ( .A1(n26789), .A2(n39250), .ZN(n39254) );
  CLKNAND2HSV4 U27502 ( .A1(n39254), .A2(n39253), .ZN(n39351) );
  XNOR2HSV4 U27503 ( .A1(n40286), .A2(n25422), .ZN(n40287) );
  CLKNAND2HSV2 U27504 ( .A1(n40285), .A2(n30779), .ZN(n25422) );
  CLKNHSV0 U27505 ( .I(n25889), .ZN(n46140) );
  INAND2HSV4 U27506 ( .A1(n46620), .B1(n59276), .ZN(n33019) );
  XOR4HSV4 U27507 ( .A1(n31316), .A2(n31315), .A3(n33019), .A4(n31314), .Z(
        n31317) );
  XNOR2HSV4 U27508 ( .A1(n39984), .A2(n39983), .ZN(n39987) );
  INHSV2 U27509 ( .I(n37864), .ZN(n25423) );
  NOR2HSV4 U27510 ( .A1(n25423), .A2(n37863), .ZN(n29632) );
  XNOR2HSV4 U27511 ( .A1(n32021), .A2(n32020), .ZN(n32023) );
  INHSV4 U27512 ( .I(n40484), .ZN(n59498) );
  NAND2HSV4 U27513 ( .A1(n26034), .A2(n26033), .ZN(n26001) );
  NAND2HSV2 U27514 ( .A1(n40278), .A2(n31225), .ZN(n39667) );
  CLKNAND2HSV4 U27515 ( .A1(n39680), .A2(n39681), .ZN(n39676) );
  INHSV4 U27516 ( .I(n39676), .ZN(n37781) );
  CLKNHSV6 U27517 ( .I(n38388), .ZN(n50929) );
  CLKNHSV0 U27518 ( .I(n38388), .ZN(n52176) );
  NOR2HSV4 U27519 ( .A1(n29774), .A2(n35034), .ZN(n57087) );
  NAND3HSV4 U27520 ( .A1(n46817), .A2(n46766), .A3(n46633), .ZN(n28761) );
  CLKNAND2HSV2 U27521 ( .A1(n28760), .A2(n28761), .ZN(n28762) );
  CLKNAND2HSV4 U27522 ( .A1(n26202), .A2(n26203), .ZN(n52734) );
  CLKNHSV6 U27523 ( .I(n51727), .ZN(n52047) );
  NAND3HSV4 U27524 ( .A1(n30991), .A2(n31005), .A3(n39741), .ZN(n30978) );
  CLKAND2HSV4 U27525 ( .A1(n30978), .A2(n52817), .Z(n29697) );
  CLKNAND2HSV2 U27526 ( .A1(n60040), .A2(n30063), .ZN(n30066) );
  NAND2HSV4 U27527 ( .A1(n30066), .A2(n30065), .ZN(n30068) );
  INHSV4 U27528 ( .I(n30088), .ZN(n25424) );
  INHSV4 U27529 ( .I(n30137), .ZN(n25425) );
  CLKNAND2HSV4 U27530 ( .A1(n25426), .A2(n32561), .ZN(n32820) );
  CLKNAND2HSV4 U27531 ( .A1(n32560), .A2(n32559), .ZN(n25426) );
  NAND3HSV4 U27532 ( .A1(n37332), .A2(n37240), .A3(n37238), .ZN(n37338) );
  BUFHSV8 U27533 ( .I(n59914), .Z(n32833) );
  INHSV4 U27534 ( .I(n30887), .ZN(n30783) );
  CLKXOR2HSV4 U27535 ( .A1(n37403), .A2(n37402), .Z(n37405) );
  XNOR2HSV2 U27536 ( .A1(n37405), .A2(n37404), .ZN(n37406) );
  DELHS1 U27537 ( .I(n59574), .Z(n25427) );
  DELHS1 U27538 ( .I(\pe1/bq[30] ), .Z(n25428) );
  CLKNAND2HSV3 U27539 ( .A1(n37101), .A2(n37100), .ZN(n37102) );
  INHSV6 U27540 ( .I(n46031), .ZN(n37040) );
  NAND2HSV4 U27541 ( .A1(n36919), .A2(n36918), .ZN(n46031) );
  NAND2HSV4 U27542 ( .A1(n25429), .A2(n30762), .ZN(n31135) );
  CLKNAND2HSV4 U27543 ( .A1(n30761), .A2(n30760), .ZN(n25429) );
  NAND2HSV4 U27544 ( .A1(n37541), .A2(n31102), .ZN(n31103) );
  NOR2HSV4 U27545 ( .A1(n31104), .A2(n31103), .ZN(n31238) );
  XNOR2HSV4 U27546 ( .A1(n25430), .A2(n46098), .ZN(n26074) );
  NAND3HSV4 U27547 ( .A1(n46081), .A2(n46079), .A3(n46080), .ZN(n25430) );
  NAND2HSV4 U27548 ( .A1(n39729), .A2(n39728), .ZN(n39740) );
  XNOR2HSV4 U27549 ( .A1(n25431), .A2(n40349), .ZN(n26826) );
  INHSV2 U27550 ( .I(n45499), .ZN(n26539) );
  CLKNHSV6 U27551 ( .I(n36309), .ZN(n36311) );
  CLKNAND2HSV8 U27552 ( .A1(n36311), .A2(n36310), .ZN(n36313) );
  NAND2HSV2 U27553 ( .A1(n25433), .A2(n39670), .ZN(n25432) );
  NOR2HSV2 U27554 ( .A1(n25435), .A2(n25434), .ZN(n25433) );
  NAND2HSV2 U27555 ( .A1(n39671), .A2(n39693), .ZN(n25434) );
  INHSV2 U27556 ( .I(n47946), .ZN(n25435) );
  XNOR2HSV4 U27557 ( .A1(n25436), .A2(n36479), .ZN(n36484) );
  XOR2HSV2 U27558 ( .A1(n36476), .A2(n36477), .Z(n25436) );
  CLKNAND2HSV2 U27559 ( .A1(n40474), .A2(n40473), .ZN(n40475) );
  NAND2HSV4 U27560 ( .A1(n40476), .A2(n40475), .ZN(n40478) );
  INHSV4 U27561 ( .I(n39664), .ZN(n39537) );
  NOR2HSV2 U27562 ( .A1(n36557), .A2(n59586), .ZN(n36472) );
  CLKNAND2HSV2 U27563 ( .A1(n59674), .A2(n41689), .ZN(n40701) );
  NOR2HSV4 U27564 ( .A1(n25438), .A2(n25437), .ZN(n39738) );
  CLKNHSV2 U27565 ( .I(n39736), .ZN(n25437) );
  CLKNAND2HSV2 U27566 ( .A1(n39737), .A2(n39735), .ZN(n25438) );
  NAND2HSV4 U27567 ( .A1(n40757), .A2(n40933), .ZN(n40650) );
  XNOR2HSV4 U27568 ( .A1(n55939), .A2(n55938), .ZN(n55943) );
  CLKNAND2HSV4 U27569 ( .A1(n26066), .A2(n26065), .ZN(n26418) );
  CLKXOR2HSV4 U27570 ( .A1(n51957), .A2(n51956), .Z(n51960) );
  CLKXOR2HSV4 U27571 ( .A1(n51527), .A2(n51526), .Z(n51529) );
  CLKNAND2HSV2 U27572 ( .A1(n59394), .A2(n40700), .ZN(n40506) );
  INHSV4 U27573 ( .I(n40506), .ZN(n40508) );
  XNOR2HSV4 U27574 ( .A1(n56257), .A2(n56256), .ZN(n56258) );
  XOR3HSV2 U27575 ( .A1(n55811), .A2(n55812), .A3(n25439), .Z(n55814) );
  CLKNHSV2 U27576 ( .I(n55813), .ZN(n25439) );
  CLKNAND2HSV4 U27577 ( .A1(n59569), .A2(n36850), .ZN(n36882) );
  NAND3HSV4 U27578 ( .A1(n36882), .A2(n36881), .A3(n29682), .ZN(n36915) );
  NAND2HSV2 U27579 ( .A1(n37298), .A2(n25787), .ZN(n42747) );
  INHSV4 U27580 ( .I(n31253), .ZN(n31369) );
  NAND2HSV2 U27581 ( .A1(n31369), .A2(\pe6/bq[28] ), .ZN(n32105) );
  INHSV4 U27582 ( .I(n37185), .ZN(n36789) );
  NAND2HSV4 U27583 ( .A1(n37012), .A2(n36955), .ZN(n36829) );
  INHSV4 U27584 ( .I(n26738), .ZN(n50111) );
  INHSV4 U27585 ( .I(n50111), .ZN(n58299) );
  BUFHSV16 U27586 ( .I(n45499), .Z(n52693) );
  NAND2HSV2 U27587 ( .A1(n52693), .A2(n48742), .ZN(n48303) );
  CLKNHSV2 U27588 ( .I(n26609), .ZN(n25440) );
  NOR2HSV2 U27589 ( .A1(n26087), .A2(n48324), .ZN(n26086) );
  CLKNAND2HSV2 U27590 ( .A1(n29735), .A2(n42316), .ZN(n26087) );
  NOR2HSV4 U27591 ( .A1(n25442), .A2(n26066), .ZN(n48162) );
  CLKNAND2HSV4 U27592 ( .A1(n45106), .A2(n44041), .ZN(n44042) );
  CLKNAND2HSV2 U27593 ( .A1(n52785), .A2(n52787), .ZN(n30775) );
  CLKXOR2HSV4 U27594 ( .A1(n50103), .A2(n50102), .Z(n50105) );
  CLKNAND2HSV2 U27595 ( .A1(n25443), .A2(n43023), .ZN(n25696) );
  AOI31HSV2 U27596 ( .A1(n43127), .A2(n43236), .A3(n36692), .B(n43022), .ZN(
        n25443) );
  CLKNAND2HSV2 U27597 ( .A1(n42928), .A2(n42927), .ZN(n42932) );
  XNOR2HSV4 U27598 ( .A1(n33253), .A2(n33252), .ZN(n25444) );
  XOR2HSV2 U27599 ( .A1(n33254), .A2(n33251), .Z(n25445) );
  OAI22HSV4 U27600 ( .A1(n36635), .A2(n36566), .B1(n36568), .B2(n36565), .ZN(
        n36567) );
  INHSV4 U27601 ( .I(n36567), .ZN(n36572) );
  INHSV6 U27602 ( .I(\pe6/ctrq ), .ZN(n31255) );
  CLKNHSV6 U27603 ( .I(n26789), .ZN(pov5[20]) );
  CLKNAND2HSV8 U27604 ( .A1(pov5[20]), .A2(n31102), .ZN(n39429) );
  BUFHSV8 U27605 ( .I(n49661), .Z(n52910) );
  MUX2NHSV4 U27606 ( .I0(n39355), .I1(n39367), .S(n29022), .ZN(n39389) );
  CLKNAND2HSV2 U27607 ( .A1(n36683), .A2(n36684), .ZN(n36688) );
  CLKNAND2HSV4 U27608 ( .A1(n36688), .A2(n36844), .ZN(n25776) );
  INHSV4 U27609 ( .I(n45783), .ZN(n25947) );
  CLKNAND2HSV4 U27610 ( .A1(n31238), .A2(n37756), .ZN(n37762) );
  CLKNAND2HSV2 U27611 ( .A1(n42046), .A2(n42045), .ZN(n42077) );
  CLKNAND2HSV4 U27612 ( .A1(n41328), .A2(n41697), .ZN(n29208) );
  NOR2HSV8 U27613 ( .A1(n34342), .A2(n34341), .ZN(n34575) );
  NAND2HSV4 U27614 ( .A1(n60009), .A2(n42335), .ZN(n40380) );
  NAND2HSV4 U27615 ( .A1(n25521), .A2(n31819), .ZN(n32033) );
  INHSV2 U27616 ( .I(n25916), .ZN(n25915) );
  INHSV4 U27617 ( .I(n36638), .ZN(n26879) );
  CLKNAND2HSV4 U27618 ( .A1(n34587), .A2(n34333), .ZN(n34334) );
  NOR2HSV4 U27619 ( .A1(n32667), .A2(n36065), .ZN(n32659) );
  CLKNHSV0 U27620 ( .I(n56059), .ZN(n56976) );
  OAI21HSV4 U27621 ( .A1(n40639), .A2(n40552), .B(n40532), .ZN(n40533) );
  INHSV4 U27622 ( .I(n40533), .ZN(n40537) );
  INHSV4 U27623 ( .I(n40590), .ZN(n40587) );
  NAND2HSV4 U27624 ( .A1(n40587), .A2(n40588), .ZN(n40592) );
  CLKNAND2HSV2 U27625 ( .A1(n48480), .A2(n36958), .ZN(n28972) );
  CLKNAND2HSV2 U27626 ( .A1(n48893), .A2(n36724), .ZN(n36745) );
  INHSV2 U27627 ( .I(n36745), .ZN(n36746) );
  BUFHSV8 U27628 ( .I(n36775), .Z(n36863) );
  NOR2HSV4 U27629 ( .A1(n36863), .A2(n37454), .ZN(n36744) );
  AOI21HSV2 U27630 ( .A1(n34587), .A2(n25447), .B(n25446), .ZN(n29709) );
  CLKNHSV2 U27631 ( .I(n34822), .ZN(n25446) );
  CLKNHSV2 U27632 ( .I(n34588), .ZN(n25447) );
  CLKNAND2HSV2 U27633 ( .A1(n36466), .A2(n36467), .ZN(n36468) );
  NAND2HSV4 U27634 ( .A1(n36723), .A2(n36722), .ZN(n25449) );
  DELHS1 U27635 ( .I(n41824), .Z(n25448) );
  INHSV4 U27636 ( .I(n40150), .ZN(n40151) );
  INHSV4 U27637 ( .I(n40149), .ZN(n40152) );
  NAND2HSV4 U27638 ( .A1(n40152), .A2(n40151), .ZN(n40153) );
  INHSV4 U27639 ( .I(n47920), .ZN(n58272) );
  NAND2HSV2 U27640 ( .A1(n58272), .A2(n57672), .ZN(n50411) );
  CLKNHSV0 U27641 ( .I(n50301), .ZN(n35033) );
  INHSV2 U27642 ( .I(n50301), .ZN(n59950) );
  XNOR2HSV4 U27643 ( .A1(n52891), .A2(n52892), .ZN(n52894) );
  BUFHSV16 U27644 ( .I(n59579), .Z(n25570) );
  NAND2HSV4 U27645 ( .A1(n26582), .A2(n32551), .ZN(n32801) );
  NAND2HSV4 U27646 ( .A1(n30991), .A2(n25450), .ZN(n37534) );
  NAND2HSV4 U27647 ( .A1(n31119), .A2(n31240), .ZN(n25450) );
  NAND2HSV4 U27648 ( .A1(n31117), .A2(n30863), .ZN(n30991) );
  CLKNAND2HSV2 U27649 ( .A1(n27578), .A2(n25451), .ZN(n27579) );
  CLKNAND2HSV2 U27650 ( .A1(n25453), .A2(n25452), .ZN(n25451) );
  CLKNHSV2 U27651 ( .I(n27577), .ZN(n25452) );
  CLKNAND2HSV2 U27652 ( .A1(n52840), .A2(n52276), .ZN(n27577) );
  CLKNHSV2 U27653 ( .I(n27576), .ZN(n25453) );
  XNOR2HSV4 U27654 ( .A1(n55283), .A2(n55282), .ZN(n55285) );
  INHSV2 U27655 ( .I(n45945), .ZN(n46073) );
  NAND2HSV2 U27656 ( .A1(n26827), .A2(n40377), .ZN(n40345) );
  AOI21HSV4 U27657 ( .A1(n30143), .A2(n30052), .B(n30090), .ZN(n30053) );
  CLKXOR2HSV4 U27658 ( .A1(n57448), .A2(n57447), .Z(n57450) );
  CLKXOR2HSV2 U27659 ( .A1(n57450), .A2(n57449), .Z(n57451) );
  CLKNAND2HSV4 U27660 ( .A1(n58104), .A2(n59663), .ZN(n27232) );
  CLKXOR2HSV2 U27661 ( .A1(n27231), .A2(n27232), .Z(n27233) );
  CLKXOR2HSV4 U27662 ( .A1(n58274), .A2(n58273), .Z(n58276) );
  CLKXOR2HSV2 U27663 ( .A1(n58276), .A2(n58275), .Z(n58277) );
  CLKNAND2HSV4 U27664 ( .A1(n58186), .A2(n47655), .ZN(n25557) );
  AOI21HSV4 U27665 ( .A1(n36916), .A2(n29701), .B(n36908), .ZN(n36912) );
  NAND2HSV4 U27666 ( .A1(n36912), .A2(n36911), .ZN(n36913) );
  NAND2HSV2 U27667 ( .A1(n39879), .A2(n59580), .ZN(n27010) );
  CLKXOR2HSV2 U27668 ( .A1(n27009), .A2(n27010), .Z(n27011) );
  CLKAND2HSV2 U27669 ( .A1(n38742), .A2(n38737), .Z(n38740) );
  CLKNAND2HSV2 U27670 ( .A1(n31368), .A2(n59278), .ZN(n31310) );
  NOR2HSV4 U27671 ( .A1(n42356), .A2(n44528), .ZN(n41907) );
  CLKNAND2HSV4 U27672 ( .A1(n25454), .A2(n33223), .ZN(n33238) );
  NAND2HSV2 U27673 ( .A1(n47903), .A2(n47567), .ZN(n52163) );
  CLKNAND2HSV4 U27674 ( .A1(n47902), .A2(n47901), .ZN(n47567) );
  INHSV4 U27675 ( .I(n30190), .ZN(n25527) );
  INHSV2 U27676 ( .I(n42316), .ZN(n42187) );
  AOI21HSV4 U27677 ( .A1(n29735), .A2(n42316), .B(n25455), .ZN(n42323) );
  CLKNAND2HSV2 U27678 ( .A1(n60104), .A2(n42484), .ZN(n25455) );
  CLKNAND2HSV4 U27679 ( .A1(n41843), .A2(n41838), .ZN(n42316) );
  XOR2HSV4 U27680 ( .A1(n31815), .A2(n31814), .Z(n25591) );
  NAND2HSV2 U27681 ( .A1(n52715), .A2(n29860), .ZN(n29861) );
  NAND2HSV4 U27682 ( .A1(n52695), .A2(n29842), .ZN(n52715) );
  XOR3HSV2 U27683 ( .A1(n25457), .A2(n30015), .A3(n25456), .Z(n30019) );
  CLKNHSV2 U27684 ( .I(n30014), .ZN(n25456) );
  XOR2HSV2 U27685 ( .A1(n30003), .A2(n30004), .Z(n25457) );
  OAI21HSV4 U27686 ( .A1(n37434), .A2(n43468), .B(n36692), .ZN(n42596) );
  INHSV2 U27687 ( .I(n47539), .ZN(n29745) );
  BUFHSV6 U27688 ( .I(n29745), .Z(n44283) );
  NOR2HSV2 U27689 ( .A1(n40016), .A2(n40160), .ZN(n40156) );
  NOR2HSV4 U27690 ( .A1(n40015), .A2(n25458), .ZN(n40160) );
  NAND2HSV2 U27691 ( .A1(n32427), .A2(n32426), .ZN(n32428) );
  CLKXOR2HSV4 U27692 ( .A1(n49600), .A2(n49599), .Z(n49601) );
  NAND3HSV4 U27693 ( .A1(n32314), .A2(n25459), .A3(n32316), .ZN(n32155) );
  NAND2HSV2 U27694 ( .A1(n29771), .A2(n59367), .ZN(n51416) );
  CLKNAND2HSV4 U27695 ( .A1(n42475), .A2(n42474), .ZN(n42483) );
  INHSV4 U27696 ( .I(n26341), .ZN(n43596) );
  CLKNAND2HSV4 U27697 ( .A1(n43899), .A2(n43596), .ZN(n43897) );
  INHSV2 U27698 ( .I(n29796), .ZN(n29795) );
  CLKNHSV6 U27699 ( .I(n31424), .ZN(n31339) );
  NAND2HSV4 U27700 ( .A1(n44807), .A2(n39007), .ZN(n38769) );
  CLKNAND2HSV4 U27701 ( .A1(n58184), .A2(n47841), .ZN(n27221) );
  NAND2HSV4 U27702 ( .A1(n43369), .A2(n43481), .ZN(n59575) );
  INHSV4 U27703 ( .I(n25570), .ZN(n58212) );
  INHSV4 U27704 ( .I(n25570), .ZN(n29752) );
  AOI21HSV4 U27705 ( .A1(n31743), .A2(n51439), .B(n32651), .ZN(n31744) );
  NAND2HSV4 U27706 ( .A1(n44182), .A2(n36654), .ZN(n44179) );
  INHSV2 U27707 ( .I(n42334), .ZN(n26282) );
  CLKNAND2HSV2 U27708 ( .A1(n48330), .A2(n48329), .ZN(n48334) );
  CLKNAND2HSV2 U27709 ( .A1(n56948), .A2(\pe3/got [17]), .ZN(n56555) );
  NAND2HSV2 U27710 ( .A1(n56173), .A2(\pe3/got [18]), .ZN(n56253) );
  XNOR2HSV1 U27711 ( .A1(n56253), .A2(n56252), .ZN(n56254) );
  XNOR2HSV4 U27712 ( .A1(n25460), .A2(n31868), .ZN(n31879) );
  CLKNAND2HSV2 U27713 ( .A1(n31958), .A2(n59022), .ZN(n25460) );
  NAND2HSV2 U27714 ( .A1(n56952), .A2(n56675), .ZN(n56333) );
  NOR2HSV4 U27715 ( .A1(n48319), .A2(n48316), .ZN(n48317) );
  CLKNAND2HSV2 U27716 ( .A1(n45113), .A2(n25461), .ZN(n45115) );
  CLKNHSV2 U27717 ( .I(n25462), .ZN(n25461) );
  CLKNAND2HSV2 U27718 ( .A1(n45112), .A2(n59979), .ZN(n25462) );
  AOI21HSV4 U27719 ( .A1(n32643), .A2(n32440), .B(n32439), .ZN(n32441) );
  BUFHSV6 U27720 ( .I(n33096), .Z(n33808) );
  INHSV4 U27721 ( .I(n33090), .ZN(n33096) );
  DELHS1 U27722 ( .I(\pe6/got [32]), .Z(n25463) );
  CLKNAND2HSV2 U27723 ( .A1(n26726), .A2(n25464), .ZN(n26725) );
  CLKNHSV2 U27724 ( .I(n27087), .ZN(n25464) );
  CLKNAND2HSV2 U27725 ( .A1(n52176), .A2(n44711), .ZN(n27087) );
  NAND2HSV2 U27726 ( .A1(n32162), .A2(n32161), .ZN(n32320) );
  CLKNAND2HSV2 U27727 ( .A1(n25553), .A2(n25552), .ZN(n25551) );
  CLKNAND2HSV2 U27728 ( .A1(n36785), .A2(n29750), .ZN(n36786) );
  CLKAND2HSV4 U27729 ( .A1(n41837), .A2(n41836), .Z(n41838) );
  NOR2HSV4 U27730 ( .A1(n26761), .A2(n35587), .ZN(n50315) );
  NAND3HSV4 U27731 ( .A1(n31291), .A2(n31292), .A3(n31290), .ZN(n31293) );
  CLKNAND2HSV4 U27732 ( .A1(n31294), .A2(n31293), .ZN(n31382) );
  NOR2HSV4 U27733 ( .A1(n39869), .A2(n25465), .ZN(n40137) );
  NOR2HSV4 U27734 ( .A1(n25467), .A2(n25466), .ZN(n25465) );
  CLKNAND2HSV2 U27735 ( .A1(n39568), .A2(n39567), .ZN(n25466) );
  CLKNHSV2 U27736 ( .I(n39872), .ZN(n25467) );
  INHSV2 U27737 ( .I(n25468), .ZN(n43350) );
  NAND2HSV2 U27738 ( .A1(n25891), .A2(n45625), .ZN(n25468) );
  XOR2HSV4 U27739 ( .A1(n32056), .A2(n32146), .Z(n52765) );
  CLKNAND2HSV2 U27740 ( .A1(n53097), .A2(n26651), .ZN(n25469) );
  INHSV2 U27741 ( .I(n25470), .ZN(n29646) );
  NAND2HSV0 U27742 ( .A1(n32035), .A2(n32047), .ZN(n25470) );
  CLKNAND2HSV2 U27743 ( .A1(n25471), .A2(n44678), .ZN(n26063) );
  NOR2HSV4 U27744 ( .A1(n48895), .A2(n44679), .ZN(n25471) );
  BUFHSV8 U27745 ( .I(n45942), .Z(n56910) );
  CLKNAND2HSV4 U27746 ( .A1(n26344), .A2(n45779), .ZN(n43595) );
  NAND2HSV2 U27747 ( .A1(n59580), .A2(n30596), .ZN(n47384) );
  NAND3HSV4 U27748 ( .A1(n25473), .A2(n45592), .A3(n45589), .ZN(n25472) );
  NOR2HSV4 U27749 ( .A1(n45595), .A2(n25474), .ZN(n25473) );
  CLKNHSV2 U27750 ( .I(n45591), .ZN(n25474) );
  XNOR2HSV4 U27751 ( .A1(n56773), .A2(n25476), .ZN(n25475) );
  XOR2HSV2 U27752 ( .A1(n56769), .A2(n56770), .Z(n25476) );
  INHSV4 U27753 ( .I(n42617), .ZN(n25477) );
  OAI21HSV2 U27754 ( .A1(n32942), .A2(n32941), .B(n32940), .ZN(n32943) );
  NOR2HSV4 U27755 ( .A1(n37770), .A2(n25478), .ZN(n39404) );
  CLKNAND2HSV2 U27756 ( .A1(n29711), .A2(n37765), .ZN(n37769) );
  NOR2HSV2 U27757 ( .A1(n53376), .A2(n53377), .ZN(n42595) );
  CLKNAND2HSV2 U27758 ( .A1(n41923), .A2(n25900), .ZN(pov1[23]) );
  NAND3HSV4 U27759 ( .A1(n42784), .A2(n25479), .A3(n42785), .ZN(n42926) );
  NOR2HSV4 U27760 ( .A1(n25815), .A2(n42791), .ZN(n25479) );
  INHSV6 U27761 ( .I(n41421), .ZN(n41239) );
  CLKNAND2HSV4 U27762 ( .A1(n47772), .A2(n26596), .ZN(n26742) );
  CLKAND2HSV4 U27763 ( .A1(n39880), .A2(\pe5/got [27]), .Z(n40127) );
  NOR2HSV2 U27764 ( .A1(n47784), .A2(n47783), .ZN(n25553) );
  XNOR2HSV4 U27765 ( .A1(n50487), .A2(n50486), .ZN(n50489) );
  NAND2HSV4 U27766 ( .A1(n40639), .A2(n46609), .ZN(n40640) );
  XNOR2HSV4 U27767 ( .A1(n52557), .A2(n52556), .ZN(n52561) );
  BUFHSV6 U27768 ( .I(n48165), .Z(n51016) );
  CLKNAND2HSV4 U27769 ( .A1(n25709), .A2(n38782), .ZN(n28544) );
  NAND2HSV2 U27770 ( .A1(n28544), .A2(n28543), .ZN(n28545) );
  CLKNAND2HSV2 U27771 ( .A1(n39699), .A2(n39698), .ZN(n59423) );
  XNOR2HSV4 U27772 ( .A1(n36423), .A2(n36422), .ZN(n36424) );
  XNOR2HSV4 U27773 ( .A1(n39365), .A2(n39228), .ZN(n39416) );
  CLKXOR2HSV4 U27774 ( .A1(n40418), .A2(n40417), .Z(n40421) );
  OAI21HSV2 U27775 ( .A1(n28510), .A2(n28511), .B(n28512), .ZN(n28513) );
  NAND2HSV2 U27776 ( .A1(n28514), .A2(n28513), .ZN(n28515) );
  AOI21HSV4 U27777 ( .A1(n29661), .A2(n25904), .B(n39719), .ZN(n39720) );
  XNOR2HSV4 U27778 ( .A1(n25481), .A2(n25480), .ZN(\pe6/poht [20]) );
  CLKNAND2HSV2 U27779 ( .A1(n58655), .A2(n59180), .ZN(n25480) );
  XNOR2HSV4 U27780 ( .A1(n58573), .A2(n58574), .ZN(n25481) );
  XNOR2HSV4 U27781 ( .A1(n51267), .A2(n51266), .ZN(n51269) );
  NAND3HSV4 U27782 ( .A1(n25903), .A2(n26500), .A3(n25902), .ZN(n26499) );
  NAND2HSV4 U27783 ( .A1(n51150), .A2(n51151), .ZN(n52558) );
  CLKNAND2HSV4 U27784 ( .A1(n51445), .A2(n31817), .ZN(n25521) );
  NAND2HSV4 U27785 ( .A1(n30062), .A2(n30074), .ZN(n26203) );
  NAND3HSV3 U27786 ( .A1(n41840), .A2(n29767), .A3(n41839), .ZN(n25900) );
  OAI21HSV4 U27787 ( .A1(n33291), .A2(n33290), .B(n26044), .ZN(n25876) );
  NOR2HSV4 U27788 ( .A1(n26051), .A2(n26050), .ZN(n33291) );
  NOR2HSV2 U27789 ( .A1(n42320), .A2(n42191), .ZN(n42192) );
  CLKNHSV6 U27790 ( .I(n50211), .ZN(n58104) );
  XNOR2HSV4 U27791 ( .A1(n25482), .A2(n42783), .ZN(n42792) );
  XNOR2HSV4 U27792 ( .A1(n42782), .A2(n42781), .ZN(n25482) );
  NAND3HSV4 U27793 ( .A1(n25483), .A2(n32959), .A3(n32958), .ZN(n32960) );
  CLKNAND2HSV4 U27794 ( .A1(n32682), .A2(n32681), .ZN(n25483) );
  CLKNAND2HSV3 U27795 ( .A1(n32157), .A2(n32059), .ZN(n32407) );
  CLKNAND2HSV4 U27796 ( .A1(n32162), .A2(n32793), .ZN(n32157) );
  CLKNHSV3 U27797 ( .I(n32061), .ZN(n59034) );
  XNOR2HSV4 U27798 ( .A1(n25488), .A2(n25484), .ZN(n32310) );
  XNOR2HSV4 U27799 ( .A1(n25487), .A2(n25485), .ZN(n25484) );
  NOR2HSV4 U27800 ( .A1(n32061), .A2(n32241), .ZN(n25487) );
  CLKNAND2HSV2 U27801 ( .A1(n32407), .A2(n35705), .ZN(n25488) );
  CLKNHSV2 U27802 ( .I(n32130), .ZN(n32165) );
  XNOR2HSV4 U27803 ( .A1(n25490), .A2(n25489), .ZN(n32223) );
  CLKNAND2HSV2 U27804 ( .A1(n32306), .A2(n59022), .ZN(n25489) );
  OAI21HSV4 U27805 ( .A1(n51443), .A2(n36055), .B(n32134), .ZN(n32306) );
  XNOR2HSV4 U27806 ( .A1(n26587), .A2(n31759), .ZN(n51443) );
  XNOR2HSV4 U27807 ( .A1(n25494), .A2(n25491), .ZN(n25490) );
  XNOR2HSV4 U27808 ( .A1(n25493), .A2(n25492), .ZN(n25491) );
  XOR2HSV2 U27809 ( .A1(n32222), .A2(n32221), .Z(n25492) );
  CLKNAND2HSV2 U27810 ( .A1(n26109), .A2(n26110), .ZN(n25493) );
  NOR2HSV4 U27811 ( .A1(n32130), .A2(n25495), .ZN(n25494) );
  CLKNHSV2 U27812 ( .I(n49665), .ZN(n25495) );
  CLKNAND2HSV2 U27813 ( .A1(n25496), .A2(n32946), .ZN(n47952) );
  CLKNAND2HSV2 U27814 ( .A1(n25496), .A2(n32804), .ZN(n32805) );
  CLKNAND2HSV4 U27815 ( .A1(n32803), .A2(n32802), .ZN(n25496) );
  CLKNHSV3 U27816 ( .I(n30020), .ZN(n30023) );
  CLKNAND2HSV4 U27817 ( .A1(n30130), .A2(n30028), .ZN(n30020) );
  CLKNAND2HSV3 U27818 ( .A1(n25498), .A2(n25497), .ZN(n30130) );
  AOI21HSV4 U27819 ( .A1(n29993), .A2(n29992), .B(n29991), .ZN(n25497) );
  CLKNAND2HSV3 U27820 ( .A1(n29997), .A2(n29998), .ZN(n25498) );
  NOR2HSV0 U27821 ( .A1(n36969), .A2(n25499), .ZN(n36880) );
  OAI21HSV2 U27822 ( .A1(n25500), .A2(n36885), .B(n43608), .ZN(n25499) );
  CLKNAND2HSV3 U27823 ( .A1(n25501), .A2(n36874), .ZN(n25500) );
  NOR2HSV3 U27824 ( .A1(n25502), .A2(n36877), .ZN(n25501) );
  CLKNHSV4 U27825 ( .I(n36847), .ZN(n25502) );
  CLKNAND2HSV4 U27826 ( .A1(n60024), .A2(n36873), .ZN(n36969) );
  CLKNAND2HSV4 U27827 ( .A1(n25909), .A2(n36892), .ZN(n60024) );
  NAND3HSV4 U27828 ( .A1(n36871), .A2(n36872), .A3(n36870), .ZN(n36892) );
  CLKNAND2HSV3 U27829 ( .A1(n36868), .A2(n36869), .ZN(n25909) );
  CLKNAND2HSV3 U27830 ( .A1(n25918), .A2(n31879), .ZN(n25504) );
  AOI21HSV4 U27831 ( .A1(n31882), .A2(n25504), .B(n25503), .ZN(n25523) );
  AOI21HSV4 U27832 ( .A1(n31881), .A2(n25504), .B(n31880), .ZN(n25503) );
  CLKNHSV4 U27833 ( .I(n32316), .ZN(n25506) );
  BUFHSV8 U27834 ( .I(n25507), .Z(n25505) );
  NOR2HSV4 U27835 ( .A1(n25506), .A2(n25505), .ZN(n26517) );
  NOR2HSV4 U27836 ( .A1(n26175), .A2(n25505), .ZN(n32336) );
  CLKNAND2HSV2 U27837 ( .A1(n25508), .A2(n31638), .ZN(n48000) );
  NAND3HSV4 U27838 ( .A1(n25508), .A2(n31638), .A3(n31261), .ZN(n31743) );
  NAND3HSV4 U27839 ( .A1(n25508), .A2(n31638), .A3(n35908), .ZN(n31636) );
  OAI21HSV4 U27840 ( .A1(n26340), .A2(n26339), .B(n26338), .ZN(n25508) );
  NOR2HSV8 U27841 ( .A1(n26547), .A2(n38375), .ZN(n53388) );
  OAI21HSV4 U27842 ( .A1(n45145), .A2(n44831), .B(n25509), .ZN(n25596) );
  AOI21HSV4 U27843 ( .A1(n45408), .A2(n44709), .B(n25510), .ZN(n25509) );
  NOR2HSV4 U27844 ( .A1(n45277), .A2(n44831), .ZN(n25510) );
  NOR2HSV4 U27845 ( .A1(n53388), .A2(n45280), .ZN(n45408) );
  NAND3HSV4 U27846 ( .A1(n25511), .A2(n26243), .A3(n26241), .ZN(n45280) );
  CLKNAND2HSV4 U27847 ( .A1(n26408), .A2(n44830), .ZN(n45145) );
  CLKNHSV2 U27848 ( .I(n25512), .ZN(n25511) );
  CLKNAND2HSV2 U27849 ( .A1(n26240), .A2(n26239), .ZN(n25512) );
  CLKNAND2HSV4 U27850 ( .A1(n32666), .A2(n32665), .ZN(n32786) );
  CLKNAND2HSV2 U27851 ( .A1(n25513), .A2(n32787), .ZN(n32788) );
  CLKNAND2HSV2 U27852 ( .A1(n32666), .A2(n25514), .ZN(n25513) );
  CLKNHSV2 U27853 ( .I(n25515), .ZN(n25514) );
  CLKNAND2HSV2 U27854 ( .A1(n32665), .A2(n29725), .ZN(n25515) );
  CLKNHSV2 U27855 ( .I(n32786), .ZN(n32800) );
  CLKNAND2HSV4 U27856 ( .A1(n58369), .A2(n46163), .ZN(n46553) );
  CLKNHSV2 U27857 ( .I(n59536), .ZN(n43136) );
  NOR2HSV4 U27858 ( .A1(n59536), .A2(n43249), .ZN(n43253) );
  AOI21HSV4 U27859 ( .A1(n59536), .A2(n43261), .B(n43260), .ZN(n25694) );
  NAND3HSV4 U27860 ( .A1(n25516), .A2(n44341), .A3(n44340), .ZN(n44349) );
  NAND3HSV3 U27861 ( .A1(n25516), .A2(n44341), .A3(n36086), .ZN(n44691) );
  CLKNAND2HSV4 U27862 ( .A1(n36079), .A2(n36078), .ZN(n25516) );
  XNOR2HSV4 U27863 ( .A1(n27429), .A2(n25517), .ZN(n27430) );
  CLKNAND2HSV2 U27864 ( .A1(n52910), .A2(\pe2/got [10]), .ZN(n25517) );
  CLKNAND2HSV2 U27865 ( .A1(n29589), .A2(n29588), .ZN(n29590) );
  XOR3HSV2 U27866 ( .A1(n54359), .A2(n25520), .A3(n25518), .Z(n29588) );
  CLKNHSV2 U27867 ( .I(n25519), .ZN(n25518) );
  CLKNAND2HSV2 U27868 ( .A1(n59521), .A2(n54716), .ZN(n25519) );
  CLKNHSV2 U27869 ( .I(n54360), .ZN(n25520) );
  OAI21HSV4 U27870 ( .A1(n32162), .A2(n32163), .B(n32055), .ZN(n32056) );
  XNOR2HSV4 U27871 ( .A1(n32033), .A2(n32035), .ZN(n32162) );
  XNOR2HSV4 U27872 ( .A1(n25523), .A2(n25522), .ZN(n32035) );
  CLKNAND2HSV2 U27873 ( .A1(n31891), .A2(n31892), .ZN(n25522) );
  CLKNAND2HSV4 U27874 ( .A1(\pe3/ti_1 ), .A2(\pe3/got [32]), .ZN(n25794) );
  XNOR2HSV4 U27875 ( .A1(n25533), .A2(n25524), .ZN(n30197) );
  NAND3HSV4 U27876 ( .A1(n25528), .A2(n25525), .A3(n29712), .ZN(n25524) );
  CLKNAND2HSV2 U27877 ( .A1(n25526), .A2(n30191), .ZN(n25525) );
  NOR2HSV0 U27878 ( .A1(n25527), .A2(n30192), .ZN(n25526) );
  CLKNAND2HSV2 U27879 ( .A1(n30195), .A2(n25529), .ZN(n25528) );
  CLKNAND2HSV2 U27880 ( .A1(n25530), .A2(n30185), .ZN(n25529) );
  AOI21HSV1 U27881 ( .A1(n30182), .A2(n25532), .B(n25531), .ZN(n25530) );
  CLKNHSV2 U27882 ( .I(n30186), .ZN(n25531) );
  CLKNHSV2 U27883 ( .I(n30187), .ZN(n25532) );
  CLKNAND2HSV2 U27884 ( .A1(n30099), .A2(n25535), .ZN(n25534) );
  CLKNHSV2 U27885 ( .I(n40142), .ZN(n25535) );
  CLKNAND2HSV2 U27886 ( .A1(n30099), .A2(n26422), .ZN(n25537) );
  OAI21HSV2 U27887 ( .A1(n37864), .A2(n53094), .B(n39007), .ZN(n37989) );
  XNOR2HSV4 U27888 ( .A1(n25539), .A2(n25538), .ZN(n37864) );
  XOR3HSV2 U27889 ( .A1(n37831), .A2(n37830), .A3(n37829), .Z(n25538) );
  OAI21HSV4 U27890 ( .A1(n37790), .A2(n37789), .B(n53092), .ZN(n25539) );
  XNOR2HSV4 U27891 ( .A1(n30565), .A2(n25540), .ZN(n30566) );
  XOR2HSV2 U27892 ( .A1(n30564), .A2(n25541), .Z(n25540) );
  XNOR2HSV4 U27893 ( .A1(n25544), .A2(n25542), .ZN(n25541) );
  XNOR2HSV4 U27894 ( .A1(n30563), .A2(n25543), .ZN(n25542) );
  XOR2HSV2 U27895 ( .A1(n30561), .A2(n30562), .Z(n25543) );
  CLKNAND2HSV2 U27896 ( .A1(n30734), .A2(n30685), .ZN(n25544) );
  XOR2HSV4 U27897 ( .A1(n37001), .A2(n25545), .Z(n25751) );
  CLKNAND2HSV3 U27898 ( .A1(\pe3/bq[31] ), .A2(\pe3/aot [32]), .ZN(n25545) );
  NAND2HSV2 U27899 ( .A1(\pe3/bq[32] ), .A2(\pe3/aot [31]), .ZN(n37001) );
  CLKNAND2HSV2 U27900 ( .A1(n47787), .A2(n25546), .ZN(n26635) );
  CLKNHSV2 U27901 ( .I(n47785), .ZN(n25546) );
  AOI21HSV4 U27902 ( .A1(n25555), .A2(n25554), .B(n25547), .ZN(n47785) );
  CLKNAND2HSV2 U27903 ( .A1(n25551), .A2(n25548), .ZN(n25547) );
  CLKNAND2HSV2 U27904 ( .A1(n25550), .A2(n25549), .ZN(n25548) );
  CLKNHSV2 U27905 ( .I(n47778), .ZN(n25549) );
  CLKNHSV2 U27906 ( .I(n47779), .ZN(n25550) );
  CLKNHSV2 U27907 ( .I(n26596), .ZN(n25552) );
  CLKNHSV2 U27908 ( .I(n47780), .ZN(n25554) );
  INAND2HSV4 U27909 ( .A1(n52847), .B1(n35011), .ZN(n47787) );
  XNOR2HSV4 U27910 ( .A1(n25557), .A2(n25556), .ZN(n52847) );
  CLKNAND2HSV2 U27911 ( .A1(n29359), .A2(n26853), .ZN(n25556) );
  CLKNAND2HSV2 U27912 ( .A1(n32232), .A2(n44519), .ZN(n32154) );
  CLKNAND2HSV2 U27913 ( .A1(n25561), .A2(n25558), .ZN(n32232) );
  NAND3HSV4 U27914 ( .A1(n25560), .A2(n25288), .A3(n25559), .ZN(n25558) );
  CLKNHSV2 U27915 ( .I(n32151), .ZN(n25559) );
  CLKNHSV2 U27916 ( .I(n32159), .ZN(n25560) );
  CLKNAND2HSV2 U27917 ( .A1(n32153), .A2(n32152), .ZN(n25561) );
  XNOR2HSV4 U27918 ( .A1(n32050), .A2(n32049), .ZN(n32153) );
  CLKNHSV1 U27919 ( .I(n29990), .ZN(n26148) );
  CLKNAND2HSV3 U27920 ( .A1(n30017), .A2(n30016), .ZN(n29889) );
  NOR2HSV4 U27921 ( .A1(n29820), .A2(n29819), .ZN(n30017) );
  AOI21HSV4 U27922 ( .A1(n29888), .A2(n25564), .B(n25563), .ZN(n25562) );
  CLKNHSV2 U27923 ( .I(n30139), .ZN(n25563) );
  NOR2HSV4 U27924 ( .A1(n29886), .A2(n30421), .ZN(n25564) );
  CLKNAND2HSV4 U27925 ( .A1(n29822), .A2(n29913), .ZN(n30016) );
  NOR2HSV8 U27926 ( .A1(n25566), .A2(n25565), .ZN(n32814) );
  CLKNAND2HSV4 U27927 ( .A1(n32230), .A2(n32229), .ZN(n25565) );
  CLKNHSV4 U27928 ( .I(n32351), .ZN(n25566) );
  XNOR2HSV4 U27929 ( .A1(n25568), .A2(n25567), .ZN(n32658) );
  NOR2HSV4 U27930 ( .A1(n32814), .A2(n31373), .ZN(n25567) );
  INAND2HSV4 U27931 ( .A1(n31971), .B1(n32833), .ZN(n25569) );
  INHSV24 U27932 ( .I(n25570), .ZN(n29774) );
  NOR2HSV4 U27933 ( .A1(n29774), .A2(n49922), .ZN(n47889) );
  CLKNAND2HSV2 U27934 ( .A1(n44661), .A2(n44525), .ZN(n26531) );
  CLKNAND2HSV2 U27935 ( .A1(n44657), .A2(n44656), .ZN(n44661) );
  CLKNAND2HSV2 U27936 ( .A1(n25576), .A2(n25580), .ZN(n44657) );
  NAND3HSV4 U27937 ( .A1(n44648), .A2(n44647), .A3(n53786), .ZN(n25574) );
  CLKNHSV2 U27938 ( .I(n55490), .ZN(n25575) );
  CLKNAND2HSV2 U27939 ( .A1(n25579), .A2(n25577), .ZN(n25576) );
  CLKNHSV2 U27940 ( .I(n48330), .ZN(n25577) );
  CLKNAND2HSV2 U27941 ( .A1(n45783), .A2(n25578), .ZN(n48330) );
  CLKNHSV2 U27942 ( .I(n45781), .ZN(n25578) );
  CLKNHSV2 U27943 ( .I(n45782), .ZN(n25579) );
  CLKNAND2HSV2 U27944 ( .A1(n25946), .A2(n25943), .ZN(n25580) );
  XNOR2HSV4 U27945 ( .A1(n43111), .A2(n43110), .ZN(n43114) );
  NAND3HSV2 U27946 ( .A1(n46817), .A2(n46766), .A3(n59031), .ZN(n28514) );
  INHSV2 U27947 ( .I(n37080), .ZN(n37084) );
  CLKNAND2HSV4 U27948 ( .A1(n40361), .A2(n26107), .ZN(n40424) );
  CLKNAND2HSV4 U27949 ( .A1(n31894), .A2(n44344), .ZN(n32041) );
  CLKNAND2HSV4 U27950 ( .A1(n32041), .A2(n31895), .ZN(n31967) );
  NOR2HSV4 U27951 ( .A1(n35583), .A2(n35587), .ZN(n35140) );
  OAI21HSV2 U27952 ( .A1(n28790), .A2(n28791), .B(n28792), .ZN(n28793) );
  INHSV4 U27953 ( .I(n35019), .ZN(n35463) );
  CLKNAND2HSV2 U27954 ( .A1(n58476), .A2(n58401), .ZN(n58349) );
  NOR2HSV8 U27955 ( .A1(n36799), .A2(n36940), .ZN(n25791) );
  CLKNHSV6 U27956 ( .I(n31898), .ZN(n31759) );
  NAND2HSV4 U27957 ( .A1(n26067), .A2(n59374), .ZN(n48449) );
  CLKXOR2HSV4 U27958 ( .A1(n37324), .A2(n37323), .Z(n37328) );
  CLKNAND2HSV4 U27959 ( .A1(n34231), .A2(n52821), .ZN(n47964) );
  INHSV2 U27960 ( .I(n47964), .ZN(n34232) );
  CLKNAND2HSV8 U27961 ( .A1(n40439), .A2(n40332), .ZN(n40362) );
  IOA22HSV4 U27962 ( .B1(n40362), .B2(n40569), .A1(n40969), .A2(\pe1/ti_7t [1]), .ZN(n41880) );
  CLKNAND2HSV4 U27963 ( .A1(n36732), .A2(n36729), .ZN(n36722) );
  CLKNAND2HSV4 U27964 ( .A1(n29737), .A2(n32348), .ZN(n31765) );
  NAND2HSV4 U27965 ( .A1(n31765), .A2(n31764), .ZN(n31874) );
  NAND2HSV4 U27966 ( .A1(n51443), .A2(n32133), .ZN(n32026) );
  NAND3HSV3 U27967 ( .A1(n46766), .A2(n53102), .A3(n49736), .ZN(n29205) );
  INHSV8 U27968 ( .I(n36718), .ZN(n36728) );
  OAI22HSV4 U27969 ( .A1(n33701), .A2(n33704), .B1(n34727), .B2(n33700), .ZN(
        n33763) );
  BUFHSV8 U27970 ( .I(\pe3/bq[31] ), .Z(n37186) );
  NAND2HSV2 U27971 ( .A1(n51726), .A2(n53093), .ZN(n28541) );
  XNOR2HSV4 U27972 ( .A1(n42312), .A2(n42311), .ZN(n42313) );
  INHSV4 U27973 ( .I(n36044), .ZN(n36043) );
  NAND2HSV4 U27974 ( .A1(n36042), .A2(n36043), .ZN(n36046) );
  CLKNAND2HSV2 U27975 ( .A1(n25860), .A2(n35808), .ZN(n35795) );
  CLKNAND2HSV2 U27976 ( .A1(n46133), .A2(\pe3/pvq [6]), .ZN(n36793) );
  BUFHSV8 U27977 ( .I(n42643), .Z(n43757) );
  CLKNAND2HSV4 U27978 ( .A1(n44662), .A2(n44663), .ZN(n40320) );
  INHSV2 U27979 ( .I(n35463), .ZN(n35469) );
  OAI21HSV4 U27980 ( .A1(n35469), .A2(n35468), .B(n35467), .ZN(n35474) );
  CLKNAND2HSV4 U27981 ( .A1(n49405), .A2(\pe3/got [29]), .ZN(n37079) );
  CLKNAND2HSV2 U27982 ( .A1(n58184), .A2(n58141), .ZN(n29148) );
  OAI21HSV2 U27983 ( .A1(n29147), .A2(n29148), .B(n29149), .ZN(n29150) );
  INHSV2 U27984 ( .I(n32157), .ZN(n32159) );
  NAND3HSV4 U27985 ( .A1(n36728), .A2(n36783), .A3(n36709), .ZN(n36693) );
  INHSV4 U27986 ( .I(n59607), .ZN(n36695) );
  AOI21HSV4 U27987 ( .A1(n25581), .A2(n25587), .B(n25586), .ZN(n31346) );
  CLKNHSV2 U27988 ( .I(n52704), .ZN(n25581) );
  OAI22HSV4 U27989 ( .A1(n52704), .A2(n25583), .B1(n25585), .B2(n25582), .ZN(
        n25584) );
  CLKNHSV2 U27990 ( .I(n25586), .ZN(n25582) );
  INAND2HSV4 U27991 ( .A1(n25585), .B1(n25587), .ZN(n25583) );
  AOI21HSV4 U27992 ( .A1(n31448), .A2(n31454), .B(n25584), .ZN(n31507) );
  CLKNHSV2 U27993 ( .I(n31449), .ZN(n25585) );
  CLKNHSV2 U27994 ( .I(n31690), .ZN(n25586) );
  CLKNHSV2 U27995 ( .I(n31345), .ZN(n25587) );
  CLKNAND2HSV2 U27996 ( .A1(n55705), .A2(n43898), .ZN(n43593) );
  CLKNAND2HSV2 U27997 ( .A1(n55705), .A2(n43234), .ZN(n45588) );
  CLKNHSV2 U27998 ( .I(n43222), .ZN(n43448) );
  XOR3HSV2 U27999 ( .A1(n25590), .A2(n25588), .A3(n43105), .Z(n43109) );
  XNOR2HSV4 U28000 ( .A1(n25589), .A2(n43104), .ZN(n25588) );
  CLKNAND2HSV2 U28001 ( .A1(n43755), .A2(n42770), .ZN(n25589) );
  INAND2HSV4 U28002 ( .A1(n42827), .B1(n59380), .ZN(n25590) );
  CLKNAND2HSV1 U28003 ( .A1(n25591), .A2(n31901), .ZN(n31897) );
  NOR2HSV2 U28004 ( .A1(n42506), .A2(n25592), .ZN(n42581) );
  INHSV1 U28005 ( .I(n37453), .ZN(n25592) );
  INAND2HSV2 U28006 ( .A1(n37451), .B1(n25593), .ZN(n37453) );
  INHSV4 U28007 ( .I(n42682), .ZN(n25593) );
  OAI21HSV4 U28008 ( .A1(n44165), .A2(n29330), .B(n44164), .ZN(n45101) );
  CLKNAND2HSV4 U28009 ( .A1(n44161), .A2(n44162), .ZN(n45102) );
  CLKNHSV2 U28010 ( .I(n44181), .ZN(n45114) );
  OAI21HSV4 U28011 ( .A1(n25596), .A2(n25595), .B(n25594), .ZN(n45132) );
  CLKNAND2HSV4 U28012 ( .A1(n35720), .A2(n25598), .ZN(n36053) );
  NAND2HSV4 U28013 ( .A1(n33088), .A2(n35717), .ZN(n25598) );
  CLKNHSV2 U28014 ( .I(n25598), .ZN(n25597) );
  CLKNAND2HSV3 U28015 ( .A1(n25649), .A2(n33075), .ZN(n25599) );
  CLKNAND2HSV4 U28016 ( .A1(n25600), .A2(n25907), .ZN(n26753) );
  CLKNAND2HSV3 U28017 ( .A1(n26779), .A2(n26777), .ZN(n25600) );
  OAI21HSV4 U28018 ( .A1(n26754), .A2(n25600), .B(n26753), .ZN(n60077) );
  NOR2HSV4 U28019 ( .A1(n35302), .A2(n25601), .ZN(n44690) );
  OAI21HSV4 U28020 ( .A1(n35301), .A2(n35313), .B(n35300), .ZN(n25601) );
  CLKNHSV2 U28021 ( .I(n25602), .ZN(n42807) );
  CLKNAND2HSV2 U28022 ( .A1(n43025), .A2(n42806), .ZN(n25602) );
  XNOR2HSV4 U28023 ( .A1(n42926), .A2(n42916), .ZN(n43025) );
  CLKNHSV2 U28024 ( .I(n38002), .ZN(n38017) );
  XNOR2HSV4 U28025 ( .A1(n25604), .A2(n25603), .ZN(n38002) );
  CLKNAND2HSV2 U28026 ( .A1(n26837), .A2(n37925), .ZN(n25603) );
  XNOR2HSV4 U28027 ( .A1(n37916), .A2(n37915), .ZN(n25604) );
  CLKNAND2HSV4 U28028 ( .A1(n25605), .A2(n35312), .ZN(n35310) );
  CLKNAND2HSV3 U28029 ( .A1(n35463), .A2(n35465), .ZN(n25605) );
  XNOR2HSV4 U28030 ( .A1(n37413), .A2(n25606), .ZN(n53377) );
  XNOR2HSV4 U28031 ( .A1(n37417), .A2(n25606), .ZN(n37433) );
  XNOR2HSV4 U28032 ( .A1(n25669), .A2(n37412), .ZN(n25606) );
  CLKNAND2HSV3 U28033 ( .A1(n31757), .A2(n31747), .ZN(n31752) );
  XNOR2HSV4 U28034 ( .A1(n25610), .A2(n25607), .ZN(n31757) );
  NOR2HSV4 U28035 ( .A1(n25609), .A2(n25608), .ZN(n25607) );
  NOR2HSV4 U28036 ( .A1(n31693), .A2(n31694), .ZN(n25608) );
  CLKNAND2HSV2 U28037 ( .A1(n26331), .A2(n31692), .ZN(n25609) );
  XNOR2HSV4 U28038 ( .A1(n25612), .A2(n25611), .ZN(n25610) );
  XNOR2HSV4 U28039 ( .A1(n31668), .A2(n31669), .ZN(n25611) );
  AOI21HSV4 U28040 ( .A1(n31675), .A2(n32822), .B(n31674), .ZN(n25612) );
  OAI21HSV4 U28041 ( .A1(n25614), .A2(n25613), .B(n33605), .ZN(n34458) );
  OAI21HSV2 U28042 ( .A1(n33699), .A2(n33597), .B(n33596), .ZN(n25613) );
  AOI21HSV4 U28043 ( .A1(n52757), .A2(n35021), .B(n33597), .ZN(n25614) );
  CLKNAND2HSV4 U28044 ( .A1(n25615), .A2(n25617), .ZN(n34867) );
  CLKNAND2HSV2 U28045 ( .A1(n60038), .A2(n25620), .ZN(n25615) );
  CLKBUFHSV2 U28046 ( .I(n34867), .Z(n25616) );
  CLKNAND2HSV0 U28047 ( .A1(n34867), .A2(\pe4/got [27]), .ZN(n33399) );
  CLKNAND2HSV2 U28048 ( .A1(n25619), .A2(n25618), .ZN(n25617) );
  CLKNHSV2 U28049 ( .I(n33340), .ZN(n25618) );
  CLKNHSV2 U28050 ( .I(n33848), .ZN(n25619) );
  CLKNHSV2 U28051 ( .I(n33339), .ZN(n25620) );
  CLKNHSV4 U28052 ( .I(n46074), .ZN(n25652) );
  INAND2HSV4 U28053 ( .A1(n25650), .B1(n45946), .ZN(n46074) );
  NOR2HSV4 U28054 ( .A1(n43913), .A2(n45941), .ZN(n45946) );
  CLKNHSV2 U28055 ( .I(n47846), .ZN(n47904) );
  OAI21HSV4 U28056 ( .A1(n35451), .A2(n25624), .B(n25621), .ZN(n35452) );
  AOI21HSV4 U28057 ( .A1(n25623), .A2(n25622), .B(n35450), .ZN(n25621) );
  NOR2HSV4 U28058 ( .A1(n35448), .A2(n34416), .ZN(n25622) );
  CLKNHSV2 U28059 ( .I(n35447), .ZN(n25623) );
  NAND3HSV4 U28060 ( .A1(n35024), .A2(n35022), .A3(n35023), .ZN(n35447) );
  CLKNAND2HSV2 U28061 ( .A1(n35446), .A2(n35445), .ZN(n25624) );
  NAND3HSV4 U28062 ( .A1(n47846), .A2(n35028), .A3(n35029), .ZN(n35284) );
  CLKNAND2HSV2 U28063 ( .A1(n35285), .A2(n35448), .ZN(n35451) );
  XNOR2HSV4 U28064 ( .A1(n35026), .A2(n35025), .ZN(n35448) );
  CLKNAND2HSV2 U28065 ( .A1(n25627), .A2(n25625), .ZN(n35285) );
  NOR2HSV4 U28066 ( .A1(n47846), .A2(n25626), .ZN(n25625) );
  CLKNHSV2 U28067 ( .I(n35028), .ZN(n25626) );
  CLKNHSV2 U28068 ( .I(n35440), .ZN(n25627) );
  CLKNHSV2 U28069 ( .I(n31424), .ZN(n25628) );
  INAND2HSV4 U28070 ( .A1(n31424), .B1(\pe6/got [28]), .ZN(n26452) );
  INAND2HSV4 U28071 ( .A1(n25629), .B1(\pe6/got [27]), .ZN(n31485) );
  INAND2HSV4 U28072 ( .A1(n31269), .B1(\pe6/got [21]), .ZN(n31788) );
  CLKNAND2HSV2 U28073 ( .A1(n46818), .A2(n25630), .ZN(n31848) );
  CLKNAND2HSV2 U28074 ( .A1(n53101), .A2(n25630), .ZN(n31993) );
  CLKNHSV2 U28075 ( .I(n25629), .ZN(n25630) );
  CLKNHSV8 U28076 ( .I(\pe4/got [32]), .ZN(n33184) );
  CLKNAND2HSV3 U28077 ( .A1(n60001), .A2(n45779), .ZN(n25631) );
  CLKNAND2HSV4 U28078 ( .A1(n25631), .A2(n47429), .ZN(n56260) );
  CLKNHSV2 U28079 ( .I(n55820), .ZN(n53279) );
  XNOR2HSV4 U28080 ( .A1(n25638), .A2(n25632), .ZN(n46439) );
  XNOR2HSV4 U28081 ( .A1(n25634), .A2(n25633), .ZN(n25632) );
  NOR2HSV4 U28082 ( .A1(n47496), .A2(n46438), .ZN(n25633) );
  XNOR2HSV4 U28083 ( .A1(n25637), .A2(n25635), .ZN(n25634) );
  XNOR2HSV4 U28084 ( .A1(n46436), .A2(n25636), .ZN(n25635) );
  CLKNHSV2 U28085 ( .I(n46437), .ZN(n25636) );
  CLKNAND2HSV2 U28086 ( .A1(n48480), .A2(n59963), .ZN(n25637) );
  CLKNAND2HSV2 U28087 ( .A1(n56260), .A2(n42815), .ZN(n25638) );
  OAI21HSV4 U28088 ( .A1(n25639), .A2(n44672), .B(n44671), .ZN(n48894) );
  CLKNHSV2 U28089 ( .I(n25640), .ZN(n29358) );
  CLKNAND2HSV2 U28090 ( .A1(n25642), .A2(n25640), .ZN(n26853) );
  NOR2HSV4 U28091 ( .A1(n44690), .A2(n25641), .ZN(n25640) );
  CLKNHSV2 U28092 ( .I(n59956), .ZN(n25641) );
  CLKNHSV2 U28093 ( .I(n29357), .ZN(n25642) );
  CLKNAND2HSV2 U28094 ( .A1(n59666), .A2(n33461), .ZN(n25643) );
  CLKNAND2HSV2 U28095 ( .A1(n25646), .A2(n25645), .ZN(n25644) );
  CLKNHSV2 U28096 ( .I(n29355), .ZN(n25645) );
  CLKNHSV2 U28097 ( .I(n29354), .ZN(n25646) );
  NAND3HSV4 U28098 ( .A1(n43909), .A2(n25647), .A3(n44674), .ZN(n43911) );
  CLKNHSV2 U28099 ( .I(n25647), .ZN(n26398) );
  CLKNHSV2 U28100 ( .I(n51451), .ZN(n25649) );
  CLKNAND2HSV3 U28101 ( .A1(n33072), .A2(n25648), .ZN(n33073) );
  CLKNAND2HSV2 U28102 ( .A1(n46075), .A2(n46074), .ZN(n46077) );
  CLKNHSV2 U28103 ( .I(n43371), .ZN(n25650) );
  NOR2HSV4 U28104 ( .A1(n26221), .A2(n26222), .ZN(n44677) );
  CLKNAND2HSV4 U28105 ( .A1(n35788), .A2(n32967), .ZN(n46588) );
  CLKNAND2HSV3 U28106 ( .A1(n32806), .A2(n32805), .ZN(n35788) );
  NOR2HSV2 U28107 ( .A1(n46588), .A2(n33063), .ZN(n33076) );
  CLKNAND2HSV2 U28108 ( .A1(n45630), .A2(n25651), .ZN(n26071) );
  CLKNAND2HSV3 U28109 ( .A1(n45945), .A2(n45944), .ZN(n45943) );
  AOI21HSV4 U28110 ( .A1(n26259), .A2(n48894), .B(n25653), .ZN(n45945) );
  XNOR2HSV4 U28111 ( .A1(n46070), .A2(n46069), .ZN(n46076) );
  NOR2HSV4 U28112 ( .A1(n45946), .A2(n43873), .ZN(n46072) );
  NOR2HSV4 U28113 ( .A1(n25655), .A2(n25654), .ZN(n25653) );
  CLKNHSV2 U28114 ( .I(\pe3/ti_7t [27]), .ZN(n25654) );
  CLKNHSV2 U28115 ( .I(n36967), .ZN(n25655) );
  CLKNAND2HSV2 U28116 ( .A1(n45942), .A2(n25656), .ZN(n45754) );
  NOR2HSV1 U28117 ( .A1(n44665), .A2(n44679), .ZN(n25656) );
  CLKNHSV2 U28118 ( .I(n43911), .ZN(n45942) );
  CLKBUFHSV2 U28119 ( .I(n25658), .Z(n25657) );
  BUFHSV8 U28120 ( .I(n25659), .Z(n25658) );
  INAND2HSV2 U28121 ( .A1(n49400), .B1(n46289), .ZN(n46290) );
  CLKNAND2HSV2 U28122 ( .A1(n25658), .A2(n32596), .ZN(n46889) );
  CLKNAND2HSV2 U28123 ( .A1(n25658), .A2(n59178), .ZN(n49908) );
  CLKNAND2HSV2 U28124 ( .A1(n25658), .A2(n59175), .ZN(n58922) );
  CLKNAND2HSV2 U28125 ( .A1(n25657), .A2(n59173), .ZN(n27460) );
  CLKNAND2HSV2 U28126 ( .A1(n25657), .A2(n59182), .ZN(n27609) );
  CLKNAND2HSV2 U28127 ( .A1(n25657), .A2(n58401), .ZN(n28746) );
  CLKNAND2HSV2 U28128 ( .A1(n25657), .A2(n36029), .ZN(n46578) );
  CLKNHSV4 U28129 ( .I(n49400), .ZN(n25659) );
  XNOR2HSV4 U28130 ( .A1(n25663), .A2(n25660), .ZN(n36224) );
  XNOR2HSV4 U28131 ( .A1(n35906), .A2(n35905), .ZN(n25661) );
  CLKNAND2HSV2 U28132 ( .A1(n59487), .A2(n59022), .ZN(n25662) );
  CLKNAND2HSV2 U28133 ( .A1(n36206), .A2(n36207), .ZN(n59487) );
  CLKNAND2HSV2 U28134 ( .A1(n36218), .A2(n25664), .ZN(n25663) );
  CLKNHSV2 U28135 ( .I(n25665), .ZN(n25664) );
  CLKNAND2HSV2 U28136 ( .A1(n36216), .A2(n35916), .ZN(n25665) );
  CLKNAND2HSV2 U28137 ( .A1(n35915), .A2(n35914), .ZN(n36216) );
  CLKNAND2HSV0 U28138 ( .A1(n35913), .A2(n35912), .ZN(n25666) );
  CLKNAND2HSV2 U28139 ( .A1(n35911), .A2(n35910), .ZN(n25667) );
  INHSV2 U28140 ( .I(n25668), .ZN(n37870) );
  CLKNAND2HSV3 U28141 ( .A1(n25668), .A2(n38025), .ZN(n37991) );
  CLKNHSV2 U28142 ( .I(n37411), .ZN(n25669) );
  XNOR2HSV4 U28143 ( .A1(n37258), .A2(n37257), .ZN(n25670) );
  CLKNHSV2 U28144 ( .I(n25670), .ZN(n52752) );
  CLKNAND2HSV3 U28145 ( .A1(n58369), .A2(n26603), .ZN(n26602) );
  CLKNAND2HSV3 U28146 ( .A1(n46157), .A2(n46552), .ZN(n25715) );
  NOR2HSV4 U28147 ( .A1(n58437), .A2(n58435), .ZN(n25672) );
  CLKNAND2HSV4 U28148 ( .A1(n25672), .A2(n48889), .ZN(n29765) );
  INHSV2 U28149 ( .I(n25973), .ZN(n25678) );
  CLKNAND2HSV4 U28150 ( .A1(n25673), .A2(n37157), .ZN(n37148) );
  NAND3HSV4 U28151 ( .A1(n25675), .A2(n25967), .A3(n25674), .ZN(n25673) );
  CLKNHSV2 U28152 ( .I(n25676), .ZN(n25674) );
  CLKNAND2HSV2 U28153 ( .A1(n25678), .A2(n25677), .ZN(n25675) );
  CLKNHSV2 U28154 ( .I(n37146), .ZN(n25676) );
  CLKNHSV2 U28155 ( .I(n25975), .ZN(n25677) );
  NOR2HSV4 U28156 ( .A1(n37150), .A2(n37246), .ZN(n25679) );
  CLKNAND2HSV4 U28157 ( .A1(n25679), .A2(n37154), .ZN(n25882) );
  CLKNAND2HSV3 U28158 ( .A1(n60030), .A2(n25680), .ZN(n26279) );
  NOR2HSV4 U28159 ( .A1(n35008), .A2(n35010), .ZN(n25680) );
  XNOR2HSV4 U28160 ( .A1(n34982), .A2(n35016), .ZN(n60030) );
  CLKNAND2HSV2 U28161 ( .A1(n35161), .A2(n35160), .ZN(n35306) );
  AOI21HSV4 U28162 ( .A1(n35008), .A2(n35015), .B(n50301), .ZN(n35160) );
  CLKNAND2HSV2 U28163 ( .A1(n25682), .A2(n35018), .ZN(n35161) );
  AOI21HSV4 U28164 ( .A1(n35014), .A2(n35013), .B(n35012), .ZN(n35154) );
  NOR2HSV4 U28165 ( .A1(n60030), .A2(n25681), .ZN(n35157) );
  CLKNAND2HSV2 U28166 ( .A1(n35014), .A2(n35021), .ZN(n25681) );
  CLKNHSV4 U28167 ( .I(n35003), .ZN(n50301) );
  CLKNAND2HSV4 U28168 ( .A1(n35008), .A2(n35283), .ZN(n25682) );
  XNOR2HSV4 U28169 ( .A1(n35006), .A2(n35005), .ZN(n35014) );
  OAI21HSV4 U28170 ( .A1(n60051), .A2(n38529), .B(n27095), .ZN(n25956) );
  XNOR2HSV4 U28171 ( .A1(n25683), .A2(n44303), .ZN(n60051) );
  XNOR2HSV4 U28172 ( .A1(n44039), .A2(n44040), .ZN(n44303) );
  XNOR2HSV4 U28173 ( .A1(n44038), .A2(n44037), .ZN(n44040) );
  OAI21HSV4 U28174 ( .A1(n44148), .A2(n43922), .B(n43921), .ZN(n44039) );
  CLKNAND2HSV2 U28175 ( .A1(n29686), .A2(n44302), .ZN(n25684) );
  OAI21HSV4 U28176 ( .A1(n44299), .A2(n44298), .B(n44297), .ZN(n25685) );
  CLKNHSV2 U28177 ( .I(n25686), .ZN(n44673) );
  CLKNAND2HSV2 U28178 ( .A1(n44668), .A2(n43896), .ZN(n25686) );
  XOR2HSV2 U28179 ( .A1(n45748), .A2(n25687), .Z(n45749) );
  XNOR2HSV4 U28180 ( .A1(n25690), .A2(n25688), .ZN(n25687) );
  NOR2HSV4 U28181 ( .A1(n48484), .A2(n25689), .ZN(n25688) );
  CLKNHSV2 U28182 ( .I(n45947), .ZN(n25689) );
  XOR2HSV2 U28183 ( .A1(n25691), .A2(n45747), .Z(n25690) );
  CLKNAND2HSV2 U28184 ( .A1(n48486), .A2(n45634), .ZN(n25691) );
  CLKNAND2HSV2 U28185 ( .A1(n43256), .A2(n43355), .ZN(n25695) );
  XNOR2HSV4 U28186 ( .A1(n25697), .A2(n25696), .ZN(n43256) );
  CLKNAND2HSV2 U28187 ( .A1(n60012), .A2(n44309), .ZN(n25698) );
  CLKNAND2HSV2 U28188 ( .A1(n25702), .A2(n25699), .ZN(n60012) );
  CLKNAND2HSV2 U28189 ( .A1(n45142), .A2(n25700), .ZN(n25699) );
  CLKNHSV2 U28190 ( .I(n25701), .ZN(n25700) );
  CLKNAND2HSV2 U28191 ( .A1(n45143), .A2(n45141), .ZN(n25701) );
  NAND3HSV4 U28192 ( .A1(n25703), .A2(n45266), .A3(n45139), .ZN(n25702) );
  CLKNHSV2 U28193 ( .I(n45264), .ZN(n25703) );
  XNOR2HSV4 U28194 ( .A1(n25707), .A2(n25706), .ZN(n25704) );
  XOR2HSV2 U28195 ( .A1(n25708), .A2(\pe3/phq [7]), .Z(n25705) );
  CLKNAND2HSV3 U28196 ( .A1(n46133), .A2(\pe3/pvq [7]), .ZN(n25706) );
  CLKNAND2HSV4 U28197 ( .A1(n42634), .A2(n59609), .ZN(n25708) );
  CLKNAND2HSV2 U28198 ( .A1(\pe3/aot [31]), .A2(\pe3/bq[31] ), .ZN(n36674) );
  CLKNAND2HSV2 U28199 ( .A1(n25709), .A2(n52922), .ZN(n25710) );
  XNOR2HSV4 U28200 ( .A1(n48160), .A2(n25712), .ZN(n25711) );
  CLKNHSV2 U28201 ( .I(n25713), .ZN(n25712) );
  NOR2HSV4 U28202 ( .A1(n51727), .A2(n25714), .ZN(n25713) );
  CLKNHSV2 U28203 ( .I(n59685), .ZN(n25714) );
  CLKNAND2HSV4 U28204 ( .A1(n59571), .A2(n43247), .ZN(n43255) );
  CLKNAND2HSV0 U28205 ( .A1(n26600), .A2(n25715), .ZN(n46300) );
  OAI21HSV4 U28206 ( .A1(n25717), .A2(n38198), .B(n25716), .ZN(n26717) );
  NOR2HSV4 U28207 ( .A1(n47981), .A2(n38180), .ZN(n25716) );
  XNOR2HSV4 U28208 ( .A1(n38175), .A2(n38174), .ZN(n47981) );
  XNOR2HSV4 U28209 ( .A1(n38103), .A2(n38102), .ZN(n38174) );
  OAI22HSV4 U28210 ( .A1(n38040), .A2(n38039), .B1(n38104), .B2(n38038), .ZN(
        n38175) );
  NOR2HSV4 U28211 ( .A1(n26718), .A2(n38109), .ZN(n38198) );
  CLKNAND2HSV2 U28212 ( .A1(n25850), .A2(n38199), .ZN(n25717) );
  CLKNAND2HSV2 U28213 ( .A1(n38012), .A2(n38109), .ZN(n25850) );
  CLKBUFHSV2 U28214 ( .I(n36861), .Z(n25718) );
  CLKNAND2HSV1 U28215 ( .A1(n25719), .A2(n36864), .ZN(n36738) );
  XNOR2HSV4 U28216 ( .A1(n52728), .A2(n25718), .ZN(n60091) );
  CLKNHSV2 U28217 ( .I(n25968), .ZN(n25974) );
  INAND2HSV4 U28218 ( .A1(n37040), .B1(n37340), .ZN(n25968) );
  CLKNAND2HSV3 U28219 ( .A1(n25720), .A2(n33201), .ZN(n33199) );
  CLKNAND2HSV3 U28220 ( .A1(n33129), .A2(n33128), .ZN(n25720) );
  CLKNAND2HSV2 U28221 ( .A1(n25720), .A2(n34571), .ZN(n26050) );
  CLKNAND2HSV2 U28222 ( .A1(n33198), .A2(n25720), .ZN(n59578) );
  INHSV2 U28223 ( .I(n25721), .ZN(n38354) );
  OAI21HSV4 U28224 ( .A1(n52749), .A2(n37930), .B(n25722), .ZN(n25723) );
  AOI21HSV4 U28225 ( .A1(n26089), .A2(n38112), .B(n26088), .ZN(n25722) );
  CLKNAND2HSV3 U28226 ( .A1(n26723), .A2(n26722), .ZN(n25724) );
  CLKNAND2HSV2 U28227 ( .A1(n25724), .A2(n25723), .ZN(n38355) );
  NOR2HSV4 U28228 ( .A1(n25724), .A2(n25723), .ZN(n25721) );
  CLKNAND2HSV4 U28229 ( .A1(n25725), .A2(n35153), .ZN(n33851) );
  CLKNHSV8 U28230 ( .I(n33795), .ZN(n25725) );
  XNOR2HSV4 U28231 ( .A1(n25785), .A2(n25781), .ZN(n25726) );
  CLKNAND2HSV2 U28232 ( .A1(n25726), .A2(n36714), .ZN(n36715) );
  XNOR2HSV4 U28233 ( .A1(n33557), .A2(n25727), .ZN(n33558) );
  XNOR2HSV4 U28234 ( .A1(n25729), .A2(n25728), .ZN(n25727) );
  XNOR2HSV4 U28235 ( .A1(n33545), .A2(n33555), .ZN(n25728) );
  XNOR2HSV4 U28236 ( .A1(n25731), .A2(n25730), .ZN(n25729) );
  CLKNAND2HSV2 U28237 ( .A1(n34285), .A2(n59369), .ZN(n25730) );
  CLKNAND2HSV2 U28238 ( .A1(n33735), .A2(\pe4/got [22]), .ZN(n25731) );
  CLKBUFHSV2 U28239 ( .I(n25733), .Z(n25732) );
  INHSV2 U28240 ( .I(n37020), .ZN(n25733) );
  CLKNAND2HSV2 U28241 ( .A1(n25733), .A2(n36788), .ZN(n36769) );
  CLKNAND2HSV2 U28242 ( .A1(n25732), .A2(n42508), .ZN(n37138) );
  CLKNAND2HSV2 U28243 ( .A1(n25732), .A2(n56335), .ZN(n42758) );
  CLKNAND2HSV2 U28244 ( .A1(n25732), .A2(\pe3/got [13]), .ZN(n43314) );
  CLKNAND2HSV3 U28245 ( .A1(n25736), .A2(n25735), .ZN(n25734) );
  CLKNHSV8 U28246 ( .I(\pe4/phq [2]), .ZN(n25735) );
  CLKNAND2HSV4 U28247 ( .A1(\pe4/got [31]), .A2(\pe4/ti_1 ), .ZN(n25736) );
  OAI21HSV4 U28248 ( .A1(n25736), .A2(n25735), .B(n25734), .ZN(n26629) );
  INHSV2 U28249 ( .I(n25740), .ZN(n25737) );
  MUX2NHSV4 U28250 ( .I0(\pe4/phq [5]), .I1(n28422), .S(n28423), .ZN(n25747)
         );
  CLKNAND2HSV2 U28251 ( .A1(n25739), .A2(n25738), .ZN(n25748) );
  IOA21HSV4 U28252 ( .A1(n33326), .A2(n57106), .B(n25737), .ZN(n25738) );
  NAND3HSV4 U28253 ( .A1(n25740), .A2(n33326), .A3(n57106), .ZN(n25739) );
  CLKNAND2HSV2 U28254 ( .A1(n59485), .A2(n33248), .ZN(n25740) );
  XOR3HSV2 U28255 ( .A1(n25748), .A2(n25745), .A3(n25741), .Z(n26645) );
  XOR2HSV2 U28256 ( .A1(n33174), .A2(n25742), .Z(n25741) );
  XNOR2HSV4 U28257 ( .A1(n25744), .A2(n25743), .ZN(n25742) );
  NOR2HSV4 U28258 ( .A1(n46618), .A2(n33564), .ZN(n25743) );
  CLKNAND2HSV2 U28259 ( .A1(n33420), .A2(\pe4/bq[31] ), .ZN(n25744) );
  XNOR2HSV4 U28260 ( .A1(n25747), .A2(n25746), .ZN(n25745) );
  CLKNAND2HSV2 U28261 ( .A1(n57254), .A2(n59523), .ZN(n25746) );
  XNOR2HSV4 U28262 ( .A1(n28198), .A2(n25749), .ZN(n28199) );
  CLKNAND2HSV2 U28263 ( .A1(n52047), .A2(n52276), .ZN(n25749) );
  CLKNAND2HSV4 U28264 ( .A1(n25750), .A2(n36972), .ZN(n36930) );
  XOR3HSV2 U28265 ( .A1(n25753), .A2(n25752), .A3(n25751), .Z(n26016) );
  AOI21HSV4 U28266 ( .A1(n26330), .A2(\pe3/phq [2]), .B(n25754), .ZN(n25752)
         );
  CLKNAND2HSV2 U28267 ( .A1(\pe3/pvq [2]), .A2(\pe3/ctrq ), .ZN(n25753) );
  NOR2HSV4 U28268 ( .A1(n25755), .A2(\pe3/phq [2]), .ZN(n25754) );
  CLKNAND2HSV2 U28269 ( .A1(\pe3/ti_1 ), .A2(\pe3/got [31]), .ZN(n25755) );
  CLKNHSV3 U28270 ( .I(\pe3/ctrq ), .ZN(n36711) );
  CLKNAND2HSV4 U28271 ( .A1(n25891), .A2(n43140), .ZN(n43493) );
  CLKNAND2HSV4 U28272 ( .A1(n43256), .A2(n43126), .ZN(n25891) );
  XNOR2HSV4 U28273 ( .A1(n25760), .A2(n25756), .ZN(n25807) );
  XNOR2HSV4 U28274 ( .A1(n25758), .A2(n25757), .ZN(n25756) );
  NOR2HSV4 U28275 ( .A1(n43494), .A2(n43867), .ZN(n25757) );
  NOR2HSV4 U28276 ( .A1(n43143), .A2(n43142), .ZN(n43494) );
  XOR2HSV2 U28277 ( .A1(n25759), .A2(n43239), .Z(n25758) );
  OAI22HSV4 U28278 ( .A1(n29643), .A2(n43237), .B1(n43344), .B2(n43238), .ZN(
        n25759) );
  BUFHSV8 U28279 ( .I(n43732), .Z(n25761) );
  CLKNAND2HSV3 U28280 ( .A1(n25762), .A2(n43728), .ZN(n43732) );
  CLKNHSV2 U28281 ( .I(n43723), .ZN(n25762) );
  CLKNHSV3 U28282 ( .I(n43732), .ZN(n29657) );
  CLKNAND2HSV2 U28283 ( .A1(n43366), .A2(n25763), .ZN(n43367) );
  OAI21HSV4 U28284 ( .A1(n25766), .A2(n25771), .B(n25764), .ZN(n26466) );
  AOI21HSV4 U28285 ( .A1(n25765), .A2(n43470), .B(n43469), .ZN(n25764) );
  CLKNAND2HSV2 U28286 ( .A1(n25805), .A2(n25804), .ZN(n43470) );
  CLKNHSV2 U28287 ( .I(n25772), .ZN(n25765) );
  CLKNAND2HSV2 U28288 ( .A1(n25802), .A2(n25803), .ZN(n43490) );
  CLKNAND2HSV3 U28289 ( .A1(n25769), .A2(n26466), .ZN(n43475) );
  CLKNAND2HSV3 U28290 ( .A1(n43472), .A2(n43471), .ZN(n25769) );
  CLKNAND2HSV2 U28291 ( .A1(n45516), .A2(n43464), .ZN(n25770) );
  NAND2HSV2 U28292 ( .A1(n25772), .A2(n43139), .ZN(n25771) );
  NAND2HSV2 U28293 ( .A1(n43256), .A2(n25773), .ZN(n25772) );
  CLKNHSV3 U28294 ( .I(n25774), .ZN(n25773) );
  CLKNAND2HSV3 U28295 ( .A1(n43126), .A2(n25775), .ZN(n25774) );
  CLKNHSV4 U28296 ( .I(n43467), .ZN(n25775) );
  NOR2HSV8 U28297 ( .A1(n25777), .A2(n25776), .ZN(n36718) );
  CLKNAND2HSV3 U28298 ( .A1(n48893), .A2(n36687), .ZN(n25777) );
  CLKNHSV3 U28299 ( .I(n25778), .ZN(n36720) );
  INAND2HSV4 U28300 ( .A1(n36721), .B1(n36718), .ZN(n25778) );
  MUX2NHSV2 U28301 ( .I0(n25780), .I1(n25779), .S(n36711), .ZN(\pe3/bqt[3] )
         );
  CLKNHSV2 U28302 ( .I(bo3[3]), .ZN(n25779) );
  CLKNHSV2 U28303 ( .I(n56529), .ZN(n25780) );
  XOR4HSV2 U28304 ( .A1(\pe3/phq [5]), .A2(n25784), .A3(n25783), .A4(n25782), 
        .Z(n25781) );
  CLKNAND2HSV2 U28305 ( .A1(n36710), .A2(n37186), .ZN(n25782) );
  NOR2HSV4 U28306 ( .A1(n45649), .A2(n59606), .ZN(n25783) );
  CLKNAND2HSV2 U28307 ( .A1(n46141), .A2(\pe3/pvq [5]), .ZN(n25784) );
  XNOR2HSV4 U28308 ( .A1(n25789), .A2(n25786), .ZN(n25785) );
  XNOR2HSV4 U28309 ( .A1(n25788), .A2(n42747), .ZN(n25786) );
  CLKNHSV2 U28310 ( .I(n36999), .ZN(n25787) );
  CLKNAND2HSV2 U28311 ( .A1(n36789), .A2(n59609), .ZN(n25788) );
  XOR2HSV2 U28312 ( .A1(n25791), .A2(n25790), .Z(n25789) );
  CLKNAND2HSV2 U28313 ( .A1(n36795), .A2(n59809), .ZN(n25790) );
  CLKNAND2HSV3 U28314 ( .A1(\pe3/bq[32] ), .A2(\pe3/aot [32]), .ZN(n25796) );
  XNOR2HSV4 U28315 ( .A1(n25795), .A2(n25792), .ZN(n49001) );
  AOI22HSV4 U28316 ( .A1(n59572), .A2(n25794), .B1(n36695), .B2(n25793), .ZN(
        n25792) );
  NOR2HSV4 U28317 ( .A1(n59611), .A2(n59572), .ZN(n25793) );
  XNOR2HSV4 U28318 ( .A1(n25797), .A2(n25796), .ZN(n25795) );
  CLKNAND2HSV2 U28319 ( .A1(\pe3/pvq [1]), .A2(\pe3/ctrq ), .ZN(n25797) );
  INHSV2 U28320 ( .I(n25798), .ZN(n29684) );
  CLKNAND2HSV2 U28321 ( .A1(n42593), .A2(n25799), .ZN(n25798) );
  CLKNAND2HSV3 U28322 ( .A1(n53377), .A2(n37435), .ZN(n25799) );
  CLKNAND2HSV2 U28323 ( .A1(n25799), .A2(n37436), .ZN(n42493) );
  INHSV2 U28324 ( .I(n25800), .ZN(n26342) );
  CLKNAND2HSV4 U28325 ( .A1(n43358), .A2(n26134), .ZN(n25800) );
  CLKNAND2HSV4 U28326 ( .A1(n25800), .A2(n43592), .ZN(n43481) );
  XNOR2HSV4 U28327 ( .A1(n43026), .A2(n43025), .ZN(n60086) );
  CLKNHSV2 U28328 ( .I(n43360), .ZN(n25801) );
  OAI22HSV2 U28329 ( .A1(n43131), .A2(n43359), .B1(n43240), .B2(n43132), .ZN(
        n25802) );
  CLKNAND2HSV1 U28330 ( .A1(n43138), .A2(n43137), .ZN(n25803) );
  CLKNAND2HSV3 U28331 ( .A1(n43494), .A2(n25890), .ZN(n25804) );
  CLKNAND2HSV3 U28332 ( .A1(n26287), .A2(n43240), .ZN(n25805) );
  XNOR2HSV4 U28333 ( .A1(n25807), .A2(n25806), .ZN(n43365) );
  AOI21HSV4 U28334 ( .A1(n25811), .A2(n26551), .B(n25809), .ZN(n25806) );
  CLKNAND2HSV3 U28335 ( .A1(n25808), .A2(n25812), .ZN(n25811) );
  NAND2HSV2 U28336 ( .A1(n43490), .A2(n43139), .ZN(n25808) );
  NOR2HSV4 U28337 ( .A1(n25810), .A2(n43487), .ZN(n25809) );
  CLKNAND2HSV2 U28338 ( .A1(n43493), .A2(n26378), .ZN(n25810) );
  CLKNHSV2 U28339 ( .I(n43744), .ZN(n25812) );
  NAND2HSV2 U28340 ( .A1(n25813), .A2(n42701), .ZN(n42616) );
  NAND3HSV4 U28341 ( .A1(n42598), .A2(n29684), .A3(n42597), .ZN(n25813) );
  NAND3HSV4 U28342 ( .A1(n25813), .A2(n42701), .A3(n42700), .ZN(n43226) );
  NAND3HSV4 U28343 ( .A1(n42617), .A2(n25814), .A3(n26691), .ZN(n42785) );
  CLKNHSV2 U28344 ( .I(n42616), .ZN(n25814) );
  CLKNAND2HSV4 U28345 ( .A1(n42789), .A2(n42613), .ZN(n25815) );
  NAND3HSV4 U28346 ( .A1(n42615), .A2(n42614), .A3(n42924), .ZN(n42789) );
  CLKNHSV2 U28347 ( .I(n25817), .ZN(n25816) );
  CLKNHSV2 U28348 ( .I(n42609), .ZN(n25818) );
  XNOR2HSV4 U28349 ( .A1(n42610), .A2(n42612), .ZN(n42617) );
  CLKNAND2HSV2 U28350 ( .A1(n25821), .A2(n25819), .ZN(n26738) );
  AOI21HSV4 U28351 ( .A1(n25820), .A2(n47784), .B(n26597), .ZN(n25819) );
  CLKNHSV2 U28352 ( .I(n26598), .ZN(n25820) );
  CLKNAND2HSV2 U28353 ( .A1(n26742), .A2(n25822), .ZN(n25821) );
  NOR2HSV4 U28354 ( .A1(n47784), .A2(n25823), .ZN(n25822) );
  CLKNHSV2 U28355 ( .I(n26740), .ZN(n25823) );
  XNOR2HSV4 U28356 ( .A1(n46563), .A2(n46564), .ZN(n47784) );
  BUFHSV4 U28357 ( .I(n38625), .Z(n25824) );
  NAND3HSV4 U28358 ( .A1(n38618), .A2(n38617), .A3(n38611), .ZN(n38625) );
  INHSV4 U28359 ( .I(n38625), .ZN(n44331) );
  INOR2HSV4 U28360 ( .A1(n44650), .B1(n44651), .ZN(n60018) );
  NAND2HSV4 U28361 ( .A1(n41705), .A2(n41704), .ZN(n42033) );
  BUFHSV8 U28362 ( .I(n45415), .Z(n59892) );
  INHSV4 U28363 ( .I(n45415), .ZN(n46976) );
  NAND2HSV4 U28364 ( .A1(n39577), .A2(n39576), .ZN(n39722) );
  NAND2HSV4 U28365 ( .A1(n39740), .A2(n40131), .ZN(n45415) );
  NOR2HSV4 U28366 ( .A1(n35166), .A2(n35165), .ZN(n45793) );
  NOR2HSV4 U28367 ( .A1(n45793), .A2(n35308), .ZN(n35302) );
  NAND2HSV0 U28368 ( .A1(n56863), .A2(n56557), .ZN(n56545) );
  NAND2HSV0 U28369 ( .A1(n56863), .A2(\pe3/got [1]), .ZN(n56879) );
  NAND2HSV0 U28370 ( .A1(n56863), .A2(n55821), .ZN(n55931) );
  NAND2HSV0 U28371 ( .A1(n56863), .A2(n46311), .ZN(n46433) );
  NAND2HSV4 U28372 ( .A1(n44166), .A2(n45114), .ZN(n44949) );
  INHSV4 U28373 ( .I(n46822), .ZN(n58447) );
  NAND2HSV4 U28374 ( .A1(n44692), .A2(n44691), .ZN(n46822) );
  INHSV4 U28375 ( .I(n58447), .ZN(n59026) );
  NAND3HSV4 U28376 ( .A1(n36060), .A2(n36059), .A3(n36058), .ZN(n36061) );
  NAND3HSV3 U28377 ( .A1(n36057), .A2(n46585), .A3(n36056), .ZN(n36058) );
  INHSV4 U28378 ( .I(n36061), .ZN(n49317) );
  CLKNHSV6 U28379 ( .I(n44326), .ZN(n52856) );
  NAND2HSV4 U28380 ( .A1(n26608), .A2(n44304), .ZN(n25825) );
  OAI21HSV2 U28381 ( .A1(n47938), .A2(n28362), .B(n28363), .ZN(n28364) );
  INHSV4 U28382 ( .I(n41846), .ZN(n25826) );
  CLKNAND2HSV4 U28383 ( .A1(n41823), .A2(n42202), .ZN(n41705) );
  CLKNAND2HSV4 U28384 ( .A1(n41607), .A2(n41608), .ZN(n41823) );
  CLKXOR2HSV4 U28385 ( .A1(n41911), .A2(n25827), .Z(n42060) );
  CLKNHSV0 U28386 ( .I(n47554), .ZN(n25828) );
  NAND2HSV0 U28387 ( .A1(n26303), .A2(n25828), .ZN(n28365) );
  INHSV2 U28388 ( .I(n44824), .ZN(n47554) );
  INHSV2 U28389 ( .I(n26303), .ZN(n26301) );
  INHSV4 U28390 ( .I(n38013), .ZN(n47997) );
  OAI21HSV0 U28391 ( .A1(n39725), .A2(n39722), .B(n37767), .ZN(n39724) );
  NOR2HSV2 U28392 ( .A1(n46620), .A2(n31487), .ZN(n26454) );
  NOR2HSV4 U28393 ( .A1(n35787), .A2(n35786), .ZN(n35793) );
  AND2HSV4 U28394 ( .A1(n35785), .A2(n35784), .Z(n35786) );
  NAND3HSV3 U28395 ( .A1(n26004), .A2(n39427), .A3(n39426), .ZN(n26555) );
  INHSV2 U28396 ( .I(n39425), .ZN(n39427) );
  INHSV4 U28397 ( .I(n50716), .ZN(n55944) );
  NAND2HSV4 U28398 ( .A1(n44349), .A2(n44348), .ZN(n47932) );
  NOR2HSV2 U28399 ( .A1(n26465), .A2(n26463), .ZN(n36067) );
  NAND2HSV2 U28400 ( .A1(n40014), .A2(n30881), .ZN(n40015) );
  BUFHSV2 U28401 ( .I(n25835), .Z(n52168) );
  INHSV4 U28402 ( .I(n26547), .ZN(n25835) );
  NAND2HSV0 U28403 ( .A1(n26415), .A2(n45388), .ZN(n45390) );
  INHSV4 U28404 ( .I(n29744), .ZN(n25830) );
  INHSV4 U28405 ( .I(n40290), .ZN(n47199) );
  INHSV4 U28406 ( .I(n52917), .ZN(n45147) );
  OAI21HSV0 U28407 ( .A1(n26464), .A2(n46575), .B(n36065), .ZN(n26463) );
  NAND2HSV2 U28408 ( .A1(n46575), .A2(n31883), .ZN(n36080) );
  NAND2HSV0 U28409 ( .A1(n26467), .A2(n59374), .ZN(n54032) );
  CLKXOR2HSV4 U28410 ( .A1(n46573), .A2(poh6[29]), .Z(po[30]) );
  INHSV4 U28411 ( .I(n54159), .ZN(n59489) );
  NOR2HSV2 U28412 ( .A1(n29761), .A2(n53190), .ZN(n53358) );
  NOR2HSV2 U28413 ( .A1(n25826), .A2(n26617), .ZN(n26616) );
  NOR2HSV2 U28414 ( .A1(n42346), .A2(n42345), .ZN(n26068) );
  OAI21HSV2 U28415 ( .A1(n41920), .A2(n42187), .B(n42318), .ZN(n42345) );
  NAND3HSV3 U28416 ( .A1(n26377), .A2(n26376), .A3(n26375), .ZN(n44952) );
  NAND2HSV4 U28417 ( .A1(n39005), .A2(n39004), .ZN(n52827) );
  NAND2HSV4 U28418 ( .A1(n39003), .A2(n39002), .ZN(n39004) );
  CLKNHSV6 U28419 ( .I(n26547), .ZN(n25834) );
  BUFHSV4 U28420 ( .I(n26415), .Z(n26414) );
  CLKNHSV6 U28421 ( .I(n26407), .ZN(n51797) );
  INHSV6 U28422 ( .I(n25834), .ZN(n26407) );
  NOR2HSV4 U28423 ( .A1(n37987), .A2(n25869), .ZN(n37873) );
  INAND2HSV2 U28424 ( .A1(n38646), .B1(n38778), .ZN(n26820) );
  INHSV4 U28425 ( .I(n38646), .ZN(n59505) );
  CLKXOR2HSV4 U28426 ( .A1(n46548), .A2(poh6[30]), .Z(po[31]) );
  NAND2HSV2 U28427 ( .A1(n47903), .A2(n51151), .ZN(n59794) );
  NAND2HSV0 U28428 ( .A1(n25834), .A2(\pe2/got [17]), .ZN(n26678) );
  NAND2HSV0 U28429 ( .A1(n25835), .A2(n26868), .ZN(n26867) );
  NAND2HSV0 U28430 ( .A1(n51797), .A2(\pe2/got [23]), .ZN(n49596) );
  NAND2HSV0 U28431 ( .A1(n51797), .A2(n52900), .ZN(n28785) );
  NAND2HSV0 U28432 ( .A1(n25834), .A2(n52276), .ZN(n52156) );
  NAND2HSV2 U28433 ( .A1(n55289), .A2(n53473), .ZN(n26276) );
  XOR3HSV2 U28434 ( .A1(n25836), .A2(n26618), .A3(n26616), .Z(n26615) );
  XNOR2HSV1 U28435 ( .A1(n41504), .A2(n41503), .ZN(n25836) );
  NAND3HSV3 U28436 ( .A1(n26523), .A2(n26522), .A3(n26521), .ZN(n26520) );
  NAND2HSV2 U28437 ( .A1(n39579), .A2(n39578), .ZN(n39714) );
  INOR2HSV2 U28438 ( .A1(n47388), .B1(n47389), .ZN(n25837) );
  CLKNAND2HSV2 U28439 ( .A1(n25837), .A2(n26871), .ZN(n53363) );
  CLKAND2HSV4 U28440 ( .A1(n39731), .A2(n30322), .Z(n29661) );
  OA21HSV4 U28441 ( .A1(n39721), .A2(n39734), .B(n39720), .Z(n25838) );
  OAI21HSV0 U28442 ( .A1(n28219), .A2(n28220), .B(n28221), .ZN(n28222) );
  NAND2HSV0 U28443 ( .A1(n28220), .A2(n28219), .ZN(n28221) );
  NAND3HSV3 U28444 ( .A1(n53511), .A2(n26524), .A3(n26520), .ZN(n54553) );
  INHSV4 U28445 ( .I(n26525), .ZN(n26524) );
  NAND2HSV4 U28446 ( .A1(n42350), .A2(n42351), .ZN(n42469) );
  NAND2HSV4 U28447 ( .A1(n42491), .A2(n42338), .ZN(n48313) );
  OR2HSV2 U28448 ( .A1(n45783), .A2(n45780), .Z(n29654) );
  INHSV4 U28449 ( .I(n48456), .ZN(n53503) );
  NAND2HSV0 U28450 ( .A1(n25831), .A2(n52415), .ZN(n52553) );
  NAND2HSV0 U28451 ( .A1(n29358), .A2(n29357), .ZN(n29359) );
  NAND2HSV4 U28452 ( .A1(n26349), .A2(n53511), .ZN(n25839) );
  CLKNAND2HSV2 U28453 ( .A1(n26349), .A2(n53511), .ZN(n25840) );
  CLKNAND2HSV2 U28454 ( .A1(n26349), .A2(n53511), .ZN(n55484) );
  NOR2HSV2 U28455 ( .A1(n44321), .A2(n44959), .ZN(n44325) );
  NAND2HSV0 U28456 ( .A1(n52163), .A2(n59685), .ZN(n51684) );
  NAND2HSV0 U28457 ( .A1(n52163), .A2(n51958), .ZN(n26712) );
  AOI21HSV0 U28458 ( .A1(n39734), .A2(n39733), .B(n37551), .ZN(n39735) );
  MUX2NHSV1 U28459 ( .I0(n39700), .I1(n26427), .S(n39701), .ZN(n39734) );
  NAND3HSV3 U28460 ( .A1(n39227), .A2(n37553), .A3(n39226), .ZN(n39365) );
  XNOR2HSV4 U28461 ( .A1(n57085), .A2(n57084), .ZN(n57088) );
  INHSV2 U28462 ( .I(n30870), .ZN(n30993) );
  XNOR2HSV4 U28463 ( .A1(n47049), .A2(n47048), .ZN(n47050) );
  XNOR2HSV4 U28464 ( .A1(n47047), .A2(n47046), .ZN(n47049) );
  NOR2HSV2 U28465 ( .A1(n58212), .A2(n33830), .ZN(n57980) );
  NOR2HSV2 U28466 ( .A1(n29774), .A2(n34460), .ZN(n50109) );
  NAND2HSV2 U28467 ( .A1(n47903), .A2(n47567), .ZN(n51961) );
  NAND2HSV2 U28468 ( .A1(n47903), .A2(n47567), .ZN(n53097) );
  XOR2HSV0 U28469 ( .A1(n47393), .A2(n25842), .Z(\pe5/poht [31]) );
  OR2HSV2 U28470 ( .A1(n45904), .A2(n51235), .Z(n25842) );
  INHSV2 U28471 ( .I(n47885), .ZN(n25843) );
  INHSV4 U28472 ( .I(n58145), .ZN(n47885) );
  NOR2HSV2 U28473 ( .A1(n39355), .A2(n26791), .ZN(n39368) );
  INHSV4 U28474 ( .I(n39355), .ZN(n39367) );
  CLKNAND2HSV4 U28475 ( .A1(n41506), .A2(n41505), .ZN(n53657) );
  NAND2HSV2 U28476 ( .A1(n55513), .A2(n54969), .ZN(n55224) );
  NAND2HSV2 U28477 ( .A1(n55513), .A2(n59750), .ZN(n29185) );
  XNOR2HSV4 U28478 ( .A1(n39388), .A2(n39387), .ZN(n39393) );
  CLKNAND2HSV2 U28479 ( .A1(n39410), .A2(n39409), .ZN(n39412) );
  NAND3HSV2 U28480 ( .A1(n25843), .A2(n47772), .A3(n47784), .ZN(n26584) );
  BUFHSV6 U28481 ( .I(n26596), .Z(n26692) );
  CLKNAND2HSV2 U28482 ( .A1(n39401), .A2(n39408), .ZN(n37775) );
  XNOR3HSV2 U28483 ( .A1(n25844), .A2(n55374), .A3(n55373), .ZN(\pe1/poht [22]) );
  XOR2HSV0 U28484 ( .A1(n55372), .A2(n26294), .Z(n25844) );
  OAI21HSV2 U28485 ( .A1(n29264), .A2(n29265), .B(n29266), .ZN(n29267) );
  AOI31HSV2 U28486 ( .A1(n45404), .A2(n45405), .A3(n26414), .B(n26139), .ZN(
        n26138) );
  XNOR2HSV4 U28487 ( .A1(n42465), .A2(n42464), .ZN(n25845) );
  NAND3HSV3 U28488 ( .A1(n52836), .A2(n40290), .A3(n30063), .ZN(n40295) );
  XNOR2HSV2 U28489 ( .A1(n51434), .A2(n51433), .ZN(n51436) );
  XOR2HSV0 U28490 ( .A1(n51246), .A2(n25846), .Z(\pe5/poht [28]) );
  XOR2HSV0 U28491 ( .A1(n51245), .A2(n51244), .Z(n25846) );
  INHSV4 U28492 ( .I(n30062), .ZN(n26201) );
  NAND2HSV4 U28493 ( .A1(n30077), .A2(n30078), .ZN(n30062) );
  NAND2HSV4 U28494 ( .A1(n26201), .A2(n30085), .ZN(n26202) );
  NAND2HSV0 U28495 ( .A1(\pe1/got [25]), .A2(n59520), .ZN(n54260) );
  NAND2HSV2 U28496 ( .A1(n26348), .A2(n26347), .ZN(n29980) );
  OAI21HSV2 U28497 ( .A1(n30197), .A2(n39222), .B(n26389), .ZN(n25984) );
  BUFHSV6 U28498 ( .I(n39880), .Z(n59893) );
  XNOR2HSV4 U28499 ( .A1(n39991), .A2(n39990), .ZN(n39994) );
  AND2HSV2 U28500 ( .A1(n37652), .A2(\pe5/got [28]), .Z(n37636) );
  NAND2HSV2 U28501 ( .A1(n53513), .A2(n55086), .ZN(n26273) );
  XOR2HSV0 U28502 ( .A1(n25847), .A2(n51357), .Z(\pe5/poht [26]) );
  XOR2HSV4 U28503 ( .A1(n51356), .A2(n51355), .Z(n25847) );
  CLKNHSV0 U28504 ( .I(n54631), .ZN(n25848) );
  INHSV4 U28505 ( .I(n58348), .ZN(n25849) );
  CLKNHSV6 U28506 ( .I(n58348), .ZN(n48888) );
  CLKNAND2HSV4 U28507 ( .A1(n29880), .A2(n29879), .ZN(n29881) );
  NOR2HSV2 U28508 ( .A1(n25833), .A2(n26676), .ZN(n26675) );
  NOR2HSV2 U28509 ( .A1(n25833), .A2(n26870), .ZN(n26869) );
  INAND2HSV2 U28510 ( .A1(n25833), .B1(n59351), .ZN(n29259) );
  INAND2HSV2 U28511 ( .A1(n45147), .B1(n52276), .ZN(n52277) );
  XOR2HSV4 U28512 ( .A1(n44816), .A2(n44815), .Z(n44819) );
  NAND2HSV4 U28513 ( .A1(n40510), .A2(n40509), .ZN(n40552) );
  CLKNHSV6 U28514 ( .I(n59338), .ZN(n59167) );
  NAND2HSV2 U28515 ( .A1(n25849), .A2(n58423), .ZN(n58350) );
  CLKNAND2HSV2 U28516 ( .A1(n40601), .A2(n26885), .ZN(n26887) );
  CLKNAND2HSV2 U28517 ( .A1(n29765), .A2(n58372), .ZN(n58476) );
  NOR2HSV2 U28518 ( .A1(n26761), .A2(n50091), .ZN(n58295) );
  NOR2HSV2 U28519 ( .A1(n26761), .A2(n50052), .ZN(n57979) );
  NOR2HSV2 U28520 ( .A1(n26761), .A2(n35488), .ZN(n57669) );
  NOR2HSV2 U28521 ( .A1(n26761), .A2(n50064), .ZN(n58213) );
  NOR2HSV2 U28522 ( .A1(n26761), .A2(n50095), .ZN(n58319) );
  CLKNHSV6 U28523 ( .I(n40346), .ZN(n40357) );
  CLKNAND2HSV4 U28524 ( .A1(n40345), .A2(n40344), .ZN(n40346) );
  INHSV4 U28525 ( .I(n40600), .ZN(n26885) );
  CLKNHSV0 U28526 ( .I(n45148), .ZN(n44713) );
  NAND2HSV4 U28527 ( .A1(n39429), .A2(n39428), .ZN(n59883) );
  INHSV4 U28528 ( .I(n40640), .ZN(n40642) );
  XNOR2HSV4 U28529 ( .A1(n50642), .A2(n50641), .ZN(n50645) );
  XNOR2HSV4 U28530 ( .A1(n50640), .A2(n50639), .ZN(n50641) );
  NAND2HSV4 U28531 ( .A1(n40813), .A2(n40812), .ZN(n41391) );
  OR2HSV2 U28532 ( .A1(n40805), .A2(n40804), .Z(n40813) );
  CLKAND2HSV2 U28533 ( .A1(n40811), .A2(n40810), .Z(n40812) );
  NAND2HSV2 U28534 ( .A1(n40635), .A2(n40482), .ZN(n40483) );
  NOR2HSV2 U28535 ( .A1(n42343), .A2(n26281), .ZN(n26280) );
  NOR2HSV2 U28536 ( .A1(n33463), .A2(n33462), .ZN(n33466) );
  CLKNAND2HSV4 U28537 ( .A1(n41840), .A2(n41839), .ZN(n41921) );
  MOAI22HSV4 U28538 ( .A1(n26284), .A2(n42197), .B1(n42197), .B2(n42198), .ZN(
        n42486) );
  BUFHSV6 U28539 ( .I(n36100), .Z(n26152) );
  XNOR2HSV4 U28540 ( .A1(n39336), .A2(n39335), .ZN(n39338) );
  XNOR2HSV4 U28541 ( .A1(n39343), .A2(n39342), .ZN(n39344) );
  XNOR2HSV4 U28542 ( .A1(n39340), .A2(n39339), .ZN(n39343) );
  NOR2HSV4 U28543 ( .A1(n25982), .A2(n25981), .ZN(n25852) );
  NOR2HSV2 U28544 ( .A1(n25982), .A2(n25981), .ZN(n25853) );
  NOR2HSV4 U28545 ( .A1(n25982), .A2(n25981), .ZN(n30252) );
  BUFHSV6 U28546 ( .I(n54683), .Z(n59934) );
  DELHS4 U28547 ( .I(n41391), .Z(n41894) );
  DELHS4 U28548 ( .I(n41391), .Z(n54115) );
  DELHS4 U28549 ( .I(n54732), .Z(n54513) );
  INHSV4 U28550 ( .I(n26020), .ZN(n26019) );
  CLKXOR2HSV4 U28551 ( .A1(n33502), .A2(n33501), .Z(n33503) );
  INHSV4 U28552 ( .I(n26026), .ZN(n26104) );
  CLKNAND2HSV2 U28553 ( .A1(n45410), .A2(n45131), .ZN(n45133) );
  BUFHSV2 U28554 ( .I(n30485), .Z(n47058) );
  NAND2HSV2 U28555 ( .A1(n30485), .A2(n39249), .ZN(n26391) );
  OR2HSV2 U28556 ( .A1(n30193), .A2(n30184), .Z(n29712) );
  NAND3HSV3 U28557 ( .A1(n26202), .A2(n26203), .A3(n30073), .ZN(n26425) );
  NAND2HSV4 U28558 ( .A1(n26425), .A2(n30138), .ZN(n25981) );
  OAI21HSV2 U28559 ( .A1(n47990), .A2(n26168), .B(n26167), .ZN(n25854) );
  INHSV4 U28560 ( .I(n33067), .ZN(n25855) );
  XOR2HSV4 U28561 ( .A1(n33071), .A2(n33070), .Z(n33067) );
  CLKNAND2HSV2 U28562 ( .A1(n38441), .A2(n38444), .ZN(n38188) );
  NAND2HSV2 U28563 ( .A1(n26802), .A2(n33575), .ZN(n33666) );
  CLKNHSV0 U28564 ( .I(n33224), .ZN(n25856) );
  CLKNHSV6 U28565 ( .I(\pe2/aot [32]), .ZN(n36240) );
  CLKNAND2HSV2 U28566 ( .A1(n29765), .A2(n58383), .ZN(n29772) );
  XNOR2HSV4 U28567 ( .A1(n40630), .A2(n40629), .ZN(n40631) );
  NAND2HSV0 U28568 ( .A1(n40341), .A2(n40340), .ZN(n25857) );
  CLKNHSV0 U28569 ( .I(n41605), .ZN(n25858) );
  INHSV4 U28570 ( .I(n47960), .ZN(n41605) );
  NAND3HSV4 U28571 ( .A1(n43950), .A2(n36399), .A3(n36398), .ZN(n36400) );
  INHSV4 U28572 ( .I(n33662), .ZN(n33514) );
  CLKNAND2HSV2 U28573 ( .A1(n36415), .A2(n36414), .ZN(n52719) );
  OAI21HSV2 U28574 ( .A1(n27774), .A2(n27775), .B(n27776), .ZN(n27777) );
  NAND2HSV2 U28575 ( .A1(n33508), .A2(n33507), .ZN(n33509) );
  OAI21HSV2 U28576 ( .A1(n29454), .A2(n29455), .B(n29456), .ZN(n29457) );
  AOI22HSV2 U28577 ( .A1(n30322), .A2(n30653), .B1(n30428), .B2(n30321), .ZN(
        n30323) );
  MUX2NHSV1 U28578 ( .I0(n30996), .I1(n30995), .S(n26043), .ZN(n30998) );
  CLKNAND2HSV2 U28579 ( .A1(n30312), .A2(n30311), .ZN(n30314) );
  INHSV4 U28580 ( .I(n30305), .ZN(n30311) );
  NAND2HSV0 U28581 ( .A1(n46169), .A2(n46553), .ZN(n46165) );
  OAI21HSV2 U28582 ( .A1(n32814), .A2(n32530), .B(n32458), .ZN(n26468) );
  CLKNHSV6 U28583 ( .I(n32458), .ZN(n32453) );
  OAI21HSV2 U28584 ( .A1(n27426), .A2(n27427), .B(n27428), .ZN(n27429) );
  NAND2HSV0 U28585 ( .A1(n27427), .A2(n27426), .ZN(n27428) );
  CLKXOR2HSV4 U28586 ( .A1(n35707), .A2(n35706), .Z(n35714) );
  NAND2HSV4 U28587 ( .A1(n59570), .A2(n36029), .ZN(n26732) );
  CLKNAND2HSV2 U28588 ( .A1(n29765), .A2(n58372), .ZN(n58655) );
  NAND3HSV3 U28589 ( .A1(n44355), .A2(n44352), .A3(n35807), .ZN(n35810) );
  CLKNHSV0 U28590 ( .I(n44352), .ZN(n44354) );
  NAND2HSV4 U28591 ( .A1(n36235), .A2(n36234), .ZN(n46151) );
  NAND3HSV3 U28592 ( .A1(n44681), .A2(n26262), .A3(n44682), .ZN(n44684) );
  CLKNAND2HSV2 U28593 ( .A1(n32661), .A2(n32660), .ZN(n32662) );
  CLKNHSV6 U28594 ( .I(n30194), .ZN(n30184) );
  INHSV4 U28595 ( .I(n33409), .ZN(n45804) );
  INHSV4 U28596 ( .I(n33575), .ZN(n33448) );
  INHSV4 U28597 ( .I(n26795), .ZN(n33602) );
  NAND2HSV2 U28598 ( .A1(n34003), .A2(n34002), .ZN(n34199) );
  BUFHSV8 U28599 ( .I(n43916), .Z(n44148) );
  OAI21HSV2 U28600 ( .A1(n31002), .A2(n37534), .B(n26681), .ZN(n26680) );
  INHSV2 U28601 ( .I(n30141), .ZN(n29663) );
  CLKNAND2HSV4 U28602 ( .A1(n44160), .A2(n44159), .ZN(n44165) );
  XNOR2HSV4 U28603 ( .A1(n26236), .A2(n45385), .ZN(n45387) );
  CLKNHSV0 U28604 ( .I(n29466), .ZN(n25859) );
  MUX2NHSV2 U28605 ( .I0(n29936), .I1(n29935), .S(n29958), .ZN(n29974) );
  CLKXOR2HSV4 U28606 ( .A1(n40759), .A2(n40758), .Z(n40760) );
  XOR2HSV4 U28607 ( .A1(n40756), .A2(n40755), .Z(n40759) );
  NAND3HSV2 U28608 ( .A1(n30307), .A2(n30313), .A3(n39733), .ZN(n30308) );
  INHSV4 U28609 ( .I(n38377), .ZN(n26790) );
  NAND2HSV2 U28610 ( .A1(n45286), .A2(n38777), .ZN(n26236) );
  NAND2HSV2 U28611 ( .A1(n45403), .A2(n25834), .ZN(n26375) );
  NAND2HSV4 U28612 ( .A1(n33279), .A2(n52731), .ZN(n33383) );
  INHSV4 U28613 ( .I(n33237), .ZN(n33239) );
  OAI21HSV4 U28614 ( .A1(n60040), .A2(n30064), .B(n30027), .ZN(n30181) );
  NAND2HSV4 U28615 ( .A1(n33244), .A2(n33243), .ZN(n52731) );
  CLKNAND2HSV2 U28616 ( .A1(n44645), .A2(n44646), .ZN(n44647) );
  XNOR2HSV4 U28617 ( .A1(n44365), .A2(n44364), .ZN(n44366) );
  CLKNAND2HSV2 U28618 ( .A1(n29738), .A2(n59599), .ZN(n33560) );
  NAND2HSV2 U28619 ( .A1(n44955), .A2(n52856), .ZN(n44965) );
  CLKNAND2HSV2 U28620 ( .A1(n31874), .A2(n31875), .ZN(n51441) );
  BUFHSV8 U28621 ( .I(n31382), .Z(n31572) );
  INHSV4 U28622 ( .I(n30334), .ZN(n52754) );
  CLKNAND2HSV2 U28623 ( .A1(n31324), .A2(n31353), .ZN(n31388) );
  INHSV8 U28624 ( .I(n40547), .ZN(n41824) );
  OAI21HSV2 U28625 ( .A1(n33085), .A2(n35704), .B(n35703), .ZN(n36100) );
  CLKNAND2HSV4 U28626 ( .A1(n60108), .A2(n41410), .ZN(n40468) );
  AOI21HSV2 U28627 ( .A1(n44379), .A2(n45788), .B(n44387), .ZN(n44386) );
  NAND2HSV2 U28628 ( .A1(n44673), .A2(n44674), .ZN(n26224) );
  INHSV2 U28629 ( .I(n29974), .ZN(n29977) );
  CLKNAND2HSV2 U28630 ( .A1(n29974), .A2(n29975), .ZN(n26347) );
  NAND2HSV0 U28631 ( .A1(n55448), .A2(n54154), .ZN(n55538) );
  NAND2HSV0 U28632 ( .A1(n53513), .A2(n55222), .ZN(n55223) );
  NAND2HSV0 U28633 ( .A1(n59520), .A2(\pe1/got [24]), .ZN(n54554) );
  NAND2HSV4 U28634 ( .A1(n46071), .A2(n46082), .ZN(n45769) );
  OAI21HSV2 U28635 ( .A1(n29582), .A2(n29583), .B(n29584), .ZN(n29585) );
  INAND2HSV2 U28636 ( .A1(n55158), .B1(n40482), .ZN(n53651) );
  NAND3HSV2 U28637 ( .A1(n29989), .A2(n29990), .A3(n29988), .ZN(n25861) );
  INAND2HSV4 U28638 ( .A1(n30325), .B1(n25983), .ZN(n25862) );
  INAND2HSV2 U28639 ( .A1(n30325), .B1(n25983), .ZN(n30304) );
  CLKNAND2HSV2 U28640 ( .A1(n45632), .A2(n45631), .ZN(n45778) );
  CLKNAND2HSV2 U28641 ( .A1(n26242), .A2(n44824), .ZN(n26241) );
  CLKNAND2HSV8 U28642 ( .A1(n40380), .A2(n40379), .ZN(n40786) );
  NAND2HSV4 U28643 ( .A1(n60051), .A2(n44309), .ZN(n26608) );
  NAND2HSV4 U28644 ( .A1(n39381), .A2(n39380), .ZN(n39576) );
  NAND2HSV2 U28645 ( .A1(n50929), .A2(n38389), .ZN(n26955) );
  NAND2HSV2 U28646 ( .A1(n26955), .A2(n26954), .ZN(n26956) );
  XNOR2HSV4 U28647 ( .A1(n45391), .A2(n45390), .ZN(n45392) );
  NAND2HSV0 U28648 ( .A1(n52416), .A2(n51485), .ZN(n45082) );
  CLKNAND2HSV4 U28649 ( .A1(n40712), .A2(n40711), .ZN(n40805) );
  NAND2HSV2 U28650 ( .A1(n38323), .A2(n38327), .ZN(n38095) );
  NAND2HSV2 U28651 ( .A1(n29930), .A2(n29931), .ZN(n60037) );
  NAND2HSV2 U28652 ( .A1(n26345), .A2(n29979), .ZN(n29981) );
  OAI22HSV0 U28653 ( .A1(n41076), .A2(n54185), .B1(n40445), .B2(n42264), .ZN(
        n40570) );
  INHSV4 U28654 ( .I(n38443), .ZN(n38452) );
  CLKNHSV4 U28655 ( .I(n38779), .ZN(n51966) );
  INHSV6 U28656 ( .I(n37346), .ZN(n37349) );
  XOR2HSV4 U28657 ( .A1(n48611), .A2(n48610), .Z(n48612) );
  DELHS4 U28658 ( .I(n38841), .Z(n59679) );
  OAI21HSV2 U28659 ( .A1(n26951), .A2(n26952), .B(n26953), .ZN(n26954) );
  CLKNAND2HSV2 U28660 ( .A1(n33296), .A2(n33300), .ZN(n33298) );
  XNOR2HSV4 U28661 ( .A1(n34230), .A2(n34229), .ZN(n34349) );
  OAI21HSV2 U28662 ( .A1(n48451), .A2(n42037), .B(n42470), .ZN(n42475) );
  NOR2HSV4 U28663 ( .A1(n38115), .A2(n38114), .ZN(n26089) );
  CLKNAND2HSV4 U28664 ( .A1(n26898), .A2(n26897), .ZN(n38115) );
  NAND2HSV0 U28665 ( .A1(n38537), .A2(\pe2/got [29]), .ZN(n38598) );
  BUFHSV6 U28666 ( .I(n38537), .Z(n59773) );
  CLKNHSV0 U28667 ( .I(n39880), .ZN(n25863) );
  INHSV2 U28668 ( .I(n25863), .ZN(n25864) );
  NAND2HSV0 U28669 ( .A1(n44145), .A2(n44780), .ZN(n36626) );
  INHSV4 U28670 ( .I(n38889), .ZN(n25865) );
  INHSV4 U28671 ( .I(n38887), .ZN(n38889) );
  CLKNAND2HSV4 U28672 ( .A1(n25941), .A2(n48619), .ZN(n36982) );
  OAI21HSV2 U28673 ( .A1(n29097), .A2(n29098), .B(n29099), .ZN(n29100) );
  NAND2HSV2 U28674 ( .A1(n44694), .A2(n37630), .ZN(n26496) );
  NAND2HSV2 U28675 ( .A1(n34994), .A2(n34419), .ZN(n35029) );
  CLKXOR2HSV2 U28676 ( .A1(n33845), .A2(n33844), .Z(n25874) );
  CLKNHSV0 U28677 ( .I(n45797), .ZN(n42811) );
  NAND3HSV4 U28678 ( .A1(n42930), .A2(n42929), .A3(n45797), .ZN(n42935) );
  NAND3HSV3 U28679 ( .A1(n25865), .A2(n52924), .A3(n44827), .ZN(n26852) );
  CLKNHSV6 U28680 ( .I(n57835), .ZN(n50211) );
  CLKNHSV0 U28681 ( .I(n31758), .ZN(n25866) );
  NAND2HSV4 U28682 ( .A1(n26658), .A2(n26656), .ZN(n31814) );
  NAND2HSV2 U28683 ( .A1(n47785), .A2(n47786), .ZN(n26634) );
  NAND2HSV2 U28684 ( .A1(n27577), .A2(n27576), .ZN(n27578) );
  AOI31HSV2 U28685 ( .A1(n29649), .A2(n44358), .A3(n44359), .B(n44357), .ZN(
        n44360) );
  OAI21HSV2 U28686 ( .A1(n29515), .A2(n29516), .B(n29517), .ZN(n29518) );
  NAND2HSV2 U28687 ( .A1(n29516), .A2(n29515), .ZN(n29517) );
  OAI21HSV2 U28688 ( .A1(n29518), .A2(n29519), .B(n29520), .ZN(n29521) );
  NAND2HSV2 U28689 ( .A1(n29519), .A2(n29518), .ZN(n29520) );
  CLKNAND2HSV4 U28690 ( .A1(n31525), .A2(n31524), .ZN(n31540) );
  XOR2HSV4 U28691 ( .A1(n56728), .A2(n56727), .Z(n56729) );
  XNOR2HSV4 U28692 ( .A1(n56726), .A2(n56725), .ZN(n56727) );
  CLKNAND2HSV8 U28693 ( .A1(n32462), .A2(n32461), .ZN(n32686) );
  INHSV4 U28694 ( .I(n41716), .ZN(n41717) );
  NOR2HSV4 U28695 ( .A1(n41908), .A2(n42031), .ZN(n41716) );
  NOR2HSV0 U28696 ( .A1(n26234), .A2(pov3[24]), .ZN(n26233) );
  CLKNAND2HSV2 U28697 ( .A1(pov3[24]), .A2(n26671), .ZN(n43730) );
  NAND2HSV4 U28698 ( .A1(n26307), .A2(n31625), .ZN(n31677) );
  NAND2HSV2 U28699 ( .A1(n38118), .A2(n38117), .ZN(n29749) );
  INHSV2 U28700 ( .I(n26838), .ZN(n26837) );
  AOI21HSV2 U28701 ( .A1(n29767), .A2(n40952), .B(n26208), .ZN(n26850) );
  NAND3HSV2 U28702 ( .A1(n52785), .A2(n52787), .A3(n26573), .ZN(n26579) );
  NAND3HSV3 U28703 ( .A1(n52785), .A2(n52787), .A3(n30757), .ZN(n30965) );
  AOI31HSV2 U28704 ( .A1(n46088), .A2(n46087), .A3(n46092), .B(n46086), .ZN(
        n46097) );
  NOR2HSV2 U28705 ( .A1(n42066), .A2(n42065), .ZN(n42081) );
  MUX2NHSV2 U28706 ( .I0(n29055), .I1(n41233), .S(n29060), .ZN(n29061) );
  AOI21HSV2 U28707 ( .A1(n41235), .A2(n41234), .B(n29053), .ZN(n29054) );
  CLKNHSV0 U28708 ( .I(n31748), .ZN(n25867) );
  INHSV2 U28709 ( .I(n25867), .ZN(n25868) );
  NAND2HSV0 U28710 ( .A1(n25848), .A2(n54033), .ZN(n54034) );
  NAND2HSV0 U28711 ( .A1(n55589), .A2(n55337), .ZN(n55083) );
  NAND2HSV0 U28712 ( .A1(n55589), .A2(n41689), .ZN(n29610) );
  NAND2HSV0 U28713 ( .A1(n55410), .A2(n54154), .ZN(n55590) );
  NAND2HSV0 U28714 ( .A1(n55145), .A2(n53513), .ZN(n55485) );
  CLKXOR2HSV2 U28715 ( .A1(n56610), .A2(n56609), .Z(n56611) );
  XNOR2HSV4 U28716 ( .A1(n56614), .A2(n56613), .ZN(n56617) );
  CLKXOR2HSV4 U28717 ( .A1(n56612), .A2(n56611), .Z(n56613) );
  CLKXOR2HSV2 U28718 ( .A1(n56849), .A2(n56848), .Z(n56850) );
  XNOR2HSV4 U28719 ( .A1(n56853), .A2(n56852), .ZN(n56858) );
  XOR2HSV4 U28720 ( .A1(n56851), .A2(n56850), .Z(n56852) );
  CLKXOR2HSV2 U28721 ( .A1(n56927), .A2(n56926), .Z(n56928) );
  XNOR2HSV4 U28722 ( .A1(n56931), .A2(n56930), .ZN(n56934) );
  XOR2HSV4 U28723 ( .A1(n56929), .A2(n56928), .Z(n56930) );
  INHSV2 U28724 ( .I(n37759), .ZN(n37761) );
  NOR2HSV4 U28725 ( .A1(n28597), .A2(n41913), .ZN(n42042) );
  NAND2HSV2 U28726 ( .A1(n40466), .A2(n41915), .ZN(n28597) );
  CLKNHSV6 U28727 ( .I(n31288), .ZN(n31291) );
  INHSV4 U28728 ( .I(n35711), .ZN(n35716) );
  INHSV2 U28729 ( .I(n46103), .ZN(n46105) );
  MUX2NHSV4 U28730 ( .I0(n47786), .I1(n47787), .S(n52848), .ZN(n26633) );
  NOR2HSV2 U28731 ( .A1(n26761), .A2(n47793), .ZN(n49962) );
  NOR2HSV2 U28732 ( .A1(n26761), .A2(n46581), .ZN(n57205) );
  NAND3HSV2 U28733 ( .A1(n30994), .A2(n30870), .A3(n26583), .ZN(n31000) );
  CLKNAND2HSV2 U28734 ( .A1(n30877), .A2(n30994), .ZN(n30878) );
  NOR2HSV4 U28735 ( .A1(n31763), .A2(n48018), .ZN(n31699) );
  OAI21HSV2 U28736 ( .A1(n31898), .A2(n31888), .B(n31887), .ZN(n31889) );
  INHSV2 U28737 ( .I(n37849), .ZN(n25869) );
  INHSV4 U28738 ( .I(n37989), .ZN(n37849) );
  INHSV4 U28739 ( .I(n42477), .ZN(n48314) );
  INHSV4 U28740 ( .I(n42476), .ZN(n44652) );
  BUFHSV4 U28741 ( .I(n37992), .Z(n25870) );
  INHSV4 U28742 ( .I(n36283), .ZN(n25871) );
  INHSV4 U28743 ( .I(n36406), .ZN(n36283) );
  INHSV2 U28744 ( .I(n41590), .ZN(n29207) );
  NAND2HSV4 U28745 ( .A1(n41708), .A2(n41411), .ZN(n41908) );
  NAND2HSV2 U28746 ( .A1(n45477), .A2(n30254), .ZN(n30145) );
  CLKNAND2HSV4 U28747 ( .A1(n26705), .A2(n26703), .ZN(n45477) );
  NOR2HSV2 U28748 ( .A1(n25852), .A2(n40130), .ZN(n26399) );
  MUX2NHSV4 U28749 ( .I0(n41696), .I1(n26847), .S(n26846), .ZN(n26845) );
  AOI21HSV2 U28750 ( .A1(n43484), .A2(n45928), .B(n45620), .ZN(n45632) );
  NOR2HSV2 U28751 ( .A1(n43592), .A2(n43591), .ZN(n26343) );
  CLKNAND2HSV4 U28752 ( .A1(n39216), .A2(n31139), .ZN(n31235) );
  INHSV2 U28753 ( .I(n31236), .ZN(n31232) );
  BUFHSV8 U28754 ( .I(n45516), .Z(n46312) );
  CLKNHSV0 U28755 ( .I(n42483), .ZN(n25872) );
  CLKNHSV0 U28756 ( .I(n25872), .ZN(n25873) );
  CLKNHSV6 U28757 ( .I(n32663), .ZN(n32674) );
  INHSV4 U28758 ( .I(n53503), .ZN(n55213) );
  INAND2HSV2 U28759 ( .A1(n26625), .B1(n42085), .ZN(n26624) );
  NAND2HSV2 U28760 ( .A1(\pe4/got [32]), .A2(\pe4/ti_1 ), .ZN(n26192) );
  CLKNAND2HSV4 U28761 ( .A1(n34094), .A2(n34095), .ZN(n34102) );
  CLKNAND2HSV4 U28762 ( .A1(n34686), .A2(n34685), .ZN(n34733) );
  BUFHSV6 U28763 ( .I(n34733), .Z(n47835) );
  INHSV4 U28764 ( .I(\pe4/ti_1 ), .ZN(n46618) );
  MUX2NHSV1 U28765 ( .I0(n29619), .I1(n46618), .S(n48068), .ZN(\pe4/ti_1t ) );
  CLKNHSV0 U28766 ( .I(n46618), .ZN(n33897) );
  CLKNAND2HSV8 U28767 ( .A1(n40154), .A2(n40153), .ZN(n52838) );
  CLKNAND2HSV2 U28768 ( .A1(n37918), .A2(n47998), .ZN(n37833) );
  NAND2HSV2 U28769 ( .A1(n29767), .A2(n41831), .ZN(n41832) );
  NAND3HSV3 U28770 ( .A1(n32812), .A2(n32813), .A3(n32811), .ZN(n35721) );
  XNOR2HSV4 U28771 ( .A1(n33846), .A2(n25874), .ZN(n33926) );
  INAND2HSV2 U28772 ( .A1(n34588), .B1(n34587), .ZN(n25875) );
  CLKNAND2HSV4 U28773 ( .A1(n33793), .A2(n33792), .ZN(n34408) );
  AOI31HSV2 U28774 ( .A1(n44964), .A2(n44962), .A3(n44963), .B(n44961), .ZN(
        n26512) );
  CLKNAND2HSV2 U28775 ( .A1(n31395), .A2(n31394), .ZN(n31396) );
  NAND2HSV4 U28776 ( .A1(n38194), .A2(n38193), .ZN(n38471) );
  OR2HSV2 U28777 ( .A1(n33999), .A2(n52797), .Z(n29667) );
  NAND2HSV2 U28778 ( .A1(n32692), .A2(n59166), .ZN(n32346) );
  INHSV6 U28779 ( .I(n30960), .ZN(n44694) );
  NAND2HSV4 U28780 ( .A1(n34451), .A2(n34450), .ZN(n34819) );
  NAND2HSV4 U28781 ( .A1(n34700), .A2(n34701), .ZN(n34340) );
  CLKNHSV3 U28782 ( .I(n50298), .ZN(n57889) );
  NAND2HSV2 U28783 ( .A1(n33345), .A2(n33344), .ZN(n26231) );
  NAND3HSV3 U28784 ( .A1(n34578), .A2(n34577), .A3(n34337), .ZN(n34698) );
  NAND2HSV2 U28785 ( .A1(n44660), .A2(n44661), .ZN(n26536) );
  CLKNHSV0 U28786 ( .I(n52820), .ZN(n25877) );
  INHSV2 U28787 ( .I(n25877), .ZN(n25878) );
  NAND2HSV4 U28788 ( .A1(n34016), .A2(n34015), .ZN(n34592) );
  INHSV4 U28789 ( .I(n33893), .ZN(n33415) );
  NAND3HSV4 U28790 ( .A1(n34001), .A2(n34000), .A3(n29667), .ZN(n25879) );
  NAND3HSV2 U28791 ( .A1(n34001), .A2(n34000), .A3(n29667), .ZN(n34229) );
  CLKNAND2HSV4 U28792 ( .A1(n33519), .A2(n33518), .ZN(n33661) );
  XNOR2HSV4 U28793 ( .A1(n33931), .A2(n33930), .ZN(n33932) );
  MUX2NHSV2 U28794 ( .I0(n33335), .I1(n33334), .S(n33333), .ZN(n25880) );
  MUX2NHSV2 U28795 ( .I0(n33335), .I1(n33334), .S(n33333), .ZN(n33336) );
  NAND3HSV3 U28796 ( .A1(n33299), .A2(n33298), .A3(n33301), .ZN(n33335) );
  NAND2HSV4 U28797 ( .A1(n33771), .A2(n33770), .ZN(n33850) );
  NAND2HSV2 U28798 ( .A1(\pe4/pvq [3]), .A2(\pe4/ctrq ), .ZN(n27824) );
  INHSV4 U28799 ( .I(n26206), .ZN(n33161) );
  XNOR2HSV4 U28800 ( .A1(n34678), .A2(n34677), .ZN(n34684) );
  NAND2HSV4 U28801 ( .A1(n33384), .A2(n33383), .ZN(n33412) );
  NAND3HSV2 U28802 ( .A1(n33384), .A2(n33383), .A3(n33382), .ZN(n45806) );
  NAND2HSV4 U28803 ( .A1(n26219), .A2(n52697), .ZN(n33157) );
  INOR2HSV4 U28804 ( .A1(n34831), .B1(n34830), .ZN(n34832) );
  INHSV2 U28805 ( .I(n35296), .ZN(n25881) );
  CLKNAND2HSV2 U28806 ( .A1(n35298), .A2(n25881), .ZN(n35166) );
  NAND3HSV4 U28807 ( .A1(n34196), .A2(n34199), .A3(n33094), .ZN(n34004) );
  NAND2HSV4 U28808 ( .A1(n35004), .A2(n35008), .ZN(n35305) );
  NOR2HSV4 U28809 ( .A1(n37833), .A2(n37832), .ZN(n37844) );
  CLKNHSV0 U28810 ( .I(n40317), .ZN(n40302) );
  NAND3HSV3 U28811 ( .A1(n33578), .A2(n33459), .A3(n33458), .ZN(n33667) );
  XNOR2HSV4 U28812 ( .A1(n32810), .A2(n32809), .ZN(n32966) );
  CLKNHSV6 U28813 ( .I(n40411), .ZN(n53411) );
  XNOR2HSV4 U28814 ( .A1(n40415), .A2(n40414), .ZN(n40423) );
  OAI21HSV2 U28815 ( .A1(n28182), .A2(n28183), .B(n28184), .ZN(n28185) );
  NAND2HSV0 U28816 ( .A1(n49661), .A2(\pe2/got [8]), .ZN(n51153) );
  NAND2HSV2 U28817 ( .A1(n40317), .A2(n40008), .ZN(n26314) );
  OAI21HSV2 U28818 ( .A1(n40404), .A2(n40403), .B(n40402), .ZN(n40405) );
  CLKNAND2HSV2 U28819 ( .A1(n34103), .A2(n34102), .ZN(n34319) );
  CLKNAND2HSV4 U28820 ( .A1(n58439), .A2(n58438), .ZN(n46306) );
  CLKNAND2HSV4 U28821 ( .A1(n32543), .A2(n32542), .ZN(n32663) );
  OAI21HSV4 U28822 ( .A1(n31709), .A2(n31708), .B(n31707), .ZN(n31745) );
  CLKNAND2HSV2 U28823 ( .A1(n40424), .A2(n26108), .ZN(n26106) );
  NOR2HSV4 U28824 ( .A1(n36082), .A2(n44339), .ZN(n36086) );
  CLKNAND2HSV4 U28825 ( .A1(n37325), .A2(n36922), .ZN(n25950) );
  NAND2HSV4 U28826 ( .A1(n47969), .A2(n47773), .ZN(n47967) );
  BUFHSV6 U28827 ( .I(n49726), .Z(n58702) );
  BUFHSV4 U28828 ( .I(n35788), .Z(n49726) );
  CLKNHSV0 U28829 ( .I(n52823), .ZN(n25883) );
  INHSV2 U28830 ( .I(n25883), .ZN(n25884) );
  CLKNAND2HSV4 U28831 ( .A1(n33164), .A2(n33163), .ZN(n33180) );
  NOR2HSV4 U28832 ( .A1(n46162), .A2(n46161), .ZN(n58437) );
  AOI21HSV2 U28833 ( .A1(n40816), .A2(n59934), .B(n40815), .ZN(n40817) );
  CLKNHSV0 U28834 ( .I(n58442), .ZN(n25885) );
  INHSV2 U28835 ( .I(n25885), .ZN(n25886) );
  NAND2HSV2 U28836 ( .A1(n47940), .A2(n36047), .ZN(n36063) );
  CLKNAND2HSV4 U28837 ( .A1(n38531), .A2(n38530), .ZN(n44043) );
  NAND3HSV4 U28838 ( .A1(n41603), .A2(n41602), .A3(n41601), .ZN(n47960) );
  NAND3HSV3 U28839 ( .A1(n41599), .A2(n41597), .A3(n41598), .ZN(n41602) );
  NAND2HSV2 U28840 ( .A1(n32943), .A2(n32967), .ZN(n32944) );
  CLKNAND2HSV2 U28841 ( .A1(n38387), .A2(n38382), .ZN(n38334) );
  INHSV2 U28842 ( .I(n38536), .ZN(n38645) );
  INHSV6 U28843 ( .I(n44826), .ZN(n44828) );
  NAND2HSV4 U28844 ( .A1(n29696), .A2(n45092), .ZN(n44824) );
  INAND2HSV2 U28845 ( .A1(n44824), .B1(n44828), .ZN(n26243) );
  NAND2HSV2 U28846 ( .A1(n58808), .A2(n59021), .ZN(n29043) );
  INHSV4 U28847 ( .I(n59338), .ZN(n59021) );
  NAND2HSV0 U28848 ( .A1(n29043), .A2(n29042), .ZN(n29044) );
  NOR2HSV4 U28849 ( .A1(n34537), .A2(n33929), .ZN(n33758) );
  NAND2HSV4 U28850 ( .A1(n41116), .A2(n41115), .ZN(n41120) );
  CLKNHSV4 U28851 ( .I(n53389), .ZN(n53792) );
  NOR2HSV4 U28852 ( .A1(n34839), .A2(n34838), .ZN(n34841) );
  OAI21HSV2 U28853 ( .A1(n28540), .A2(n28541), .B(n28542), .ZN(n28543) );
  NAND2HSV0 U28854 ( .A1(n28541), .A2(n28540), .ZN(n28542) );
  NAND2HSV0 U28855 ( .A1(n45410), .A2(n45409), .ZN(n26136) );
  NAND2HSV4 U28856 ( .A1(n25900), .A2(n40541), .ZN(n42082) );
  NAND2HSV4 U28857 ( .A1(n34710), .A2(n34709), .ZN(n34842) );
  BUFHSV4 U28858 ( .I(n35569), .Z(n49966) );
  OAI21HSV4 U28859 ( .A1(n33857), .A2(n33856), .B(n33855), .ZN(n35569) );
  NOR2HSV4 U28860 ( .A1(n45929), .A2(n45928), .ZN(n45935) );
  NOR2HSV0 U28861 ( .A1(n31535), .A2(n32057), .ZN(n31526) );
  INHSV4 U28862 ( .I(n39682), .ZN(n39675) );
  INHSV4 U28863 ( .I(n37085), .ZN(n37325) );
  AOI22HSV4 U28864 ( .A1(n32678), .A2(n32794), .B1(n32786), .B2(n32677), .ZN(
        n32679) );
  XNOR2HSV4 U28865 ( .A1(n47383), .A2(n47382), .ZN(n25887) );
  NAND2HSV4 U28866 ( .A1(n51230), .A2(n51229), .ZN(n52668) );
  NOR2HSV2 U28867 ( .A1(n30440), .A2(n31122), .ZN(n30306) );
  INAND2HSV2 U28868 ( .A1(n30421), .B1(n30780), .ZN(n30507) );
  NAND2HSV0 U28869 ( .A1(n53198), .A2(n53197), .ZN(n53209) );
  NAND2HSV0 U28870 ( .A1(n53198), .A2(n51200), .ZN(n51271) );
  XNOR2HSV2 U28871 ( .A1(n39575), .A2(n39574), .ZN(n39715) );
  CLKNHSV0 U28872 ( .I(n39574), .ZN(n39243) );
  CLKNAND2HSV2 U28873 ( .A1(n44662), .A2(n44663), .ZN(n51411) );
  MUX2NHSV2 U28874 ( .I0(n29847), .I1(n28446), .S(n28450), .ZN(n29945) );
  MUX2NHSV1 U28875 ( .I0(n28447), .I1(n29876), .S(n28449), .ZN(n28450) );
  NAND2HSV4 U28876 ( .A1(n45777), .A2(n45776), .ZN(n45930) );
  NAND2HSV0 U28877 ( .A1(n58145), .A2(n28877), .ZN(n26598) );
  AOI21HSV2 U28878 ( .A1(n45783), .A2(n45782), .B(n45781), .ZN(n53519) );
  INHSV4 U28879 ( .I(n55226), .ZN(n54159) );
  OAI21HSV2 U28880 ( .A1(n28327), .A2(n28328), .B(n28329), .ZN(n28330) );
  NAND2HSV0 U28881 ( .A1(n28328), .A2(n28327), .ZN(n28329) );
  INHSV4 U28882 ( .I(n53791), .ZN(n55593) );
  INHSV6 U28883 ( .I(n59732), .ZN(n53791) );
  OAI21HSV2 U28884 ( .A1(n28199), .A2(n28200), .B(n28201), .ZN(n28202) );
  NAND2HSV0 U28885 ( .A1(n28200), .A2(n28199), .ZN(n28201) );
  XNOR2HSV4 U28886 ( .A1(n26074), .A2(n26073), .ZN(n25888) );
  INHSV2 U28887 ( .I(\pe3/ctrq ), .ZN(n25889) );
  NOR2HSV4 U28888 ( .A1(n36730), .A2(n36720), .ZN(n36723) );
  CLKNAND2HSV2 U28889 ( .A1(n46095), .A2(n46094), .ZN(n46096) );
  INHSV4 U28890 ( .I(n36751), .ZN(n59347) );
  CLKNAND2HSV4 U28891 ( .A1(n44680), .A2(n45506), .ZN(n44674) );
  NOR2HSV2 U28892 ( .A1(n56420), .A2(n25993), .ZN(n25992) );
  CLKNAND2HSV4 U28893 ( .A1(n26071), .A2(n45935), .ZN(n46118) );
  XNOR2HSV1 U28894 ( .A1(n26288), .A2(n26287), .ZN(n29474) );
  INAND2HSV2 U28895 ( .A1(n43372), .B1(n26119), .ZN(n26118) );
  CLKXOR2HSV4 U28896 ( .A1(n43118), .A2(n43117), .Z(n25890) );
  NAND2HSV2 U28897 ( .A1(n43236), .A2(n29750), .ZN(n43117) );
  INHSV2 U28898 ( .I(n43133), .ZN(n46532) );
  CLKNAND2HSV4 U28899 ( .A1(n43028), .A2(n43027), .ZN(n43621) );
  INHSV4 U28900 ( .I(n43129), .ZN(n43142) );
  XNOR2HSV1 U28901 ( .A1(n25942), .A2(n25941), .ZN(pov3[9]) );
  NAND3HSV4 U28902 ( .A1(n29641), .A2(n37167), .A3(n37414), .ZN(n37261) );
  NOR2HSV2 U28903 ( .A1(n36858), .A2(n37454), .ZN(n36776) );
  XNOR2HSV2 U28904 ( .A1(n36884), .A2(n36883), .ZN(n36909) );
  INHSV2 U28905 ( .I(n45769), .ZN(n45767) );
  NOR2HSV4 U28906 ( .A1(n43245), .A2(n43244), .ZN(n43358) );
  CLKNHSV0 U28907 ( .I(n43453), .ZN(n25892) );
  INHSV2 U28908 ( .I(n25892), .ZN(n25893) );
  CLKBUFHSV2 U28909 ( .I(n57188), .Z(n25894) );
  CLKNAND2HSV2 U28910 ( .A1(n25894), .A2(n58102), .ZN(n57749) );
  CLKNAND2HSV2 U28911 ( .A1(n25894), .A2(n57413), .ZN(n50385) );
  CLKNAND2HSV2 U28912 ( .A1(n25894), .A2(n58314), .ZN(n57887) );
  CLKNAND2HSV0 U28913 ( .A1(n25894), .A2(n58298), .ZN(n28672) );
  CLKNHSV2 U28914 ( .I(n48892), .ZN(n57188) );
  CLKNHSV2 U28915 ( .I(n42797), .ZN(n52792) );
  NOR2HSV4 U28916 ( .A1(n25896), .A2(n25895), .ZN(n42803) );
  NOR2HSV4 U28917 ( .A1(n42802), .A2(n43361), .ZN(n25895) );
  CLKNAND2HSV2 U28918 ( .A1(n42601), .A2(n42617), .ZN(n42607) );
  CLKNAND2HSV2 U28919 ( .A1(n25897), .A2(n42801), .ZN(n25896) );
  NOR2HSV4 U28920 ( .A1(n52791), .A2(n29720), .ZN(n25898) );
  CLKNHSV3 U28921 ( .I(n25901), .ZN(n40000) );
  XNOR2HSV4 U28922 ( .A1(n39994), .A2(n39993), .ZN(n25901) );
  CLKNAND2HSV1 U28923 ( .A1(n25901), .A2(n39998), .ZN(n26769) );
  CLKNAND2HSV2 U28924 ( .A1(n25903), .A2(n25902), .ZN(n25904) );
  CLKNAND2HSV2 U28925 ( .A1(n39700), .A2(n39701), .ZN(n25902) );
  CLKNAND2HSV2 U28926 ( .A1(n25905), .A2(n26501), .ZN(n25903) );
  CLKNHSV4 U28927 ( .I(n39701), .ZN(n25905) );
  XNOR2HSV4 U28928 ( .A1(n25906), .A2(n25904), .ZN(n27808) );
  CLKNHSV2 U28929 ( .I(n27807), .ZN(n25906) );
  NAND2HSV3 U28930 ( .A1(n26755), .A2(n26782), .ZN(n25907) );
  INHSV2 U28931 ( .I(n25909), .ZN(n25908) );
  INHSV2 U28932 ( .I(n25911), .ZN(n25912) );
  CLKNHSV2 U28933 ( .I(n47996), .ZN(n25911) );
  AOI21HSV4 U28934 ( .A1(n25915), .A2(n25914), .B(n25913), .ZN(n31881) );
  MUX2NHSV2 U28935 ( .I0(n31872), .I1(n31871), .S(n31879), .ZN(n25913) );
  CLKNHSV2 U28936 ( .I(n31879), .ZN(n25914) );
  CLKNAND2HSV2 U28937 ( .A1(n47996), .A2(n25917), .ZN(n25916) );
  CLKNHSV2 U28938 ( .I(n32444), .ZN(n25917) );
  CLKNHSV2 U28939 ( .I(n31897), .ZN(n25918) );
  XNOR2HSV4 U28940 ( .A1(n31815), .A2(n31814), .ZN(n47996) );
  AOI31HSV2 U28941 ( .A1(n38635), .A2(n38624), .A3(n25926), .B(n25924), .ZN(
        n25919) );
  NOR2HSV4 U28942 ( .A1(n52815), .A2(n38756), .ZN(n25920) );
  CLKNHSV2 U28943 ( .I(n25922), .ZN(n25921) );
  NOR2HSV4 U28944 ( .A1(n38756), .A2(n38757), .ZN(n38876) );
  XNOR2HSV4 U28945 ( .A1(n38634), .A2(n38633), .ZN(n52815) );
  NOR2HSV4 U28946 ( .A1(n25824), .A2(n52813), .ZN(n38756) );
  CLKNAND2HSV2 U28947 ( .A1(n52812), .A2(n25923), .ZN(n25922) );
  CLKNHSV2 U28948 ( .I(n38757), .ZN(n25923) );
  CLKNHSV2 U28949 ( .I(n25925), .ZN(n25924) );
  CLKNAND2HSV2 U28950 ( .A1(n25927), .A2(n44322), .ZN(n25925) );
  CLKNHSV2 U28951 ( .I(n25928), .ZN(n25926) );
  CLKNHSV2 U28952 ( .I(n38622), .ZN(n25927) );
  CLKNHSV2 U28953 ( .I(n44322), .ZN(n25928) );
  CLKNAND2HSV3 U28954 ( .A1(n59504), .A2(n40972), .ZN(n40673) );
  CLKNAND2HSV4 U28955 ( .A1(n26887), .A2(n26886), .ZN(n59504) );
  INHSV2 U28956 ( .I(n25929), .ZN(n40674) );
  CLKNAND2HSV2 U28957 ( .A1(n40673), .A2(n25930), .ZN(n25929) );
  NOR2HSV4 U28958 ( .A1(n40672), .A2(n40671), .ZN(n25930) );
  XNOR2HSV4 U28959 ( .A1(n40666), .A2(n40665), .ZN(n40672) );
  OAI21HSV4 U28960 ( .A1(n29746), .A2(n45276), .B(n25934), .ZN(n25931) );
  CLKNAND2HSV2 U28961 ( .A1(n47539), .A2(n25933), .ZN(n25932) );
  CLKNHSV2 U28962 ( .I(n38874), .ZN(n25933) );
  OAI22HSV4 U28963 ( .A1(n38870), .A2(n38869), .B1(n38868), .B2(n38867), .ZN(
        n25934) );
  XNOR2HSV4 U28964 ( .A1(n25938), .A2(n25935), .ZN(n32458) );
  OAI21HSV4 U28965 ( .A1(n25937), .A2(n25936), .B(n32411), .ZN(n25935) );
  CLKNAND2HSV2 U28966 ( .A1(n32512), .A2(n32513), .ZN(n25936) );
  CLKBUFHSV2 U28967 ( .I(n25940), .Z(n25939) );
  CLKNAND2HSV3 U28968 ( .A1(n38118), .A2(n38117), .ZN(n39080) );
  CLKNAND2HSV3 U28969 ( .A1(n38113), .A2(n52749), .ZN(n38118) );
  BUFHSV8 U28970 ( .I(n39080), .Z(n25940) );
  CLKNHSV2 U28971 ( .I(n29279), .ZN(n25942) );
  CLKNAND2HSV3 U28972 ( .A1(n25945), .A2(n25944), .ZN(n25943) );
  INHSV2 U28973 ( .I(n44655), .ZN(n25944) );
  INHSV2 U28974 ( .I(n44654), .ZN(n25945) );
  CLKNAND2HSV3 U28975 ( .A1(n48328), .A2(n25948), .ZN(n25946) );
  CLKNHSV4 U28976 ( .I(n40335), .ZN(n25948) );
  INHSV2 U28977 ( .I(n45781), .ZN(n25949) );
  CLKNAND2HSV3 U28978 ( .A1(n25950), .A2(n36982), .ZN(n37104) );
  NAND3HSV4 U28979 ( .A1(n25950), .A2(n36982), .A3(n36981), .ZN(n37101) );
  CLKNAND2HSV4 U28980 ( .A1(n25951), .A2(n36859), .ZN(n42682) );
  NAND3HSV4 U28981 ( .A1(n25882), .A2(n37267), .A3(n42509), .ZN(n25951) );
  CLKNAND2HSV2 U28982 ( .A1(n25951), .A2(n42694), .ZN(n37412) );
  XNOR2HSV1 U28983 ( .A1(n25954), .A2(n25952), .ZN(n33331) );
  CLKNAND2HSV3 U28984 ( .A1(n46611), .A2(n33461), .ZN(n25952) );
  CLKNAND2HSV4 U28985 ( .A1(n25953), .A2(n33201), .ZN(n46611) );
  CLKNAND2HSV3 U28986 ( .A1(n59578), .A2(n34220), .ZN(n25953) );
  XOR3HSV4 U28987 ( .A1(n33329), .A2(n25955), .A3(n33330), .Z(n25954) );
  CLKNHSV2 U28988 ( .I(n45094), .ZN(n45096) );
  XOR2HSV2 U28989 ( .A1(n25958), .A2(n45090), .Z(n25957) );
  XNOR2HSV4 U28990 ( .A1(n45088), .A2(n45087), .ZN(n25958) );
  CLKNAND2HSV4 U28991 ( .A1(n25959), .A2(n43352), .ZN(n43348) );
  NAND3HSV4 U28992 ( .A1(n25959), .A2(n43352), .A3(n43351), .ZN(n43356) );
  NAND3HSV4 U28993 ( .A1(n25960), .A2(n43751), .A3(n43750), .ZN(n45584) );
  NAND2HSV3 U28994 ( .A1(n25960), .A2(n43751), .ZN(pov3[24]) );
  CLKNAND2HSV4 U28995 ( .A1(n26128), .A2(n26124), .ZN(n25961) );
  CLKNAND2HSV2 U28996 ( .A1(n25961), .A2(n43593), .ZN(n43597) );
  CLKNAND2HSV2 U28997 ( .A1(n25962), .A2(n25973), .ZN(n25969) );
  CLKNHSV2 U28998 ( .I(n37147), .ZN(n25972) );
  CLKNAND2HSV2 U28999 ( .A1(n25971), .A2(n25963), .ZN(n25970) );
  OAI21HSV4 U29000 ( .A1(n25975), .A2(n25972), .B(n25964), .ZN(n25963) );
  CLKNAND2HSV2 U29001 ( .A1(n25975), .A2(n37146), .ZN(n25964) );
  CLKNHSV4 U29002 ( .I(n26188), .ZN(n25975) );
  NAND3HSV4 U29003 ( .A1(n25966), .A2(n37147), .A3(n25965), .ZN(n37157) );
  CLKNAND2HSV2 U29004 ( .A1(n25973), .A2(n25974), .ZN(n25965) );
  INAND2HSV4 U29005 ( .A1(n25973), .B1(n25975), .ZN(n25966) );
  CLKNAND2HSV2 U29006 ( .A1(n25968), .A2(n25973), .ZN(n25967) );
  CLKNAND2HSV2 U29007 ( .A1(n25970), .A2(n25969), .ZN(n37162) );
  CLKNHSV2 U29008 ( .I(n25973), .ZN(n25971) );
  CLKNAND2HSV4 U29009 ( .A1(n37106), .A2(n37272), .ZN(n25973) );
  CLKNHSV3 U29010 ( .I(n25979), .ZN(n25976) );
  CLKNHSV0 U29011 ( .I(n36930), .ZN(n36779) );
  OAI21HSV4 U29012 ( .A1(n25980), .A2(n36930), .B(n25977), .ZN(n36857) );
  AOI21HSV4 U29013 ( .A1(n36928), .A2(n25978), .B(n36781), .ZN(n25977) );
  NOR2HSV4 U29014 ( .A1(n36925), .A2(n43880), .ZN(n25978) );
  XNOR2HSV4 U29015 ( .A1(n36750), .A2(n36749), .ZN(n36925) );
  CLKNHSV2 U29016 ( .I(n36747), .ZN(n25979) );
  CLKNAND2HSV2 U29017 ( .A1(n59508), .A2(n56620), .ZN(n50796) );
  CLKNAND2HSV0 U29018 ( .A1(n59508), .A2(\pe3/got [1]), .ZN(n26200) );
  INHSV2 U29019 ( .I(n56682), .ZN(n59508) );
  CLKNHSV3 U29020 ( .I(n30197), .ZN(n26388) );
  AOI21HSV4 U29021 ( .A1(n25985), .A2(n26388), .B(n25984), .ZN(n25983) );
  CLKNAND2HSV2 U29022 ( .A1(n29714), .A2(n30138), .ZN(n30140) );
  NOR2HSV4 U29023 ( .A1(n25853), .A2(n25986), .ZN(n30325) );
  CLKNAND2HSV2 U29024 ( .A1(n30197), .A2(n30196), .ZN(n25986) );
  INHSV2 U29025 ( .I(n27094), .ZN(n25987) );
  NOR2HSV4 U29026 ( .A1(n25987), .A2(n25988), .ZN(n38513) );
  NOR2HSV2 U29027 ( .A1(n27093), .A2(n27092), .ZN(n25988) );
  XNOR2HSV4 U29028 ( .A1(n38614), .A2(n38513), .ZN(n28461) );
  BUFHSV8 U29029 ( .I(n56780), .Z(n25989) );
  CLKNHSV4 U29030 ( .I(n56420), .ZN(n56173) );
  CLKNHSV2 U29031 ( .I(n56780), .ZN(n49403) );
  XNOR2HSV4 U29032 ( .A1(n25991), .A2(n25990), .ZN(n56165) );
  CLKNAND2HSV2 U29033 ( .A1(n25989), .A2(n56171), .ZN(n25990) );
  XOR2HSV2 U29034 ( .A1(n56163), .A2(n25992), .Z(n25991) );
  CLKNHSV2 U29035 ( .I(\pe3/got [20]), .ZN(n25993) );
  NAND3HSV4 U29036 ( .A1(n25994), .A2(n37245), .A3(n37155), .ZN(n37153) );
  CLKNAND2HSV2 U29037 ( .A1(n37151), .A2(n37152), .ZN(n25994) );
  NOR2HSV4 U29038 ( .A1(n25995), .A2(n36782), .ZN(n36787) );
  INHSV4 U29039 ( .I(n36728), .ZN(n25995) );
  XOR3HSV2 U29040 ( .A1(n25999), .A2(n25996), .A3(n36800), .Z(n36801) );
  XNOR2HSV4 U29041 ( .A1(n36790), .A2(\pe3/phq [6]), .ZN(n25998) );
  XNOR2HSV4 U29042 ( .A1(n36798), .A2(n26000), .ZN(n25999) );
  XNOR2HSV4 U29043 ( .A1(n36792), .A2(n36793), .ZN(n26000) );
  NOR2HSV4 U29044 ( .A1(n26001), .A2(n29698), .ZN(n26070) );
  CLKNHSV2 U29045 ( .I(n26002), .ZN(n26003) );
  XNOR2HSV4 U29046 ( .A1(n26184), .A2(n26183), .ZN(n26002) );
  CLKNAND2HSV2 U29047 ( .A1(n26002), .A2(n26822), .ZN(n52697) );
  OAI22HSV4 U29048 ( .A1(n26002), .A2(n26181), .B1(n26180), .B2(n26179), .ZN(
        n26821) );
  XOR2HSV2 U29049 ( .A1(n48016), .A2(n26003), .Z(n60083) );
  CLKNAND2HSV3 U29050 ( .A1(n39426), .A2(n26004), .ZN(n39424) );
  CLKNAND2HSV3 U29051 ( .A1(n39412), .A2(n39411), .ZN(n26004) );
  NAND3HSV1 U29052 ( .A1(n48469), .A2(n48467), .A3(n48468), .ZN(n26354) );
  CLKNAND2HSV2 U29053 ( .A1(n26005), .A2(n26007), .ZN(n48467) );
  CLKNAND2HSV4 U29054 ( .A1(n26006), .A2(n48466), .ZN(n48469) );
  CLKNAND2HSV2 U29055 ( .A1(n38459), .A2(n26008), .ZN(n38463) );
  CLKNHSV2 U29056 ( .I(n38460), .ZN(n26008) );
  XNOR2HSV4 U29057 ( .A1(n26009), .A2(n26963), .ZN(n38460) );
  CLKNHSV2 U29058 ( .I(n26767), .ZN(n26009) );
  CLKNAND2HSV3 U29059 ( .A1(n29513), .A2(n26010), .ZN(n26012) );
  CLKNAND2HSV3 U29060 ( .A1(n26011), .A2(n26013), .ZN(n26010) );
  INHSV1 U29061 ( .I(n29512), .ZN(n26011) );
  XNOR2HSV4 U29062 ( .A1(n29514), .A2(n26012), .ZN(n29515) );
  CLKNHSV2 U29063 ( .I(n29511), .ZN(n26013) );
  XNOR2HSV4 U29064 ( .A1(n27322), .A2(n26014), .ZN(n45593) );
  CLKNAND2HSV2 U29065 ( .A1(n48486), .A2(n45947), .ZN(n26014) );
  CLKNAND2HSV4 U29066 ( .A1(n37349), .A2(n37420), .ZN(n26015) );
  CLKNHSV2 U29067 ( .I(n26015), .ZN(n37435) );
  CLKNHSV4 U29068 ( .I(n45621), .ZN(n37238) );
  XNOR2HSV4 U29069 ( .A1(n26017), .A2(n26016), .ZN(n48893) );
  AOI21HSV4 U29070 ( .A1(n49001), .A2(n37238), .B(n26630), .ZN(n26017) );
  CLKBUFHSV2 U29071 ( .I(n26218), .Z(n26018) );
  MUX2NHSV4 U29072 ( .I0(n26021), .I1(n26019), .S(n33127), .ZN(n33128) );
  CLKNAND2HSV3 U29073 ( .A1(n26218), .A2(n33694), .ZN(n26020) );
  CLKNAND2HSV3 U29074 ( .A1(n26218), .A2(n35274), .ZN(n26021) );
  AOI21HSV4 U29075 ( .A1(n26018), .A2(n26024), .B(n26022), .ZN(n33129) );
  CLKNHSV2 U29076 ( .I(n33109), .ZN(n26023) );
  CLKNHSV2 U29077 ( .I(n26025), .ZN(n26024) );
  CLKNAND2HSV2 U29078 ( .A1(n33108), .A2(n34419), .ZN(n26025) );
  CLKNHSV2 U29079 ( .I(n31816), .ZN(n26027) );
  CLKNHSV2 U29080 ( .I(n26028), .ZN(n40164) );
  CLKNAND2HSV2 U29081 ( .A1(n40166), .A2(n26028), .ZN(n40167) );
  CLKNAND2HSV2 U29082 ( .A1(n40320), .A2(n48741), .ZN(n26028) );
  XNOR2HSV4 U29083 ( .A1(n26031), .A2(n26029), .ZN(n33211) );
  XNOR2HSV4 U29084 ( .A1(n33208), .A2(n26030), .ZN(n26029) );
  CLKNAND2HSV2 U29085 ( .A1(n33897), .A2(n33748), .ZN(n26030) );
  NOR2HSV8 U29086 ( .A1(n26326), .A2(n26032), .ZN(n29698) );
  CLKNHSV4 U29087 ( .I(n26327), .ZN(n26032) );
  CLKNAND2HSV3 U29088 ( .A1(n45584), .A2(n43864), .ZN(n26033) );
  INHSV2 U29089 ( .I(n26035), .ZN(n26802) );
  NAND2HSV4 U29090 ( .A1(n33573), .A2(n33458), .ZN(n26035) );
  CLKNAND2HSV2 U29091 ( .A1(n26035), .A2(n26807), .ZN(n26806) );
  CLKNAND2HSV3 U29092 ( .A1(n26037), .A2(n26036), .ZN(n26038) );
  INHSV2 U29093 ( .I(n42491), .ZN(n26036) );
  NOR2HSV4 U29094 ( .A1(n42331), .A2(n44651), .ZN(n42338) );
  CLKNAND2HSV3 U29095 ( .A1(n26040), .A2(n26039), .ZN(n42336) );
  AOI31HSV2 U29096 ( .A1(n26087), .A2(n60104), .A3(n48312), .B(n42319), .ZN(
        n26039) );
  CLKNAND2HSV3 U29097 ( .A1(n26086), .A2(n26085), .ZN(n26040) );
  XNOR2HSV4 U29098 ( .A1(n42337), .A2(n42336), .ZN(n42491) );
  XNOR2HSV4 U29099 ( .A1(n42201), .A2(n26041), .ZN(n42337) );
  XOR2HSV2 U29100 ( .A1(n42313), .A2(n42314), .Z(n26041) );
  CLKNAND2HSV4 U29101 ( .A1(n42330), .A2(n42326), .ZN(n44650) );
  XNOR2HSV4 U29102 ( .A1(n30587), .A2(n30588), .ZN(n26043) );
  OAI21HSV4 U29103 ( .A1(n33196), .A2(n33195), .B(n25876), .ZN(n33224) );
  NOR2HSV4 U29104 ( .A1(n26048), .A2(n26047), .ZN(n26044) );
  CLKNAND2HSV2 U29105 ( .A1(n26045), .A2(n26046), .ZN(n33195) );
  AOI31HSV2 U29106 ( .A1(n26055), .A2(n26053), .A3(n26054), .B(n26052), .ZN(
        n26045) );
  OAI21HSV4 U29107 ( .A1(n26057), .A2(n26056), .B(n29740), .ZN(n26046) );
  INHSV2 U29108 ( .I(n33292), .ZN(n26055) );
  CLKNAND2HSV2 U29109 ( .A1(n26049), .A2(n33192), .ZN(n26048) );
  CLKNAND2HSV2 U29110 ( .A1(n33194), .A2(n26054), .ZN(n26049) );
  CLKNHSV2 U29111 ( .I(n33198), .ZN(n26051) );
  CLKNHSV2 U29112 ( .I(n33187), .ZN(n26052) );
  CLKNHSV2 U29113 ( .I(n33171), .ZN(n26053) );
  XNOR2HSV4 U29114 ( .A1(n26644), .A2(n33179), .ZN(n26054) );
  CLKNHSV2 U29115 ( .I(n33182), .ZN(n26056) );
  CLKNHSV2 U29116 ( .I(n33183), .ZN(n26057) );
  NOR2HSV4 U29117 ( .A1(n26060), .A2(n26059), .ZN(n26058) );
  CLKNHSV2 U29118 ( .I(n40873), .ZN(n26059) );
  CLKNHSV2 U29119 ( .I(n54729), .ZN(n26060) );
  CLKNHSV2 U29120 ( .I(n26061), .ZN(n37422) );
  AOI21HSV2 U29121 ( .A1(n26062), .A2(n46087), .B(n45756), .ZN(n43914) );
  CLKNHSV2 U29122 ( .I(n45758), .ZN(n26062) );
  INHSV2 U29123 ( .I(n45143), .ZN(n26064) );
  NOR2HSV8 U29124 ( .A1(n45140), .A2(n38344), .ZN(n45264) );
  XOR2HSV4 U29125 ( .A1(n53387), .A2(n45389), .Z(n45140) );
  MUX2NHSV2 U29126 ( .I0(n45271), .I1(n45266), .S(n45264), .ZN(n45410) );
  CLKNHSV2 U29127 ( .I(n45143), .ZN(n45266) );
  NOR2HSV4 U29128 ( .A1(n26064), .A2(n45099), .ZN(n45271) );
  CLKNHSV0 U29129 ( .I(n26066), .ZN(n52841) );
  CLKNHSV2 U29130 ( .I(n26419), .ZN(n26065) );
  CLKBUFHSV2 U29131 ( .I(n54729), .Z(n26067) );
  OAI21HSV4 U29132 ( .A1(n42347), .A2(n26069), .B(n26068), .ZN(n54729) );
  CLKNHSV2 U29133 ( .I(n29760), .ZN(n26069) );
  CLKNAND2HSV2 U29134 ( .A1(n54729), .A2(n59994), .ZN(n26699) );
  XNOR2HSV4 U29135 ( .A1(n46118), .A2(n46116), .ZN(n46560) );
  XNOR2HSV4 U29136 ( .A1(n26074), .A2(n26073), .ZN(n46561) );
  NAND3HSV4 U29137 ( .A1(n46111), .A2(n46110), .A3(n46109), .ZN(n26073) );
  XNOR2HSV4 U29138 ( .A1(n26078), .A2(n26075), .ZN(n42324) );
  XOR3HSV2 U29139 ( .A1(n26077), .A2(n26076), .A3(n42185), .Z(n26075) );
  XNOR2HSV4 U29140 ( .A1(n42184), .A2(n42183), .ZN(n26076) );
  CLKNAND2HSV2 U29141 ( .A1(n59377), .A2(\pe1/got [28]), .ZN(n26077) );
  CLKNHSV2 U29142 ( .I(n26737), .ZN(n26079) );
  CLKNHSV2 U29143 ( .I(n26081), .ZN(n26080) );
  CLKNAND2HSV2 U29144 ( .A1(n31364), .A2(n32783), .ZN(n26081) );
  NAND3HSV4 U29145 ( .A1(n31365), .A2(n29670), .A3(n26082), .ZN(n31579) );
  NAND3HSV4 U29146 ( .A1(n31392), .A2(n31348), .A3(n31358), .ZN(n26082) );
  CLKNAND2HSV2 U29147 ( .A1(n38607), .A2(n38890), .ZN(n26083) );
  XNOR2HSV4 U29148 ( .A1(n38464), .A2(n26084), .ZN(n38607) );
  AOI21HSV4 U29149 ( .A1(n38453), .A2(n38452), .B(n38451), .ZN(n38464) );
  CLKNAND2HSV3 U29150 ( .A1(n29760), .A2(n42315), .ZN(n26085) );
  CLKNHSV2 U29151 ( .I(n44827), .ZN(n26088) );
  CLKNHSV2 U29152 ( .I(n54037), .ZN(n55229) );
  XNOR2HSV4 U29153 ( .A1(n26096), .A2(n26090), .ZN(n42058) );
  XNOR2HSV4 U29154 ( .A1(n26095), .A2(n26091), .ZN(n26090) );
  XNOR2HSV4 U29155 ( .A1(n26094), .A2(n26092), .ZN(n26091) );
  XNOR2HSV4 U29156 ( .A1(n26093), .A2(n42027), .ZN(n26092) );
  CLKNHSV2 U29157 ( .I(n42028), .ZN(n26093) );
  CLKNAND2HSV2 U29158 ( .A1(n53768), .A2(\pe1/got [25]), .ZN(n26094) );
  INAND2HSV4 U29159 ( .A1(n54037), .B1(n41689), .ZN(n26095) );
  CLKNAND2HSV2 U29160 ( .A1(n48336), .A2(n59374), .ZN(n26096) );
  CLKNAND2HSV2 U29161 ( .A1(n53656), .A2(n53655), .ZN(n48336) );
  CLKNAND2HSV2 U29162 ( .A1(pov1[23]), .A2(n42202), .ZN(n53656) );
  CLKNAND2HSV3 U29163 ( .A1(n60020), .A2(n38383), .ZN(n26099) );
  INAND2HSV4 U29164 ( .A1(n45091), .B1(n38383), .ZN(n26097) );
  BUFHSV8 U29165 ( .I(n38903), .Z(n26098) );
  CLKNAND2HSV4 U29166 ( .A1(n26099), .A2(n38470), .ZN(n38903) );
  XNOR2HSV4 U29167 ( .A1(n26101), .A2(n26100), .ZN(n51445) );
  NAND3HSV4 U29168 ( .A1(n26102), .A2(n26251), .A3(n26250), .ZN(n26100) );
  XNOR2HSV4 U29169 ( .A1(n26105), .A2(n26104), .ZN(n26101) );
  XNOR2HSV4 U29170 ( .A1(n26249), .A2(n26248), .ZN(n26105) );
  INHSV2 U29171 ( .I(n26106), .ZN(n40336) );
  AOI21HSV4 U29172 ( .A1(n26268), .A2(n26267), .B(n26272), .ZN(n26107) );
  CLKNAND2HSV4 U29173 ( .A1(n26271), .A2(n26270), .ZN(n40361) );
  INHSV1 U29174 ( .I(n40424), .ZN(n40567) );
  CLKNHSV2 U29175 ( .I(n40393), .ZN(n26108) );
  CLKNHSV4 U29176 ( .I(n31970), .ZN(n26109) );
  INHSV2 U29177 ( .I(n32166), .ZN(n26110) );
  CLKNHSV2 U29178 ( .I(n31970), .ZN(n26114) );
  INAND2HSV4 U29179 ( .A1(n31970), .B1(n26111), .ZN(n32021) );
  CLKNHSV2 U29180 ( .I(n31971), .ZN(n26111) );
  CLKNAND2HSV2 U29181 ( .A1(n26114), .A2(n26112), .ZN(n32303) );
  CLKNHSV2 U29182 ( .I(n46750), .ZN(n26112) );
  CLKNAND2HSV2 U29183 ( .A1(n26114), .A2(n26113), .ZN(n32398) );
  CLKNHSV2 U29184 ( .I(n32631), .ZN(n26113) );
  CLKNAND2HSV2 U29185 ( .A1(n26114), .A2(\pe6/got [7]), .ZN(n27377) );
  CLKNHSV4 U29186 ( .I(n44668), .ZN(n45508) );
  XNOR2HSV4 U29187 ( .A1(n43903), .A2(n43906), .ZN(n44668) );
  XNOR2HSV4 U29188 ( .A1(n26118), .A2(n26115), .ZN(n43465) );
  XNOR2HSV4 U29189 ( .A1(n26117), .A2(n26116), .ZN(n26115) );
  CLKNAND2HSV2 U29190 ( .A1(n43463), .A2(n42936), .ZN(n26116) );
  XNOR2HSV4 U29191 ( .A1(n43462), .A2(n43461), .ZN(n26117) );
  CLKNHSV2 U29192 ( .I(n43371), .ZN(n26119) );
  NOR2HSV4 U29193 ( .A1(n43143), .A2(n43142), .ZN(n43372) );
  CLKNHSV2 U29194 ( .I(n26213), .ZN(n26120) );
  NAND2HSV2 U29195 ( .A1(n45794), .A2(n26122), .ZN(n26132) );
  NOR2HSV4 U29196 ( .A1(n26213), .A2(n26133), .ZN(n26122) );
  CLKNAND2HSV2 U29197 ( .A1(n45794), .A2(n26123), .ZN(n26129) );
  CLKNHSV2 U29198 ( .I(n26209), .ZN(n26123) );
  AOI22HSV4 U29199 ( .A1(n26127), .A2(n26211), .B1(n26126), .B2(n26125), .ZN(
        n26124) );
  CLKNHSV2 U29200 ( .I(n26209), .ZN(n26125) );
  CLKNAND2HSV2 U29201 ( .A1(n45794), .A2(n43868), .ZN(n26127) );
  OAI21HSV4 U29202 ( .A1(n26131), .A2(n26130), .B(n26129), .ZN(n26128) );
  NOR2HSV4 U29203 ( .A1(n26216), .A2(n26213), .ZN(n26130) );
  CLKNHSV2 U29204 ( .I(n26132), .ZN(n26131) );
  CLKNHSV2 U29205 ( .I(n43868), .ZN(n26133) );
  CLKNAND2HSV3 U29206 ( .A1(n43350), .A2(n43349), .ZN(n26134) );
  CLKNAND2HSV3 U29207 ( .A1(n41330), .A2(n41329), .ZN(n41508) );
  CLKNAND2HSV3 U29208 ( .A1(n60107), .A2(n44649), .ZN(n41330) );
  CLKNAND2HSV2 U29209 ( .A1(n26135), .A2(\pe3/got [22]), .ZN(n29514) );
  CLKNAND2HSV2 U29210 ( .A1(n26135), .A2(n56675), .ZN(n29434) );
  CLKNAND2HSV0 U29211 ( .A1(n26135), .A2(n45755), .ZN(n28357) );
  CLKNHSV2 U29212 ( .I(n49403), .ZN(n26135) );
  CLKNAND2HSV1 U29213 ( .A1(n45406), .A2(n36562), .ZN(n26139) );
  CLKNAND2HSV3 U29214 ( .A1(n26143), .A2(n26140), .ZN(n29989) );
  NOR2HSV4 U29215 ( .A1(n26142), .A2(n26141), .ZN(n26140) );
  CLKNAND2HSV2 U29216 ( .A1(n30016), .A2(n30139), .ZN(n26142) );
  CLKNAND2HSV2 U29217 ( .A1(n29885), .A2(n29884), .ZN(n26143) );
  CLKNAND2HSV3 U29218 ( .A1(n29989), .A2(n26145), .ZN(n26144) );
  NOR2HSV3 U29219 ( .A1(n26147), .A2(n26146), .ZN(n26145) );
  INHSV2 U29220 ( .I(n39398), .ZN(n26146) );
  INHSV2 U29221 ( .I(n29988), .ZN(n26147) );
  CLKNHSV2 U29222 ( .I(n44526), .ZN(n26532) );
  CLKNAND2HSV2 U29223 ( .A1(n26150), .A2(n48326), .ZN(n44526) );
  XNOR2HSV4 U29224 ( .A1(n42483), .A2(n48329), .ZN(n60015) );
  CLKNHSV2 U29225 ( .I(n44523), .ZN(n26149) );
  NOR2HSV4 U29226 ( .A1(n48325), .A2(n44521), .ZN(n26150) );
  XNOR2HSV4 U29227 ( .A1(n42486), .A2(n42485), .ZN(n48325) );
  CLKNAND2HSV2 U29228 ( .A1(n26151), .A2(\pe3/got [24]), .ZN(n55935) );
  CLKNAND2HSV2 U29229 ( .A1(n26151), .A2(n56421), .ZN(n56549) );
  CLKNAND2HSV2 U29230 ( .A1(n26151), .A2(n56618), .ZN(n56670) );
  CLKNAND2HSV0 U29231 ( .A1(n26151), .A2(n56342), .ZN(n53278) );
  CLKNHSV2 U29232 ( .I(n26152), .ZN(n44330) );
  CLKNAND2HSV2 U29233 ( .A1(n26152), .A2(n46289), .ZN(n36021) );
  CLKNHSV2 U29234 ( .I(n40338), .ZN(n41720) );
  NOR2HSV4 U29235 ( .A1(n40338), .A2(\pe1/ti_7t [1]), .ZN(n40339) );
  CLKNHSV2 U29236 ( .I(n30085), .ZN(n30074) );
  CLKNAND2HSV1 U29237 ( .A1(n30085), .A2(n30083), .ZN(n30076) );
  XNOR2HSV4 U29238 ( .A1(n29987), .A2(n29986), .ZN(n30085) );
  INHSV24 U29239 ( .I(n26163), .ZN(n26153) );
  INHSV24 U29240 ( .I(n30331), .ZN(n26154) );
  XNOR2HSV4 U29241 ( .A1(n26393), .A2(n26390), .ZN(n47988) );
  NAND3HSV4 U29242 ( .A1(n26158), .A2(n26156), .A3(n26155), .ZN(n26167) );
  CLKNAND2HSV2 U29243 ( .A1(n30329), .A2(n26162), .ZN(n26155) );
  CLKNHSV2 U29244 ( .I(n26157), .ZN(n26156) );
  MOAI22HSV4 U29245 ( .A1(n30328), .A2(n26165), .B1(n26154), .B2(n26153), .ZN(
        n26157) );
  CLKNAND2HSV1 U29246 ( .A1(n47988), .A2(n30330), .ZN(n26168) );
  NOR3HSV4 U29247 ( .A1(n26160), .A2(n30329), .A3(n26159), .ZN(n47990) );
  CLKNHSV2 U29248 ( .I(n26161), .ZN(n26159) );
  NOR2HSV4 U29249 ( .A1(n30328), .A2(n30051), .ZN(n26160) );
  CLKNHSV2 U29250 ( .I(n26164), .ZN(n26161) );
  CLKNHSV2 U29251 ( .I(n30331), .ZN(n26162) );
  NOR2HSV4 U29252 ( .A1(n26164), .A2(n39245), .ZN(n26163) );
  NOR2HSV4 U29253 ( .A1(n30327), .A2(n39733), .ZN(n26164) );
  CLKNHSV2 U29254 ( .I(n26166), .ZN(n26165) );
  NOR2HSV4 U29255 ( .A1(n30331), .A2(n30051), .ZN(n26166) );
  OAI21HSV4 U29256 ( .A1(n47990), .A2(n26168), .B(n26167), .ZN(n30780) );
  CLKNAND2HSV4 U29257 ( .A1(n43741), .A2(n43740), .ZN(n26169) );
  AOI21HSV4 U29258 ( .A1(n43738), .A2(n26169), .B(n43486), .ZN(n43903) );
  NAND2HSV2 U29259 ( .A1(\pe1/bq[29] ), .A2(\pe1/aot [32]), .ZN(n26170) );
  CLKNHSV2 U29260 ( .I(n40558), .ZN(n40342) );
  INAND2HSV4 U29261 ( .A1(n40558), .B1(n26171), .ZN(n40413) );
  CLKNHSV2 U29262 ( .I(n40787), .ZN(n26171) );
  XNOR2HSV4 U29263 ( .A1(n26173), .A2(n26172), .ZN(n40326) );
  XNOR2HSV4 U29264 ( .A1(n40413), .A2(n26174), .ZN(n26173) );
  CLKNHSV2 U29265 ( .I(n40787), .ZN(n40488) );
  CLKNHSV2 U29266 ( .I(n33564), .ZN(n33263) );
  CLKNHSV4 U29267 ( .I(n32314), .ZN(n26175) );
  CLKNAND2HSV4 U29268 ( .A1(n32336), .A2(n29647), .ZN(n32514) );
  AND2HSV8 U29269 ( .A1(n32316), .A2(n32315), .Z(n29647) );
  CLKNAND2HSV3 U29270 ( .A1(n31969), .A2(n32407), .ZN(n32316) );
  CLKNHSV0 U29271 ( .I(n32314), .ZN(n47974) );
  AOI21HSV4 U29272 ( .A1(n25288), .A2(n26176), .B(n32153), .ZN(n32335) );
  CLKNHSV2 U29273 ( .I(n32051), .ZN(n26176) );
  CLKNAND2HSV3 U29274 ( .A1(n26177), .A2(n26178), .ZN(n33198) );
  INHSV2 U29275 ( .I(n33129), .ZN(n26177) );
  INHSV2 U29276 ( .I(n33128), .ZN(n26178) );
  CLKNHSV2 U29277 ( .I(\pe4/ti_7t [2]), .ZN(n26179) );
  CLKNHSV2 U29278 ( .I(n59997), .ZN(n26180) );
  CLKNHSV2 U29279 ( .I(n33095), .ZN(n26182) );
  XNOR2HSV4 U29280 ( .A1(n33092), .A2(n33091), .ZN(n33153) );
  XOR2HSV2 U29281 ( .A1(n26627), .A2(n26628), .Z(n26183) );
  XNOR2HSV4 U29282 ( .A1(n26629), .A2(n33946), .ZN(n26184) );
  NOR2HSV4 U29283 ( .A1(n26186), .A2(n26185), .ZN(n32926) );
  CLKNHSV2 U29284 ( .I(n32925), .ZN(n26185) );
  CLKNHSV2 U29285 ( .I(n26187), .ZN(n26186) );
  NOR2HSV0 U29286 ( .A1(n26187), .A2(n32047), .ZN(n51447) );
  OAI21HSV4 U29287 ( .A1(n26187), .A2(n32949), .B(n32925), .ZN(n46592) );
  CLKNAND2HSV4 U29288 ( .A1(n32690), .A2(n32691), .ZN(n26187) );
  CLKNHSV2 U29289 ( .I(n25968), .ZN(n26188) );
  CLKNAND2HSV2 U29290 ( .A1(n32684), .A2(n32683), .ZN(n32959) );
  OAI21HSV4 U29291 ( .A1(n35781), .A2(n35784), .B(n26189), .ZN(n35787) );
  MUX2NHSV2 U29292 ( .I0(n35780), .I1(n31903), .S(n35779), .ZN(n26189) );
  XNOR2HSV4 U29293 ( .A1(n26190), .A2(n35776), .ZN(n35779) );
  CLKNAND2HSV2 U29294 ( .A1(n36102), .A2(n32354), .ZN(n26190) );
  CLKNAND2HSV2 U29295 ( .A1(n47951), .A2(n33089), .ZN(n35784) );
  CLKNHSV2 U29296 ( .I(\pe4/ti_1 ), .ZN(n33118) );
  XNOR2HSV4 U29297 ( .A1(n33092), .A2(n33091), .ZN(n29766) );
  MUX2NHSV2 U29298 ( .I0(n28876), .I1(\pe4/phq [1]), .S(n26191), .ZN(n33091)
         );
  XNOR2HSV4 U29299 ( .A1(n26193), .A2(n26192), .ZN(n33092) );
  NOR2HSV4 U29300 ( .A1(n33090), .A2(n26194), .ZN(n26193) );
  CLKNHSV2 U29301 ( .I(\pe4/pvq [1]), .ZN(n26194) );
  CLKNAND2HSV3 U29302 ( .A1(n41472), .A2(n40873), .ZN(n26196) );
  CLKNAND2HSV2 U29303 ( .A1(n40552), .A2(n40636), .ZN(n26195) );
  XNOR2HSV4 U29304 ( .A1(n40578), .A2(n40577), .ZN(n26197) );
  CLKNAND2HSV2 U29305 ( .A1(n59441), .A2(n56176), .ZN(n56732) );
  CLKNAND2HSV2 U29306 ( .A1(n56817), .A2(n56888), .ZN(n56890) );
  CLKNAND2HSV2 U29307 ( .A1(n56058), .A2(n56908), .ZN(n56978) );
  CLKNAND2HSV0 U29308 ( .A1(n59441), .A2(n55940), .ZN(n55941) );
  CLKNHSV2 U29309 ( .I(n56854), .ZN(n59441) );
  XOR2HSV2 U29310 ( .A1(n56947), .A2(n26198), .Z(n56951) );
  XOR3HSV2 U29311 ( .A1(n56946), .A2(n26200), .A3(n26199), .Z(n26198) );
  CLKNAND2HSV2 U29312 ( .A1(n48480), .A2(n56908), .ZN(n26199) );
  CLKNAND2HSV4 U29313 ( .A1(n60105), .A2(n41410), .ZN(n41708) );
  MUX2NHSV4 U29314 ( .I0(n41590), .I1(n29207), .S(n29209), .ZN(n60105) );
  CLKNHSV2 U29315 ( .I(n26204), .ZN(n41922) );
  XNOR2HSV4 U29316 ( .A1(n41830), .A2(n41829), .ZN(n26204) );
  AOI21HSV4 U29317 ( .A1(n26204), .A2(n41917), .B(n41916), .ZN(n42041) );
  XNOR2HSV4 U29318 ( .A1(n26205), .A2(n29442), .ZN(n29443) );
  NOR2HSV4 U29319 ( .A1(n33155), .A2(n33154), .ZN(n26206) );
  OAI21HSV4 U29320 ( .A1(n29766), .A2(n33339), .B(n33152), .ZN(n33154) );
  XNOR2HSV4 U29321 ( .A1(n26207), .A2(n33106), .ZN(n33155) );
  XNOR2HSV4 U29322 ( .A1(n33102), .A2(n33101), .ZN(n26207) );
  CLKNHSV2 U29323 ( .I(n42044), .ZN(n26208) );
  CLKNHSV4 U29324 ( .I(n46588), .ZN(n33070) );
  XNOR2HSV4 U29325 ( .A1(n33071), .A2(n33070), .ZN(n33084) );
  CLKNHSV2 U29326 ( .I(n26215), .ZN(n26216) );
  CLKNAND2HSV2 U29327 ( .A1(n56265), .A2(n26210), .ZN(n26215) );
  CLKNHSV2 U29328 ( .I(n26217), .ZN(n26210) );
  NOR2HSV4 U29329 ( .A1(n26215), .A2(n26212), .ZN(n26211) );
  XNOR2HSV4 U29330 ( .A1(n43589), .A2(n26214), .ZN(n26213) );
  CLKNHSV2 U29331 ( .I(n43590), .ZN(n26214) );
  CLKNAND2HSV2 U29332 ( .A1(n26215), .A2(n43868), .ZN(n26209) );
  CLKNHSV2 U29333 ( .I(n37169), .ZN(n26217) );
  BUFHSV8 U29334 ( .I(n33157), .Z(n26218) );
  INHSV2 U29335 ( .I(n26821), .ZN(n26219) );
  CLKNHSV4 U29336 ( .I(n32157), .ZN(n29757) );
  CLKNAND2HSV4 U29337 ( .A1(n32325), .A2(n26220), .ZN(n32158) );
  CLKNHSV2 U29338 ( .I(n26518), .ZN(n26220) );
  XNOR2HSV4 U29339 ( .A1(n32050), .A2(n32049), .ZN(n32314) );
  CLKNHSV2 U29340 ( .I(n33157), .ZN(n33172) );
  XNOR2HSV4 U29341 ( .A1(n33155), .A2(n33107), .ZN(n33108) );
  CLKNHSV2 U29342 ( .I(n44675), .ZN(n26221) );
  CLKNAND2HSV2 U29343 ( .A1(n44676), .A2(n26223), .ZN(n26222) );
  CLKNHSV2 U29344 ( .I(n36980), .ZN(n26223) );
  NAND2HSV2 U29345 ( .A1(n43902), .A2(n43903), .ZN(n26225) );
  XNOR2HSV4 U29346 ( .A1(n26230), .A2(n26226), .ZN(n33442) );
  XNOR2HSV4 U29347 ( .A1(n33441), .A2(n26227), .ZN(n26226) );
  XNOR2HSV4 U29348 ( .A1(n26229), .A2(n26228), .ZN(n26227) );
  CLKNAND2HSV2 U29349 ( .A1(n46611), .A2(n33748), .ZN(n26228) );
  XOR3HSV2 U29350 ( .A1(n33440), .A2(n33439), .A3(n33438), .Z(n26229) );
  CLKNAND2HSV2 U29351 ( .A1(n33413), .A2(n57208), .ZN(n26230) );
  NAND3HSV4 U29352 ( .A1(n26232), .A2(n33346), .A3(n26231), .ZN(n33413) );
  CLKNHSV2 U29353 ( .I(n33343), .ZN(n26232) );
  CLKNAND2HSV2 U29354 ( .A1(n25761), .A2(n26233), .ZN(n43735) );
  CLKNHSV2 U29355 ( .I(n43734), .ZN(n26234) );
  CLKNHSV2 U29356 ( .I(n39679), .ZN(n39686) );
  XOR2HSV2 U29357 ( .A1(n39678), .A2(n39393), .Z(n39679) );
  CLKNAND2HSV2 U29358 ( .A1(n39401), .A2(n39408), .ZN(n39678) );
  NOR2HSV4 U29359 ( .A1(n39404), .A2(n29724), .ZN(n39401) );
  NAND3HSV2 U29360 ( .A1(n44949), .A2(n45108), .A3(n45092), .ZN(n45286) );
  CLKNAND2HSV3 U29361 ( .A1(n44173), .A2(n45113), .ZN(n45092) );
  CLKNAND2HSV2 U29362 ( .A1(n44709), .A2(n44824), .ZN(n26245) );
  CLKNHSV2 U29363 ( .I(n26237), .ZN(n44822) );
  CLKNAND2HSV2 U29364 ( .A1(n26243), .A2(n26239), .ZN(n26237) );
  CLKNHSV2 U29365 ( .I(n26238), .ZN(n44823) );
  CLKNAND2HSV2 U29366 ( .A1(n26241), .A2(n26240), .ZN(n26238) );
  CLKNHSV2 U29367 ( .I(n44821), .ZN(n26239) );
  INAND2HSV4 U29368 ( .A1(n26244), .B1(n44828), .ZN(n26240) );
  NOR2HSV4 U29369 ( .A1(n44828), .A2(n26246), .ZN(n26242) );
  CLKNHSV2 U29370 ( .I(n26245), .ZN(n44829) );
  CLKNHSV2 U29371 ( .I(n45280), .ZN(n45282) );
  CLKNHSV2 U29372 ( .I(n36320), .ZN(n26244) );
  CLKNHSV2 U29373 ( .I(n44709), .ZN(n26246) );
  INAND2HSV4 U29374 ( .A1(n31903), .B1(n26247), .ZN(n31880) );
  INAND2HSV4 U29375 ( .A1(n31904), .B1(n26247), .ZN(n31962) );
  CLKNAND2HSV2 U29376 ( .A1(n26109), .A2(n59292), .ZN(n58890) );
  CLKNAND2HSV0 U29377 ( .A1(n26247), .A2(n58724), .ZN(n58778) );
  CLKNHSV8 U29378 ( .I(n31970), .ZN(n26247) );
  NAND2HSV2 U29379 ( .A1(n47996), .A2(n26255), .ZN(n26253) );
  CLKXOR2HSV4 U29380 ( .A1(n31813), .A2(n31812), .Z(n26248) );
  AOI21HSV4 U29381 ( .A1(n51441), .A2(n31876), .B(n31767), .ZN(n26249) );
  CLKNAND2HSV2 U29382 ( .A1(n26255), .A2(n26257), .ZN(n26250) );
  CLKNAND2HSV2 U29383 ( .A1(n31898), .A2(n26252), .ZN(n26251) );
  CLKNHSV2 U29384 ( .I(n26253), .ZN(n26252) );
  CLKNHSV2 U29385 ( .I(n26256), .ZN(n26255) );
  NOR2HSV4 U29386 ( .A1(n31761), .A2(n32685), .ZN(n26256) );
  CLKNHSV2 U29387 ( .I(n31760), .ZN(n26257) );
  INAND2HSV4 U29388 ( .A1(n26260), .B1(n44665), .ZN(n26258) );
  CLKNHSV2 U29389 ( .I(n44664), .ZN(n26260) );
  CLKNAND2HSV2 U29390 ( .A1(n36222), .A2(n26261), .ZN(n36223) );
  CLKNAND2HSV1 U29391 ( .A1(n26261), .A2(n46568), .ZN(n36235) );
  XNOR2HSV4 U29392 ( .A1(n44375), .A2(n47933), .ZN(n26261) );
  CLKNHSV2 U29393 ( .I(n59504), .ZN(n40594) );
  CLKNAND2HSV2 U29394 ( .A1(n59504), .A2(n41134), .ZN(n40718) );
  CLKNHSV4 U29395 ( .I(n39002), .ZN(n26263) );
  NOR2HSV2 U29396 ( .A1(n52827), .A2(n44156), .ZN(n44158) );
  NOR2HSV8 U29397 ( .A1(n26266), .A2(n26265), .ZN(n26413) );
  CLKNAND2HSV4 U29398 ( .A1(n26637), .A2(n26636), .ZN(n26265) );
  CLKNHSV4 U29399 ( .I(n26632), .ZN(n26266) );
  AOI21HSV4 U29400 ( .A1(n40367), .A2(n40365), .B(n26605), .ZN(n26267) );
  NOR3HSV4 U29401 ( .A1(n40363), .A2(n26606), .A3(n40362), .ZN(n26268) );
  CLKNHSV2 U29402 ( .I(n40424), .ZN(n26269) );
  NAND3HSV3 U29403 ( .A1(n60110), .A2(n51113), .A3(n40331), .ZN(n26270) );
  CLKNHSV3 U29404 ( .I(n40334), .ZN(n26271) );
  CLKNHSV2 U29405 ( .I(n26607), .ZN(n26272) );
  XOR3HSV2 U29406 ( .A1(n26274), .A2(n55338), .A3(n26273), .Z(\pe1/poht [19])
         );
  XNOR2HSV4 U29407 ( .A1(n55336), .A2(n26275), .ZN(n26274) );
  XOR2HSV2 U29408 ( .A1(n26277), .A2(n26276), .Z(n26275) );
  XNOR2HSV4 U29409 ( .A1(n55333), .A2(n26278), .ZN(n26277) );
  XOR2HSV2 U29410 ( .A1(n55335), .A2(n55334), .Z(n26278) );
  CLKNHSV2 U29411 ( .I(n42343), .ZN(n47936) );
  NAND3HSV4 U29412 ( .A1(n53368), .A2(n60015), .A3(n42484), .ZN(n44527) );
  XNOR2HSV4 U29413 ( .A1(n42486), .A2(n42485), .ZN(n53368) );
  AOI21HSV4 U29414 ( .A1(n26283), .A2(n26282), .B(n26280), .ZN(n42485) );
  CLKNAND2HSV0 U29415 ( .A1(n42489), .A2(n42327), .ZN(n26281) );
  CLKNHSV2 U29416 ( .I(n42199), .ZN(n26284) );
  INHSV2 U29417 ( .I(n26286), .ZN(n39697) );
  XNOR2HSV4 U29418 ( .A1(n39715), .A2(n39714), .ZN(n26286) );
  NAND3HSV4 U29419 ( .A1(n26286), .A2(n39580), .A3(n39581), .ZN(n39698) );
  INAND2HSV4 U29420 ( .A1(n39697), .B1(n39732), .ZN(n39736) );
  NOR2HSV4 U29421 ( .A1(n43372), .A2(n36721), .ZN(n26287) );
  CLKNHSV2 U29422 ( .I(n25890), .ZN(n26288) );
  CLKNHSV2 U29423 ( .I(n29746), .ZN(n52534) );
  XNOR2HSV4 U29424 ( .A1(n26291), .A2(n26289), .ZN(n44024) );
  XNOR2HSV4 U29425 ( .A1(n44021), .A2(n26290), .ZN(n26289) );
  INAND2HSV4 U29426 ( .A1(n29746), .B1(n38723), .ZN(n26290) );
  CLKNAND2HSV2 U29427 ( .A1(n51687), .A2(n38327), .ZN(n26291) );
  INAND2HSV4 U29428 ( .A1(n26293), .B1(n26292), .ZN(n51687) );
  CLKNAND2HSV2 U29429 ( .A1(n60021), .A2(n44309), .ZN(n26292) );
  CLKNHSV2 U29430 ( .I(n43923), .ZN(n26293) );
  INHSV2 U29431 ( .I(n54635), .ZN(n55576) );
  XOR2HSV2 U29432 ( .A1(n26298), .A2(n26295), .Z(n26294) );
  XNOR2HSV4 U29433 ( .A1(n26297), .A2(n26296), .ZN(n26295) );
  XNOR2HSV4 U29434 ( .A1(n55371), .A2(n55370), .ZN(n26296) );
  CLKNAND2HSV2 U29435 ( .A1(n55332), .A2(n55448), .ZN(n26297) );
  NOR2HSV2 U29436 ( .A1(n54635), .A2(n26299), .ZN(n26298) );
  CLKNHSV2 U29437 ( .I(n59750), .ZN(n26299) );
  AOI31HSV2 U29438 ( .A1(n44823), .A2(n44822), .A3(n26301), .B(n26300), .ZN(
        n26302) );
  CLKNHSV2 U29439 ( .I(n26306), .ZN(n26300) );
  CLKNHSV2 U29440 ( .I(n38375), .ZN(n26303) );
  NAND2HSV2 U29441 ( .A1(n26407), .A2(n26305), .ZN(n26304) );
  CLKNHSV2 U29442 ( .I(n45280), .ZN(n26305) );
  CLKNHSV2 U29443 ( .I(n45146), .ZN(n26306) );
  CLKNHSV2 U29444 ( .I(\pe4/got [31]), .ZN(n33189) );
  CLKNHSV4 U29445 ( .I(n26339), .ZN(n29668) );
  CLKNAND2HSV4 U29446 ( .A1(n31677), .A2(n26308), .ZN(n26339) );
  CLKNAND2HSV4 U29447 ( .A1(n31627), .A2(n31628), .ZN(n31625) );
  CLKNHSV2 U29448 ( .I(n26309), .ZN(n26308) );
  INHSV24 U29449 ( .I(n31533), .ZN(n26309) );
  XNOR2HSV4 U29450 ( .A1(n26314), .A2(n26310), .ZN(n40166) );
  XNOR2HSV4 U29451 ( .A1(n26311), .A2(n39865), .ZN(n26310) );
  XNOR2HSV4 U29452 ( .A1(n26313), .A2(n26312), .ZN(n26311) );
  XNOR2HSV4 U29453 ( .A1(n39863), .A2(n39864), .ZN(n26312) );
  CLKNAND2HSV2 U29454 ( .A1(n45499), .A2(\pe5/got [28]), .ZN(n26313) );
  AOI22HSV4 U29455 ( .A1(\pe5/ti_7t [28]), .A2(n40007), .B1(n40010), .B2(
        n40006), .ZN(n40294) );
  CLKNHSV2 U29456 ( .I(n30441), .ZN(n30515) );
  CLKNAND2HSV2 U29457 ( .A1(n26316), .A2(n26315), .ZN(n30246) );
  MUX2NHSV2 U29458 ( .I0(n30208), .I1(n30209), .S(n26318), .ZN(n26315) );
  MUX2NHSV2 U29459 ( .I0(n30205), .I1(n26320), .S(n26317), .ZN(n26316) );
  CLKNHSV2 U29460 ( .I(n26318), .ZN(n26317) );
  NOR2HSV4 U29461 ( .A1(n30441), .A2(n26319), .ZN(n26318) );
  CLKNHSV2 U29462 ( .I(n30254), .ZN(n26319) );
  CLKNHSV2 U29463 ( .I(n26321), .ZN(n26320) );
  CLKNAND2HSV2 U29464 ( .A1(n60074), .A2(n30299), .ZN(n26321) );
  XNOR2HSV4 U29465 ( .A1(n30068), .A2(n30067), .ZN(n60074) );
  CLKNAND2HSV3 U29466 ( .A1(n60060), .A2(n26322), .ZN(n45925) );
  NOR2HSV2 U29467 ( .A1(n45626), .A2(n45621), .ZN(n26322) );
  CLKNAND2HSV4 U29468 ( .A1(n44689), .A2(n44688), .ZN(n60060) );
  XNOR2HSV4 U29469 ( .A1(n29810), .A2(n26323), .ZN(n29824) );
  XNOR2HSV4 U29470 ( .A1(n26325), .A2(n26324), .ZN(n26323) );
  CLKNAND2HSV2 U29471 ( .A1(n30925), .A2(\pe5/pvq [8]), .ZN(n26324) );
  XNOR2HSV4 U29472 ( .A1(n29809), .A2(\pe5/phq [8]), .ZN(n26325) );
  CLKNAND2HSV3 U29473 ( .A1(n26329), .A2(n26328), .ZN(n26326) );
  CLKNAND2HSV3 U29474 ( .A1(n49253), .A2(n43877), .ZN(n26328) );
  CLKNAND2HSV1 U29475 ( .A1(n43876), .A2(n43875), .ZN(n26329) );
  CLKNAND2HSV2 U29476 ( .A1(\pe3/ti_1 ), .A2(\pe3/got [31]), .ZN(n26330) );
  NOR2HSV4 U29477 ( .A1(n31757), .A2(n48010), .ZN(n31762) );
  NAND3HSV4 U29478 ( .A1(n31694), .A2(n26333), .A3(n26332), .ZN(n26331) );
  CLKNHSV2 U29479 ( .I(n36055), .ZN(n26332) );
  CLKNAND2HSV2 U29480 ( .A1(n31679), .A2(n31680), .ZN(n26333) );
  CLKNAND2HSV0 U29481 ( .A1(\pe3/bq[30] ), .A2(\pe3/aot [32]), .ZN(n36675) );
  CLKNAND2HSV3 U29482 ( .A1(n31470), .A2(n31471), .ZN(n26334) );
  OAI21HSV4 U29483 ( .A1(n26336), .A2(n26337), .B(n26335), .ZN(n31676) );
  CLKNAND2HSV2 U29484 ( .A1(n31470), .A2(n31471), .ZN(n26336) );
  AOI21HSV4 U29485 ( .A1(n31677), .A2(n31531), .B(n31676), .ZN(n26338) );
  CLKNHSV2 U29486 ( .I(n31536), .ZN(n26340) );
  AOI21HSV4 U29487 ( .A1(n26343), .A2(n26342), .B(n43478), .ZN(n43594) );
  CLKNHSV2 U29488 ( .I(n43481), .ZN(n26344) );
  NAND4HSV4 U29489 ( .A1(n26348), .A2(n26345), .A3(n26347), .A4(n29979), .ZN(
        n29982) );
  NAND3HSV4 U29490 ( .A1(n29930), .A2(n29931), .A3(n26346), .ZN(n26345) );
  CLKNHSV2 U29491 ( .I(n37766), .ZN(n26346) );
  CLKNAND2HSV3 U29492 ( .A1(n29977), .A2(n29976), .ZN(n26348) );
  CLKNAND2HSV0 U29493 ( .A1(n55484), .A2(n59756), .ZN(n55603) );
  CLKNAND2HSV3 U29494 ( .A1(n60036), .A2(n41727), .ZN(n26349) );
  CLKNAND2HSV3 U29495 ( .A1(n26535), .A2(n26534), .ZN(n60036) );
  NOR2HSV4 U29496 ( .A1(n26353), .A2(n26350), .ZN(n54631) );
  CLKNAND2HSV2 U29497 ( .A1(n26352), .A2(n26351), .ZN(n26350) );
  CLKNAND2HSV2 U29498 ( .A1(n41242), .A2(\pe1/ti_7t [31]), .ZN(n26351) );
  CLKNAND2HSV2 U29499 ( .A1(n48470), .A2(n48471), .ZN(n26352) );
  MUX2NHSV2 U29500 ( .I0(n26355), .I1(n26354), .S(n60036), .ZN(n26353) );
  CLKNAND2HSV2 U29501 ( .A1(n48470), .A2(n40654), .ZN(n26355) );
  CLKNAND2HSV2 U29502 ( .A1(n48467), .A2(n48469), .ZN(n48470) );
  CLKNAND2HSV3 U29503 ( .A1(n26356), .A2(n29805), .ZN(n29811) );
  INHSV2 U29504 ( .I(n29803), .ZN(n26356) );
  CLKNAND2HSV3 U29505 ( .A1(n26358), .A2(n26357), .ZN(n29803) );
  INHSV1 U29506 ( .I(n29801), .ZN(n26357) );
  CLKNAND2HSV4 U29507 ( .A1(n31510), .A2(n31472), .ZN(n32697) );
  CLKNAND2HSV4 U29508 ( .A1(n31458), .A2(n31457), .ZN(n31510) );
  CLKNAND2HSV4 U29509 ( .A1(n31507), .A2(n31506), .ZN(n31472) );
  XNOR2HSV4 U29510 ( .A1(n26365), .A2(n26359), .ZN(n31664) );
  XNOR2HSV4 U29511 ( .A1(n26361), .A2(n26360), .ZN(n26359) );
  XOR2HSV2 U29512 ( .A1(n31661), .A2(n31662), .Z(n26360) );
  XNOR2HSV4 U29513 ( .A1(n26363), .A2(n26362), .ZN(n26361) );
  XNOR2HSV4 U29514 ( .A1(n31660), .A2(n31659), .ZN(n26362) );
  NOR2HSV4 U29515 ( .A1(n31434), .A2(n26364), .ZN(n26363) );
  CLKNHSV2 U29516 ( .I(n31710), .ZN(n26364) );
  CLKNAND2HSV2 U29517 ( .A1(n32697), .A2(\pe6/got [27]), .ZN(n26365) );
  CLKNAND2HSV2 U29518 ( .A1(n26367), .A2(n26366), .ZN(n26510) );
  CLKNHSV2 U29519 ( .I(n44966), .ZN(n26366) );
  CLKNHSV2 U29520 ( .I(n44965), .ZN(n26367) );
  CLKBUFHSV2 U29521 ( .I(n59775), .Z(n26368) );
  INAND2HSV4 U29522 ( .A1(n26369), .B1(n26368), .ZN(n52262) );
  CLKNHSV2 U29523 ( .I(n59354), .ZN(n26369) );
  INAND2HSV4 U29524 ( .A1(n26370), .B1(n26368), .ZN(n52143) );
  CLKNHSV2 U29525 ( .I(n52051), .ZN(n26370) );
  INAND2HSV4 U29526 ( .A1(n26371), .B1(n26368), .ZN(n47638) );
  CLKNHSV2 U29527 ( .I(n52172), .ZN(n26371) );
  INAND2HSV4 U29528 ( .A1(n26372), .B1(n26368), .ZN(n49583) );
  CLKNHSV2 U29529 ( .I(n51796), .ZN(n26372) );
  INAND2HSV4 U29530 ( .A1(n26373), .B1(n26368), .ZN(n48145) );
  CLKNHSV2 U29531 ( .I(n49493), .ZN(n26373) );
  INAND2HSV4 U29532 ( .A1(n26374), .B1(n26368), .ZN(n51002) );
  CLKNHSV2 U29533 ( .I(n52418), .ZN(n26374) );
  CLKNHSV2 U29534 ( .I(n26548), .ZN(n26376) );
  CLKNAND2HSV2 U29535 ( .A1(n45400), .A2(n26549), .ZN(n26377) );
  CLKNHSV2 U29536 ( .I(n26550), .ZN(n26378) );
  CLKNAND2HSV2 U29537 ( .A1(n40964), .A2(n26379), .ZN(n26382) );
  CLKNHSV2 U29538 ( .I(n26383), .ZN(n26379) );
  INHSV2 U29539 ( .I(n26380), .ZN(n26381) );
  CLKNHSV2 U29540 ( .I(n52763), .ZN(n26380) );
  XNOR2HSV4 U29541 ( .A1(n40960), .A2(n40945), .ZN(n52763) );
  IOA22HSV4 U29542 ( .B1(n40967), .B2(n26381), .A1(n51114), .A2(n41117), .ZN(
        n52760) );
  NAND3HSV4 U29543 ( .A1(n26385), .A2(n26384), .A3(n26382), .ZN(n41117) );
  CLKNHSV2 U29544 ( .I(n40963), .ZN(n26383) );
  AOI22HSV4 U29545 ( .A1(n40962), .A2(\pe1/ti_7t [14]), .B1(n40961), .B2(
        n40960), .ZN(n26384) );
  CLKNAND2HSV2 U29546 ( .A1(n40956), .A2(n40964), .ZN(n26385) );
  NAND3HSV4 U29547 ( .A1(n26388), .A2(n26387), .A3(n26386), .ZN(n30328) );
  CLKNAND2HSV2 U29548 ( .A1(n30140), .A2(n39222), .ZN(n26386) );
  CLKNAND2HSV0 U29549 ( .A1(n30141), .A2(n39222), .ZN(n26387) );
  CLKNHSV2 U29550 ( .I(n30197), .ZN(n47994) );
  CLKNHSV2 U29551 ( .I(n30198), .ZN(n26389) );
  XNOR2HSV4 U29552 ( .A1(n26392), .A2(n26391), .ZN(n26390) );
  XNOR2HSV4 U29553 ( .A1(n30135), .A2(n30136), .ZN(n26392) );
  NOR2HSV4 U29554 ( .A1(n30252), .A2(n40293), .ZN(n26393) );
  CLKNAND2HSV2 U29555 ( .A1(n45605), .A2(n45606), .ZN(n45603) );
  AOI22HSV4 U29556 ( .A1(n45506), .A2(n26394), .B1(n45508), .B2(n45507), .ZN(
        n45606) );
  NOR2HSV4 U29557 ( .A1(n26396), .A2(n26395), .ZN(n26394) );
  CLKNHSV2 U29558 ( .I(n45505), .ZN(n26395) );
  CLKNHSV2 U29559 ( .I(n46090), .ZN(n26397) );
  CLKNAND2HSV2 U29560 ( .A1(n30138), .A2(n26424), .ZN(n30339) );
  XNOR2HSV4 U29561 ( .A1(n26400), .A2(n26399), .ZN(n30305) );
  XNOR2HSV4 U29562 ( .A1(n26401), .A2(n29662), .ZN(n26400) );
  INHSV4 U29563 ( .I(n42810), .ZN(n42917) );
  NOR2HSV4 U29564 ( .A1(n26402), .A2(n42908), .ZN(n42909) );
  XOR2HSV2 U29565 ( .A1(n26403), .A2(n42906), .Z(n26402) );
  NOR2HSV4 U29566 ( .A1(n43025), .A2(n59998), .ZN(n42906) );
  NOR2HSV4 U29567 ( .A1(n42810), .A2(n26404), .ZN(n26403) );
  CLKNHSV2 U29568 ( .I(n43905), .ZN(n26404) );
  XNOR2HSV4 U29569 ( .A1(n26405), .A2(n31477), .ZN(n31478) );
  XNOR2HSV4 U29570 ( .A1(n31318), .A2(n31317), .ZN(n31477) );
  CLKNAND2HSV2 U29571 ( .A1(n31475), .A2(n31476), .ZN(n26406) );
  INHSV2 U29572 ( .I(n26409), .ZN(n40353) );
  NAND2HSV2 U29573 ( .A1(n40347), .A2(n26411), .ZN(n26409) );
  CLKBUFHSV2 U29574 ( .I(n26412), .Z(n26410) );
  CLKNHSV2 U29575 ( .I(n59999), .ZN(n26411) );
  CLKNAND2HSV3 U29576 ( .A1(n26412), .A2(n40427), .ZN(n40391) );
  CLKNAND2HSV2 U29577 ( .A1(n26410), .A2(n55087), .ZN(n41767) );
  CLKNAND2HSV2 U29578 ( .A1(n26410), .A2(n54970), .ZN(n41883) );
  CLKNAND2HSV2 U29579 ( .A1(n26410), .A2(n53473), .ZN(n41458) );
  CLKNAND2HSV2 U29580 ( .A1(n26410), .A2(n44605), .ZN(n42144) );
  INHSV2 U29581 ( .I(n40347), .ZN(n26412) );
  NAND2HSV2 U29582 ( .A1(n45275), .A2(n26415), .ZN(n26823) );
  NAND3HSV2 U29583 ( .A1(n44707), .A2(n44708), .A3(n44706), .ZN(n26415) );
  CLKNAND2HSV0 U29584 ( .A1(n52918), .A2(n59371), .ZN(n51523) );
  CLKNAND2HSV2 U29585 ( .A1(n26414), .A2(n59354), .ZN(n28535) );
  CLKNAND2HSV4 U29586 ( .A1(n42693), .A2(n42692), .ZN(n26416) );
  NAND2HSV3 U29587 ( .A1(n26416), .A2(n42703), .ZN(n42705) );
  CLKNAND2HSV2 U29588 ( .A1(n26417), .A2(n59629), .ZN(n58106) );
  CLKNAND2HSV2 U29589 ( .A1(n26417), .A2(\pe4/got [27]), .ZN(n57085) );
  CLKNAND2HSV2 U29590 ( .A1(n51961), .A2(n51796), .ZN(n49663) );
  CLKNHSV2 U29591 ( .I(n45399), .ZN(n26419) );
  NOR2HSV4 U29592 ( .A1(n48162), .A2(n48161), .ZN(n47903) );
  CLKNAND2HSV4 U29593 ( .A1(n26420), .A2(n26421), .ZN(n45794) );
  CLKNAND2HSV3 U29594 ( .A1(n43488), .A2(n43487), .ZN(n26421) );
  NAND2HSV3 U29595 ( .A1(n30081), .A2(n30082), .ZN(n30138) );
  CLKNHSV2 U29596 ( .I(n40142), .ZN(n26422) );
  XNOR2HSV4 U29597 ( .A1(n30179), .A2(n30180), .ZN(n26423) );
  CLKNHSV2 U29598 ( .I(n39722), .ZN(n26433) );
  CLKNHSV2 U29599 ( .I(n39700), .ZN(n26434) );
  CLKNAND2HSV2 U29600 ( .A1(n39701), .A2(n26443), .ZN(n26441) );
  XNOR2HSV4 U29601 ( .A1(n26438), .A2(n26437), .ZN(n39701) );
  CLKNHSV2 U29602 ( .I(n26428), .ZN(n26427) );
  INAND2HSV4 U29603 ( .A1(n26443), .B1(n39722), .ZN(n26428) );
  NOR2HSV4 U29604 ( .A1(n26430), .A2(n26429), .ZN(n26435) );
  CLKNHSV2 U29605 ( .I(n26436), .ZN(n26429) );
  CLKNHSV2 U29606 ( .I(n26441), .ZN(n26430) );
  NOR2HSV2 U29607 ( .A1(n26432), .A2(n26431), .ZN(n26437) );
  CLKNAND2HSV2 U29608 ( .A1(n39690), .A2(n39689), .ZN(n26431) );
  CLKNHSV2 U29609 ( .I(n39691), .ZN(n26432) );
  MUX2NHSV2 U29610 ( .I0(n26434), .I1(n26433), .S(n39701), .ZN(n26442) );
  CLKNAND2HSV2 U29611 ( .A1(n26435), .A2(n26442), .ZN(n26440) );
  CLKNHSV2 U29612 ( .I(n52767), .ZN(n26436) );
  CLKNAND2HSV4 U29613 ( .A1(n39722), .A2(n26439), .ZN(n39700) );
  XNOR2HSV4 U29614 ( .A1(n39674), .A2(n39673), .ZN(n26438) );
  INHSV2 U29615 ( .I(n26443), .ZN(n26439) );
  NAND3HSV3 U29616 ( .A1(n60068), .A2(n26440), .A3(n39718), .ZN(n39719) );
  CLKNHSV2 U29617 ( .I(n26444), .ZN(n26443) );
  XNOR2HSV4 U29618 ( .A1(n39726), .A2(n39717), .ZN(n60068) );
  CLKNHSV2 U29619 ( .I(n26506), .ZN(n26444) );
  XNOR2HSV4 U29620 ( .A1(n26450), .A2(n26445), .ZN(n31372) );
  XNOR2HSV4 U29621 ( .A1(n26447), .A2(n26446), .ZN(n26445) );
  XOR2HSV2 U29622 ( .A1(n31370), .A2(\pe6/phq [5]), .Z(n26446) );
  XNOR2HSV4 U29623 ( .A1(n26449), .A2(n26448), .ZN(n26447) );
  CLKNAND2HSV2 U29624 ( .A1(n31491), .A2(\pe6/bq[31] ), .ZN(n26448) );
  CLKNAND2HSV2 U29625 ( .A1(n31593), .A2(\pe6/pvq [5]), .ZN(n26449) );
  XNOR2HSV4 U29626 ( .A1(n26453), .A2(n26451), .ZN(n26450) );
  XNOR2HSV4 U29627 ( .A1(n46179), .A2(n26452), .ZN(n26451) );
  CLKNAND2HSV2 U29628 ( .A1(n31368), .A2(n31367), .ZN(n46179) );
  XOR2HSV2 U29629 ( .A1(n26454), .A2(n32105), .Z(n26453) );
  XNOR2HSV4 U29630 ( .A1(n26456), .A2(n26455), .ZN(n31499) );
  XOR2HSV2 U29631 ( .A1(n31490), .A2(n31496), .Z(n26455) );
  XNOR2HSV4 U29632 ( .A1(n26458), .A2(n26457), .ZN(n26456) );
  XNOR2HSV4 U29633 ( .A1(n31486), .A2(n31485), .ZN(n26457) );
  XNOR2HSV4 U29634 ( .A1(n26459), .A2(n31495), .ZN(n26458) );
  XNOR2HSV4 U29635 ( .A1(n26460), .A2(\pe6/phq [6]), .ZN(n26459) );
  CLKNAND2HSV3 U29636 ( .A1(n44389), .A2(n44346), .ZN(n26465) );
  CLKNAND2HSV2 U29637 ( .A1(n26461), .A2(n46575), .ZN(n44346) );
  XNOR2HSV4 U29638 ( .A1(n36028), .A2(n36027), .ZN(n46575) );
  NOR2HSV4 U29639 ( .A1(n44342), .A2(n36066), .ZN(n26461) );
  XOR2HSV4 U29640 ( .A1(n35918), .A2(n36035), .Z(n44342) );
  CLKBUFHSV2 U29641 ( .I(n46575), .Z(n26462) );
  NOR2HSV4 U29642 ( .A1(n44342), .A2(n46159), .ZN(n26464) );
  CLKBUFHSV2 U29643 ( .I(n59732), .Z(n26467) );
  CLKNAND2HSV3 U29644 ( .A1(n42487), .A2(n44527), .ZN(n59732) );
  CLKNAND2HSV2 U29645 ( .A1(n32459), .A2(n26470), .ZN(n26469) );
  CLKNHSV2 U29646 ( .I(n32457), .ZN(n26470) );
  NOR2HSV4 U29647 ( .A1(n26472), .A2(n26471), .ZN(n32832) );
  CLKNHSV2 U29648 ( .I(n33061), .ZN(n26471) );
  CLKNHSV2 U29649 ( .I(n41240), .ZN(n41241) );
  CLKNAND2HSV4 U29650 ( .A1(n60026), .A2(n42488), .ZN(n41506) );
  CLKXOR2HSV4 U29651 ( .A1(n26473), .A2(n41240), .Z(n60026) );
  CLKNAND2HSV1 U29652 ( .A1(n41239), .A2(n41328), .ZN(n26473) );
  AOI21HSV4 U29653 ( .A1(n26474), .A2(n60030), .B(n59950), .ZN(n35454) );
  NOR2HSV4 U29654 ( .A1(n35014), .A2(n47777), .ZN(n26474) );
  CLKNHSV2 U29655 ( .I(n59883), .ZN(n52567) );
  XNOR2HSV4 U29656 ( .A1(n39214), .A2(n26475), .ZN(n39238) );
  XNOR2HSV4 U29657 ( .A1(n26479), .A2(n26476), .ZN(n26475) );
  XOR2HSV2 U29658 ( .A1(n39212), .A2(n26477), .Z(n26476) );
  XNOR2HSV4 U29659 ( .A1(n39213), .A2(n26478), .ZN(n26477) );
  XNOR2HSV4 U29660 ( .A1(n39210), .A2(n39211), .ZN(n26478) );
  INAND2HSV4 U29661 ( .A1(n37635), .B1(n59883), .ZN(n26479) );
  INAND2HSV4 U29662 ( .A1(n26482), .B1(n26480), .ZN(n42606) );
  CLKNHSV2 U29663 ( .I(n26481), .ZN(n26480) );
  XNOR2HSV4 U29664 ( .A1(n26481), .A2(n26482), .ZN(n42797) );
  XNOR2HSV4 U29665 ( .A1(n42588), .A2(n42587), .ZN(n26481) );
  CLKNHSV4 U29666 ( .I(n31256), .ZN(n26489) );
  NAND2HSV3 U29667 ( .A1(n26484), .A2(n26483), .ZN(n31283) );
  CLKNAND2HSV2 U29668 ( .A1(n31369), .A2(n31418), .ZN(n26483) );
  CLKNAND2HSV2 U29669 ( .A1(n32881), .A2(\pe6/pvq [1]), .ZN(n26484) );
  BUFHSV8 U29670 ( .I(n31257), .Z(n26485) );
  CLKNAND2HSV3 U29671 ( .A1(n26488), .A2(n26486), .ZN(n31260) );
  OAI21HSV4 U29672 ( .A1(n31256), .A2(n31424), .B(n26487), .ZN(n26486) );
  CLKNHSV2 U29673 ( .I(\pe6/phq [1]), .ZN(n26487) );
  NAND3HSV4 U29674 ( .A1(n31339), .A2(n26489), .A3(\pe6/phq [1]), .ZN(n26488)
         );
  CLKNHSV2 U29675 ( .I(n31260), .ZN(n31257) );
  NAND3HSV4 U29676 ( .A1(n26490), .A2(n31257), .A3(n31261), .ZN(n31259) );
  CLKNAND2HSV2 U29677 ( .A1(n31284), .A2(n31283), .ZN(n26490) );
  NAND3HSV4 U29678 ( .A1(n26515), .A2(n26513), .A3(n26491), .ZN(n31284) );
  NOR2HSV4 U29679 ( .A1(n26514), .A2(n31253), .ZN(n26491) );
  XNOR2HSV4 U29680 ( .A1(n26494), .A2(n26492), .ZN(n37637) );
  NOR2HSV4 U29681 ( .A1(n39664), .A2(n37635), .ZN(n26492) );
  AOI21HSV4 U29682 ( .A1(n31144), .A2(n31145), .B(n26493), .ZN(n39664) );
  XNOR2HSV4 U29683 ( .A1(n37634), .A2(n26495), .ZN(n26494) );
  XOR3HSV2 U29684 ( .A1(n37633), .A2(n26496), .A3(n37632), .Z(n26495) );
  CLKNHSV2 U29685 ( .I(n26497), .ZN(n39666) );
  CLKNAND2HSV2 U29686 ( .A1(n59883), .A2(n26498), .ZN(n26497) );
  CLKNHSV2 U29687 ( .I(n31081), .ZN(n26498) );
  NOR2HSV4 U29688 ( .A1(n39731), .A2(n26499), .ZN(n26505) );
  XNOR2HSV4 U29689 ( .A1(n39715), .A2(n39714), .ZN(n39731) );
  CLKNHSV2 U29690 ( .I(n40309), .ZN(n26500) );
  CLKNHSV2 U29691 ( .I(n26503), .ZN(n26502) );
  CLKNHSV2 U29692 ( .I(n26506), .ZN(n26503) );
  CLKNHSV2 U29693 ( .I(n39722), .ZN(n26504) );
  NOR2HSV4 U29694 ( .A1(n40285), .A2(n26505), .ZN(n39737) );
  INHSV2 U29695 ( .I(n39692), .ZN(n26506) );
  CLKNHSV3 U29696 ( .I(n35305), .ZN(n35307) );
  CLKNHSV4 U29697 ( .I(n60030), .ZN(n35004) );
  XNOR2HSV4 U29698 ( .A1(n35006), .A2(n35005), .ZN(n35008) );
  OAI21HSV4 U29699 ( .A1(n26509), .A2(n26508), .B(n26507), .ZN(n45143) );
  CLKNAND2HSV2 U29700 ( .A1(n26512), .A2(n26546), .ZN(n26508) );
  CLKNHSV2 U29701 ( .I(n26510), .ZN(n26509) );
  CLKNHSV2 U29702 ( .I(n31255), .ZN(n26513) );
  CLKNHSV2 U29703 ( .I(\pe6/bq[32] ), .ZN(n26514) );
  CLKNHSV2 U29704 ( .I(n31254), .ZN(n26515) );
  CLKBUFHSV4 U29705 ( .I(n26596), .Z(n26516) );
  CLKNAND2HSV2 U29706 ( .A1(n26516), .A2(n57574), .ZN(n50414) );
  CLKNAND2HSV2 U29707 ( .A1(n26516), .A2(n35318), .ZN(n57577) );
  CLKNAND2HSV2 U29708 ( .A1(n26516), .A2(n58137), .ZN(n58249) );
  CLKNAND2HSV2 U29709 ( .A1(n26516), .A2(n57672), .ZN(n50310) );
  CLKNAND2HSV2 U29710 ( .A1(n26516), .A2(n59350), .ZN(n57449) );
  CLKNAND2HSV2 U29711 ( .A1(n32421), .A2(n26517), .ZN(n32233) );
  CLKAND2HSV4 U29712 ( .A1(n32314), .A2(n32315), .Z(n32421) );
  CLKNHSV2 U29713 ( .I(n32044), .ZN(n26518) );
  OAI21HSV2 U29714 ( .A1(n26538), .A2(n26537), .B(n26536), .ZN(n26534) );
  CLKNAND2HSV2 U29715 ( .A1(n44527), .A2(n44525), .ZN(n26537) );
  CLKNHSV2 U29716 ( .I(n44526), .ZN(n26538) );
  CLKNHSV2 U29717 ( .I(n26531), .ZN(n26519) );
  NOR2HSV4 U29718 ( .A1(n26531), .A2(n26533), .ZN(n26521) );
  CLKNHSV2 U29719 ( .I(n26532), .ZN(n26522) );
  AOI21HSV4 U29720 ( .A1(n26529), .A2(n26528), .B(n26526), .ZN(n26525) );
  CLKNHSV2 U29721 ( .I(n26533), .ZN(n26527) );
  CLKNHSV2 U29722 ( .I(n26538), .ZN(n26528) );
  CLKNHSV2 U29723 ( .I(n26537), .ZN(n26529) );
  CLKNHSV2 U29724 ( .I(n41727), .ZN(n26533) );
  NOR2HSV8 U29725 ( .A1(n25838), .A2(n39738), .ZN(n39739) );
  CLKNAND2HSV3 U29726 ( .A1(n39739), .A2(n40017), .ZN(n40290) );
  CLKNAND2HSV4 U29727 ( .A1(n39711), .A2(n39712), .ZN(n40017) );
  OAI22HSV4 U29728 ( .A1(n26541), .A2(n26540), .B1(n26545), .B2(n26539), .ZN(
        n26544) );
  CLKNHSV2 U29729 ( .I(n40289), .ZN(n26540) );
  CLKNHSV2 U29730 ( .I(n26542), .ZN(n26541) );
  CLKNAND2HSV2 U29731 ( .A1(n45499), .A2(n26543), .ZN(n26542) );
  CLKNHSV2 U29732 ( .I(n40288), .ZN(n26543) );
  OAI21HSV1 U29733 ( .A1(n40318), .A2(n29914), .B(n40317), .ZN(n40304) );
  CLKNAND2HSV2 U29734 ( .A1(n40287), .A2(n30142), .ZN(n26545) );
  CLKNAND2HSV2 U29735 ( .A1(n26417), .A2(n57753), .ZN(n57978) );
  CLKNAND2HSV2 U29736 ( .A1(n26417), .A2(n58153), .ZN(n58188) );
  CLKNAND2HSV2 U29737 ( .A1(n26417), .A2(n58137), .ZN(n50123) );
  CLKNAND2HSV2 U29738 ( .A1(n26417), .A2(n58246), .ZN(n58211) );
  CLKNAND2HSV2 U29739 ( .A1(n26417), .A2(n58216), .ZN(n58252) );
  CLKNAND2HSV2 U29740 ( .A1(n26417), .A2(n58258), .ZN(n58278) );
  CLKNAND2HSV2 U29741 ( .A1(n26417), .A2(n58314), .ZN(n58293) );
  CLKNHSV2 U29742 ( .I(n45405), .ZN(n26548) );
  AND3HSV8 U29743 ( .A1(n44707), .A2(n44708), .A3(n44706), .Z(n26547) );
  CLKNHSV2 U29744 ( .I(n27236), .ZN(n26549) );
  CLKNAND2HSV0 U29745 ( .A1(n26552), .A2(n36671), .ZN(n26550) );
  CLKNHSV2 U29746 ( .I(n43488), .ZN(n47949) );
  CLKNAND2HSV2 U29747 ( .A1(n25891), .A2(n43140), .ZN(n45516) );
  NOR2HSV4 U29748 ( .A1(n43470), .A2(n43130), .ZN(n43487) );
  CLKNHSV2 U29749 ( .I(n43466), .ZN(n26552) );
  MUX2NHSV2 U29750 ( .I0(n26553), .I1(n26554), .S(n40398), .ZN(n40404) );
  XNOR2HSV4 U29751 ( .A1(n40392), .A2(n40391), .ZN(n40398) );
  CLKNHSV2 U29752 ( .I(n40394), .ZN(n26554) );
  CLKNAND2HSV3 U29753 ( .A1(n39424), .A2(n39425), .ZN(n26556) );
  CLKNAND2HSV4 U29754 ( .A1(n26556), .A2(n26555), .ZN(n39557) );
  XNOR2HSV4 U29755 ( .A1(n39557), .A2(n39556), .ZN(n39717) );
  AOI31HSV2 U29756 ( .A1(n36630), .A2(n44780), .A3(n36521), .B(n36520), .ZN(
        n26557) );
  CLKNHSV8 U29757 ( .I(n48896), .ZN(n37791) );
  CLKNAND2HSV3 U29758 ( .A1(n26558), .A2(n26557), .ZN(n48896) );
  CLKNAND2HSV1 U29759 ( .A1(n36518), .A2(n36629), .ZN(n26558) );
  CLKNHSV2 U29760 ( .I(n38455), .ZN(n26559) );
  CLKNAND2HSV2 U29761 ( .A1(n52286), .A2(n38723), .ZN(n38724) );
  CLKNAND2HSV2 U29762 ( .A1(n52286), .A2(n44711), .ZN(n26819) );
  CLKNAND2HSV2 U29763 ( .A1(n52286), .A2(n38778), .ZN(n38864) );
  CLKNAND2HSV2 U29764 ( .A1(n52286), .A2(n52922), .ZN(n44278) );
  CLKNAND2HSV0 U29765 ( .A1(n52286), .A2(n38390), .ZN(n44802) );
  NOR2HSV4 U29766 ( .A1(n26563), .A2(n26561), .ZN(n26566) );
  CLKNHSV2 U29767 ( .I(n26567), .ZN(n26562) );
  CLKNHSV2 U29768 ( .I(n42607), .ZN(n52791) );
  AOI21HSV4 U29769 ( .A1(n26566), .A2(n42606), .B(n42799), .ZN(n42608) );
  CLKNHSV2 U29770 ( .I(n42590), .ZN(n26567) );
  XNOR2HSV4 U29771 ( .A1(n38464), .A2(n26569), .ZN(n38519) );
  CLKNAND2HSV2 U29772 ( .A1(n38462), .A2(n38463), .ZN(n26569) );
  CLKNAND2HSV3 U29773 ( .A1(n38458), .A2(n38604), .ZN(n38518) );
  CLKNHSV4 U29774 ( .I(n38606), .ZN(n26571) );
  INHSV2 U29775 ( .I(n26579), .ZN(n26572) );
  NAND3HSV4 U29776 ( .A1(n31085), .A2(n31087), .A3(n30681), .ZN(n26578) );
  CLKNHSV2 U29777 ( .I(n26574), .ZN(n26573) );
  INAND2HSV4 U29778 ( .A1(n40169), .B1(n30757), .ZN(n26574) );
  IOA21HSV4 U29779 ( .A1(n31140), .A2(n26572), .B(n26575), .ZN(n30997) );
  NOR2HSV4 U29780 ( .A1(n26577), .A2(n26576), .ZN(n26575) );
  CLKNHSV2 U29781 ( .I(n30759), .ZN(n26576) );
  NOR2HSV4 U29782 ( .A1(n26578), .A2(n31140), .ZN(n26577) );
  XNOR2HSV4 U29783 ( .A1(n30750), .A2(n30749), .ZN(n31140) );
  CLKNAND2HSV2 U29784 ( .A1(n43226), .A2(n42697), .ZN(n26580) );
  XNOR2HSV4 U29785 ( .A1(n26686), .A2(n26687), .ZN(n26581) );
  AOI31HSV2 U29786 ( .A1(n42925), .A2(n42926), .A3(n42924), .B(n42923), .ZN(
        n42927) );
  CLKNAND2HSV2 U29787 ( .A1(n26582), .A2(n32675), .ZN(n32676) );
  OAI21HSV4 U29788 ( .A1(n32686), .A2(n32674), .B(n32673), .ZN(n26582) );
  CLKNHSV2 U29789 ( .I(n39733), .ZN(n26583) );
  CLKXOR2HSV4 U29790 ( .A1(n52800), .A2(n30862), .Z(n30870) );
  NOR2HSV4 U29791 ( .A1(n31121), .A2(n31123), .ZN(n30994) );
  OAI21HSV4 U29792 ( .A1(n30859), .A2(n30860), .B(n31102), .ZN(n31123) );
  NOR2HSV4 U29793 ( .A1(n30861), .A2(n31091), .ZN(n31121) );
  OAI21HSV4 U29794 ( .A1(pov4[29]), .A2(n28669), .B(n47779), .ZN(n52848) );
  CLKNAND2HSV2 U29795 ( .A1(n31897), .A2(n31896), .ZN(n26587) );
  XOR4HSV2 U29796 ( .A1(n42651), .A2(n26593), .A3(n26591), .A4(n26588), .Z(
        n36700) );
  XNOR2HSV4 U29797 ( .A1(n26590), .A2(n26589), .ZN(n26588) );
  CLKNAND2HSV2 U29798 ( .A1(n36795), .A2(n36710), .ZN(n26590) );
  XOR2HSV2 U29799 ( .A1(n26595), .A2(n26594), .Z(n26593) );
  CLKNAND2HSV2 U29800 ( .A1(n59609), .A2(\pe3/bq[31] ), .ZN(n26594) );
  CLKNAND2HSV2 U29801 ( .A1(n37298), .A2(n59614), .ZN(n26595) );
  AOI21HSV4 U29802 ( .A1(n36861), .A2(n36901), .B(n36839), .ZN(n36964) );
  BUFHSV8 U29803 ( .I(n58145), .Z(n26596) );
  CLKNHSV2 U29804 ( .I(n26739), .ZN(n26597) );
  XNOR2HSV4 U29805 ( .A1(n26599), .A2(n27149), .ZN(n27150) );
  CLKNAND2HSV2 U29806 ( .A1(n59021), .A2(n49665), .ZN(n26599) );
  CLKNHSV2 U29807 ( .I(n26601), .ZN(n26600) );
  CLKNAND2HSV2 U29808 ( .A1(n26602), .A2(n46587), .ZN(n26601) );
  CLKNHSV2 U29809 ( .I(n46158), .ZN(n26603) );
  INHSV24 U29810 ( .I(n47935), .ZN(n26604) );
  CLKNHSV2 U29811 ( .I(n40493), .ZN(n53530) );
  CLKNHSV2 U29812 ( .I(n47935), .ZN(n40331) );
  NOR2HSV4 U29813 ( .A1(n26604), .A2(n59376), .ZN(n26605) );
  INOR2HSV2 U29814 ( .A1(n40443), .B1(n40568), .ZN(n40363) );
  INHSV2 U29815 ( .I(n51112), .ZN(n26606) );
  CLKNHSV4 U29816 ( .I(n40520), .ZN(n40365) );
  CLKNHSV8 U29817 ( .I(n40371), .ZN(n26607) );
  NOR2HSV8 U29818 ( .A1(n40598), .A2(n40327), .ZN(n40371) );
  CLKNHSV2 U29819 ( .I(n44321), .ZN(n44326) );
  CLKNAND2HSV2 U29820 ( .A1(n26610), .A2(n46082), .ZN(n36752) );
  CLKNHSV2 U29821 ( .I(n36729), .ZN(n26609) );
  XNOR2HSV4 U29822 ( .A1(n26615), .A2(n26611), .ZN(n41843) );
  CLKNAND2HSV2 U29823 ( .A1(n42355), .A2(n42200), .ZN(n26611) );
  OAI21HSV4 U29824 ( .A1(n26614), .A2(n26613), .B(n26612), .ZN(n42355) );
  AOI22HSV4 U29825 ( .A1(n41720), .A2(\pe1/ti_7t [22]), .B1(n26613), .B2(
        n41711), .ZN(n26612) );
  CLKNHSV2 U29826 ( .I(n41703), .ZN(n26614) );
  CLKNHSV2 U29827 ( .I(n42084), .ZN(n26617) );
  CLKNAND2HSV2 U29828 ( .A1(n59391), .A2(\pe1/got [28]), .ZN(n26618) );
  CLKNAND2HSV0 U29829 ( .A1(n52924), .A2(n38026), .ZN(n38534) );
  CLKNAND2HSV2 U29830 ( .A1(n52924), .A2(n38327), .ZN(n39099) );
  CLKNAND2HSV2 U29831 ( .A1(n44970), .A2(n53086), .ZN(n44020) );
  CLKNAND2HSV2 U29832 ( .A1(n44970), .A2(n59584), .ZN(n44282) );
  AOI21HSV4 U29833 ( .A1(n38890), .A2(n52924), .B(n38889), .ZN(n38895) );
  CLKNAND2HSV4 U29834 ( .A1(n38531), .A2(n38530), .ZN(n52924) );
  CLKNAND2HSV2 U29835 ( .A1(n26622), .A2(n26624), .ZN(n26619) );
  CLKNHSV2 U29836 ( .I(n26624), .ZN(n26623) );
  CLKNHSV2 U29837 ( .I(n42471), .ZN(n26625) );
  CLKNAND2HSV2 U29838 ( .A1(n33096), .A2(\pe4/pvq [2]), .ZN(n26627) );
  NOR2HSV4 U29839 ( .A1(n36692), .A2(n36670), .ZN(n36696) );
  NOR2HSV4 U29840 ( .A1(n36692), .A2(n26631), .ZN(n26630) );
  INAND2HSV4 U29841 ( .A1(n36670), .B1(n59962), .ZN(n26631) );
  CLKNAND2HSV3 U29842 ( .A1(n26633), .A2(n47775), .ZN(n26632) );
  NAND3HSV4 U29843 ( .A1(n26635), .A2(n26634), .A3(n60077), .ZN(n26637) );
  CLKNHSV2 U29844 ( .I(n47789), .ZN(n26636) );
  XNOR2HSV1 U29845 ( .A1(n26638), .A2(n27575), .ZN(n27576) );
  NAND2HSV3 U29846 ( .A1(n27574), .A2(n26639), .ZN(n26638) );
  INHSV2 U29847 ( .I(n26640), .ZN(n26639) );
  NOR2HSV2 U29848 ( .A1(n27572), .A2(n27573), .ZN(n26640) );
  XNOR2HSV4 U29849 ( .A1(n26641), .A2(n49662), .ZN(n49664) );
  XNOR2HSV4 U29850 ( .A1(n49660), .A2(n26642), .ZN(n26641) );
  XOR3HSV2 U29851 ( .A1(n49659), .A2(n26700), .A3(n26701), .Z(n26642) );
  CLKNAND2HSV4 U29852 ( .A1(n26643), .A2(n33801), .ZN(n33179) );
  CLKNHSV4 U29853 ( .I(n33172), .ZN(n26643) );
  CLKNHSV2 U29854 ( .I(n33172), .ZN(n33173) );
  XNOR2HSV4 U29855 ( .A1(n26646), .A2(n26645), .ZN(n33178) );
  NOR2HSV4 U29856 ( .A1(n33177), .A2(n33176), .ZN(n26646) );
  CLKNAND2HSV4 U29857 ( .A1(n26647), .A2(n33169), .ZN(n33292) );
  CLKNAND2HSV3 U29858 ( .A1(n33168), .A2(n26666), .ZN(n26647) );
  INHSV2 U29859 ( .I(n26649), .ZN(n26648) );
  CLKNAND2HSV4 U29860 ( .A1(n39553), .A2(n39554), .ZN(n39872) );
  CLKNHSV2 U29861 ( .I(n39567), .ZN(n26649) );
  AOI21HSV4 U29862 ( .A1(n39570), .A2(n39246), .B(n39245), .ZN(n26650) );
  CLKNAND2HSV4 U29863 ( .A1(n26685), .A2(n26684), .ZN(n39570) );
  CLKNHSV2 U29864 ( .I(n49000), .ZN(n26651) );
  XNOR2HSV4 U29865 ( .A1(n26653), .A2(n48999), .ZN(n26652) );
  XOR2HSV2 U29866 ( .A1(n26654), .A2(n48998), .Z(n26653) );
  NAND2HSV2 U29867 ( .A1(n31752), .A2(n31751), .ZN(n26658) );
  XNOR2HSV4 U29868 ( .A1(n31744), .A2(n26655), .ZN(n26660) );
  NAND3HSV4 U29869 ( .A1(n26657), .A2(n31757), .A3(n31756), .ZN(n26656) );
  CLKNHSV2 U29870 ( .I(n26659), .ZN(n26657) );
  XNOR2HSV4 U29871 ( .A1(n26661), .A2(n26660), .ZN(n31815) );
  NOR2HSV4 U29872 ( .A1(n31705), .A2(n52705), .ZN(n26661) );
  CLKNHSV2 U29873 ( .I(n34043), .ZN(n35501) );
  XNOR2HSV1 U29874 ( .A1(n26664), .A2(n26662), .ZN(n33165) );
  XNOR2HSV1 U29875 ( .A1(n26663), .A2(n33131), .ZN(n26662) );
  NAND2HSV2 U29876 ( .A1(n33173), .A2(n59350), .ZN(n26663) );
  XNOR2HSV2 U29877 ( .A1(n26665), .A2(n33150), .ZN(n26664) );
  CLKNAND2HSV3 U29878 ( .A1(n34043), .A2(n33263), .ZN(n26665) );
  CLKNAND2HSV4 U29879 ( .A1(n26667), .A2(n26666), .ZN(n34043) );
  CLKNHSV4 U29880 ( .I(n33180), .ZN(n26666) );
  CLKNAND2HSV3 U29881 ( .A1(n33181), .A2(n29650), .ZN(n26667) );
  BUFHSV8 U29882 ( .I(n43614), .Z(n26668) );
  OAI21HSV4 U29883 ( .A1(n26668), .A2(n26670), .B(n26669), .ZN(n43729) );
  AOI21HSV4 U29884 ( .A1(n26668), .A2(n43620), .B(n43619), .ZN(n26669) );
  CLKNHSV2 U29885 ( .I(n43615), .ZN(n26670) );
  AOI21HSV4 U29886 ( .A1(n26668), .A2(n26673), .B(n26672), .ZN(n26671) );
  CLKNHSV2 U29887 ( .I(n43616), .ZN(n26672) );
  CLKNHSV2 U29888 ( .I(n43867), .ZN(n26673) );
  XNOR2HSV4 U29889 ( .A1(n52041), .A2(n26674), .ZN(n52044) );
  XNOR2HSV4 U29890 ( .A1(n26677), .A2(n26675), .ZN(n26674) );
  CLKNHSV2 U29891 ( .I(n52050), .ZN(n26676) );
  XNOR2HSV4 U29892 ( .A1(n26678), .A2(n52040), .ZN(n26677) );
  CLKNAND2HSV3 U29893 ( .A1(n37533), .A2(n39693), .ZN(n26679) );
  XNOR2HSV4 U29894 ( .A1(n30998), .A2(n30997), .ZN(n37533) );
  CLKNAND2HSV3 U29895 ( .A1(n26679), .A2(n31001), .ZN(n26681) );
  CLKNHSV2 U29896 ( .I(n31000), .ZN(n37532) );
  CLKNAND2HSV4 U29897 ( .A1(n26682), .A2(n26680), .ZN(n39542) );
  CLKNAND2HSV2 U29898 ( .A1(n37536), .A2(n30999), .ZN(n26682) );
  BUFHSV8 U29899 ( .I(n39570), .Z(n26683) );
  CLKNAND2HSV1 U29900 ( .A1(n39575), .A2(n39574), .ZN(n26684) );
  NAND2HSV2 U29901 ( .A1(n39243), .A2(n39244), .ZN(n26685) );
  CLKNHSV2 U29902 ( .I(n39570), .ZN(n39866) );
  XNOR2HSV4 U29903 ( .A1(n37526), .A2(n37525), .ZN(n42612) );
  NAND3HSV4 U29904 ( .A1(n37450), .A2(n37448), .A3(n37449), .ZN(n42610) );
  XNOR2HSV4 U29905 ( .A1(n42688), .A2(n42687), .ZN(n26686) );
  NOR2HSV4 U29906 ( .A1(n26690), .A2(n26689), .ZN(n26688) );
  CLKNHSV2 U29907 ( .I(n42695), .ZN(n26689) );
  CLKNHSV2 U29908 ( .I(n42689), .ZN(n26691) );
  OAI21HSV4 U29909 ( .A1(n35486), .A2(n47930), .B(n35485), .ZN(n58145) );
  OAI21HSV4 U29910 ( .A1(n35477), .A2(n35478), .B(n35476), .ZN(n35485) );
  NAND3HSV4 U29911 ( .A1(n35458), .A2(n35461), .A3(n35459), .ZN(n47930) );
  CLKNHSV2 U29912 ( .I(n35455), .ZN(n26693) );
  CLKNHSV2 U29913 ( .I(n35462), .ZN(n26694) );
  CLKNHSV2 U29914 ( .I(n35457), .ZN(n26695) );
  CLKNHSV2 U29915 ( .I(n54729), .ZN(n53389) );
  XNOR2HSV4 U29916 ( .A1(n26699), .A2(n26696), .ZN(n42197) );
  XNOR2HSV4 U29917 ( .A1(n42058), .A2(n26697), .ZN(n26696) );
  NOR2HSV4 U29918 ( .A1(n55144), .A2(n26698), .ZN(n26697) );
  CLKNHSV2 U29919 ( .I(n41731), .ZN(n26698) );
  CLKNHSV2 U29920 ( .I(n45147), .ZN(n52048) );
  CLKNAND2HSV1 U29921 ( .A1(n51797), .A2(n52172), .ZN(n26700) );
  NOR2HSV2 U29922 ( .A1(n25833), .A2(n26702), .ZN(n26701) );
  INHSV2 U29923 ( .I(n59375), .ZN(n26702) );
  NAND3HSV4 U29924 ( .A1(n26704), .A2(n29642), .A3(n29846), .ZN(n26703) );
  CLKNHSV2 U29925 ( .I(n29666), .ZN(n26704) );
  CLKNAND2HSV2 U29926 ( .A1(n29864), .A2(n29863), .ZN(n26705) );
  CLKNAND2HSV3 U29927 ( .A1(n45477), .A2(n30028), .ZN(n26711) );
  XNOR2HSV4 U29928 ( .A1(n26711), .A2(n26706), .ZN(n30050) );
  XNOR3HSV2 U29929 ( .A1(n26710), .A2(n26707), .A3(n30047), .ZN(n26706) );
  XNOR2HSV4 U29930 ( .A1(n26709), .A2(n26708), .ZN(n26707) );
  XNOR2HSV4 U29931 ( .A1(n30042), .A2(n30045), .ZN(n26708) );
  XNOR2HSV4 U29932 ( .A1(n30044), .A2(n30043), .ZN(n26709) );
  NOR2HSV4 U29933 ( .A1(n30106), .A2(n30595), .ZN(n26710) );
  XNOR2HSV4 U29934 ( .A1(n26715), .A2(n26714), .ZN(n26713) );
  XNOR2HSV4 U29935 ( .A1(n26716), .A2(n51606), .ZN(n26715) );
  XNOR2HSV4 U29936 ( .A1(n51604), .A2(n51605), .ZN(n26716) );
  CLKNAND2HSV2 U29937 ( .A1(n26719), .A2(n26717), .ZN(n38181) );
  CLKNAND2HSV2 U29938 ( .A1(n38167), .A2(n38108), .ZN(n26718) );
  AOI31HSV2 U29939 ( .A1(n47981), .A2(n26720), .A3(n25851), .B(n44156), .ZN(
        n26719) );
  CLKNAND2HSV2 U29940 ( .A1(n38000), .A2(n37999), .ZN(n26722) );
  CLKNAND2HSV3 U29941 ( .A1(n37997), .A2(n37998), .ZN(n26723) );
  XNOR2HSV4 U29942 ( .A1(n26724), .A2(n27089), .ZN(n27090) );
  CLKNAND2HSV2 U29943 ( .A1(n26725), .A2(n27088), .ZN(n26724) );
  CLKNHSV2 U29944 ( .I(n27086), .ZN(n26726) );
  XNOR2HSV4 U29945 ( .A1(n36300), .A2(n36301), .ZN(n36315) );
  XNOR2HSV4 U29946 ( .A1(n26727), .A2(n36292), .ZN(n36301) );
  XNOR2HSV4 U29947 ( .A1(n36290), .A2(n36291), .ZN(n26727) );
  XNOR2HSV4 U29948 ( .A1(n26731), .A2(n26728), .ZN(n36300) );
  NOR2HSV4 U29949 ( .A1(n26730), .A2(n26729), .ZN(n26728) );
  CLKNHSV2 U29950 ( .I(n45008), .ZN(n26729) );
  CLKNHSV2 U29951 ( .I(n38742), .ZN(n26730) );
  OAI21HSV4 U29952 ( .A1(n36297), .A2(n36296), .B(n36295), .ZN(n26731) );
  BUFHSV8 U29953 ( .I(\pe5/ctrq ), .Z(n26734) );
  NAND3HSV4 U29954 ( .A1(n26734), .A2(n26733), .A3(\pe5/pvq [2]), .ZN(n26736)
         );
  CLKNAND2HSV2 U29955 ( .A1(n41921), .A2(n41922), .ZN(n26737) );
  CLKNHSV2 U29956 ( .I(n26741), .ZN(n26739) );
  CLKNHSV2 U29957 ( .I(n34221), .ZN(n26740) );
  CLKNHSV2 U29958 ( .I(n46566), .ZN(n26741) );
  OAI21HSV4 U29959 ( .A1(n37539), .A2(n37538), .B(n37537), .ZN(n60054) );
  CLKNAND2HSV3 U29960 ( .A1(n60054), .A2(n40008), .ZN(n26744) );
  XNOR2HSV4 U29961 ( .A1(n37759), .A2(n26743), .ZN(n37545) );
  XNOR2HSV4 U29962 ( .A1(n37531), .A2(n26744), .ZN(n26743) );
  XNOR2HSV4 U29963 ( .A1(n31095), .A2(n31096), .ZN(n37531) );
  NAND3HSV4 U29964 ( .A1(n37541), .A2(n37550), .A3(n37540), .ZN(n39116) );
  CLKNAND2HSV3 U29965 ( .A1(n52816), .A2(n31242), .ZN(n37541) );
  CLKNAND2HSV4 U29966 ( .A1(n31099), .A2(n31100), .ZN(n37550) );
  CLKNHSV2 U29967 ( .I(n45259), .ZN(n45258) );
  XNOR2HSV4 U29968 ( .A1(n26745), .A2(n45256), .ZN(n45259) );
  XOR2HSV2 U29969 ( .A1(n26746), .A2(n45255), .Z(n26745) );
  XOR2HSV2 U29970 ( .A1(n45254), .A2(n45253), .Z(n26746) );
  INOR2HSV4 U29971 ( .A1(n26779), .B1(n26747), .ZN(n26750) );
  CLKNAND2HSV2 U29972 ( .A1(n26777), .A2(n26748), .ZN(n26747) );
  CLKNHSV2 U29973 ( .I(n26752), .ZN(n26748) );
  OAI21HSV4 U29974 ( .A1(n26753), .A2(n26752), .B(n26749), .ZN(n59579) );
  AOI21HSV4 U29975 ( .A1(n26751), .A2(n26750), .B(n29728), .ZN(n26749) );
  CLKNHSV2 U29976 ( .I(n26754), .ZN(n26751) );
  CLKNHSV2 U29977 ( .I(n35604), .ZN(n26752) );
  CLKNAND2HSV2 U29978 ( .A1(n26782), .A2(n26755), .ZN(n26754) );
  INHSV2 U29979 ( .I(n26785), .ZN(n26756) );
  CLKNHSV2 U29980 ( .I(n26757), .ZN(n39672) );
  CLKNHSV2 U29981 ( .I(n39693), .ZN(n26758) );
  OAI21HSV4 U29982 ( .A1(n39415), .A2(n39669), .B(n39416), .ZN(n47947) );
  CLKNAND2HSV2 U29983 ( .A1(n39413), .A2(n39414), .ZN(n39669) );
  CLKNHSV2 U29984 ( .I(n26759), .ZN(n47565) );
  NOR2HSV4 U29985 ( .A1(n47564), .A2(n47563), .ZN(n26759) );
  CLKNAND2HSV2 U29986 ( .A1(n25709), .A2(n51796), .ZN(n47563) );
  XNOR2HSV4 U29987 ( .A1(n26760), .A2(n47562), .ZN(n47564) );
  XNOR2HSV4 U29988 ( .A1(n47560), .A2(n47561), .ZN(n26760) );
  NOR2HSV4 U29989 ( .A1(n36331), .A2(n26762), .ZN(n36333) );
  CLKNHSV2 U29990 ( .I(n38108), .ZN(n26762) );
  NOR2HSV4 U29991 ( .A1(n36315), .A2(n38603), .ZN(n36331) );
  CLKNHSV2 U29992 ( .I(n36665), .ZN(n36250) );
  CLKNHSV2 U29993 ( .I(n36443), .ZN(n45303) );
  OAI21HSV4 U29994 ( .A1(n26766), .A2(n26765), .B(n26763), .ZN(n36260) );
  OAI21HSV4 U29995 ( .A1(n36443), .A2(n26764), .B(n36249), .ZN(n26763) );
  CLKNHSV2 U29996 ( .I(\pe2/got [32]), .ZN(n26764) );
  CLKNHSV2 U29997 ( .I(n45008), .ZN(n26765) );
  INAND2HSV4 U29998 ( .A1(n36665), .B1(\pe2/phq [1]), .ZN(n26766) );
  NAND3HSV4 U29999 ( .A1(n40003), .A2(n40002), .A3(n39878), .ZN(n26768) );
  CLKNAND2HSV2 U30000 ( .A1(n40137), .A2(n39870), .ZN(n40002) );
  NAND3HSV4 U30001 ( .A1(n39875), .A2(n40141), .A3(n39876), .ZN(n40003) );
  XNOR2HSV4 U30002 ( .A1(n26768), .A2(n40004), .ZN(n40014) );
  CLKNAND2HSV3 U30003 ( .A1(n26770), .A2(n26769), .ZN(n40004) );
  CLKNAND2HSV3 U30004 ( .A1(n40000), .A2(n39999), .ZN(n26770) );
  CLKNHSV2 U30005 ( .I(n44264), .ZN(n52120) );
  NOR2HSV4 U30006 ( .A1(n44264), .A2(n26772), .ZN(n26771) );
  CLKNHSV2 U30007 ( .I(n38512), .ZN(n26772) );
  XNOR2HSV4 U30008 ( .A1(n26774), .A2(n38325), .ZN(n26773) );
  CLKNAND2HSV2 U30009 ( .A1(n38510), .A2(n38324), .ZN(n26774) );
  CLKNAND2HSV3 U30010 ( .A1(n26776), .A2(n26775), .ZN(n38736) );
  CLKNAND2HSV2 U30011 ( .A1(n38522), .A2(n38525), .ZN(n26775) );
  CLKNAND2HSV2 U30012 ( .A1(n38521), .A2(n52808), .ZN(n26776) );
  CLKNHSV3 U30013 ( .I(n35603), .ZN(n26780) );
  NAND2HSV2 U30014 ( .A1(n35479), .A2(n46566), .ZN(n26786) );
  CLKNAND2HSV2 U30015 ( .A1(n26778), .A2(n58186), .ZN(n26777) );
  NOR2HSV4 U30016 ( .A1(n35603), .A2(n26788), .ZN(n26778) );
  CLKNHSV2 U30017 ( .I(n26788), .ZN(n26781) );
  AOI21HSV4 U30018 ( .A1(n35480), .A2(n26784), .B(n26783), .ZN(n26782) );
  CLKNHSV2 U30019 ( .I(n26787), .ZN(n26783) );
  CLKNHSV2 U30020 ( .I(n26786), .ZN(n26784) );
  CLKNHSV2 U30021 ( .I(n46565), .ZN(n26785) );
  CLKNHSV2 U30022 ( .I(n35484), .ZN(n26787) );
  CLKNHSV2 U30023 ( .I(n52755), .ZN(n26788) );
  CLKNAND2HSV0 U30024 ( .A1(n52778), .A2(n38885), .ZN(n38378) );
  NOR2HSV4 U30025 ( .A1(n38361), .A2(n38362), .ZN(n38371) );
  OAI21HSV4 U30026 ( .A1(n26794), .A2(n26792), .B(n39366), .ZN(n26791) );
  NAND3HSV4 U30027 ( .A1(n37553), .A2(n39226), .A3(n26793), .ZN(n26792) );
  CLKNHSV2 U30028 ( .I(n39414), .ZN(n26793) );
  CLKNHSV2 U30029 ( .I(n39227), .ZN(n26794) );
  XNOR2HSV4 U30030 ( .A1(n37644), .A2(n37643), .ZN(n39355) );
  CLKNHSV4 U30031 ( .I(n46602), .ZN(n26798) );
  CLKNAND2HSV4 U30032 ( .A1(n26796), .A2(n26795), .ZN(n46602) );
  INHSV2 U30033 ( .I(n33697), .ZN(n26796) );
  INHSV24 U30034 ( .I(n33702), .ZN(n26797) );
  NOR2HSV4 U30035 ( .A1(n26798), .A2(n26797), .ZN(n33679) );
  BUFHSV8 U30036 ( .I(n44313), .Z(n26799) );
  CLKNHSV2 U30037 ( .I(n26799), .ZN(n47938) );
  XNOR2HSV4 U30038 ( .A1(n44306), .A2(n44305), .ZN(n44313) );
  NOR2HSV4 U30039 ( .A1(n60028), .A2(n26799), .ZN(n44294) );
  NOR2HSV4 U30040 ( .A1(n44180), .A2(n26801), .ZN(n26800) );
  OAI21HSV4 U30041 ( .A1(n44179), .A2(n44178), .B(n44177), .ZN(n26801) );
  NOR2HSV4 U30042 ( .A1(n44168), .A2(n45089), .ZN(n44180) );
  CLKNAND2HSV4 U30043 ( .A1(n33408), .A2(n33407), .ZN(n33573) );
  NAND3HSV4 U30044 ( .A1(n33447), .A2(n33446), .A3(n33192), .ZN(n33575) );
  CLKNAND2HSV2 U30045 ( .A1(n26806), .A2(n26803), .ZN(n33460) );
  NAND3HSV1 U30046 ( .A1(n33447), .A2(n33446), .A3(n26804), .ZN(n26803) );
  CLKNHSV2 U30047 ( .I(n26805), .ZN(n26804) );
  CLKNAND2HSV2 U30048 ( .A1(n33192), .A2(n26807), .ZN(n26805) );
  CLKNHSV2 U30049 ( .I(n33457), .ZN(n26807) );
  XOR2HSV2 U30050 ( .A1(n28527), .A2(n26808), .Z(n28528) );
  AOI21HSV4 U30051 ( .A1(n26813), .A2(n26810), .B(n26809), .ZN(n26808) );
  NOR2HSV4 U30052 ( .A1(n26810), .A2(n26813), .ZN(n26809) );
  XNOR2HSV4 U30053 ( .A1(n26812), .A2(n26811), .ZN(n26810) );
  CLKNHSV2 U30054 ( .I(n28526), .ZN(n26811) );
  CLKNAND2HSV2 U30055 ( .A1(n53288), .A2(n51228), .ZN(n26812) );
  NOR2HSV4 U30056 ( .A1(n47139), .A2(n47140), .ZN(n26813) );
  NOR2HSV3 U30057 ( .A1(n38471), .A2(n38337), .ZN(n38338) );
  NAND3HSV3 U30058 ( .A1(n38355), .A2(n38354), .A3(n38183), .ZN(n38337) );
  CLKNHSV0 U30059 ( .I(n38338), .ZN(n52774) );
  NOR2HSV4 U30060 ( .A1(n26816), .A2(n26814), .ZN(n39096) );
  CLKNHSV2 U30061 ( .I(n26815), .ZN(n26814) );
  CLKNAND2HSV2 U30062 ( .A1(n45071), .A2(n26817), .ZN(n26815) );
  MUX2NHSV2 U30063 ( .I0(n26820), .I1(n53086), .S(n26817), .ZN(n26816) );
  XNOR2HSV4 U30064 ( .A1(n26819), .A2(n26818), .ZN(n26817) );
  CLKNHSV2 U30065 ( .I(n39094), .ZN(n26818) );
  AOI21HSV4 U30066 ( .A1(n29766), .A2(n34203), .B(n33849), .ZN(n26822) );
  CLKNHSV0 U30067 ( .I(n40424), .ZN(n40347) );
  XNOR2HSV4 U30068 ( .A1(n26826), .A2(n26824), .ZN(n40377) );
  XOR2HSV2 U30069 ( .A1(n40350), .A2(n40348), .Z(n26824) );
  CLKNAND2HSV2 U30070 ( .A1(n40342), .A2(n26825), .ZN(n40350) );
  CLKNHSV2 U30071 ( .I(n40556), .ZN(n26825) );
  CLKNHSV2 U30072 ( .I(n26828), .ZN(n26827) );
  CLKNAND2HSV2 U30073 ( .A1(n40424), .A2(n41225), .ZN(n26828) );
  XNOR2HSV4 U30074 ( .A1(n40505), .A2(n26829), .ZN(n40528) );
  CLKNHSV2 U30075 ( .I(n26830), .ZN(n26829) );
  CLKNAND2HSV2 U30076 ( .A1(n40786), .A2(n40636), .ZN(n26830) );
  XNOR2HSV4 U30077 ( .A1(n40502), .A2(n40503), .ZN(n40505) );
  CLKNAND2HSV2 U30078 ( .A1(n27835), .A2(n26831), .ZN(n40503) );
  CLKNAND2HSV2 U30079 ( .A1(n26833), .A2(n26832), .ZN(n26831) );
  NOR2HSV4 U30080 ( .A1(n27834), .A2(n44528), .ZN(n26832) );
  CLKNHSV2 U30081 ( .I(n26269), .ZN(n26833) );
  CLKNAND2HSV3 U30082 ( .A1(n30397), .A2(n30396), .ZN(n30568) );
  NOR2HSV4 U30083 ( .A1(n30251), .A2(n26835), .ZN(n26834) );
  CLKNHSV2 U30084 ( .I(n30396), .ZN(n26835) );
  XNOR2HSV4 U30085 ( .A1(n30405), .A2(n30404), .ZN(n30251) );
  XNOR2HSV4 U30086 ( .A1(n30250), .A2(n30249), .ZN(n30404) );
  CLKNHSV2 U30087 ( .I(n38002), .ZN(n26836) );
  OAI21HSV1 U30088 ( .A1(n37927), .A2(n37926), .B(n37924), .ZN(n26838) );
  OAI21HSV4 U30089 ( .A1(n60019), .A2(n44821), .B(n37875), .ZN(n37928) );
  XNOR2HSV4 U30090 ( .A1(n38023), .A2(n36669), .ZN(n60019) );
  BUFHSV8 U30091 ( .I(n41412), .Z(n26839) );
  CLKNHSV2 U30092 ( .I(n44529), .ZN(n55091) );
  XNOR2HSV4 U30093 ( .A1(n26845), .A2(n26840), .ZN(n41707) );
  CLKNAND2HSV2 U30094 ( .A1(n26842), .A2(n26841), .ZN(n26840) );
  AOI31HSV2 U30095 ( .A1(n41699), .A2(n26839), .A3(n42484), .B(n41698), .ZN(
        n26841) );
  CLKNAND2HSV2 U30096 ( .A1(n26844), .A2(n26843), .ZN(n26842) );
  NOR2HSV0 U30097 ( .A1(n41699), .A2(n25448), .ZN(n26843) );
  CLKNAND2HSV2 U30098 ( .A1(n26851), .A2(n44523), .ZN(n26844) );
  XNOR2HSV4 U30099 ( .A1(n41695), .A2(n41694), .ZN(n26846) );
  NOR2HSV4 U30100 ( .A1(n44529), .A2(n26848), .ZN(n26847) );
  CLKNHSV2 U30101 ( .I(n42084), .ZN(n26848) );
  NOR2HSV4 U30102 ( .A1(n29774), .A2(n26849), .ZN(n47791) );
  CLKNHSV2 U30103 ( .I(n58314), .ZN(n26849) );
  INHSV2 U30104 ( .I(n41412), .ZN(n44529) );
  BUFHSV4 U30105 ( .I(n41412), .Z(n26851) );
  CLKNAND2HSV2 U30106 ( .A1(n41415), .A2(n26851), .ZN(n41416) );
  AOI21HSV4 U30107 ( .A1(n38770), .A2(n26852), .B(n38769), .ZN(n52823) );
  CLKNAND2HSV2 U30108 ( .A1(n52847), .A2(n35011), .ZN(n47786) );
  MUX2NHSV2 U30109 ( .I0(n26855), .I1(n26854), .S(n55512), .ZN(n48319) );
  CLKNHSV2 U30110 ( .I(n26858), .ZN(n26854) );
  CLKNHSV2 U30111 ( .I(n26856), .ZN(n26855) );
  CLKNAND2HSV2 U30112 ( .A1(n26858), .A2(n26857), .ZN(n26856) );
  CLKNHSV2 U30113 ( .I(n48310), .ZN(n26857) );
  CLKNAND2HSV2 U30114 ( .A1(n48311), .A2(n48312), .ZN(n26858) );
  NAND2HSV2 U30115 ( .A1(n29776), .A2(n30142), .ZN(n26861) );
  NAND2HSV3 U30116 ( .A1(n47141), .A2(n47052), .ZN(n48309) );
  CLKNAND2HSV4 U30117 ( .A1(pov5[31]), .A2(n44520), .ZN(n47141) );
  XNOR2HSV4 U30118 ( .A1(n26863), .A2(n26860), .ZN(n26859) );
  XNOR2HSV4 U30119 ( .A1(n26862), .A2(n26861), .ZN(n26860) );
  XNOR2HSV4 U30120 ( .A1(n48307), .A2(n48308), .ZN(n26862) );
  CLKNAND2HSV2 U30121 ( .A1(n52668), .A2(n48740), .ZN(n26863) );
  CLKNAND2HSV2 U30122 ( .A1(n48309), .A2(n52799), .ZN(n26864) );
  CLKNHSV4 U30123 ( .I(n33393), .ZN(n33395) );
  CLKNAND2HSV4 U30124 ( .A1(n33412), .A2(n33277), .ZN(n33393) );
  CLKNAND2HSV4 U30125 ( .A1(n33284), .A2(n33283), .ZN(n33384) );
  XOR2HSV2 U30126 ( .A1(n26869), .A2(n26866), .Z(n26865) );
  XNOR2HSV4 U30127 ( .A1(n26867), .A2(n53091), .ZN(n26866) );
  CLKNHSV2 U30128 ( .I(n44710), .ZN(n26868) );
  CLKNHSV2 U30129 ( .I(n52916), .ZN(n26870) );
  OAI21HSV4 U30130 ( .A1(n40315), .A2(n40316), .B(n40314), .ZN(n47388) );
  NAND2HSV3 U30131 ( .A1(n26871), .A2(n47388), .ZN(pov5[31]) );
  CLKNAND2HSV4 U30132 ( .A1(n47392), .A2(n47391), .ZN(n26871) );
  INHSV2 U30133 ( .I(pov5[31]), .ZN(n47196) );
  CLKNAND2HSV4 U30134 ( .A1(n40713), .A2(n40805), .ZN(n40810) );
  CLKNHSV4 U30135 ( .I(n39112), .ZN(n39113) );
  CLKNHSV4 U30136 ( .I(n39110), .ZN(n43917) );
  NAND2HSV4 U30137 ( .A1(n37837), .A2(n36662), .ZN(n37847) );
  NAND3HSV4 U30138 ( .A1(n36325), .A2(n36324), .A3(n36323), .ZN(n36429) );
  AOI21HSV0 U30139 ( .A1(\pe5/ctrq ), .A2(\pe5/pvq [1]), .B(\pe5/phq [1]), 
        .ZN(n29801) );
  CLKNAND2HSV4 U30140 ( .A1(n36401), .A2(n36400), .ZN(n36421) );
  CLKNAND2HSV2 U30141 ( .A1(n60002), .A2(n36414), .ZN(n39106) );
  CLKNAND2HSV4 U30142 ( .A1(n40941), .A2(n40940), .ZN(n40946) );
  NAND3HSV4 U30143 ( .A1(n48007), .A2(n40537), .A3(n40536), .ZN(n40648) );
  CLKNHSV4 U30144 ( .I(n47885), .ZN(n58186) );
  CLKNAND2HSV2 U30145 ( .A1(n38345), .A2(n38108), .ZN(n26872) );
  NAND2HSV2 U30146 ( .A1(n38346), .A2(n26873), .ZN(n38348) );
  CLKNHSV2 U30147 ( .I(n26872), .ZN(n26873) );
  INHSV4 U30148 ( .I(n36570), .ZN(n26874) );
  NAND2HSV2 U30149 ( .A1(n36363), .A2(n36362), .ZN(n60102) );
  NOR2HSV4 U30150 ( .A1(n38339), .A2(n38338), .ZN(n38346) );
  INHSV6 U30151 ( .I(n36577), .ZN(n36570) );
  INOR2HSV2 U30152 ( .A1(n44181), .B1(n44172), .ZN(n44173) );
  NAND2HSV4 U30153 ( .A1(n30752), .A2(n30751), .ZN(n52785) );
  OAI21HSV4 U30154 ( .A1(n31086), .A2(n29133), .B(n30060), .ZN(n39121) );
  CLKAND2HSV4 U30155 ( .A1(n25825), .A2(n44953), .Z(n29680) );
  CLKNAND2HSV4 U30156 ( .A1(n36585), .A2(n36659), .ZN(n37789) );
  INHSV4 U30157 ( .I(n37789), .ZN(n36586) );
  NAND2HSV2 U30158 ( .A1(n38169), .A2(n38168), .ZN(n26877) );
  CLKNAND2HSV4 U30159 ( .A1(n26875), .A2(n26876), .ZN(n26878) );
  NAND2HSV4 U30160 ( .A1(n26877), .A2(n26878), .ZN(n38171) );
  CLKNHSV2 U30161 ( .I(n38169), .ZN(n26875) );
  INHSV4 U30162 ( .I(n38168), .ZN(n26876) );
  CLKNAND2HSV2 U30163 ( .A1(n36638), .A2(n36639), .ZN(n26881) );
  CLKNAND2HSV8 U30164 ( .A1(n26881), .A2(n26882), .ZN(n36647) );
  CLKNHSV2 U30165 ( .I(n36639), .ZN(n26880) );
  NAND2HSV2 U30166 ( .A1(n38166), .A2(n38165), .ZN(n38169) );
  CLKNAND2HSV2 U30167 ( .A1(n36280), .A2(n36279), .ZN(n36287) );
  NAND2HSV4 U30168 ( .A1(n36411), .A2(n36410), .ZN(n36422) );
  NOR2HSV4 U30169 ( .A1(n38471), .A2(n38196), .ZN(n27217) );
  CLKNAND2HSV4 U30170 ( .A1(n40468), .A2(n40467), .ZN(n40700) );
  CLKNAND2HSV4 U30171 ( .A1(n40947), .A2(n40946), .ZN(n40954) );
  INHSV6 U30172 ( .I(n36269), .ZN(n36376) );
  CLKNAND2HSV2 U30173 ( .A1(n40599), .A2(n40600), .ZN(n26886) );
  CLKAND2HSV2 U30174 ( .A1(n41921), .A2(n41922), .Z(n26888) );
  INHSV4 U30175 ( .I(n38468), .ZN(n38469) );
  NAND2HSV0 U30176 ( .A1(n25284), .A2(n59601), .ZN(n34547) );
  CLKNHSV6 U30177 ( .I(n36269), .ZN(n36341) );
  INHSV8 U30178 ( .I(\pe2/ti_1 ), .ZN(n36350) );
  CLKXOR2HSV4 U30179 ( .A1(n48996), .A2(n48995), .Z(n48997) );
  CLKNAND2HSV2 U30180 ( .A1(n33791), .A2(n33790), .ZN(n33792) );
  CLKNAND2HSV2 U30181 ( .A1(n34232), .A2(n47965), .ZN(n34578) );
  CLKNAND2HSV4 U30182 ( .A1(n45135), .A2(n45134), .ZN(n45136) );
  CLKNAND2HSV2 U30183 ( .A1(n35143), .A2(n59955), .ZN(n35005) );
  CLKNAND2HSV4 U30184 ( .A1(n34350), .A2(n34349), .ZN(n34685) );
  CLKNAND2HSV2 U30185 ( .A1(n45262), .A2(n45261), .ZN(n45413) );
  NAND2HSV2 U30186 ( .A1(n41915), .A2(n41914), .ZN(n41917) );
  OAI21HSV2 U30187 ( .A1(n41049), .A2(n41240), .B(n41048), .ZN(n41060) );
  NAND2HSV2 U30188 ( .A1(n40357), .A2(n40356), .ZN(n40354) );
  INHSV4 U30189 ( .I(n45133), .ZN(n45134) );
  CLKNAND2HSV4 U30190 ( .A1(n36433), .A2(n36293), .ZN(n36297) );
  CLKNHSV6 U30191 ( .I(n36299), .ZN(n36269) );
  AND3HSV4 U30192 ( .A1(n40511), .A2(n40526), .A3(n40646), .Z(n29688) );
  CLKNAND2HSV4 U30193 ( .A1(n41051), .A2(n41050), .ZN(n40971) );
  NAND2HSV2 U30194 ( .A1(n36619), .A2(n36661), .ZN(n36463) );
  NAND2HSV0 U30195 ( .A1(n38613), .A2(n38616), .ZN(n26891) );
  INHSV2 U30196 ( .I(n38616), .ZN(n26890) );
  AOI31HSV0 U30197 ( .A1(n38355), .A2(n38354), .A3(n44316), .B(n38353), .ZN(
        n38356) );
  CLKNAND2HSV4 U30198 ( .A1(n26790), .A2(n38457), .ZN(n38606) );
  INHSV2 U30199 ( .I(n36656), .ZN(n36657) );
  NAND2HSV2 U30200 ( .A1(n38097), .A2(n38096), .ZN(n26895) );
  NAND2HSV4 U30201 ( .A1(n26893), .A2(n26894), .ZN(n26896) );
  CLKNAND2HSV4 U30202 ( .A1(n26895), .A2(n26896), .ZN(n38103) );
  CLKNHSV2 U30203 ( .I(n38096), .ZN(n26894) );
  CLKXOR2HSV4 U30204 ( .A1(n38095), .A2(n38094), .Z(n38097) );
  OAI21HSV2 U30205 ( .A1(n26960), .A2(n26961), .B(n26962), .ZN(n26963) );
  OAI21HSV2 U30206 ( .A1(n26957), .A2(n26958), .B(n26959), .ZN(n26960) );
  NAND2HSV2 U30207 ( .A1(n26958), .A2(n26957), .ZN(n26959) );
  OAI21HSV2 U30208 ( .A1(n26954), .A2(n26955), .B(n26956), .ZN(n26957) );
  NAND2HSV2 U30209 ( .A1(n52718), .A2(n29743), .ZN(n36416) );
  NAND2HSV2 U30210 ( .A1(n37928), .A2(n38002), .ZN(n26897) );
  INHSV4 U30211 ( .I(n38115), .ZN(n52749) );
  OAI22HSV2 U30212 ( .A1(n36644), .A2(n36643), .B1(n36642), .B2(n36641), .ZN(
        n36649) );
  NAND3HSV3 U30213 ( .A1(n44176), .A2(n44175), .A3(n44174), .ZN(n45089) );
  NOR2HSV4 U30214 ( .A1(n38515), .A2(n45099), .ZN(n38457) );
  NAND2HSV4 U30215 ( .A1(n37975), .A2(n37846), .ZN(n37927) );
  NAND3HSV2 U30216 ( .A1(n44176), .A2(n44175), .A3(n44174), .ZN(n44817) );
  NAND3HSV4 U30217 ( .A1(n44155), .A2(n29769), .A3(n44312), .ZN(n44175) );
  INHSV6 U30218 ( .I(n38206), .ZN(n38388) );
  NAND2HSV4 U30219 ( .A1(n37978), .A2(n38026), .ZN(n37863) );
  CLKNAND2HSV2 U30220 ( .A1(n38445), .A2(n38447), .ZN(n38197) );
  NOR2HSV2 U30221 ( .A1(n26879), .A2(n36523), .ZN(n36643) );
  NAND2HSV4 U30222 ( .A1(n36470), .A2(n36471), .ZN(n44780) );
  BUFHSV8 U30223 ( .I(n34447), .Z(n34099) );
  NAND2HSV4 U30224 ( .A1(n34700), .A2(n34701), .ZN(n34451) );
  NOR2HSV2 U30225 ( .A1(n30425), .A2(n30424), .ZN(n30508) );
  XNOR4HSV2 U30226 ( .A1(n36681), .A2(n36680), .A3(n36679), .A4(n36678), .ZN(
        n36683) );
  NAND2HSV2 U30227 ( .A1(n30780), .A2(n39249), .ZN(n30395) );
  NAND2HSV2 U30228 ( .A1(n31279), .A2(n31288), .ZN(n31280) );
  INHSV2 U30229 ( .I(n31088), .ZN(n31145) );
  INAND2HSV2 U30230 ( .A1(n42692), .B1(n42691), .ZN(n42696) );
  INHSV2 U30231 ( .I(n37156), .ZN(n37150) );
  NAND2HSV2 U30232 ( .A1(n38461), .A2(n38460), .ZN(n38462) );
  NAND2HSV0 U30233 ( .A1(n36639), .A2(n38183), .ZN(n36523) );
  NOR2HSV2 U30234 ( .A1(n40677), .A2(n41056), .ZN(n40669) );
  INHSV4 U30235 ( .I(\pe2/got [29]), .ZN(n36458) );
  NAND2HSV2 U30236 ( .A1(n46824), .A2(n46760), .ZN(n44363) );
  NAND2HSV2 U30237 ( .A1(n40528), .A2(n40527), .ZN(n40511) );
  NAND2HSV2 U30238 ( .A1(n33224), .A2(n33461), .ZN(n33441) );
  CLKNAND2HSV2 U30239 ( .A1(n40775), .A2(n40774), .ZN(n40780) );
  INHSV2 U30240 ( .I(n40777), .ZN(n40774) );
  INHSV4 U30241 ( .I(n47987), .ZN(n40777) );
  NAND2HSV2 U30242 ( .A1(n40810), .A2(n40714), .ZN(n40715) );
  NAND2HSV2 U30243 ( .A1(n40934), .A2(n40933), .ZN(n40938) );
  NAND2HSV2 U30244 ( .A1(n35457), .A2(n59955), .ZN(n35152) );
  INHSV2 U30245 ( .I(n44294), .ZN(n44954) );
  NAND2HSV2 U30246 ( .A1(n60013), .A2(n52745), .ZN(n47901) );
  NAND2HSV0 U30247 ( .A1(n36557), .A2(n38382), .ZN(n36558) );
  NOR2HSV2 U30248 ( .A1(n37870), .A2(n37869), .ZN(n37987) );
  NAND2HSV2 U30249 ( .A1(n38379), .A2(n38537), .ZN(n38380) );
  INHSV4 U30250 ( .I(n40552), .ZN(n40785) );
  INHSV4 U30251 ( .I(n40534), .ZN(n40639) );
  XOR2HSV0 U30252 ( .A1(n40135), .A2(n40134), .Z(n40148) );
  CLKNAND2HSV2 U30253 ( .A1(n32426), .A2(n32234), .ZN(n32522) );
  OAI21HSV2 U30254 ( .A1(n27675), .A2(n27676), .B(n27677), .ZN(n27678) );
  NAND2HSV2 U30255 ( .A1(n41604), .A2(n47960), .ZN(n41608) );
  NAND2HSV0 U30256 ( .A1(n35915), .A2(n44519), .ZN(n35913) );
  INHSV2 U30257 ( .I(n38368), .ZN(n38861) );
  NAND2HSV2 U30258 ( .A1(n38105), .A2(n38104), .ZN(n38107) );
  NAND2HSV2 U30259 ( .A1(n29749), .A2(n38382), .ZN(n38170) );
  CLKNAND2HSV2 U30260 ( .A1(n37975), .A2(n37848), .ZN(n37855) );
  INAND2HSV2 U30261 ( .A1(n37835), .B1(n37834), .ZN(n37836) );
  CLKNAND2HSV2 U30262 ( .A1(n34847), .A2(n34987), .ZN(n34848) );
  NAND2HSV2 U30263 ( .A1(n57166), .A2(n33190), .ZN(n33194) );
  NAND2HSV2 U30264 ( .A1(n40165), .A2(n40164), .ZN(n40168) );
  NAND2HSV2 U30265 ( .A1(n53524), .A2(n40873), .ZN(n40632) );
  NAND2HSV0 U30266 ( .A1(n41243), .A2(n41212), .ZN(n41046) );
  NAND2HSV2 U30267 ( .A1(n32790), .A2(n29725), .ZN(n32791) );
  OAI21HSV2 U30268 ( .A1(n42346), .A2(n42345), .B(n59394), .ZN(n42351) );
  INHSV4 U30269 ( .I(n34343), .ZN(n34104) );
  MUX2NHSV1 U30270 ( .I0(n28459), .I1(n38616), .S(n28462), .ZN(n38626) );
  NAND2HSV2 U30271 ( .A1(n38537), .A2(n36398), .ZN(n38538) );
  CLKXOR2HSV2 U30272 ( .A1(n40705), .A2(n40704), .Z(n40706) );
  NOR2HSV2 U30273 ( .A1(n26269), .A2(n41228), .ZN(n40425) );
  NAND2HSV4 U30274 ( .A1(n45128), .A2(n45127), .ZN(n53387) );
  NAND3HSV2 U30275 ( .A1(n45126), .A2(n45125), .A3(n45124), .ZN(n45127) );
  NAND2HSV2 U30276 ( .A1(n45126), .A2(n45124), .ZN(n45122) );
  CLKNAND2HSV2 U30277 ( .A1(n45110), .A2(n45109), .ZN(n45121) );
  NAND2HSV2 U30278 ( .A1(n40317), .A2(n37554), .ZN(n40319) );
  INHSV4 U30279 ( .I(\pe4/got [11]), .ZN(n34460) );
  INHSV4 U30280 ( .I(\pe3/got [14]), .ZN(n46042) );
  INHSV2 U30281 ( .I(n39675), .ZN(n37779) );
  NAND2HSV2 U30282 ( .A1(n55513), .A2(n54965), .ZN(n54967) );
  INAND2HSV2 U30283 ( .A1(n55158), .B1(\pe1/got [18]), .ZN(n54966) );
  NAND2HSV2 U30284 ( .A1(n55513), .A2(n54452), .ZN(n54450) );
  NAND2HSV2 U30285 ( .A1(n55537), .A2(\pe1/got [23]), .ZN(n54555) );
  NAND2HSV2 U30286 ( .A1(n55537), .A2(n55331), .ZN(n55374) );
  NAND2HSV4 U30287 ( .A1(n32560), .A2(n32559), .ZN(n32690) );
  NAND2HSV2 U30288 ( .A1(n52697), .A2(n35604), .ZN(n33159) );
  NAND2HSV0 U30289 ( .A1(n36475), .A2(n45005), .ZN(n36442) );
  NOR2HSV2 U30290 ( .A1(n36443), .A2(n38472), .ZN(n36444) );
  NAND3HSV2 U30291 ( .A1(n52756), .A2(n60031), .A3(n34436), .ZN(n33672) );
  INHSV2 U30292 ( .I(n42049), .ZN(n42075) );
  INHSV4 U30293 ( .I(\pe4/aot [17]), .ZN(n35175) );
  XNOR2HSV1 U30294 ( .A1(n33115), .A2(\pe4/phq [4]), .ZN(n33116) );
  NAND2HSV2 U30295 ( .A1(n33306), .A2(n35370), .ZN(n33251) );
  NAND2HSV2 U30296 ( .A1(n33621), .A2(n59523), .ZN(n33252) );
  NAND2HSV0 U30297 ( .A1(n57327), .A2(n35075), .ZN(n33254) );
  INHSV2 U30298 ( .I(\pe2/aot [17]), .ZN(n38946) );
  INHSV2 U30299 ( .I(\pe2/aot [19]), .ZN(n52080) );
  NOR2HSV2 U30300 ( .A1(n44095), .A2(n37953), .ZN(n36482) );
  NAND2HSV2 U30301 ( .A1(n40553), .A2(n40488), .ZN(n40489) );
  INHSV4 U30302 ( .I(n39713), .ZN(n39732) );
  NAND3HSV3 U30303 ( .A1(n35285), .A2(n35284), .A3(n35283), .ZN(n35288) );
  OAI21HSV2 U30304 ( .A1(n35433), .A2(n35432), .B(n35431), .ZN(n35444) );
  NAND2HSV2 U30305 ( .A1(n35432), .A2(n35433), .ZN(n35431) );
  NAND2HSV2 U30306 ( .A1(n33307), .A2(n33263), .ZN(n33264) );
  NAND2HSV4 U30307 ( .A1(pov4[16]), .A2(n33848), .ZN(n34016) );
  AND3HSV2 U30308 ( .A1(n38442), .A2(n38340), .A3(n38441), .Z(n38453) );
  NAND2HSV2 U30309 ( .A1(n38446), .A2(n38445), .ZN(n38450) );
  INAND2HSV2 U30310 ( .A1(n38729), .B1(n38728), .ZN(n38731) );
  INAND2HSV2 U30311 ( .A1(n34854), .B1(n34853), .ZN(n34863) );
  NOR2HSV2 U30312 ( .A1(n34852), .A2(n33098), .ZN(n34853) );
  OAI21HSV2 U30313 ( .A1(n40419), .A2(n40413), .B(n40386), .ZN(n40388) );
  INHSV4 U30314 ( .I(n43236), .ZN(n43344) );
  NAND2HSV2 U30315 ( .A1(\pe2/bq[32] ), .A2(n52449), .ZN(n36275) );
  NAND2HSV4 U30316 ( .A1(n36656), .A2(n36655), .ZN(n36582) );
  NOR2HSV2 U30317 ( .A1(n36513), .A2(n36512), .ZN(n36509) );
  NOR2HSV2 U30318 ( .A1(n45235), .A2(n49000), .ZN(n38868) );
  NAND2HSV0 U30319 ( .A1(n45101), .A2(n45100), .ZN(n45104) );
  INHSV2 U30320 ( .I(n44956), .ZN(n44958) );
  CLKNHSV0 U30321 ( .I(n41117), .ZN(n41118) );
  NAND2HSV2 U30322 ( .A1(n41111), .A2(n41217), .ZN(n41112) );
  NAND3HSV3 U30323 ( .A1(n34996), .A2(n34995), .A3(n34993), .ZN(n35434) );
  INHSV4 U30324 ( .I(\pe4/bq[20] ), .ZN(n48023) );
  NOR2HSV2 U30325 ( .A1(n38371), .A2(n44821), .ZN(n38372) );
  NOR2HSV2 U30326 ( .A1(n36418), .A2(n36417), .ZN(n36420) );
  OAI21HSV2 U30327 ( .A1(n52718), .A2(n29743), .B(n37846), .ZN(n36418) );
  CLKNAND2HSV2 U30328 ( .A1(n40942), .A2(n29653), .ZN(n40861) );
  NAND2HSV4 U30329 ( .A1(n32155), .A2(n32238), .ZN(n52780) );
  NOR2HSV2 U30330 ( .A1(n29774), .A2(n35488), .ZN(n50062) );
  NOR2HSV2 U30331 ( .A1(n29774), .A2(n33749), .ZN(n57582) );
  NOR2HSV2 U30332 ( .A1(n29774), .A2(n35587), .ZN(n50419) );
  NOR2HSV2 U30333 ( .A1(n29774), .A2(n50064), .ZN(n50125) );
  AND2HSV2 U30334 ( .A1(n37765), .A2(n37764), .Z(n37773) );
  NAND2HSV2 U30335 ( .A1(n38036), .A2(n37860), .ZN(n37861) );
  INHSV4 U30336 ( .I(\pe1/got [12]), .ZN(n54879) );
  NAND3HSV2 U30337 ( .A1(n43742), .A2(n43741), .A3(n43740), .ZN(n43878) );
  AOI21HSV2 U30338 ( .A1(n29940), .A2(n52714), .B(n29939), .ZN(n29957) );
  NAND2HSV2 U30339 ( .A1(n40519), .A2(n40518), .ZN(n40538) );
  CLKNAND2HSV2 U30340 ( .A1(n40487), .A2(n40523), .ZN(n40504) );
  CLKNAND2HSV2 U30341 ( .A1(n39716), .A2(n47927), .ZN(n39726) );
  NAND2HSV4 U30342 ( .A1(n44036), .A2(n44035), .ZN(n45083) );
  INHSV4 U30343 ( .I(\pe4/aot [18]), .ZN(n57025) );
  INHSV4 U30344 ( .I(\pe3/aot [19]), .ZN(n42835) );
  NAND2HSV2 U30345 ( .A1(n52856), .A2(n52895), .ZN(n52881) );
  INHSV2 U30346 ( .I(\pe1/aot [27]), .ZN(n41074) );
  NAND2HSV2 U30347 ( .A1(n31135), .A2(n31107), .ZN(n52819) );
  CLKNAND2HSV2 U30348 ( .A1(n33161), .A2(n33160), .ZN(n52699) );
  CLKNAND2HSV2 U30349 ( .A1(n29781), .A2(n34428), .ZN(n52730) );
  NAND2HSV2 U30350 ( .A1(n34008), .A2(n35570), .ZN(n52795) );
  NAND2HSV4 U30351 ( .A1(n38036), .A2(n38004), .ZN(n53386) );
  NOR2HSV2 U30352 ( .A1(n29632), .A2(n44307), .ZN(n37872) );
  CLKNAND2HSV2 U30353 ( .A1(n38363), .A2(n38271), .ZN(n52777) );
  NAND2HSV2 U30354 ( .A1(n41591), .A2(n41590), .ZN(n41603) );
  BUFHSV2 U30355 ( .I(n47957), .Z(n47958) );
  NAND2HSV2 U30356 ( .A1(n29862), .A2(n52717), .ZN(n29863) );
  NAND2HSV2 U30357 ( .A1(n29856), .A2(n29855), .ZN(n29857) );
  NAND2HSV2 U30358 ( .A1(n49381), .A2(n32418), .ZN(n32644) );
  INHSV2 U30359 ( .I(n34339), .ZN(n34583) );
  NAND2HSV2 U30360 ( .A1(n39234), .A2(n39389), .ZN(n39682) );
  NAND2HSV2 U30361 ( .A1(n25849), .A2(n58401), .ZN(n58374) );
  NAND2HSV2 U30362 ( .A1(n55484), .A2(n59755), .ZN(n55610) );
  NAND2HSV2 U30363 ( .A1(n50318), .A2(n57974), .ZN(n47860) );
  XOR2HSV0 U30364 ( .A1(n26899), .A2(n47192), .Z(n47193) );
  XOR2HSV0 U30365 ( .A1(n47191), .A2(n47190), .Z(n26899) );
  XOR2HSV0 U30366 ( .A1(n47189), .A2(n26900), .Z(n47190) );
  XOR2HSV0 U30367 ( .A1(n47188), .A2(n47187), .Z(n26900) );
  XOR2HSV0 U30368 ( .A1(n47186), .A2(n26901), .Z(n47188) );
  XOR2HSV0 U30369 ( .A1(n47185), .A2(n47184), .Z(n26901) );
  NAND2HSV0 U30370 ( .A1(n55589), .A2(n59755), .ZN(n53187) );
  NAND2HSV2 U30371 ( .A1(n43879), .A2(n43878), .ZN(n59515) );
  NOR2HSV2 U30372 ( .A1(n40375), .A2(n40374), .ZN(n40376) );
  NAND2HSV2 U30373 ( .A1(n39697), .A2(n39696), .ZN(n39699) );
  NAND2HSV2 U30374 ( .A1(n39872), .A2(n39580), .ZN(n39696) );
  INHSV4 U30375 ( .I(n51894), .ZN(n59790) );
  XNOR2HSV2 U30376 ( .A1(n51415), .A2(n51414), .ZN(n51417) );
  NOR2HSV2 U30377 ( .A1(n29774), .A2(n50207), .ZN(n50209) );
  NOR2HSV2 U30378 ( .A1(n29774), .A2(n49954), .ZN(n58191) );
  NOR2HSV2 U30379 ( .A1(n58212), .A2(n50214), .ZN(n58214) );
  NOR2HSV2 U30380 ( .A1(n29774), .A2(n50091), .ZN(n58320) );
  INHSV6 U30381 ( .I(n58294), .ZN(n58298) );
  NAND2HSV0 U30382 ( .A1(n56965), .A2(\pe3/got [18]), .ZN(n56336) );
  NOR2HSV2 U30383 ( .A1(n37423), .A2(n42689), .ZN(n42691) );
  NAND2HSV2 U30384 ( .A1(n29866), .A2(n39430), .ZN(n29867) );
  NAND2HSV0 U30385 ( .A1(n30165), .A2(n30029), .ZN(n30030) );
  AOI21HSV2 U30386 ( .A1(n30280), .A2(n59936), .B(n30279), .ZN(n30296) );
  NAND2HSV0 U30387 ( .A1(n30401), .A2(n30684), .ZN(n30402) );
  NAND2HSV0 U30388 ( .A1(n30422), .A2(n52754), .ZN(n30425) );
  NAND3HSV2 U30389 ( .A1(n31087), .A2(n31086), .A3(n31085), .ZN(n31088) );
  AOI21HSV2 U30390 ( .A1(n31145), .A2(n52788), .B(n31090), .ZN(n31092) );
  CLKNAND2HSV2 U30391 ( .A1(n31107), .A2(n31240), .ZN(n31113) );
  NAND2HSV2 U30392 ( .A1(n39537), .A2(n30046), .ZN(n31231) );
  IOA22HSV1 U30393 ( .B1(n31560), .B2(n32589), .A1(n31776), .A2(n31491), .ZN(
        n31492) );
  NAND2HSV0 U30394 ( .A1(n43780), .A2(n59614), .ZN(n36797) );
  NAND3HSV3 U30395 ( .A1(n59364), .A2(n37082), .A3(n37081), .ZN(n37083) );
  NAND2HSV2 U30396 ( .A1(n37174), .A2(n37173), .ZN(n37227) );
  NAND3HSV2 U30397 ( .A1(n39396), .A2(n39680), .A3(n39682), .ZN(n39397) );
  NOR2HSV2 U30398 ( .A1(n43106), .A2(n43231), .ZN(n43108) );
  NAND2HSV2 U30399 ( .A1(n43237), .A2(n43234), .ZN(n43238) );
  NOR2HSV0 U30400 ( .A1(n43871), .A2(n43361), .ZN(n43362) );
  NAND3HSV2 U30401 ( .A1(n31291), .A2(n31290), .A3(n31292), .ZN(n31281) );
  NAND3HSV2 U30402 ( .A1(n42505), .A2(n42504), .A3(n42503), .ZN(n42588) );
  NAND3HSV2 U30403 ( .A1(n42581), .A2(n42580), .A3(n29717), .ZN(n42582) );
  OAI21HSV2 U30404 ( .A1(n36907), .A2(n37089), .B(n36906), .ZN(n36908) );
  NOR2HSV0 U30405 ( .A1(n36984), .A2(n36983), .ZN(n36985) );
  NAND2HSV2 U30406 ( .A1(n37237), .A2(n37236), .ZN(n37240) );
  AOI21HSV2 U30407 ( .A1(n37756), .A2(n40006), .B(n37755), .ZN(n37757) );
  NAND2HSV2 U30408 ( .A1(n29835), .A2(n29877), .ZN(n29839) );
  NAND2HSV2 U30409 ( .A1(n42583), .A2(n42582), .ZN(n42586) );
  NOR2HSV2 U30410 ( .A1(n31123), .A2(n31122), .ZN(n31124) );
  NOR2HSV0 U30411 ( .A1(n42925), .A2(n42919), .ZN(n42920) );
  NAND2HSV2 U30412 ( .A1(n32426), .A2(n29652), .ZN(n32313) );
  NAND2HSV2 U30413 ( .A1(n31389), .A2(n31450), .ZN(n31447) );
  NAND2HSV2 U30414 ( .A1(\pe6/bq[31] ), .A2(\pe6/aot [31]), .ZN(n31330) );
  NAND2HSV2 U30415 ( .A1(n31302), .A2(n31261), .ZN(n31263) );
  NAND2HSV2 U30416 ( .A1(n37325), .A2(n37161), .ZN(n37086) );
  NAND2HSV0 U30417 ( .A1(n36795), .A2(n55987), .ZN(n36796) );
  NAND2HSV2 U30418 ( .A1(n37762), .A2(n37764), .ZN(n37530) );
  XNOR2HSV1 U30419 ( .A1(n31809), .A2(n31808), .ZN(n31810) );
  NOR2HSV2 U30420 ( .A1(n30426), .A2(n30319), .ZN(n30315) );
  NAND2HSV2 U30421 ( .A1(n37420), .A2(n43360), .ZN(n37421) );
  NAND2HSV2 U30422 ( .A1(n30985), .A2(n30984), .ZN(n30986) );
  NAND2HSV2 U30423 ( .A1(n42921), .A2(n42920), .ZN(n42928) );
  NAND2HSV0 U30424 ( .A1(n30288), .A2(n30029), .ZN(n30005) );
  NAND2HSV2 U30425 ( .A1(n31106), .A2(n29697), .ZN(n30979) );
  BUFHSV2 U30426 ( .I(n36783), .Z(n36784) );
  AOI21HSV0 U30427 ( .A1(n33326), .A2(n59661), .B(n34145), .ZN(n26902) );
  AO31HSV2 U30428 ( .A1(n33326), .A2(n59661), .A3(n34145), .B(n26902), .Z(
        n26903) );
  NAND2HSV0 U30429 ( .A1(n33556), .A2(n35370), .ZN(n26904) );
  NAND2HSV2 U30430 ( .A1(n26904), .A2(n26903), .ZN(n26905) );
  OAI21HSV2 U30431 ( .A1(n26903), .A2(n26904), .B(n26905), .ZN(n26906) );
  NAND2HSV0 U30432 ( .A1(n34030), .A2(n57242), .ZN(n26907) );
  NAND2HSV2 U30433 ( .A1(n26907), .A2(n26906), .ZN(n26908) );
  OAI21HSV2 U30434 ( .A1(n26906), .A2(n26907), .B(n26908), .ZN(n33327) );
  NAND2HSV0 U30435 ( .A1(\pe4/bq[20] ), .A2(n35347), .ZN(n26909) );
  NAND2HSV0 U30436 ( .A1(n33711), .A2(n57585), .ZN(n26910) );
  NAND2HSV0 U30437 ( .A1(n26910), .A2(n26909), .ZN(n26911) );
  OAI21HSV2 U30438 ( .A1(n26909), .A2(n26910), .B(n26911), .ZN(n26912) );
  NAND2HSV0 U30439 ( .A1(n33716), .A2(\pe4/bq[12] ), .ZN(n26913) );
  NAND2HSV2 U30440 ( .A1(n26913), .A2(n26912), .ZN(n26914) );
  OAI21HSV2 U30441 ( .A1(n26912), .A2(n26913), .B(n26914), .ZN(n26915) );
  NAND2HSV0 U30442 ( .A1(n57460), .A2(n57504), .ZN(n26916) );
  NAND2HSV2 U30443 ( .A1(n26916), .A2(n26915), .ZN(n26917) );
  OAI21HSV2 U30444 ( .A1(n26915), .A2(n26916), .B(n26917), .ZN(n35540) );
  CLKNAND2HSV0 U30445 ( .A1(n36183), .A2(n44393), .ZN(n26918) );
  CLKNAND2HSV0 U30446 ( .A1(n26918), .A2(n36184), .ZN(n26919) );
  OAI21HSV0 U30447 ( .A1(n36184), .A2(n26918), .B(n26919), .ZN(n26920) );
  NAND2HSV0 U30448 ( .A1(n44477), .A2(n32167), .ZN(n26921) );
  CLKNAND2HSV0 U30449 ( .A1(n26921), .A2(n26920), .ZN(n26922) );
  OAI21HSV0 U30450 ( .A1(n26920), .A2(n26921), .B(n26922), .ZN(n26923) );
  CLKNAND2HSV0 U30451 ( .A1(n36107), .A2(n59180), .ZN(n26924) );
  CLKNAND2HSV0 U30452 ( .A1(n26924), .A2(n26923), .ZN(n26925) );
  OAI21HSV0 U30453 ( .A1(n26923), .A2(n26924), .B(n26925), .ZN(n26926) );
  NAND2HSV0 U30454 ( .A1(n36185), .A2(n58711), .ZN(n26927) );
  CLKNAND2HSV0 U30455 ( .A1(n26927), .A2(n26926), .ZN(n26928) );
  OAI21HSV0 U30456 ( .A1(n26926), .A2(n26927), .B(n26928), .ZN(n26929) );
  CLKNAND2HSV0 U30457 ( .A1(n49319), .A2(\pe6/got [14]), .ZN(n26930) );
  CLKNAND2HSV0 U30458 ( .A1(n26930), .A2(n26929), .ZN(n26931) );
  OAI21HSV0 U30459 ( .A1(n26929), .A2(n26930), .B(n26931), .ZN(n26932) );
  NAND2HSV0 U30460 ( .A1(n49829), .A2(\pe6/got [15]), .ZN(n26933) );
  CLKNAND2HSV0 U30461 ( .A1(n26933), .A2(n26932), .ZN(n26934) );
  OAI21HSV0 U30462 ( .A1(n26932), .A2(n26933), .B(n26934), .ZN(n26935) );
  NAND2HSV0 U30463 ( .A1(n35722), .A2(n36106), .ZN(n26936) );
  CLKNAND2HSV0 U30464 ( .A1(n26936), .A2(n26935), .ZN(n26937) );
  OAI21HSV0 U30465 ( .A1(n26935), .A2(n26936), .B(n26937), .ZN(n26938) );
  CLKNAND2HSV0 U30466 ( .A1(n44392), .A2(n49098), .ZN(n26939) );
  CLKNAND2HSV0 U30467 ( .A1(n26939), .A2(n26938), .ZN(n26940) );
  OAI21HSV0 U30468 ( .A1(n26938), .A2(n26939), .B(n26940), .ZN(n26941) );
  NAND2HSV0 U30469 ( .A1(n36105), .A2(n36104), .ZN(n26942) );
  CLKNAND2HSV0 U30470 ( .A1(n26942), .A2(n26941), .ZN(n26943) );
  OAI21HSV0 U30471 ( .A1(n26941), .A2(n26942), .B(n26943), .ZN(n26944) );
  NAND2HSV0 U30472 ( .A1(n35922), .A2(n46632), .ZN(n26945) );
  CLKNAND2HSV0 U30473 ( .A1(n26945), .A2(n26944), .ZN(n26946) );
  OAI21HSV2 U30474 ( .A1(n26944), .A2(n26945), .B(n26946), .ZN(n36187) );
  NOR2HSV2 U30475 ( .A1(n41700), .A2(n26947), .ZN(n41725) );
  XOR2HSV0 U30476 ( .A1(n38439), .A2(n38438), .Z(n26948) );
  NAND2HSV0 U30477 ( .A1(n39008), .A2(n38510), .ZN(n26949) );
  CLKNAND2HSV0 U30478 ( .A1(n26949), .A2(n26948), .ZN(n26950) );
  OAI21HSV0 U30479 ( .A1(n26948), .A2(n26949), .B(n26950), .ZN(n26951) );
  NAND2HSV0 U30480 ( .A1(n44711), .A2(n52120), .ZN(n26952) );
  CLKNAND2HSV0 U30481 ( .A1(n26952), .A2(n26951), .ZN(n26953) );
  NAND2HSV0 U30482 ( .A1(\pe2/got [27]), .A2(n59583), .ZN(n26958) );
  NAND2HSV0 U30483 ( .A1(n36623), .A2(n29749), .ZN(n26961) );
  CLKNAND2HSV0 U30484 ( .A1(n26961), .A2(n26960), .ZN(n26962) );
  NOR2HSV0 U30485 ( .A1(n43896), .A2(n37268), .ZN(n26964) );
  OAI21HSV0 U30486 ( .A1(\pe2/ti_7t [27]), .A2(n44315), .B(n44314), .ZN(n26965) );
  AOI21HSV2 U30487 ( .A1(n44313), .A2(n44316), .B(n26965), .ZN(n44960) );
  NAND2HSV0 U30488 ( .A1(n33245), .A2(n33507), .ZN(n26966) );
  XOR2HSV0 U30489 ( .A1(n57749), .A2(n57751), .Z(n26967) );
  XOR2HSV0 U30490 ( .A1(n57750), .A2(n26967), .Z(n26968) );
  NAND2HSV0 U30491 ( .A1(n57675), .A2(n58111), .ZN(n26969) );
  CLKNAND2HSV0 U30492 ( .A1(n26969), .A2(n26968), .ZN(n26970) );
  OAI21HSV0 U30493 ( .A1(n26968), .A2(n26969), .B(n26970), .ZN(n26971) );
  NAND2HSV0 U30494 ( .A1(n57818), .A2(n57547), .ZN(n26972) );
  CLKNAND2HSV0 U30495 ( .A1(n26972), .A2(n26971), .ZN(n26973) );
  OAI21HSV0 U30496 ( .A1(n26971), .A2(n26972), .B(n26973), .ZN(n26974) );
  NAND2HSV0 U30497 ( .A1(\pe4/got [10]), .A2(n57550), .ZN(n26975) );
  CLKNAND2HSV0 U30498 ( .A1(n26975), .A2(n26974), .ZN(n26976) );
  OAI21HSV0 U30499 ( .A1(n26974), .A2(n26975), .B(n26976), .ZN(n26977) );
  NAND2HSV0 U30500 ( .A1(n58153), .A2(n57817), .ZN(n26978) );
  CLKNAND2HSV0 U30501 ( .A1(n26978), .A2(n26977), .ZN(n26979) );
  OAI21HSV0 U30502 ( .A1(n26977), .A2(n26978), .B(n26979), .ZN(n26980) );
  NAND2HSV0 U30503 ( .A1(n47657), .A2(n57308), .ZN(n26981) );
  CLKNAND2HSV0 U30504 ( .A1(n26981), .A2(n26980), .ZN(n26982) );
  OAI21HSV0 U30505 ( .A1(n26980), .A2(n26981), .B(n26982), .ZN(n26983) );
  NAND2HSV0 U30506 ( .A1(n58097), .A2(n50189), .ZN(n26984) );
  CLKNAND2HSV0 U30507 ( .A1(n26984), .A2(n26983), .ZN(n26985) );
  OAI21HSV0 U30508 ( .A1(n26983), .A2(n26984), .B(n26985), .ZN(n26986) );
  CLKNAND2HSV0 U30509 ( .A1(n57674), .A2(n58154), .ZN(n26987) );
  CLKNAND2HSV0 U30510 ( .A1(n26987), .A2(n26986), .ZN(n26988) );
  OAI21HSV0 U30511 ( .A1(n26986), .A2(n26987), .B(n26988), .ZN(n26989) );
  CLKNAND2HSV0 U30512 ( .A1(n57974), .A2(n57819), .ZN(n26990) );
  CLKNAND2HSV0 U30513 ( .A1(n26990), .A2(n26989), .ZN(n26991) );
  OAI21HSV2 U30514 ( .A1(n26989), .A2(n26990), .B(n26991), .ZN(n26992) );
  CLKNAND2HSV0 U30515 ( .A1(n57752), .A2(n57960), .ZN(n26993) );
  CLKNAND2HSV0 U30516 ( .A1(n26993), .A2(n26992), .ZN(n26994) );
  OAI21HSV2 U30517 ( .A1(n26992), .A2(n26993), .B(n26994), .ZN(n26995) );
  CLKNAND2HSV0 U30518 ( .A1(n57753), .A2(n58220), .ZN(n26996) );
  CLKNAND2HSV0 U30519 ( .A1(n26996), .A2(n26995), .ZN(n26997) );
  OAI21HSV0 U30520 ( .A1(n26995), .A2(n26996), .B(n26997), .ZN(n26998) );
  CLKNAND2HSV0 U30521 ( .A1(n57755), .A2(n57754), .ZN(n26999) );
  CLKNAND2HSV0 U30522 ( .A1(n26999), .A2(n26998), .ZN(n27000) );
  OAI21HSV0 U30523 ( .A1(n26998), .A2(n26999), .B(n27000), .ZN(n57756) );
  XOR2HSV0 U30524 ( .A1(n45502), .A2(n45501), .Z(n27001) );
  AOI21HSV0 U30525 ( .A1(\pe5/got [25]), .A2(n51272), .B(n27001), .ZN(n27002)
         );
  AO31HSV2 U30526 ( .A1(\pe5/got [25]), .A2(n51272), .A3(n27001), .B(n27002), 
        .Z(n27003) );
  NAND2HSV0 U30527 ( .A1(n51155), .A2(n48742), .ZN(n27004) );
  CLKNAND2HSV0 U30528 ( .A1(n27004), .A2(n27003), .ZN(n27005) );
  OAI21HSV0 U30529 ( .A1(n27003), .A2(n27004), .B(n27005), .ZN(n27006) );
  NAND2HSV0 U30530 ( .A1(n29775), .A2(\pe5/got [27]), .ZN(n27007) );
  CLKNAND2HSV0 U30531 ( .A1(n27007), .A2(n27006), .ZN(n27008) );
  OAI21HSV0 U30532 ( .A1(n27006), .A2(n27007), .B(n27008), .ZN(n27009) );
  NAND2HSV0 U30533 ( .A1(n52562), .A2(n30142), .ZN(n27012) );
  CLKNAND2HSV0 U30534 ( .A1(n27012), .A2(n27011), .ZN(n27013) );
  OAI21HSV0 U30535 ( .A1(n27011), .A2(n27012), .B(n27013), .ZN(\pe5/poht [3])
         );
  NAND2HSV0 U30536 ( .A1(n59260), .A2(n58360), .ZN(n27014) );
  AOI21HSV0 U30537 ( .A1(\pe6/aot [1]), .A2(n58339), .B(n27014), .ZN(n27015)
         );
  AO31HSV2 U30538 ( .A1(\pe6/aot [1]), .A2(n58339), .A3(n27014), .B(n27015), 
        .Z(n27016) );
  NAND2HSV0 U30539 ( .A1(n58336), .A2(n58353), .ZN(n27017) );
  CLKNAND2HSV0 U30540 ( .A1(n27017), .A2(n27016), .ZN(n27018) );
  OAI21HSV0 U30541 ( .A1(n27016), .A2(n27017), .B(n27018), .ZN(n27019) );
  NAND2HSV0 U30542 ( .A1(\pe6/got [1]), .A2(n59024), .ZN(n27020) );
  CLKNAND2HSV0 U30543 ( .A1(n27020), .A2(n27019), .ZN(n27021) );
  OAI21HSV0 U30544 ( .A1(n27019), .A2(n27020), .B(n27021), .ZN(n27022) );
  NAND2HSV0 U30545 ( .A1(n48888), .A2(n58331), .ZN(n27023) );
  CLKNAND2HSV0 U30546 ( .A1(n27023), .A2(n27022), .ZN(n27024) );
  OAI21HSV2 U30547 ( .A1(n27022), .A2(n27023), .B(n27024), .ZN(n27025) );
  CLKNAND2HSV0 U30548 ( .A1(n59023), .A2(n48891), .ZN(n27026) );
  CLKNAND2HSV0 U30549 ( .A1(n27026), .A2(n27025), .ZN(n27027) );
  OAI21HSV0 U30550 ( .A1(n27025), .A2(n27026), .B(n27027), .ZN(\pe6/poht [29])
         );
  OAI22HSV0 U30551 ( .A1(n34479), .A2(n50129), .B1(n50134), .B2(n35043), .ZN(
        n27028) );
  OAI21HSV0 U30552 ( .A1(n34355), .A2(n34248), .B(n27028), .ZN(n27029) );
  NAND2HSV0 U30553 ( .A1(n27029), .A2(n50339), .ZN(n27030) );
  OAI21HSV2 U30554 ( .A1(n27029), .A2(n50339), .B(n27030), .ZN(n33722) );
  XOR2HSV0 U30555 ( .A1(n35756), .A2(n35757), .Z(n27031) );
  XOR2HSV0 U30556 ( .A1(n35749), .A2(n35748), .Z(n27032) );
  XOR2HSV0 U30557 ( .A1(n27031), .A2(n27032), .Z(n27033) );
  XOR2HSV0 U30558 ( .A1(n35771), .A2(n35772), .Z(n27034) );
  XOR2HSV0 U30559 ( .A1(n35765), .A2(n35764), .Z(n27035) );
  XOR2HSV0 U30560 ( .A1(n27034), .A2(n27035), .Z(n27036) );
  XOR2HSV0 U30561 ( .A1(n35737), .A2(n35738), .Z(n27037) );
  XOR2HSV0 U30562 ( .A1(n35731), .A2(n35730), .Z(n27038) );
  XOR2HSV0 U30563 ( .A1(n27037), .A2(n27038), .Z(n27039) );
  CLKNHSV0 U30564 ( .I(n58859), .ZN(n27040) );
  CLKNHSV0 U30565 ( .I(n35739), .ZN(n27041) );
  MUX2NHSV0 U30566 ( .I0(n27041), .I1(n35739), .S(n35741), .ZN(n27042) );
  MUX2NHSV0 U30567 ( .I0(n58859), .I1(n27040), .S(n27042), .ZN(n27043) );
  XOR2HSV0 U30568 ( .A1(n27039), .A2(n35742), .Z(n27044) );
  XOR2HSV0 U30569 ( .A1(n27043), .A2(n27044), .Z(n27045) );
  NAND2HSV0 U30570 ( .A1(n58525), .A2(n35725), .ZN(n27046) );
  CLKNAND2HSV0 U30571 ( .A1(n27046), .A2(n27045), .ZN(n27047) );
  OAI21HSV0 U30572 ( .A1(n27045), .A2(n27046), .B(n27047), .ZN(n27048) );
  XOR2HSV0 U30573 ( .A1(n27033), .A2(n27036), .Z(n27049) );
  XOR2HSV0 U30574 ( .A1(n27048), .A2(n27049), .Z(n27050) );
  NAND2HSV0 U30575 ( .A1(n44393), .A2(n32286), .ZN(n27051) );
  CLKNAND2HSV0 U30576 ( .A1(n27051), .A2(n27050), .ZN(n27052) );
  OAI21HSV0 U30577 ( .A1(n27050), .A2(n27051), .B(n27052), .ZN(n27053) );
  NAND2HSV0 U30578 ( .A1(n35724), .A2(n44477), .ZN(n27054) );
  CLKNAND2HSV0 U30579 ( .A1(n27054), .A2(n27053), .ZN(n27055) );
  OAI21HSV0 U30580 ( .A1(n27053), .A2(n27054), .B(n27055), .ZN(n27056) );
  NAND2HSV0 U30581 ( .A1(n58719), .A2(n59121), .ZN(n27057) );
  CLKNAND2HSV0 U30582 ( .A1(n27057), .A2(n27056), .ZN(n27058) );
  OAI21HSV0 U30583 ( .A1(n27056), .A2(n27057), .B(n27058), .ZN(n27059) );
  NAND2HSV0 U30584 ( .A1(n58811), .A2(n36183), .ZN(n27060) );
  CLKNAND2HSV0 U30585 ( .A1(n27060), .A2(n27059), .ZN(n27061) );
  OAI21HSV0 U30586 ( .A1(n27059), .A2(n27060), .B(n27061), .ZN(n27062) );
  NAND2HSV0 U30587 ( .A1(n58713), .A2(n35813), .ZN(n27063) );
  CLKNAND2HSV0 U30588 ( .A1(n27063), .A2(n27062), .ZN(n27064) );
  OAI21HSV0 U30589 ( .A1(n27062), .A2(n27063), .B(n27064), .ZN(n27065) );
  NAND2HSV0 U30590 ( .A1(n36107), .A2(\pe6/got [15]), .ZN(n27066) );
  CLKNAND2HSV0 U30591 ( .A1(n27066), .A2(n27065), .ZN(n27067) );
  OAI21HSV0 U30592 ( .A1(n27065), .A2(n27066), .B(n27067), .ZN(n27068) );
  CLKNAND2HSV0 U30593 ( .A1(n36106), .A2(n36185), .ZN(n27069) );
  CLKNAND2HSV0 U30594 ( .A1(n27069), .A2(n27068), .ZN(n27070) );
  OAI21HSV2 U30595 ( .A1(n27068), .A2(n27069), .B(n27070), .ZN(n35773) );
  NAND2HSV0 U30596 ( .A1(n34594), .A2(n34405), .ZN(n27071) );
  CLKNAND2HSV0 U30597 ( .A1(n27071), .A2(n34406), .ZN(n27072) );
  OAI21HSV0 U30598 ( .A1(n34406), .A2(n27071), .B(n27072), .ZN(n27073) );
  NAND2HSV0 U30599 ( .A1(n34351), .A2(n34459), .ZN(n27074) );
  CLKNAND2HSV0 U30600 ( .A1(n27074), .A2(n27073), .ZN(n27075) );
  OAI21HSV0 U30601 ( .A1(n27073), .A2(n27074), .B(n27075), .ZN(n27076) );
  NAND2HSV0 U30602 ( .A1(n34239), .A2(n46601), .ZN(n27077) );
  CLKNAND2HSV0 U30603 ( .A1(n27077), .A2(n27076), .ZN(n27078) );
  OAI21HSV0 U30604 ( .A1(n27076), .A2(n27077), .B(n27078), .ZN(n27079) );
  NAND2HSV0 U30605 ( .A1(n59603), .A2(n25894), .ZN(n27080) );
  NAND2HSV0 U30606 ( .A1(n27080), .A2(n27079), .ZN(n27081) );
  OAI21HSV2 U30607 ( .A1(n27079), .A2(n27080), .B(n27081), .ZN(n34407) );
  INHSV4 U30608 ( .I(n25940), .ZN(n27082) );
  XOR2HSV0 U30609 ( .A1(n38509), .A2(n38508), .Z(n27083) );
  XOR2HSV0 U30610 ( .A1(n38511), .A2(n27083), .Z(n27084) );
  AOI21HSV0 U30611 ( .A1(n52120), .A2(n39008), .B(n27084), .ZN(n27085) );
  AO31HSV0 U30612 ( .A1(n52120), .A2(n39008), .A3(n27084), .B(n27085), .Z(
        n27086) );
  CLKNAND2HSV0 U30613 ( .A1(n27087), .A2(n27086), .ZN(n27088) );
  NAND2HSV0 U30614 ( .A1(n38512), .A2(n59583), .ZN(n27089) );
  OAI21HSV0 U30615 ( .A1(n38472), .A2(n27082), .B(n27090), .ZN(n27091) );
  OAI31HSV2 U30616 ( .A1(n38472), .A2(n27090), .A3(n27082), .B(n27091), .ZN(
        n27092) );
  CLKNAND2HSV2 U30617 ( .A1(n51802), .A2(\pe2/got [28]), .ZN(n27093) );
  NAND2HSV2 U30618 ( .A1(n27093), .A2(n27092), .ZN(n27094) );
  NOR2HSV0 U30619 ( .A1(n49000), .A2(n44967), .ZN(n27095) );
  XOR2HSV0 U30620 ( .A1(n49949), .A2(n49950), .Z(n27096) );
  XOR2HSV0 U30621 ( .A1(n49928), .A2(n49927), .Z(n27097) );
  XOR2HSV0 U30622 ( .A1(n27096), .A2(n27097), .Z(n27098) );
  XOR2HSV0 U30623 ( .A1(n49936), .A2(n27098), .Z(n27099) );
  NAND2HSV0 U30624 ( .A1(n58282), .A2(n59526), .ZN(n27100) );
  CLKNAND2HSV0 U30625 ( .A1(n27100), .A2(n27099), .ZN(n27101) );
  OAI21HSV0 U30626 ( .A1(n27099), .A2(n27100), .B(n27101), .ZN(n27102) );
  NAND2HSV0 U30627 ( .A1(n57427), .A2(\pe4/got [2]), .ZN(n27103) );
  CLKNAND2HSV0 U30628 ( .A1(n27103), .A2(n27102), .ZN(n27104) );
  OAI21HSV0 U30629 ( .A1(n27102), .A2(n27103), .B(n27104), .ZN(n27105) );
  NAND2HSV0 U30630 ( .A1(n58258), .A2(n58029), .ZN(n27106) );
  CLKNAND2HSV0 U30631 ( .A1(n27106), .A2(n27105), .ZN(n27107) );
  OAI21HSV0 U30632 ( .A1(n27105), .A2(n27106), .B(n27107), .ZN(n27108) );
  NAND2HSV0 U30633 ( .A1(n58097), .A2(n58298), .ZN(n27109) );
  CLKNAND2HSV0 U30634 ( .A1(n27109), .A2(n27108), .ZN(n27110) );
  OAI21HSV0 U30635 ( .A1(n27108), .A2(n27109), .B(n27110), .ZN(n27111) );
  NAND2HSV0 U30636 ( .A1(n57951), .A2(n50213), .ZN(n27112) );
  CLKNAND2HSV0 U30637 ( .A1(n27112), .A2(n27111), .ZN(n27113) );
  OAI21HSV0 U30638 ( .A1(n27111), .A2(n27112), .B(n27113), .ZN(n27114) );
  CLKNAND2HSV0 U30639 ( .A1(n58216), .A2(n58183), .ZN(n27115) );
  CLKNAND2HSV0 U30640 ( .A1(n27115), .A2(n27114), .ZN(n27116) );
  OAI21HSV2 U30641 ( .A1(n27114), .A2(n27115), .B(n27116), .ZN(n27117) );
  NAND2HSV0 U30642 ( .A1(n58184), .A2(n58037), .ZN(n27118) );
  CLKNAND2HSV0 U30643 ( .A1(n27118), .A2(n27117), .ZN(n27119) );
  OAI21HSV2 U30644 ( .A1(n27117), .A2(n27118), .B(n27119), .ZN(n27120) );
  NAND2HSV0 U30645 ( .A1(n58111), .A2(n58103), .ZN(n27121) );
  CLKNAND2HSV0 U30646 ( .A1(n27121), .A2(n27120), .ZN(n27122) );
  OAI21HSV2 U30647 ( .A1(n27120), .A2(n27121), .B(n27122), .ZN(n27123) );
  NAND2HSV0 U30648 ( .A1(n58140), .A2(n58185), .ZN(n27124) );
  CLKNAND2HSV0 U30649 ( .A1(n27124), .A2(n27123), .ZN(n27125) );
  OAI21HSV0 U30650 ( .A1(n27123), .A2(n27124), .B(n27125), .ZN(n49952) );
  CLKNHSV0 U30651 ( .I(n47933), .ZN(n27126) );
  NAND2HSV0 U30652 ( .A1(n47932), .A2(n27126), .ZN(n27127) );
  OAI211HSV1 U30653 ( .A1(n27126), .A2(n47932), .B(n27127), .C(n48013), .ZN(
        n27128) );
  NAND2HSV0 U30654 ( .A1(n27128), .A2(poh6[28]), .ZN(n27129) );
  OAI21HSV2 U30655 ( .A1(poh6[28]), .A2(n27128), .B(n27129), .ZN(po[29]) );
  XOR2HSV0 U30656 ( .A1(n59019), .A2(n59018), .Z(n27130) );
  XOR2HSV0 U30657 ( .A1(n59020), .A2(n27130), .Z(n27131) );
  NAND2HSV0 U30658 ( .A1(n59028), .A2(n59328), .ZN(n27132) );
  CLKNAND2HSV0 U30659 ( .A1(n27132), .A2(n27131), .ZN(n27133) );
  OAI21HSV0 U30660 ( .A1(n27131), .A2(n27132), .B(n27133), .ZN(n27134) );
  NAND2HSV0 U30661 ( .A1(n58934), .A2(n59175), .ZN(n27135) );
  CLKNAND2HSV0 U30662 ( .A1(n27135), .A2(n27134), .ZN(n27136) );
  OAI21HSV0 U30663 ( .A1(n27134), .A2(n27135), .B(n27136), .ZN(n27137) );
  NAND2HSV0 U30664 ( .A1(n59528), .A2(n59027), .ZN(n27138) );
  CLKNAND2HSV0 U30665 ( .A1(n27138), .A2(n27137), .ZN(n27139) );
  OAI21HSV0 U30666 ( .A1(n27137), .A2(n27138), .B(n27139), .ZN(n27140) );
  NAND2HSV0 U30667 ( .A1(n59026), .A2(n32970), .ZN(n27141) );
  CLKNAND2HSV0 U30668 ( .A1(n27141), .A2(n27140), .ZN(n27142) );
  OAI21HSV0 U30669 ( .A1(n27140), .A2(n27141), .B(n27142), .ZN(n27143) );
  CLKNAND2HSV0 U30670 ( .A1(n59170), .A2(n59173), .ZN(n27144) );
  CLKNAND2HSV0 U30671 ( .A1(n27144), .A2(n27143), .ZN(n27145) );
  OAI21HSV0 U30672 ( .A1(n27143), .A2(n27144), .B(n27145), .ZN(n27146) );
  NAND2HSV0 U30673 ( .A1(n32354), .A2(n59024), .ZN(n27147) );
  CLKNAND2HSV0 U30674 ( .A1(n27147), .A2(n27146), .ZN(n27148) );
  OAI21HSV0 U30675 ( .A1(n27146), .A2(n27147), .B(n27148), .ZN(n27149) );
  NAND2HSV0 U30676 ( .A1(n59022), .A2(n29772), .ZN(n27151) );
  CLKNAND2HSV0 U30677 ( .A1(n27151), .A2(n27150), .ZN(n27152) );
  NAND2HSV0 U30678 ( .A1(n34743), .A2(n33611), .ZN(n27153) );
  AOI21HSV0 U30679 ( .A1(n33969), .A2(n33960), .B(n27153), .ZN(n27154) );
  AO31HSV2 U30680 ( .A1(n33969), .A2(n33960), .A3(n27153), .B(n27154), .Z(
        n27155) );
  NAND2HSV0 U30681 ( .A1(n34598), .A2(n33726), .ZN(n27156) );
  NAND2HSV2 U30682 ( .A1(n27156), .A2(n27155), .ZN(n27157) );
  OAI21HSV2 U30683 ( .A1(n27155), .A2(n27156), .B(n27157), .ZN(n27158) );
  NAND2HSV0 U30684 ( .A1(n33934), .A2(n57859), .ZN(n27159) );
  NAND2HSV2 U30685 ( .A1(n27159), .A2(n27158), .ZN(n27160) );
  OAI21HSV2 U30686 ( .A1(n27158), .A2(n27159), .B(n27160), .ZN(n33734) );
  CLKNHSV0 U30687 ( .I(n35495), .ZN(n27161) );
  CLKNHSV0 U30688 ( .I(n35494), .ZN(n27162) );
  NAND2HSV0 U30689 ( .A1(n57234), .A2(n57929), .ZN(n27163) );
  CLKNAND2HSV0 U30690 ( .A1(n27163), .A2(n57105), .ZN(n27164) );
  OAI21HSV2 U30691 ( .A1(n57105), .A2(n27163), .B(n27164), .ZN(n27165) );
  MUX2NHSV1 U30692 ( .I0(n27162), .I1(n35494), .S(n27165), .ZN(n27166) );
  MUX2NHSV1 U30693 ( .I0(n27161), .I1(n35495), .S(n27166), .ZN(n35496) );
  NAND2HSV0 U30694 ( .A1(\pe4/got [20]), .A2(n34396), .ZN(n27167) );
  CLKAND2HSV4 U30695 ( .A1(n59602), .A2(n34868), .Z(n27168) );
  XOR2HSV0 U30696 ( .A1(n34073), .A2(n34072), .Z(n27169) );
  CLKXOR2HSV2 U30697 ( .A1(n34074), .A2(n27169), .Z(n27170) );
  XOR2HSV4 U30698 ( .A1(n27168), .A2(n27170), .Z(n27171) );
  XOR2HSV4 U30699 ( .A1(n27167), .A2(n27171), .Z(n27172) );
  NAND2HSV0 U30700 ( .A1(n34594), .A2(n57530), .ZN(n27173) );
  XOR2HSV4 U30701 ( .A1(n27172), .A2(n27173), .Z(n34076) );
  NAND2HSV0 U30702 ( .A1(n34593), .A2(n57190), .ZN(n27174) );
  CLKNAND2HSV0 U30703 ( .A1(n27174), .A2(n34407), .ZN(n27175) );
  OAI21HSV0 U30704 ( .A1(n34407), .A2(n27174), .B(n27175), .ZN(n27176) );
  NAND2HSV0 U30705 ( .A1(n47771), .A2(n34007), .ZN(n27177) );
  NAND2HSV0 U30706 ( .A1(n27177), .A2(n27176), .ZN(n27178) );
  OAI21HSV0 U30707 ( .A1(n27176), .A2(n27177), .B(n27178), .ZN(n34413) );
  NAND2HSV0 U30708 ( .A1(n51362), .A2(n30783), .ZN(n27179) );
  CLKNAND2HSV0 U30709 ( .A1(n27179), .A2(n45478), .ZN(n27180) );
  OAI21HSV0 U30710 ( .A1(n45478), .A2(n27179), .B(n27180), .ZN(n27181) );
  NAND2HSV0 U30711 ( .A1(n48169), .A2(n51161), .ZN(n27182) );
  CLKNAND2HSV0 U30712 ( .A1(n27182), .A2(n27181), .ZN(n27183) );
  OAI21HSV0 U30713 ( .A1(n27181), .A2(n27182), .B(n27183), .ZN(n27184) );
  CLKNAND2HSV0 U30714 ( .A1(n51331), .A2(n37659), .ZN(n27185) );
  CLKNAND2HSV0 U30715 ( .A1(n27185), .A2(n27184), .ZN(n27186) );
  OAI21HSV0 U30716 ( .A1(n27184), .A2(n27185), .B(n27186), .ZN(n27187) );
  CLKNAND2HSV0 U30717 ( .A1(n48750), .A2(n51302), .ZN(n27188) );
  CLKNAND2HSV0 U30718 ( .A1(n27188), .A2(n27187), .ZN(n27189) );
  OAI21HSV0 U30719 ( .A1(n27187), .A2(n27188), .B(n27189), .ZN(n27190) );
  CLKNAND2HSV0 U30720 ( .A1(n48841), .A2(n47338), .ZN(n27191) );
  CLKNAND2HSV0 U30721 ( .A1(n27191), .A2(n27190), .ZN(n27192) );
  OAI21HSV0 U30722 ( .A1(n27190), .A2(n27191), .B(n27192), .ZN(n27193) );
  NAND2HSV0 U30723 ( .A1(n52580), .A2(n51200), .ZN(n27194) );
  CLKNAND2HSV0 U30724 ( .A1(n27194), .A2(n27193), .ZN(n27195) );
  OAI21HSV0 U30725 ( .A1(n27193), .A2(n27194), .B(n27195), .ZN(n27196) );
  NAND2HSV0 U30726 ( .A1(n51159), .A2(n51162), .ZN(n27197) );
  CLKNAND2HSV0 U30727 ( .A1(n27197), .A2(n27196), .ZN(n27198) );
  OAI21HSV0 U30728 ( .A1(n27196), .A2(n27197), .B(n27198), .ZN(n27199) );
  NAND2HSV0 U30729 ( .A1(n29770), .A2(n50698), .ZN(n27200) );
  CLKNAND2HSV0 U30730 ( .A1(n27200), .A2(n27199), .ZN(n27201) );
  OAI21HSV0 U30731 ( .A1(n27199), .A2(n27200), .B(n27201), .ZN(n27202) );
  NAND2HSV0 U30732 ( .A1(n52641), .A2(n48748), .ZN(n27203) );
  CLKNAND2HSV0 U30733 ( .A1(n27203), .A2(n27202), .ZN(n27204) );
  OAI21HSV0 U30734 ( .A1(n27202), .A2(n27203), .B(n27204), .ZN(n27205) );
  CLKNAND2HSV0 U30735 ( .A1(n52574), .A2(n52571), .ZN(n27206) );
  CLKNAND2HSV0 U30736 ( .A1(n27206), .A2(n27205), .ZN(n27207) );
  OAI21HSV0 U30737 ( .A1(n27205), .A2(n27206), .B(n27207), .ZN(n27208) );
  CLKNAND2HSV0 U30738 ( .A1(n48749), .A2(n51160), .ZN(n27209) );
  CLKNAND2HSV0 U30739 ( .A1(n27209), .A2(n27208), .ZN(n27210) );
  OAI21HSV0 U30740 ( .A1(n27208), .A2(n27209), .B(n27210), .ZN(n27211) );
  NAND2HSV0 U30741 ( .A1(n48167), .A2(n44694), .ZN(n27212) );
  CLKNAND2HSV0 U30742 ( .A1(n27212), .A2(n27211), .ZN(n27213) );
  OAI21HSV0 U30743 ( .A1(n27211), .A2(n27212), .B(n27213), .ZN(n27214) );
  CLKNAND2HSV0 U30744 ( .A1(n52568), .A2(n52572), .ZN(n27215) );
  CLKNAND2HSV0 U30745 ( .A1(n27215), .A2(n27214), .ZN(n27216) );
  OAI21HSV0 U30746 ( .A1(n27214), .A2(n27215), .B(n27216), .ZN(n45480) );
  AOI21HSV2 U30747 ( .A1(n27217), .A2(n38337), .B(n38899), .ZN(n38445) );
  NAND2HSV0 U30748 ( .A1(\pe4/got [11]), .A2(n58272), .ZN(n27218) );
  CLKNAND2HSV0 U30749 ( .A1(n59837), .A2(n58140), .ZN(n27219) );
  NAND2HSV0 U30750 ( .A1(n58103), .A2(n58102), .ZN(n27220) );
  CLKNHSV0 U30751 ( .I(n58101), .ZN(n27222) );
  NAND2HSV0 U30752 ( .A1(n34967), .A2(n58030), .ZN(n27223) );
  MUX2NHSV0 U30753 ( .I0(n58101), .I1(n27222), .S(n27223), .ZN(n27224) );
  XOR2HSV0 U30754 ( .A1(n27221), .A2(n27224), .Z(n27225) );
  NAND2HSV0 U30755 ( .A1(n59672), .A2(n58246), .ZN(n27226) );
  XOR2HSV0 U30756 ( .A1(n27225), .A2(n27226), .Z(n27227) );
  XOR2HSV0 U30757 ( .A1(n27220), .A2(n27227), .Z(n27228) );
  NAND2HSV0 U30758 ( .A1(n58111), .A2(n58185), .ZN(n27229) );
  XOR2HSV0 U30759 ( .A1(n27228), .A2(n27229), .Z(n27230) );
  XOR2HSV0 U30760 ( .A1(n27219), .A2(n27230), .Z(n27231) );
  XOR2HSV0 U30761 ( .A1(n27218), .A2(n27233), .Z(n27234) );
  CLKNAND2HSV0 U30762 ( .A1(n26516), .A2(n58110), .ZN(n27235) );
  XOR2HSV0 U30763 ( .A1(n27234), .A2(n27235), .Z(n58105) );
  CLKNHSV0 U30764 ( .I(n45401), .ZN(n27236) );
  NAND2HSV0 U30765 ( .A1(n58448), .A2(n46587), .ZN(n27237) );
  CLKNHSV0 U30766 ( .I(n46590), .ZN(n27238) );
  CLKNHSV0 U30767 ( .I(n46588), .ZN(n27239) );
  MUX2NHSV0 U30768 ( .I0(n27239), .I1(n46588), .S(n46589), .ZN(n27240) );
  MUX2NHSV0 U30769 ( .I0(n27238), .I1(n46590), .S(n27240), .ZN(n27241) );
  NAND2HSV0 U30770 ( .A1(n27241), .A2(n27237), .ZN(n27242) );
  OAI211HSV1 U30771 ( .A1(n27237), .A2(n27241), .B(n27242), .C(n48013), .ZN(
        n27243) );
  NAND2HSV0 U30772 ( .A1(n27243), .A2(poh6[23]), .ZN(n27244) );
  OAI21HSV2 U30773 ( .A1(poh6[23]), .A2(n27243), .B(n27244), .ZN(po[24]) );
  XOR2HSV0 U30774 ( .A1(n47266), .A2(n47265), .Z(n27245) );
  AOI21HSV0 U30775 ( .A1(n31149), .A2(n47268), .B(n27245), .ZN(n27246) );
  AO31HSV2 U30776 ( .A1(n31149), .A2(n47268), .A3(n27245), .B(n27246), .Z(
        n27247) );
  NAND2HSV0 U30777 ( .A1(n59535), .A2(n47267), .ZN(n27248) );
  CLKNAND2HSV0 U30778 ( .A1(n27248), .A2(n27247), .ZN(n27249) );
  OAI21HSV0 U30779 ( .A1(n27247), .A2(n27248), .B(n27249), .ZN(n27250) );
  CLKNAND2HSV0 U30780 ( .A1(n52564), .A2(n47200), .ZN(n27251) );
  CLKNAND2HSV0 U30781 ( .A1(n27251), .A2(n27250), .ZN(n27252) );
  OAI21HSV0 U30782 ( .A1(n27250), .A2(n27251), .B(n27252), .ZN(n27253) );
  NAND2HSV0 U30783 ( .A1(n52563), .A2(n37654), .ZN(n27254) );
  CLKNAND2HSV0 U30784 ( .A1(n27254), .A2(n27253), .ZN(n27255) );
  OAI21HSV0 U30785 ( .A1(n27253), .A2(n27254), .B(n27255), .ZN(n27256) );
  NAND2HSV0 U30786 ( .A1(n29777), .A2(n37630), .ZN(n27257) );
  CLKNAND2HSV0 U30787 ( .A1(n27257), .A2(n27256), .ZN(n27258) );
  OAI21HSV0 U30788 ( .A1(n27256), .A2(n27257), .B(n27258), .ZN(n27259) );
  NAND2HSV0 U30789 ( .A1(n59580), .A2(n48742), .ZN(n27260) );
  CLKNAND2HSV0 U30790 ( .A1(n27260), .A2(n27259), .ZN(n27261) );
  OAI21HSV0 U30791 ( .A1(n27259), .A2(n27260), .B(n27261), .ZN(n27262) );
  NAND2HSV0 U30792 ( .A1(n59421), .A2(n31225), .ZN(n27263) );
  CLKNAND2HSV0 U30793 ( .A1(n27263), .A2(n27262), .ZN(n27264) );
  OAI21HSV0 U30794 ( .A1(n27262), .A2(n27263), .B(n27264), .ZN(\pe5/poht [5])
         );
  CLKNHSV0 U30795 ( .I(n58395), .ZN(n27265) );
  MUX2NHSV0 U30796 ( .I0(n27265), .I1(n58395), .S(n58396), .ZN(n27266) );
  XOR2HSV0 U30797 ( .A1(n58397), .A2(n27266), .Z(n27267) );
  NAND2HSV0 U30798 ( .A1(n58402), .A2(n58403), .ZN(n27268) );
  CLKNAND2HSV0 U30799 ( .A1(n27268), .A2(n27267), .ZN(n27269) );
  OAI21HSV0 U30800 ( .A1(n27267), .A2(n27268), .B(n27269), .ZN(n27270) );
  NAND2HSV0 U30801 ( .A1(n29753), .A2(n58816), .ZN(n27271) );
  CLKNAND2HSV0 U30802 ( .A1(n27271), .A2(n27270), .ZN(n27272) );
  OAI21HSV0 U30803 ( .A1(n27270), .A2(n27271), .B(n27272), .ZN(n27273) );
  NAND2HSV0 U30804 ( .A1(n58423), .A2(n58385), .ZN(n27274) );
  CLKNAND2HSV0 U30805 ( .A1(n27274), .A2(n27273), .ZN(n27275) );
  OAI21HSV0 U30806 ( .A1(n27273), .A2(n27274), .B(n27275), .ZN(n27276) );
  NAND2HSV0 U30807 ( .A1(n58656), .A2(n58401), .ZN(n27277) );
  CLKNAND2HSV0 U30808 ( .A1(n27277), .A2(n27276), .ZN(n27278) );
  OAI21HSV0 U30809 ( .A1(n27276), .A2(n27277), .B(n27278), .ZN(n27279) );
  NAND2HSV0 U30810 ( .A1(n58384), .A2(n59169), .ZN(n27280) );
  CLKNAND2HSV0 U30811 ( .A1(n27280), .A2(n27279), .ZN(n27281) );
  OAI21HSV0 U30812 ( .A1(n27279), .A2(n27280), .B(n27281), .ZN(n27282) );
  NAND2HSV0 U30813 ( .A1(n58398), .A2(n48888), .ZN(n27283) );
  CLKNAND2HSV0 U30814 ( .A1(n27283), .A2(n27282), .ZN(n27284) );
  OAI21HSV2 U30815 ( .A1(n27282), .A2(n27283), .B(n27284), .ZN(n27285) );
  NAND2HSV0 U30816 ( .A1(n36109), .A2(n59340), .ZN(n27286) );
  CLKNAND2HSV0 U30817 ( .A1(n27286), .A2(n27285), .ZN(n27287) );
  OAI21HSV0 U30818 ( .A1(n27285), .A2(n27286), .B(n27287), .ZN(\pe6/poht [25])
         );
  XOR2HSV0 U30819 ( .A1(n33353), .A2(n33354), .Z(n27288) );
  XOR2HSV0 U30820 ( .A1(n33352), .A2(n33351), .Z(n27289) );
  XOR2HSV0 U30821 ( .A1(n27288), .A2(n27289), .Z(n27290) );
  CLKNHSV0 U30822 ( .I(n33812), .ZN(n27291) );
  CLKNHSV0 U30823 ( .I(n34148), .ZN(n27292) );
  MUX2NHSV0 U30824 ( .I0(n27292), .I1(n34148), .S(n33349), .ZN(n27293) );
  MUX2NHSV0 U30825 ( .I0(n27291), .I1(n33812), .S(n27293), .ZN(n27294) );
  XOR2HSV0 U30826 ( .A1(n27294), .A2(\pe4/phq [15]), .Z(n27295) );
  XOR2HSV0 U30827 ( .A1(n27290), .A2(n33347), .Z(n27296) );
  XOR2HSV0 U30828 ( .A1(n27295), .A2(n27296), .Z(n27297) );
  NAND2HSV0 U30829 ( .A1(n33831), .A2(n57359), .ZN(n27298) );
  NAND2HSV0 U30830 ( .A1(n27298), .A2(n27297), .ZN(n27299) );
  OAI21HSV2 U30831 ( .A1(n27297), .A2(n27298), .B(n27299), .ZN(n33373) );
  XOR2HSV0 U30832 ( .A1(n45580), .A2(n45578), .Z(n27300) );
  XOR2HSV0 U30833 ( .A1(n45577), .A2(n45579), .Z(n27301) );
  XOR2HSV0 U30834 ( .A1(n27300), .A2(n27301), .Z(n27302) );
  AOI21HSV0 U30835 ( .A1(n59965), .A2(n45732), .B(n27302), .ZN(n27303) );
  AO31HSV2 U30836 ( .A1(n59965), .A2(n45732), .A3(n27302), .B(n27303), .Z(
        n27304) );
  NAND2HSV0 U30837 ( .A1(n45636), .A2(n55945), .ZN(n27305) );
  CLKNAND2HSV0 U30838 ( .A1(n27305), .A2(n27304), .ZN(n27306) );
  OAI21HSV0 U30839 ( .A1(n27304), .A2(n27305), .B(n27306), .ZN(n27307) );
  NAND2HSV0 U30840 ( .A1(n46052), .A2(n45581), .ZN(n27308) );
  CLKNAND2HSV0 U30841 ( .A1(n27308), .A2(n27307), .ZN(n27309) );
  OAI21HSV0 U30842 ( .A1(n27307), .A2(n27308), .B(n27309), .ZN(n27310) );
  NAND2HSV0 U30843 ( .A1(n45582), .A2(n48483), .ZN(n27311) );
  CLKNAND2HSV0 U30844 ( .A1(n27311), .A2(n27310), .ZN(n27312) );
  OAI21HSV0 U30845 ( .A1(n27310), .A2(n27311), .B(n27312), .ZN(n27313) );
  CLKNAND2HSV0 U30846 ( .A1(n56624), .A2(n55821), .ZN(n27314) );
  CLKNAND2HSV0 U30847 ( .A1(n27314), .A2(n27313), .ZN(n27315) );
  OAI21HSV0 U30848 ( .A1(n27313), .A2(n27314), .B(n27315), .ZN(n27316) );
  NAND2HSV0 U30849 ( .A1(n56066), .A2(n59617), .ZN(n27317) );
  CLKNAND2HSV0 U30850 ( .A1(n27317), .A2(n27316), .ZN(n27318) );
  OAI21HSV0 U30851 ( .A1(n27316), .A2(n27317), .B(n27318), .ZN(n27319) );
  CLKNAND2HSV0 U30852 ( .A1(n45634), .A2(n46312), .ZN(n27320) );
  CLKNAND2HSV0 U30853 ( .A1(n27320), .A2(n27319), .ZN(n27321) );
  OAI21HSV0 U30854 ( .A1(n27319), .A2(n27320), .B(n27321), .ZN(n27322) );
  AOI21HSV0 U30855 ( .A1(n34003), .A2(n33998), .B(n33696), .ZN(n27323) );
  NAND2HSV0 U30856 ( .A1(n34196), .A2(n27323), .ZN(n33999) );
  INOR2HSV1 U30857 ( .A1(n38387), .B1(n52772), .ZN(n38269) );
  INOR2HSV0 U30858 ( .A1(n46121), .B1(n38886), .ZN(n38604) );
  NAND2HSV0 U30859 ( .A1(n44715), .A2(n38781), .ZN(n27324) );
  CLKNAND2HSV0 U30860 ( .A1(n27324), .A2(n38589), .ZN(n27325) );
  OAI21HSV0 U30861 ( .A1(n38589), .A2(n27324), .B(n27325), .ZN(n27326) );
  NAND2HSV0 U30862 ( .A1(n38702), .A2(\pe2/got [19]), .ZN(n27327) );
  CLKNAND2HSV0 U30863 ( .A1(n27327), .A2(n27326), .ZN(n27328) );
  OAI21HSV0 U30864 ( .A1(n27326), .A2(n27327), .B(n27328), .ZN(n27329) );
  NAND2HSV0 U30865 ( .A1(n39010), .A2(n45290), .ZN(n27330) );
  CLKNAND2HSV0 U30866 ( .A1(n27330), .A2(n27329), .ZN(n27331) );
  OAI21HSV0 U30867 ( .A1(n27329), .A2(n27330), .B(n27331), .ZN(n27332) );
  NAND2HSV0 U30868 ( .A1(n39011), .A2(n52167), .ZN(n27333) );
  CLKNAND2HSV0 U30869 ( .A1(n27333), .A2(n27332), .ZN(n27334) );
  OAI21HSV0 U30870 ( .A1(n27332), .A2(n27333), .B(n27334), .ZN(n27335) );
  NAND2HSV0 U30871 ( .A1(n52367), .A2(n43925), .ZN(n27336) );
  CLKNAND2HSV0 U30872 ( .A1(n27336), .A2(n27335), .ZN(n27337) );
  OAI21HSV0 U30873 ( .A1(n27335), .A2(n27336), .B(n27337), .ZN(n27338) );
  NAND2HSV0 U30874 ( .A1(n45218), .A2(n43924), .ZN(n27339) );
  CLKNAND2HSV0 U30875 ( .A1(n27339), .A2(n27338), .ZN(n27340) );
  OAI21HSV0 U30876 ( .A1(n27338), .A2(n27339), .B(n27340), .ZN(n27341) );
  NAND2HSV0 U30877 ( .A1(\pe2/got [24]), .A2(n38780), .ZN(n27342) );
  CLKNAND2HSV0 U30878 ( .A1(n27342), .A2(n27341), .ZN(n27343) );
  OAI21HSV2 U30879 ( .A1(n27341), .A2(n27342), .B(n27343), .ZN(n38591) );
  XOR2HSV0 U30880 ( .A1(n49678), .A2(n49679), .Z(n27344) );
  XOR2HSV0 U30881 ( .A1(n49673), .A2(n49672), .Z(n27345) );
  XOR2HSV0 U30882 ( .A1(n27344), .A2(n27345), .Z(n27346) );
  CLKNHSV0 U30883 ( .I(n49683), .ZN(n27347) );
  CLKNHSV0 U30884 ( .I(n49685), .ZN(n27348) );
  CLKNHSV0 U30885 ( .I(n59188), .ZN(n27349) );
  MUX2NHSV0 U30886 ( .I0(n27349), .I1(n59188), .S(n49684), .ZN(n27350) );
  MUX2NHSV0 U30887 ( .I0(n27348), .I1(n49685), .S(n27350), .ZN(n27351) );
  MUX2NHSV0 U30888 ( .I0(n27347), .I1(n49683), .S(n27351), .ZN(n27352) );
  XOR2HSV0 U30889 ( .A1(n49698), .A2(n49690), .Z(n27353) );
  XOR2HSV0 U30890 ( .A1(n27352), .A2(n49691), .Z(n27354) );
  XOR2HSV0 U30891 ( .A1(n27353), .A2(n27354), .Z(n27355) );
  XOR2HSV0 U30892 ( .A1(n27355), .A2(n49712), .Z(n27356) );
  XOR2HSV0 U30893 ( .A1(n27346), .A2(n49713), .Z(n27357) );
  XOR2HSV0 U30894 ( .A1(n27356), .A2(n27357), .Z(n27358) );
  NAND2HSV0 U30895 ( .A1(n58817), .A2(n59594), .ZN(n27359) );
  CLKNAND2HSV0 U30896 ( .A1(n27359), .A2(n27358), .ZN(n27360) );
  OAI21HSV0 U30897 ( .A1(n27358), .A2(n27359), .B(n27360), .ZN(n27361) );
  NAND2HSV0 U30898 ( .A1(n59039), .A2(n59121), .ZN(n27362) );
  CLKNAND2HSV0 U30899 ( .A1(n27362), .A2(n27361), .ZN(n27363) );
  OAI21HSV0 U30900 ( .A1(n27361), .A2(n27362), .B(n27363), .ZN(n27364) );
  CLKNAND2HSV0 U30901 ( .A1(n58423), .A2(n59295), .ZN(n27365) );
  CLKNAND2HSV0 U30902 ( .A1(n27365), .A2(n27364), .ZN(n27366) );
  OAI21HSV0 U30903 ( .A1(n27364), .A2(n27365), .B(n27366), .ZN(n27367) );
  NAND2HSV0 U30904 ( .A1(\pe6/got [4]), .A2(n59183), .ZN(n27368) );
  CLKNAND2HSV0 U30905 ( .A1(n27368), .A2(n27367), .ZN(n27369) );
  OAI21HSV0 U30906 ( .A1(n27367), .A2(n27368), .B(n27369), .ZN(n27370) );
  CLKNAND2HSV0 U30907 ( .A1(n58661), .A2(n59678), .ZN(n27371) );
  CLKNAND2HSV0 U30908 ( .A1(n27371), .A2(n27370), .ZN(n27372) );
  OAI21HSV0 U30909 ( .A1(n27370), .A2(n27371), .B(n27372), .ZN(n27373) );
  NAND2HSV0 U30910 ( .A1(n58723), .A2(n59917), .ZN(n27374) );
  CLKNAND2HSV0 U30911 ( .A1(n27374), .A2(n27373), .ZN(n27375) );
  OAI21HSV0 U30912 ( .A1(n27373), .A2(n27374), .B(n27375), .ZN(n27376) );
  CLKNAND2HSV0 U30913 ( .A1(n27377), .A2(n27376), .ZN(n27378) );
  OAI21HSV0 U30914 ( .A1(n27376), .A2(n27377), .B(n27378), .ZN(n27379) );
  NAND2HSV0 U30915 ( .A1(n58526), .A2(n58815), .ZN(n27380) );
  CLKNAND2HSV0 U30916 ( .A1(n27380), .A2(n27379), .ZN(n27381) );
  OAI21HSV0 U30917 ( .A1(n27379), .A2(n27380), .B(n27381), .ZN(n27382) );
  NAND2HSV0 U30918 ( .A1(n59037), .A2(n59036), .ZN(n27383) );
  CLKNAND2HSV0 U30919 ( .A1(n27383), .A2(n27382), .ZN(n27384) );
  OAI21HSV0 U30920 ( .A1(n27382), .A2(n27383), .B(n27384), .ZN(n27385) );
  NAND2HSV0 U30921 ( .A1(\pe6/got [10]), .A2(n44392), .ZN(n27386) );
  CLKNAND2HSV0 U30922 ( .A1(n27386), .A2(n27385), .ZN(n27387) );
  OAI21HSV0 U30923 ( .A1(n27385), .A2(n27386), .B(n27387), .ZN(n27388) );
  NAND2HSV0 U30924 ( .A1(n59033), .A2(n59181), .ZN(n27389) );
  CLKNAND2HSV0 U30925 ( .A1(n27389), .A2(n27388), .ZN(n27390) );
  OAI21HSV0 U30926 ( .A1(n27388), .A2(n27389), .B(n27390), .ZN(n49714) );
  CLKNHSV0 U30927 ( .I(n57231), .ZN(n27391) );
  MUX2NHSV0 U30928 ( .I0(n27391), .I1(n57231), .S(n47906), .ZN(n27392) );
  XOR2HSV0 U30929 ( .A1(n47919), .A2(n27392), .Z(n27393) );
  XOR2HSV0 U30930 ( .A1(n47918), .A2(n47917), .Z(n27394) );
  XOR2HSV0 U30931 ( .A1(n27393), .A2(n27394), .Z(n27395) );
  NAND2HSV0 U30932 ( .A1(n58300), .A2(n58183), .ZN(n27396) );
  CLKNAND2HSV0 U30933 ( .A1(n27396), .A2(n27395), .ZN(n27397) );
  OAI21HSV0 U30934 ( .A1(n27395), .A2(n27396), .B(n27397), .ZN(n27398) );
  NAND2HSV0 U30935 ( .A1(n58314), .A2(n47904), .ZN(n27399) );
  CLKNAND2HSV0 U30936 ( .A1(n27399), .A2(n27398), .ZN(n27400) );
  OAI21HSV0 U30937 ( .A1(n27398), .A2(n27399), .B(n27400), .ZN(n27401) );
  NAND2HSV0 U30938 ( .A1(\pe4/got [3]), .A2(n35033), .ZN(n27402) );
  CLKNAND2HSV0 U30939 ( .A1(n27402), .A2(n27401), .ZN(n27403) );
  OAI21HSV0 U30940 ( .A1(n27401), .A2(n27402), .B(n27403), .ZN(n27404) );
  NAND2HSV0 U30941 ( .A1(n58193), .A2(n58258), .ZN(n27405) );
  CLKNAND2HSV0 U30942 ( .A1(n27405), .A2(n27404), .ZN(n27406) );
  OAI21HSV0 U30943 ( .A1(n27404), .A2(n27405), .B(n27406), .ZN(n27407) );
  NAND2HSV0 U30944 ( .A1(n58246), .A2(n58104), .ZN(n27408) );
  CLKNAND2HSV0 U30945 ( .A1(n27408), .A2(n27407), .ZN(n27409) );
  OAI21HSV2 U30946 ( .A1(n27407), .A2(n27408), .B(n27409), .ZN(n27410) );
  NAND2HSV0 U30947 ( .A1(n58272), .A2(n58184), .ZN(n27411) );
  NAND2HSV2 U30948 ( .A1(n27411), .A2(n27410), .ZN(n27412) );
  OAI21HSV2 U30949 ( .A1(n27410), .A2(n27411), .B(n27412), .ZN(n27413) );
  NAND2HSV0 U30950 ( .A1(n58216), .A2(n58207), .ZN(n27414) );
  CLKNAND2HSV0 U30951 ( .A1(n27414), .A2(n27413), .ZN(n27415) );
  OAI21HSV2 U30952 ( .A1(n27413), .A2(n27414), .B(n27415), .ZN(n47921) );
  NAND2HSV0 U30953 ( .A1(n47950), .A2(n47951), .ZN(n27416) );
  NAND2HSV0 U30954 ( .A1(n27416), .A2(poh6[21]), .ZN(n27417) );
  OAI21HSV2 U30955 ( .A1(poh6[21]), .A2(n27416), .B(n27417), .ZN(po[22]) );
  NAND2HSV0 U30956 ( .A1(n48013), .A2(n47961), .ZN(n27418) );
  NAND2HSV0 U30957 ( .A1(n27418), .A2(poh6[19]), .ZN(n27419) );
  OAI21HSV2 U30958 ( .A1(poh6[19]), .A2(n27418), .B(n27419), .ZN(po[20]) );
  XOR2HSV0 U30959 ( .A1(n51483), .A2(n51482), .Z(n27420) );
  XOR2HSV0 U30960 ( .A1(n51484), .A2(n27420), .Z(n27421) );
  AOI21HSV0 U30961 ( .A1(n25834), .A2(n52890), .B(n27421), .ZN(n27422) );
  AO31HSV2 U30962 ( .A1(n51797), .A2(n52890), .A3(n27421), .B(n27422), .Z(
        n27423) );
  NAND2HSV0 U30963 ( .A1(n52048), .A2(n59371), .ZN(n27424) );
  CLKNAND2HSV0 U30964 ( .A1(n27424), .A2(n27423), .ZN(n27425) );
  OAI21HSV0 U30965 ( .A1(n27423), .A2(n27424), .B(n27425), .ZN(n27426) );
  NAND2HSV0 U30966 ( .A1(n52414), .A2(n52052), .ZN(n27427) );
  NAND2HSV0 U30967 ( .A1(n51892), .A2(n59794), .ZN(n27431) );
  CLKNAND2HSV0 U30968 ( .A1(n27431), .A2(n27430), .ZN(n27432) );
  OAI21HSV0 U30969 ( .A1(n27430), .A2(n27431), .B(n27432), .ZN(\pe2/poht [21])
         );
  XOR2HSV0 U30970 ( .A1(n45899), .A2(n45898), .Z(n27433) );
  NAND2HSV0 U30971 ( .A1(n53290), .A2(n39433), .ZN(n27434) );
  CLKNAND2HSV0 U30972 ( .A1(n27434), .A2(n27433), .ZN(n27435) );
  OAI21HSV0 U30973 ( .A1(n27433), .A2(n27434), .B(n27435), .ZN(n27436) );
  NAND2HSV0 U30974 ( .A1(n52693), .A2(n47056), .ZN(n27437) );
  CLKNAND2HSV0 U30975 ( .A1(n27437), .A2(n27436), .ZN(n27438) );
  OAI21HSV0 U30976 ( .A1(n27436), .A2(n27437), .B(n27438), .ZN(n27439) );
  NAND2HSV0 U30977 ( .A1(n53288), .A2(n45816), .ZN(n27440) );
  CLKNAND2HSV0 U30978 ( .A1(n27440), .A2(n27439), .ZN(n27441) );
  OAI21HSV0 U30979 ( .A1(n27439), .A2(n27440), .B(n27441), .ZN(n27442) );
  NAND2HSV0 U30980 ( .A1(n53287), .A2(n40170), .ZN(n27443) );
  CLKNAND2HSV0 U30981 ( .A1(n27443), .A2(n27442), .ZN(n27444) );
  OAI21HSV0 U30982 ( .A1(n27442), .A2(n27443), .B(n27444), .ZN(n27445) );
  NAND2HSV0 U30983 ( .A1(n48744), .A2(n29779), .ZN(n27446) );
  CLKNAND2HSV0 U30984 ( .A1(n27446), .A2(n27445), .ZN(n27447) );
  OAI21HSV0 U30985 ( .A1(n27445), .A2(n27446), .B(n27447), .ZN(n27448) );
  NAND2HSV0 U30986 ( .A1(n59580), .A2(\pe5/got [23]), .ZN(n27449) );
  CLKNAND2HSV0 U30987 ( .A1(n27449), .A2(n27448), .ZN(n27450) );
  CLKNAND2HSV0 U30988 ( .A1(n48309), .A2(\pe5/got [24]), .ZN(n27452) );
  OAI21HSV0 U30989 ( .A1(n27451), .A2(n27452), .B(n27453), .ZN(\pe5/poht [8])
         );
  NAND2HSV0 U30990 ( .A1(n59028), .A2(n59027), .ZN(n27454) );
  CLKNAND2HSV0 U30991 ( .A1(n27454), .A2(n59164), .ZN(n27455) );
  OAI21HSV0 U30992 ( .A1(n59164), .A2(n27454), .B(n27455), .ZN(n27456) );
  NAND2HSV0 U30993 ( .A1(n58934), .A2(n59165), .ZN(n27457) );
  CLKNAND2HSV0 U30994 ( .A1(n27457), .A2(n27456), .ZN(n27458) );
  OAI21HSV0 U30995 ( .A1(n27456), .A2(n27457), .B(n27458), .ZN(n27459) );
  CLKNAND2HSV0 U30996 ( .A1(n27460), .A2(n27459), .ZN(n27461) );
  OAI21HSV0 U30997 ( .A1(n27459), .A2(n27460), .B(n27461), .ZN(n27462) );
  NAND2HSV0 U30998 ( .A1(n59026), .A2(n59025), .ZN(n27463) );
  CLKNAND2HSV0 U30999 ( .A1(n27463), .A2(n27462), .ZN(n27464) );
  OAI21HSV0 U31000 ( .A1(n27462), .A2(n27463), .B(n27464), .ZN(n27465) );
  NAND2HSV0 U31001 ( .A1(n59170), .A2(n32815), .ZN(n27466) );
  CLKNAND2HSV0 U31002 ( .A1(n27466), .A2(n27465), .ZN(n27467) );
  OAI21HSV0 U31003 ( .A1(n27465), .A2(n27466), .B(n27467), .ZN(n27468) );
  CLKNAND2HSV0 U31004 ( .A1(n33061), .A2(n59024), .ZN(n27469) );
  CLKNAND2HSV0 U31005 ( .A1(n27469), .A2(n27468), .ZN(n27470) );
  OAI21HSV0 U31006 ( .A1(n27468), .A2(n27469), .B(n27470), .ZN(n27471) );
  NAND2HSV0 U31007 ( .A1(n59167), .A2(n59166), .ZN(n27472) );
  CLKNAND2HSV0 U31008 ( .A1(n27472), .A2(n27471), .ZN(n27473) );
  OAI21HSV0 U31009 ( .A1(n27471), .A2(n27472), .B(n27473), .ZN(n27474) );
  NAND2HSV0 U31010 ( .A1(n59168), .A2(n59340), .ZN(n27475) );
  CLKNAND2HSV0 U31011 ( .A1(n27475), .A2(n27474), .ZN(n27476) );
  OAI21HSV0 U31012 ( .A1(n27474), .A2(n27475), .B(n27476), .ZN(\pe6/poht [2])
         );
  OAI22HSV0 U31013 ( .A1(n57026), .A2(n48024), .B1(n57326), .B2(n47809), .ZN(
        n27477) );
  OAI21HSV0 U31014 ( .A1(n34919), .A2(n57708), .B(n27477), .ZN(n27478) );
  CLKNAND2HSV0 U31015 ( .A1(n27478), .A2(n57112), .ZN(n27479) );
  OAI21HSV0 U31016 ( .A1(n27478), .A2(n57112), .B(n27479), .ZN(n34774) );
  AOI22HSV0 U31017 ( .A1(n44750), .A2(\pe2/bq[16] ), .B1(n38792), .B2(n59588), 
        .ZN(n27480) );
  AOI21HSV0 U31018 ( .A1(n52938), .A2(n44729), .B(n27480), .ZN(n27481) );
  AOI21HSV0 U31019 ( .A1(\pe2/pvq [17]), .A2(n59497), .B(\pe2/phq [17]), .ZN(
        n27482) );
  AO31HSV2 U31020 ( .A1(\pe2/pvq [17]), .A2(n59497), .A3(\pe2/phq [17]), .B(
        n27482), .Z(n27483) );
  XOR2HSV0 U31021 ( .A1(n27481), .A2(n27483), .Z(n38399) );
  CLKNAND2HSV0 U31022 ( .A1(n40890), .A2(n54824), .ZN(n27484) );
  AOI21HSV0 U31023 ( .A1(n40889), .A2(n59385), .B(n27484), .ZN(n27485) );
  AO31HSV2 U31024 ( .A1(n40889), .A2(n59385), .A3(n27484), .B(n27485), .Z(
        n40894) );
  NAND2HSV4 U31025 ( .A1(n36584), .A2(n36583), .ZN(n36659) );
  CLKNHSV0 U31026 ( .I(n47310), .ZN(n27486) );
  MUX2NHSV0 U31027 ( .I0(n27486), .I1(n47310), .S(n47239), .ZN(n27487) );
  XOR2HSV0 U31028 ( .A1(n47228), .A2(n47229), .Z(n27488) );
  XOR2HSV0 U31029 ( .A1(n47215), .A2(n47214), .Z(n27489) );
  XOR2HSV0 U31030 ( .A1(n27488), .A2(n27489), .Z(n27490) );
  XOR2HSV0 U31031 ( .A1(n27490), .A2(n27487), .Z(n27491) );
  XOR2HSV0 U31032 ( .A1(n47235), .A2(n47240), .Z(n27492) );
  XOR2HSV0 U31033 ( .A1(n27491), .A2(n27492), .Z(n27493) );
  CLKNHSV0 U31034 ( .I(n47314), .ZN(n27494) );
  MUX2NHSV0 U31035 ( .I0(n47314), .I1(n27494), .S(n50510), .ZN(n27495) );
  XOR2HSV0 U31036 ( .A1(n47243), .A2(n27493), .Z(n27496) );
  XOR2HSV0 U31037 ( .A1(n27495), .A2(n27496), .Z(n27497) );
  NAND2HSV0 U31038 ( .A1(n51362), .A2(n37659), .ZN(n27498) );
  CLKNAND2HSV0 U31039 ( .A1(n27498), .A2(n27497), .ZN(n27499) );
  OAI21HSV0 U31040 ( .A1(n27497), .A2(n27498), .B(n27499), .ZN(n27500) );
  NAND2HSV0 U31041 ( .A1(n39654), .A2(n51161), .ZN(n27501) );
  CLKNAND2HSV0 U31042 ( .A1(n27501), .A2(n27500), .ZN(n27502) );
  OAI21HSV0 U31043 ( .A1(n27500), .A2(n27501), .B(n27502), .ZN(n27503) );
  CLKNAND2HSV0 U31044 ( .A1(n52579), .A2(n47338), .ZN(n27504) );
  CLKNAND2HSV0 U31045 ( .A1(n27504), .A2(n27503), .ZN(n27505) );
  OAI21HSV0 U31046 ( .A1(n27503), .A2(n27504), .B(n27505), .ZN(n27506) );
  NAND2HSV0 U31047 ( .A1(n52580), .A2(n52577), .ZN(n27507) );
  CLKNAND2HSV0 U31048 ( .A1(n27507), .A2(n27506), .ZN(n27508) );
  OAI21HSV0 U31049 ( .A1(n27506), .A2(n27507), .B(n27508), .ZN(n27509) );
  NAND2HSV0 U31050 ( .A1(n51334), .A2(n52578), .ZN(n27510) );
  CLKNAND2HSV0 U31051 ( .A1(n27510), .A2(n27509), .ZN(n27511) );
  OAI21HSV0 U31052 ( .A1(n27509), .A2(n27510), .B(n27511), .ZN(n27512) );
  NAND2HSV0 U31053 ( .A1(n29770), .A2(n51200), .ZN(n27513) );
  CLKNAND2HSV0 U31054 ( .A1(n27513), .A2(n27512), .ZN(n27514) );
  OAI21HSV2 U31055 ( .A1(n27512), .A2(n27513), .B(n27514), .ZN(n27515) );
  NAND2HSV0 U31056 ( .A1(n52575), .A2(n52573), .ZN(n27516) );
  NAND2HSV2 U31057 ( .A1(n27516), .A2(n27515), .ZN(n27517) );
  OAI21HSV2 U31058 ( .A1(n27515), .A2(n27516), .B(n27517), .ZN(n27518) );
  NAND2HSV0 U31059 ( .A1(n52574), .A2(n50698), .ZN(n27519) );
  CLKNAND2HSV0 U31060 ( .A1(n27519), .A2(n27518), .ZN(n27520) );
  OAI21HSV0 U31061 ( .A1(n27518), .A2(n27519), .B(n27520), .ZN(n47244) );
  AOI21HSV2 U31062 ( .A1(n45623), .A2(n43891), .B(n45624), .ZN(n27521) );
  INOR2HSV0 U31063 ( .A1(\pe2/ti_7t [15]), .B1(n44309), .ZN(n38270) );
  XOR2HSV0 U31064 ( .A1(n33060), .A2(n33059), .Z(n27522) );
  NAND2HSV0 U31065 ( .A1(n46172), .A2(n35812), .ZN(n27523) );
  CLKNAND2HSV0 U31066 ( .A1(n27523), .A2(n27522), .ZN(n27524) );
  OAI21HSV0 U31067 ( .A1(n27522), .A2(n27523), .B(n27524), .ZN(n27525) );
  NAND2HSV0 U31068 ( .A1(n59032), .A2(n32970), .ZN(n27526) );
  CLKNAND2HSV0 U31069 ( .A1(n27526), .A2(n27525), .ZN(n27527) );
  OAI21HSV0 U31070 ( .A1(n27525), .A2(n27526), .B(n27527), .ZN(n27528) );
  NAND2HSV0 U31071 ( .A1(n59144), .A2(n31710), .ZN(n27529) );
  CLKNAND2HSV0 U31072 ( .A1(n27529), .A2(n27528), .ZN(n27530) );
  OAI21HSV0 U31073 ( .A1(n27528), .A2(n27529), .B(n27530), .ZN(n27531) );
  CLKNAND2HSV0 U31074 ( .A1(n35775), .A2(\pe6/got [26]), .ZN(n27532) );
  CLKNAND2HSV0 U31075 ( .A1(n27532), .A2(n27531), .ZN(n27533) );
  OAI21HSV2 U31076 ( .A1(n27531), .A2(n27532), .B(n27533), .ZN(n27534) );
  NAND2HSV0 U31077 ( .A1(n35721), .A2(n32815), .ZN(n27535) );
  NAND2HSV0 U31078 ( .A1(n27535), .A2(n27534), .ZN(n27536) );
  OAI21HSV2 U31079 ( .A1(n27534), .A2(n27535), .B(n27536), .ZN(n27537) );
  NAND2HSV2 U31080 ( .A1(n36102), .A2(n33061), .ZN(n27538) );
  NAND2HSV2 U31081 ( .A1(n27538), .A2(n27537), .ZN(n27539) );
  OAI21HSV2 U31082 ( .A1(n27537), .A2(n27538), .B(n27539), .ZN(n27540) );
  CLKNAND2HSV0 U31083 ( .A1(n46170), .A2(n35705), .ZN(n27541) );
  NAND2HSV2 U31084 ( .A1(n27541), .A2(n27540), .ZN(n27542) );
  OAI21HSV2 U31085 ( .A1(n27540), .A2(n27541), .B(n27542), .ZN(n46589) );
  INOR2HSV0 U31086 ( .A1(\pe4/ti_7t [22]), .B1(n35011), .ZN(n34860) );
  XOR2HSV0 U31087 ( .A1(n56660), .A2(n56661), .Z(n27543) );
  XOR2HSV0 U31088 ( .A1(n56639), .A2(n56638), .Z(n27544) );
  XOR2HSV0 U31089 ( .A1(n27543), .A2(n27544), .Z(n27545) );
  CLKNAND2HSV0 U31090 ( .A1(n59821), .A2(n56862), .ZN(n27546) );
  CLKNAND2HSV0 U31091 ( .A1(n27546), .A2(n27545), .ZN(n27547) );
  OAI21HSV0 U31092 ( .A1(n27545), .A2(n27546), .B(n27547), .ZN(n27548) );
  NAND2HSV0 U31093 ( .A1(n59811), .A2(\pe3/got [1]), .ZN(n27549) );
  CLKNAND2HSV0 U31094 ( .A1(n27549), .A2(n27548), .ZN(n27550) );
  OAI21HSV0 U31095 ( .A1(n27548), .A2(n27549), .B(n27550), .ZN(n27551) );
  NAND2HSV0 U31096 ( .A1(n56624), .A2(n56735), .ZN(n27552) );
  CLKNAND2HSV0 U31097 ( .A1(n27552), .A2(n27551), .ZN(n27553) );
  OAI21HSV0 U31098 ( .A1(n27551), .A2(n27552), .B(n27553), .ZN(n27554) );
  NAND2HSV0 U31099 ( .A1(n56662), .A2(n56684), .ZN(n27555) );
  CLKNAND2HSV0 U31100 ( .A1(n27555), .A2(n27554), .ZN(n27556) );
  OAI21HSV0 U31101 ( .A1(n27554), .A2(n27555), .B(n27556), .ZN(n27557) );
  NAND2HSV0 U31102 ( .A1(n56685), .A2(n56623), .ZN(n27558) );
  CLKNAND2HSV0 U31103 ( .A1(n27558), .A2(n27557), .ZN(n27559) );
  OAI21HSV0 U31104 ( .A1(n27557), .A2(n27558), .B(n27559), .ZN(n27560) );
  NAND2HSV0 U31105 ( .A1(n56779), .A2(n56737), .ZN(n27561) );
  CLKNAND2HSV0 U31106 ( .A1(n27561), .A2(n27560), .ZN(n27562) );
  OAI21HSV0 U31107 ( .A1(n27560), .A2(n27561), .B(n27562), .ZN(n27563) );
  CLKNAND2HSV0 U31108 ( .A1(n56622), .A2(n56266), .ZN(n27564) );
  CLKNAND2HSV0 U31109 ( .A1(n27564), .A2(n27563), .ZN(n27565) );
  OAI21HSV2 U31110 ( .A1(n27563), .A2(n27564), .B(n27565), .ZN(n27566) );
  NAND2HSV0 U31111 ( .A1(n56736), .A2(n56855), .ZN(n27567) );
  CLKNAND2HSV0 U31112 ( .A1(n27567), .A2(n27566), .ZN(n27568) );
  OAI21HSV0 U31113 ( .A1(n27566), .A2(n27567), .B(n27568), .ZN(n56663) );
  XOR2HSV0 U31114 ( .A1(n47647), .A2(n47646), .Z(n27569) );
  XOR2HSV0 U31115 ( .A1(n47649), .A2(n27569), .Z(n27570) );
  AOI21HSV0 U31116 ( .A1(n51889), .A2(n51797), .B(n27570), .ZN(n27571) );
  AO31HSV2 U31117 ( .A1(n51889), .A2(n51797), .A3(n27570), .B(n27571), .Z(
        n27572) );
  NAND2HSV0 U31118 ( .A1(n51120), .A2(n59685), .ZN(n27573) );
  CLKNAND2HSV0 U31119 ( .A1(n27573), .A2(n27572), .ZN(n27574) );
  NAND2HSV0 U31120 ( .A1(n52854), .A2(n52922), .ZN(n27575) );
  NAND2HSV0 U31121 ( .A1(n53097), .A2(n43924), .ZN(n27580) );
  CLKNAND2HSV0 U31122 ( .A1(n27580), .A2(n27579), .ZN(n27581) );
  OAI21HSV0 U31123 ( .A1(n27579), .A2(n27580), .B(n27581), .ZN(\pe2/poht [9])
         );
  XOR2HSV0 U31124 ( .A1(n46973), .A2(n46972), .Z(n27582) );
  AOI21HSV0 U31125 ( .A1(n51224), .A2(n59892), .B(n27582), .ZN(n27583) );
  AO31HSV2 U31126 ( .A1(n51224), .A2(n59892), .A3(n27582), .B(n27583), .Z(
        n27584) );
  NAND2HSV0 U31127 ( .A1(n52693), .A2(n46974), .ZN(n27585) );
  CLKNAND2HSV0 U31128 ( .A1(n27585), .A2(n27584), .ZN(n27586) );
  OAI21HSV0 U31129 ( .A1(n27584), .A2(n27585), .B(n27586), .ZN(n27587) );
  NAND2HSV0 U31130 ( .A1(n53288), .A2(n39433), .ZN(n27588) );
  CLKNAND2HSV0 U31131 ( .A1(n27588), .A2(n27587), .ZN(n27589) );
  OAI21HSV0 U31132 ( .A1(n27587), .A2(n27588), .B(n27589), .ZN(n27590) );
  NAND2HSV0 U31133 ( .A1(n53287), .A2(n47056), .ZN(n27591) );
  CLKNAND2HSV0 U31134 ( .A1(n27591), .A2(n27590), .ZN(n27592) );
  OAI21HSV0 U31135 ( .A1(n27590), .A2(n27591), .B(n27592), .ZN(n27593) );
  NAND2HSV0 U31136 ( .A1(n29775), .A2(\pe5/got [20]), .ZN(n27594) );
  CLKNAND2HSV0 U31137 ( .A1(n27594), .A2(n27593), .ZN(n27595) );
  OAI21HSV0 U31138 ( .A1(n27593), .A2(n27594), .B(n27595), .ZN(n27596) );
  NAND2HSV0 U31139 ( .A1(n59580), .A2(n40170), .ZN(n27597) );
  CLKNAND2HSV0 U31140 ( .A1(n27597), .A2(n27596), .ZN(n27598) );
  OAI21HSV0 U31141 ( .A1(n27596), .A2(n27597), .B(n27598), .ZN(n27599) );
  NAND2HSV0 U31142 ( .A1(n59421), .A2(n47267), .ZN(n27600) );
  CLKNAND2HSV0 U31143 ( .A1(n27600), .A2(n27599), .ZN(n27601) );
  OAI21HSV0 U31144 ( .A1(n27599), .A2(n27600), .B(n27601), .ZN(\pe5/poht [10])
         );
  XOR2HSV0 U31145 ( .A1(n58610), .A2(n58609), .Z(n27602) );
  NAND2HSV0 U31146 ( .A1(n58611), .A2(n58659), .ZN(n27603) );
  CLKNAND2HSV0 U31147 ( .A1(n27603), .A2(n27602), .ZN(n27604) );
  OAI21HSV0 U31148 ( .A1(n27602), .A2(n27603), .B(n27604), .ZN(n27605) );
  CLKNAND2HSV0 U31149 ( .A1(n53109), .A2(n58709), .ZN(n27606) );
  CLKNAND2HSV0 U31150 ( .A1(n27606), .A2(n27605), .ZN(n27607) );
  OAI21HSV0 U31151 ( .A1(n27605), .A2(n27606), .B(n27607), .ZN(n27608) );
  CLKNAND2HSV0 U31152 ( .A1(n27609), .A2(n27608), .ZN(n27610) );
  OAI21HSV0 U31153 ( .A1(n27608), .A2(n27609), .B(n27610), .ZN(n27611) );
  CLKNAND2HSV0 U31154 ( .A1(n58657), .A2(\pe6/got [9]), .ZN(n27612) );
  CLKNAND2HSV0 U31155 ( .A1(n27612), .A2(n27611), .ZN(n27613) );
  OAI21HSV0 U31156 ( .A1(n27611), .A2(n27612), .B(n27613), .ZN(n27614) );
  NAND2HSV0 U31157 ( .A1(n58576), .A2(n58812), .ZN(n27615) );
  CLKNAND2HSV0 U31158 ( .A1(n27615), .A2(n27614), .ZN(n27616) );
  OAI21HSV0 U31159 ( .A1(n27614), .A2(n27615), .B(n27616), .ZN(n27617) );
  CLKNAND2HSV0 U31160 ( .A1(n58720), .A2(n58575), .ZN(n27618) );
  CLKNAND2HSV0 U31161 ( .A1(n27618), .A2(n27617), .ZN(n27619) );
  OAI21HSV0 U31162 ( .A1(n27617), .A2(n27618), .B(n27619), .ZN(n27620) );
  NAND2HSV0 U31163 ( .A1(n48888), .A2(\pe6/got [12]), .ZN(n27621) );
  CLKNAND2HSV0 U31164 ( .A1(n27621), .A2(n27620), .ZN(n27622) );
  OAI21HSV0 U31165 ( .A1(n27620), .A2(n27621), .B(n27622), .ZN(n27623) );
  CLKNAND2HSV0 U31166 ( .A1(n27623), .A2(n27624), .ZN(n27625) );
  OAI21HSV0 U31167 ( .A1(n27623), .A2(n27624), .B(n27625), .ZN(\pe6/poht [19])
         );
  XOR2HSV0 U31168 ( .A1(n45530), .A2(n45531), .Z(n27626) );
  XOR2HSV0 U31169 ( .A1(n45524), .A2(n45523), .Z(n27627) );
  XOR2HSV0 U31170 ( .A1(n27626), .A2(n27627), .Z(n27628) );
  CLKNAND2HSV0 U31171 ( .A1(n59648), .A2(n59799), .ZN(n27629) );
  CLKNAND2HSV0 U31172 ( .A1(n27629), .A2(n27628), .ZN(n27630) );
  OAI21HSV0 U31173 ( .A1(n27628), .A2(n27629), .B(n27630), .ZN(n27631) );
  XOR2HSV0 U31174 ( .A1(n45574), .A2(n45575), .Z(n27632) );
  XOR2HSV0 U31175 ( .A1(n45571), .A2(n45570), .Z(n27633) );
  XOR2HSV0 U31176 ( .A1(n27632), .A2(n27633), .Z(n27634) );
  XOR2HSV0 U31177 ( .A1(n27634), .A2(n45562), .Z(n27635) );
  XOR2HSV0 U31178 ( .A1(n27631), .A2(n45563), .Z(n27636) );
  XOR2HSV0 U31179 ( .A1(n27635), .A2(n27636), .Z(n27637) );
  NAND2HSV0 U31180 ( .A1(n59647), .A2(n48511), .ZN(n27638) );
  CLKNAND2HSV0 U31181 ( .A1(n27638), .A2(n27637), .ZN(n27639) );
  OAI21HSV0 U31182 ( .A1(n27637), .A2(n27638), .B(n27639), .ZN(n27640) );
  NAND2HSV0 U31183 ( .A1(n45950), .A2(n48487), .ZN(n27641) );
  CLKNAND2HSV0 U31184 ( .A1(n27641), .A2(n27640), .ZN(n27642) );
  OAI21HSV0 U31185 ( .A1(n27640), .A2(n27641), .B(n27642), .ZN(n27643) );
  NAND2HSV0 U31186 ( .A1(n56855), .A2(n37316), .ZN(n27644) );
  CLKNAND2HSV0 U31187 ( .A1(n27644), .A2(n27643), .ZN(n27645) );
  OAI21HSV0 U31188 ( .A1(n27643), .A2(n27644), .B(n27645), .ZN(n27646) );
  NAND2HSV0 U31189 ( .A1(n59645), .A2(n42938), .ZN(n27647) );
  CLKNAND2HSV0 U31190 ( .A1(n27647), .A2(n27646), .ZN(n27648) );
  OAI21HSV0 U31191 ( .A1(n27646), .A2(n27647), .B(n27648), .ZN(n27649) );
  NAND2HSV0 U31192 ( .A1(n56619), .A2(n55707), .ZN(n27650) );
  CLKNAND2HSV0 U31193 ( .A1(n27650), .A2(n27649), .ZN(n27651) );
  OAI21HSV0 U31194 ( .A1(n27649), .A2(n27650), .B(n27651), .ZN(n27652) );
  NAND2HSV0 U31195 ( .A1(n46313), .A2(n59967), .ZN(n27653) );
  CLKNAND2HSV0 U31196 ( .A1(n27653), .A2(n27652), .ZN(n27654) );
  OAI21HSV0 U31197 ( .A1(n27652), .A2(n27653), .B(n27654), .ZN(n27655) );
  NAND2HSV0 U31198 ( .A1(n55895), .A2(n56494), .ZN(n27656) );
  CLKNAND2HSV0 U31199 ( .A1(n27656), .A2(n27655), .ZN(n27657) );
  OAI21HSV0 U31200 ( .A1(n27655), .A2(n27656), .B(n27657), .ZN(n27658) );
  NAND2HSV0 U31201 ( .A1(n55706), .A2(n56421), .ZN(n27659) );
  CLKNAND2HSV0 U31202 ( .A1(n27659), .A2(n27658), .ZN(n27660) );
  OAI21HSV0 U31203 ( .A1(n27658), .A2(n27659), .B(n27660), .ZN(n27661) );
  NAND2HSV0 U31204 ( .A1(n56493), .A2(n49255), .ZN(n27662) );
  CLKNAND2HSV0 U31205 ( .A1(n27662), .A2(n27661), .ZN(n27663) );
  OAI21HSV0 U31206 ( .A1(n27661), .A2(n27662), .B(n27663), .ZN(n27664) );
  CLKNAND2HSV0 U31207 ( .A1(n45518), .A2(n55948), .ZN(n27665) );
  CLKNAND2HSV0 U31208 ( .A1(n27665), .A2(n27664), .ZN(n27666) );
  OAI21HSV0 U31209 ( .A1(n27664), .A2(n27665), .B(n27666), .ZN(n45579) );
  XOR2HSV0 U31210 ( .A1(n33824), .A2(n33825), .Z(n27667) );
  XOR2HSV0 U31211 ( .A1(n33823), .A2(n33822), .Z(n27668) );
  XOR2HSV0 U31212 ( .A1(n27667), .A2(n27668), .Z(n27669) );
  XOR2HSV0 U31213 ( .A1(n33828), .A2(n33829), .Z(n27670) );
  XOR2HSV0 U31214 ( .A1(n33827), .A2(n33826), .Z(n27671) );
  XOR2HSV0 U31215 ( .A1(n27670), .A2(n27671), .Z(n27672) );
  XOR2HSV0 U31216 ( .A1(n33820), .A2(n33821), .Z(n27673) );
  CLKXOR2HSV2 U31217 ( .A1(n33815), .A2(n33814), .Z(n27674) );
  XOR2HSV4 U31218 ( .A1(n27673), .A2(n27674), .Z(n27675) );
  NAND2HSV0 U31219 ( .A1(n34042), .A2(n33976), .ZN(n27676) );
  NAND2HSV2 U31220 ( .A1(n27676), .A2(n27675), .ZN(n27677) );
  XOR2HSV0 U31221 ( .A1(n27669), .A2(n27672), .Z(n27679) );
  CLKXOR2HSV4 U31222 ( .A1(n27678), .A2(n27679), .Z(n27680) );
  NAND2HSV0 U31223 ( .A1(n35321), .A2(n57359), .ZN(n27681) );
  NAND2HSV2 U31224 ( .A1(n27681), .A2(n27680), .ZN(n27682) );
  OAI21HSV2 U31225 ( .A1(n27680), .A2(n27681), .B(n27682), .ZN(n27683) );
  NAND2HSV0 U31226 ( .A1(n57285), .A2(n33831), .ZN(n27684) );
  CLKNAND2HSV0 U31227 ( .A1(n27684), .A2(n27683), .ZN(n27685) );
  OAI21HSV0 U31228 ( .A1(n27683), .A2(n27684), .B(n27685), .ZN(n33832) );
  CLKNHSV0 U31229 ( .I(n36205), .ZN(n27686) );
  MUX2NHSV2 U31230 ( .I0(n27686), .I1(n36205), .S(n36204), .ZN(n44362) );
  NAND2HSV0 U31231 ( .A1(n34593), .A2(n47771), .ZN(n27687) );
  CLKNAND2HSV0 U31232 ( .A1(n27687), .A2(n34310), .ZN(n27688) );
  OAI21HSV0 U31233 ( .A1(n34310), .A2(n27687), .B(n27688), .ZN(n27689) );
  NAND2HSV0 U31234 ( .A1(n59350), .A2(n57547), .ZN(n27690) );
  NAND2HSV0 U31235 ( .A1(n27690), .A2(n27689), .ZN(n27691) );
  OAI21HSV0 U31236 ( .A1(n27689), .A2(n27690), .B(n27691), .ZN(n34313) );
  OAI21HSV0 U31237 ( .A1(\pe3/ti_7t [29]), .A2(n45625), .B(n45624), .ZN(n27692) );
  IAO21HSV2 U31238 ( .A1(n45623), .A2(n45622), .B(n27692), .ZN(n46108) );
  IOA21HSV4 U31239 ( .A1(n59509), .A2(n38627), .B(n36501), .ZN(n44906) );
  XOR2HSV0 U31240 ( .A1(n59017), .A2(n59016), .Z(n27693) );
  NAND2HSV0 U31241 ( .A1(n59292), .A2(n59917), .ZN(n27694) );
  CLKNAND2HSV0 U31242 ( .A1(n27694), .A2(n27693), .ZN(n27695) );
  OAI21HSV0 U31243 ( .A1(n27693), .A2(n27694), .B(n27695), .ZN(n27696) );
  CLKNAND2HSV0 U31244 ( .A1(n58723), .A2(n58939), .ZN(n27697) );
  CLKNAND2HSV0 U31245 ( .A1(n27697), .A2(n27696), .ZN(n27698) );
  OAI21HSV0 U31246 ( .A1(n27696), .A2(n27697), .B(n27698), .ZN(n27699) );
  CLKNAND2HSV0 U31247 ( .A1(\pe6/got [7]), .A2(n32165), .ZN(n27700) );
  CLKNAND2HSV0 U31248 ( .A1(n27700), .A2(n27699), .ZN(n27701) );
  OAI21HSV0 U31249 ( .A1(n27699), .A2(n27700), .B(n27701), .ZN(n27702) );
  NAND2HSV0 U31250 ( .A1(n59182), .A2(n59036), .ZN(n27703) );
  CLKNAND2HSV0 U31251 ( .A1(n27703), .A2(n27702), .ZN(n27704) );
  OAI21HSV0 U31252 ( .A1(n27702), .A2(n27703), .B(n27704), .ZN(n27705) );
  CLKNAND2HSV0 U31253 ( .A1(n59037), .A2(n59420), .ZN(n27706) );
  CLKNAND2HSV0 U31254 ( .A1(n27706), .A2(n27705), .ZN(n27707) );
  OAI21HSV0 U31255 ( .A1(n27705), .A2(n27706), .B(n27707), .ZN(n27708) );
  NAND2HSV0 U31256 ( .A1(\pe6/got [10]), .A2(n36105), .ZN(n27709) );
  CLKNAND2HSV0 U31257 ( .A1(n27709), .A2(n27708), .ZN(n27710) );
  OAI21HSV0 U31258 ( .A1(n27708), .A2(n27709), .B(n27710), .ZN(n27711) );
  CLKNAND2HSV0 U31259 ( .A1(n59181), .A2(n58722), .ZN(n27712) );
  CLKNAND2HSV0 U31260 ( .A1(n27712), .A2(n27711), .ZN(n27713) );
  OAI21HSV0 U31261 ( .A1(n27711), .A2(n27712), .B(n27713), .ZN(n27714) );
  CLKNAND2HSV0 U31262 ( .A1(n33039), .A2(n59317), .ZN(n27715) );
  CLKNAND2HSV0 U31263 ( .A1(n27715), .A2(n27714), .ZN(n27716) );
  OAI21HSV0 U31264 ( .A1(n27714), .A2(n27715), .B(n27716), .ZN(n27717) );
  NAND2HSV0 U31265 ( .A1(n58811), .A2(n35775), .ZN(n27718) );
  CLKNAND2HSV0 U31266 ( .A1(n27718), .A2(n27717), .ZN(n27719) );
  OAI21HSV0 U31267 ( .A1(n27717), .A2(n27718), .B(n27719), .ZN(n27720) );
  CLKNAND2HSV0 U31268 ( .A1(n58938), .A2(n49741), .ZN(n27721) );
  CLKNAND2HSV0 U31269 ( .A1(n27721), .A2(n27720), .ZN(n27722) );
  OAI21HSV0 U31270 ( .A1(n27720), .A2(n27721), .B(n27722), .ZN(n27723) );
  NAND2HSV0 U31271 ( .A1(\pe6/got [15]), .A2(n59916), .ZN(n27724) );
  CLKNAND2HSV0 U31272 ( .A1(n27724), .A2(n27723), .ZN(n27725) );
  OAI21HSV0 U31273 ( .A1(n27723), .A2(n27724), .B(n27725), .ZN(n27726) );
  NAND2HSV0 U31274 ( .A1(n59177), .A2(n58937), .ZN(n27727) );
  CLKNAND2HSV0 U31275 ( .A1(n27727), .A2(n27726), .ZN(n27728) );
  OAI21HSV0 U31276 ( .A1(n27726), .A2(n27727), .B(n27728), .ZN(n27729) );
  NAND2HSV0 U31277 ( .A1(n49098), .A2(n49726), .ZN(n27730) );
  CLKNAND2HSV0 U31278 ( .A1(n27730), .A2(n27729), .ZN(n27731) );
  OAI21HSV0 U31279 ( .A1(n27729), .A2(n27730), .B(n27731), .ZN(n27732) );
  CLKNAND2HSV0 U31280 ( .A1(\pe6/got [18]), .A2(n58936), .ZN(n27733) );
  CLKNAND2HSV0 U31281 ( .A1(n27733), .A2(n27732), .ZN(n27734) );
  OAI21HSV0 U31282 ( .A1(n27732), .A2(n27733), .B(n27734), .ZN(n59018) );
  XOR2HSV0 U31283 ( .A1(n58125), .A2(n58121), .Z(n27735) );
  XOR2HSV0 U31284 ( .A1(n58119), .A2(n58122), .Z(n27736) );
  XOR2HSV0 U31285 ( .A1(n27735), .A2(n27736), .Z(n27737) );
  CLKNHSV0 U31286 ( .I(n58136), .ZN(n27738) );
  XOR2HSV0 U31287 ( .A1(n58134), .A2(n58133), .Z(n27739) );
  XOR2HSV0 U31288 ( .A1(n58135), .A2(n27739), .Z(n27740) );
  MUX2NHSV0 U31289 ( .I0(n58136), .I1(n27738), .S(n27740), .ZN(n27741) );
  XOR2HSV0 U31290 ( .A1(n58120), .A2(n27737), .Z(n27742) );
  XOR2HSV0 U31291 ( .A1(n27741), .A2(n27742), .Z(n27743) );
  NAND2HSV0 U31292 ( .A1(n58096), .A2(\pe4/got [2]), .ZN(n27744) );
  CLKNAND2HSV0 U31293 ( .A1(n27744), .A2(n27743), .ZN(n27745) );
  OAI21HSV0 U31294 ( .A1(n27743), .A2(n27744), .B(n27745), .ZN(n27746) );
  NAND2HSV0 U31295 ( .A1(n59935), .A2(n58300), .ZN(n27747) );
  CLKNAND2HSV0 U31296 ( .A1(n27747), .A2(n27746), .ZN(n27748) );
  OAI21HSV0 U31297 ( .A1(n27746), .A2(n27747), .B(n27748), .ZN(n27749) );
  NAND2HSV0 U31298 ( .A1(n58112), .A2(n58298), .ZN(n27750) );
  CLKNAND2HSV0 U31299 ( .A1(n27750), .A2(n27749), .ZN(n27751) );
  OAI21HSV0 U31300 ( .A1(n27749), .A2(n27750), .B(n27751), .ZN(n27752) );
  NAND2HSV0 U31301 ( .A1(n58246), .A2(n47841), .ZN(n27753) );
  CLKNAND2HSV0 U31302 ( .A1(n27753), .A2(n27752), .ZN(n27754) );
  OAI21HSV2 U31303 ( .A1(n27752), .A2(n27753), .B(n27754), .ZN(n27755) );
  NAND2HSV0 U31304 ( .A1(n58030), .A2(n59672), .ZN(n27756) );
  NAND2HSV2 U31305 ( .A1(n27756), .A2(n27755), .ZN(n27757) );
  OAI21HSV2 U31306 ( .A1(n27755), .A2(n27756), .B(n27757), .ZN(n27758) );
  NAND2HSV0 U31307 ( .A1(n58220), .A2(n58137), .ZN(n27759) );
  NAND2HSV2 U31308 ( .A1(n27759), .A2(n27758), .ZN(n27760) );
  OAI21HSV2 U31309 ( .A1(n27758), .A2(n27759), .B(n27760), .ZN(n27761) );
  NAND2HSV0 U31310 ( .A1(n58185), .A2(n58216), .ZN(n27762) );
  NAND2HSV2 U31311 ( .A1(n27762), .A2(n27761), .ZN(n27763) );
  OAI21HSV2 U31312 ( .A1(n27761), .A2(n27762), .B(n27763), .ZN(n58138) );
  AND2HSV2 U31313 ( .A1(n44662), .A2(n44663), .Z(n45924) );
  OAI21HSV0 U31314 ( .A1(n52710), .A2(n33085), .B(poh6[22]), .ZN(n27764) );
  OAI31HSV0 U31315 ( .A1(n52710), .A2(poh6[22]), .A3(n33085), .B(n27764), .ZN(
        po[23]) );
  AO21HSV1 U31316 ( .A1(n60037), .A2(n39417), .B(n29991), .Z(n30255) );
  NAND2HSV0 U31317 ( .A1(n51893), .A2(n52125), .ZN(n27765) );
  CLKNAND2HSV0 U31318 ( .A1(n27765), .A2(n51725), .ZN(n27766) );
  OAI21HSV0 U31319 ( .A1(n51725), .A2(n27765), .B(n27766), .ZN(n27767) );
  XOR2HSV0 U31320 ( .A1(n51724), .A2(n27767), .Z(n27768) );
  NAND2HSV0 U31321 ( .A1(n52052), .A2(n51797), .ZN(n27769) );
  CLKNAND2HSV0 U31322 ( .A1(n27769), .A2(n27768), .ZN(n27770) );
  OAI21HSV0 U31323 ( .A1(n27768), .A2(n27769), .B(n27770), .ZN(n27771) );
  NAND2HSV0 U31324 ( .A1(n25831), .A2(\pe2/got [10]), .ZN(n27772) );
  CLKNAND2HSV0 U31325 ( .A1(n27772), .A2(n27771), .ZN(n27773) );
  OAI21HSV0 U31326 ( .A1(n27771), .A2(n27772), .B(n27773), .ZN(n27774) );
  NAND2HSV0 U31327 ( .A1(n51892), .A2(n52414), .ZN(n27775) );
  CLKNAND2HSV0 U31328 ( .A1(n27775), .A2(n27774), .ZN(n27776) );
  NAND2HSV0 U31329 ( .A1(n52418), .A2(n51961), .ZN(n27781) );
  XOR2HSV0 U31330 ( .A1(n59337), .A2(n59336), .Z(n27783) );
  NAND2HSV0 U31331 ( .A1(n58717), .A2(n59173), .ZN(n27784) );
  CLKNAND2HSV0 U31332 ( .A1(n27784), .A2(n27783), .ZN(n27785) );
  OAI21HSV0 U31333 ( .A1(n27783), .A2(n27784), .B(n27785), .ZN(n27786) );
  NAND2HSV0 U31334 ( .A1(n58716), .A2(\pe6/got [26]), .ZN(n27787) );
  CLKNAND2HSV0 U31335 ( .A1(n27787), .A2(n27786), .ZN(n27788) );
  OAI21HSV0 U31336 ( .A1(n27786), .A2(n27787), .B(n27788), .ZN(n27789) );
  NAND2HSV0 U31337 ( .A1(n59528), .A2(n49665), .ZN(n27790) );
  CLKNAND2HSV0 U31338 ( .A1(n27790), .A2(n27789), .ZN(n27791) );
  OAI21HSV0 U31339 ( .A1(n27789), .A2(n27790), .B(n27791), .ZN(n27792) );
  CLKNAND2HSV0 U31340 ( .A1(n59172), .A2(n59171), .ZN(n27793) );
  CLKNAND2HSV0 U31341 ( .A1(n27793), .A2(n27792), .ZN(n27794) );
  OAI21HSV0 U31342 ( .A1(n27792), .A2(n27793), .B(n27794), .ZN(n27795) );
  NAND2HSV0 U31343 ( .A1(n59170), .A2(n35705), .ZN(n27796) );
  CLKNAND2HSV0 U31344 ( .A1(n27796), .A2(n27795), .ZN(n27797) );
  OAI21HSV0 U31345 ( .A1(n27795), .A2(n27796), .B(n27797), .ZN(n27798) );
  NAND2HSV0 U31346 ( .A1(n32967), .A2(n59169), .ZN(n27799) );
  CLKNAND2HSV0 U31347 ( .A1(n27799), .A2(n27798), .ZN(n27800) );
  OAI21HSV0 U31348 ( .A1(n27798), .A2(n27799), .B(n27800), .ZN(n27801) );
  NAND2HSV0 U31349 ( .A1(n48888), .A2(n59339), .ZN(n27802) );
  CLKNAND2HSV0 U31350 ( .A1(n27802), .A2(n27801), .ZN(n27803) );
  OAI21HSV0 U31351 ( .A1(n27801), .A2(n27802), .B(n27803), .ZN(n27804) );
  NAND2HSV0 U31352 ( .A1(n32783), .A2(n59340), .ZN(n27805) );
  CLKNAND2HSV0 U31353 ( .A1(n27805), .A2(n27804), .ZN(n27806) );
  OAI21HSV0 U31354 ( .A1(n27804), .A2(n27805), .B(n27806), .ZN(po6) );
  NAND2HSV0 U31355 ( .A1(n59892), .A2(n48741), .ZN(n27807) );
  NAND2HSV0 U31356 ( .A1(n47927), .A2(n51404), .ZN(n27809) );
  NAND2HSV0 U31357 ( .A1(n27809), .A2(n27808), .ZN(n27810) );
  OAI21HSV0 U31358 ( .A1(n27808), .A2(n27809), .B(n27810), .ZN(pov5[27]) );
  CLKNHSV0 U31359 ( .I(n34248), .ZN(n27811) );
  NAND2HSV0 U31360 ( .A1(n35491), .A2(n57846), .ZN(n27812) );
  NAND2HSV0 U31361 ( .A1(n27812), .A2(n34633), .ZN(n27813) );
  OAI21HSV0 U31362 ( .A1(n34633), .A2(n27812), .B(n27813), .ZN(n27814) );
  NAND2HSV0 U31363 ( .A1(n47658), .A2(n34359), .ZN(n27815) );
  NAND2HSV0 U31364 ( .A1(n27815), .A2(n27814), .ZN(n27816) );
  OAI21HSV0 U31365 ( .A1(n27814), .A2(n27815), .B(n27816), .ZN(n27817) );
  MUX2NHSV0 U31366 ( .I0(n27811), .I1(n34248), .S(n27817), .ZN(n34250) );
  CLKNHSV0 U31367 ( .I(n52938), .ZN(n27818) );
  NAND2HSV0 U31368 ( .A1(\pe2/pvq [14]), .A2(n53014), .ZN(n27819) );
  NAND2HSV0 U31369 ( .A1(n27819), .A2(\pe2/phq [14]), .ZN(n27820) );
  OAI21HSV2 U31370 ( .A1(\pe2/phq [14]), .A2(n27819), .B(n27820), .ZN(n27821)
         );
  MUX2NHSV1 U31371 ( .I0(n52938), .I1(n27818), .S(n27821), .ZN(n37961) );
  CLKNAND2HSV0 U31372 ( .A1(n38542), .A2(n59970), .ZN(n27822) );
  OAI21HSV0 U31373 ( .A1(n38973), .A2(n38213), .B(n27822), .ZN(n27823) );
  OAI31HSV0 U31374 ( .A1(n38973), .A2(n27822), .A3(n38213), .B(n27823), .ZN(
        n38130) );
  NAND2HSV0 U31375 ( .A1(n27824), .A2(\pe4/phq [3]), .ZN(n27825) );
  OAI21HSV2 U31376 ( .A1(\pe4/phq [3]), .A2(n27824), .B(n27825), .ZN(n33101)
         );
  NAND2HSV0 U31377 ( .A1(n42373), .A2(n44566), .ZN(n27826) );
  NAND2HSV0 U31378 ( .A1(n41877), .A2(n41645), .ZN(n27827) );
  CLKNAND2HSV0 U31379 ( .A1(n27827), .A2(n27826), .ZN(n27828) );
  OAI21HSV0 U31380 ( .A1(n27826), .A2(n27827), .B(n27828), .ZN(n27829) );
  NAND2HSV0 U31381 ( .A1(n42155), .A2(n41522), .ZN(n27830) );
  NAND2HSV0 U31382 ( .A1(n27830), .A2(n27829), .ZN(n27831) );
  OAI21HSV0 U31383 ( .A1(n27829), .A2(n27830), .B(n27831), .ZN(n41523) );
  NAND2HSV0 U31384 ( .A1(n40683), .A2(n53411), .ZN(n27832) );
  CLKNAND2HSV0 U31385 ( .A1(n27832), .A2(n41270), .ZN(n27833) );
  OAI21HSV0 U31386 ( .A1(n41270), .A2(n27832), .B(n27833), .ZN(n27834) );
  OAI21HSV0 U31387 ( .A1(n26269), .A2(n44528), .B(n27834), .ZN(n27835) );
  NAND2HSV0 U31388 ( .A1(n44392), .A2(n46171), .ZN(n27836) );
  CLKNAND2HSV0 U31389 ( .A1(n27836), .A2(n35897), .ZN(n27837) );
  OAI21HSV0 U31390 ( .A1(n35897), .A2(n27836), .B(n27837), .ZN(n27838) );
  NAND2HSV0 U31391 ( .A1(n36105), .A2(n49098), .ZN(n27839) );
  CLKNAND2HSV0 U31392 ( .A1(n27839), .A2(n27838), .ZN(n27840) );
  OAI21HSV0 U31393 ( .A1(n27838), .A2(n27839), .B(n27840), .ZN(n27841) );
  NAND2HSV0 U31394 ( .A1(n58722), .A2(n36104), .ZN(n27842) );
  CLKNAND2HSV0 U31395 ( .A1(n27842), .A2(n27841), .ZN(n27843) );
  OAI21HSV0 U31396 ( .A1(n27841), .A2(n27842), .B(n27843), .ZN(n27844) );
  NAND2HSV0 U31397 ( .A1(n59144), .A2(n35922), .ZN(n27845) );
  CLKNAND2HSV0 U31398 ( .A1(n27845), .A2(n27844), .ZN(n27846) );
  OAI21HSV0 U31399 ( .A1(n27844), .A2(n27845), .B(n27846), .ZN(n27847) );
  NAND2HSV0 U31400 ( .A1(n59676), .A2(n59176), .ZN(n27848) );
  CLKNAND2HSV0 U31401 ( .A1(n27848), .A2(n27847), .ZN(n27849) );
  OAI21HSV0 U31402 ( .A1(n27847), .A2(n27848), .B(n27849), .ZN(n27850) );
  NAND2HSV0 U31403 ( .A1(n58664), .A2(\pe6/got [21]), .ZN(n27851) );
  CLKNAND2HSV0 U31404 ( .A1(n27851), .A2(n27850), .ZN(n27852) );
  OAI21HSV0 U31405 ( .A1(n27850), .A2(n27851), .B(n27852), .ZN(n27853) );
  NAND2HSV0 U31406 ( .A1(n58663), .A2(n58714), .ZN(n27854) );
  CLKNAND2HSV0 U31407 ( .A1(n27854), .A2(n27853), .ZN(n27855) );
  OAI21HSV0 U31408 ( .A1(n27853), .A2(n27854), .B(n27855), .ZN(n27856) );
  CLKNAND2HSV0 U31409 ( .A1(n35812), .A2(n44390), .ZN(n27857) );
  CLKNAND2HSV0 U31410 ( .A1(n27857), .A2(n27856), .ZN(n27858) );
  OAI21HSV0 U31411 ( .A1(n27856), .A2(n27857), .B(n27858), .ZN(n27859) );
  NAND2HSV0 U31412 ( .A1(\pe6/got [24]), .A2(n36196), .ZN(n27860) );
  CLKNAND2HSV0 U31413 ( .A1(n27860), .A2(n27859), .ZN(n27861) );
  OAI21HSV0 U31414 ( .A1(n27859), .A2(n27860), .B(n27861), .ZN(n35899) );
  AOI21HSV0 U31415 ( .A1(n44027), .A2(n38886), .B(n44831), .ZN(n27862) );
  OAI21HSV4 U31416 ( .A1(n60095), .A2(n37931), .B(n27862), .ZN(n39003) );
  XOR2HSV0 U31417 ( .A1(n50120), .A2(n50121), .Z(n27863) );
  XOR2HSV0 U31418 ( .A1(n50119), .A2(n50118), .Z(n27864) );
  XOR2HSV0 U31419 ( .A1(n27863), .A2(n27864), .Z(n27865) );
  XOR2HSV0 U31420 ( .A1(n27865), .A2(n50117), .Z(n27866) );
  XOR2HSV0 U31421 ( .A1(n50113), .A2(n50112), .Z(n27867) );
  XOR2HSV0 U31422 ( .A1(n27866), .A2(n27867), .Z(n27868) );
  NAND2HSV0 U31423 ( .A1(n58300), .A2(n59950), .ZN(n27869) );
  CLKNAND2HSV0 U31424 ( .A1(n27869), .A2(n27868), .ZN(n27870) );
  OAI21HSV0 U31425 ( .A1(n27868), .A2(n27869), .B(n27870), .ZN(n27871) );
  NAND2HSV0 U31426 ( .A1(n58193), .A2(n58314), .ZN(n27872) );
  CLKNAND2HSV0 U31427 ( .A1(n27872), .A2(n27871), .ZN(n27873) );
  OAI21HSV0 U31428 ( .A1(n27871), .A2(n27872), .B(n27873), .ZN(n27874) );
  NAND2HSV0 U31429 ( .A1(n58104), .A2(n58298), .ZN(n27875) );
  CLKNAND2HSV0 U31430 ( .A1(n27875), .A2(n27874), .ZN(n27876) );
  OAI21HSV0 U31431 ( .A1(n27874), .A2(n27875), .B(n27876), .ZN(n27877) );
  NAND2HSV0 U31432 ( .A1(n58272), .A2(n58258), .ZN(n27878) );
  CLKNAND2HSV0 U31433 ( .A1(n27878), .A2(n27877), .ZN(n27879) );
  OAI21HSV0 U31434 ( .A1(n27877), .A2(n27878), .B(n27879), .ZN(n27880) );
  NAND2HSV0 U31435 ( .A1(n58246), .A2(n58207), .ZN(n27881) );
  NAND2HSV0 U31436 ( .A1(n27881), .A2(n27880), .ZN(n27882) );
  OAI21HSV2 U31437 ( .A1(n27880), .A2(n27881), .B(n27882), .ZN(n50122) );
  XOR2HSV0 U31438 ( .A1(n56474), .A2(n56473), .Z(n27883) );
  XOR2HSV0 U31439 ( .A1(n56476), .A2(n27883), .Z(n27884) );
  NAND2HSV0 U31440 ( .A1(n59810), .A2(n59356), .ZN(n27885) );
  CLKNAND2HSV0 U31441 ( .A1(n27885), .A2(n27884), .ZN(n27886) );
  OAI21HSV0 U31442 ( .A1(n27884), .A2(n27885), .B(n27886), .ZN(n27887) );
  NAND2HSV0 U31443 ( .A1(n55824), .A2(n56734), .ZN(n27888) );
  CLKNAND2HSV0 U31444 ( .A1(n27888), .A2(n27887), .ZN(n27889) );
  OAI21HSV0 U31445 ( .A1(n27887), .A2(n27888), .B(n27889), .ZN(n27890) );
  NAND2HSV0 U31446 ( .A1(n59811), .A2(n56781), .ZN(n27891) );
  CLKNAND2HSV0 U31447 ( .A1(n27891), .A2(n27890), .ZN(n27892) );
  OAI21HSV0 U31448 ( .A1(n27890), .A2(n27891), .B(n27892), .ZN(n27893) );
  NAND2HSV0 U31449 ( .A1(n56624), .A2(n56560), .ZN(n27894) );
  CLKNAND2HSV0 U31450 ( .A1(n27894), .A2(n27893), .ZN(n27895) );
  OAI21HSV0 U31451 ( .A1(n27893), .A2(n27894), .B(n27895), .ZN(n27896) );
  NAND2HSV0 U31452 ( .A1(n56888), .A2(n43463), .ZN(n27897) );
  CLKNAND2HSV0 U31453 ( .A1(n27897), .A2(n27896), .ZN(n27898) );
  OAI21HSV0 U31454 ( .A1(n27896), .A2(n27897), .B(n27898), .ZN(n27899) );
  NAND2HSV0 U31455 ( .A1(n56685), .A2(\pe3/got [8]), .ZN(n27900) );
  CLKNAND2HSV0 U31456 ( .A1(n27900), .A2(n27899), .ZN(n27901) );
  OAI21HSV0 U31457 ( .A1(n27899), .A2(n27900), .B(n27901), .ZN(n27902) );
  NAND2HSV0 U31458 ( .A1(n56559), .A2(n56737), .ZN(n27903) );
  CLKNAND2HSV0 U31459 ( .A1(n27903), .A2(n27902), .ZN(n27904) );
  OAI21HSV0 U31460 ( .A1(n27902), .A2(n27903), .B(n27904), .ZN(n27905) );
  NAND2HSV0 U31461 ( .A1(n56561), .A2(n56495), .ZN(n27906) );
  CLKNAND2HSV0 U31462 ( .A1(n27906), .A2(n27905), .ZN(n27907) );
  OAI21HSV2 U31463 ( .A1(n27905), .A2(n27906), .B(n27907), .ZN(n27908) );
  NAND2HSV0 U31464 ( .A1(n56736), .A2(n56557), .ZN(n27909) );
  NAND2HSV2 U31465 ( .A1(n27909), .A2(n27908), .ZN(n27910) );
  OAI21HSV2 U31466 ( .A1(n27908), .A2(n27909), .B(n27910), .ZN(n56477) );
  CLKNAND2HSV0 U31467 ( .A1(n57209), .A2(n57888), .ZN(n27911) );
  CLKNAND2HSV0 U31468 ( .A1(n27911), .A2(n57187), .ZN(n27912) );
  OAI21HSV0 U31469 ( .A1(n57187), .A2(n27911), .B(n27912), .ZN(n27913) );
  NAND2HSV0 U31470 ( .A1(n57820), .A2(n57324), .ZN(n27914) );
  CLKNAND2HSV0 U31471 ( .A1(n27914), .A2(n27913), .ZN(n27915) );
  OAI21HSV0 U31472 ( .A1(n27913), .A2(n27914), .B(n27915), .ZN(n27916) );
  NAND2HSV0 U31473 ( .A1(n57424), .A2(n57188), .ZN(n27917) );
  CLKNAND2HSV0 U31474 ( .A1(n27917), .A2(n27916), .ZN(n27918) );
  OAI21HSV0 U31475 ( .A1(n27916), .A2(n27917), .B(n27918), .ZN(n27919) );
  NAND2HSV0 U31476 ( .A1(n57675), .A2(n57307), .ZN(n27920) );
  CLKNAND2HSV0 U31477 ( .A1(n27920), .A2(n27919), .ZN(n27921) );
  OAI21HSV0 U31478 ( .A1(n27919), .A2(n27920), .B(n27921), .ZN(n27922) );
  NAND2HSV0 U31479 ( .A1(n57189), .A2(n25284), .ZN(n27923) );
  CLKNAND2HSV0 U31480 ( .A1(n27923), .A2(n27922), .ZN(n27924) );
  OAI21HSV0 U31481 ( .A1(n27922), .A2(n27923), .B(n27924), .ZN(n27925) );
  CLKNAND2HSV0 U31482 ( .A1(n57457), .A2(n34409), .ZN(n27926) );
  CLKNAND2HSV0 U31483 ( .A1(n27926), .A2(n27925), .ZN(n27927) );
  OAI21HSV0 U31484 ( .A1(n27925), .A2(n27926), .B(n27927), .ZN(n27928) );
  CLKNAND2HSV0 U31485 ( .A1(n57427), .A2(n57834), .ZN(n27929) );
  CLKNAND2HSV0 U31486 ( .A1(n27929), .A2(n27928), .ZN(n27930) );
  OAI21HSV0 U31487 ( .A1(n27928), .A2(n27929), .B(n27930), .ZN(n27931) );
  NAND2HSV0 U31488 ( .A1(n57564), .A2(n58029), .ZN(n27932) );
  CLKNAND2HSV0 U31489 ( .A1(n27932), .A2(n27931), .ZN(n27933) );
  OAI21HSV0 U31490 ( .A1(n27931), .A2(n27932), .B(n27933), .ZN(n27934) );
  CLKNAND2HSV0 U31491 ( .A1(n57554), .A2(n50404), .ZN(n27935) );
  CLKNAND2HSV0 U31492 ( .A1(n27935), .A2(n27934), .ZN(n27936) );
  OAI21HSV0 U31493 ( .A1(n27934), .A2(n27935), .B(n27936), .ZN(n27937) );
  CLKNAND2HSV0 U31494 ( .A1(n58112), .A2(n57760), .ZN(n27938) );
  CLKNAND2HSV0 U31495 ( .A1(n27938), .A2(n27937), .ZN(n27939) );
  OAI21HSV0 U31496 ( .A1(n27937), .A2(n27938), .B(n27939), .ZN(n27940) );
  CLKNAND2HSV0 U31497 ( .A1(n57819), .A2(\pe4/got [23]), .ZN(n27941) );
  CLKNAND2HSV0 U31498 ( .A1(n27941), .A2(n27940), .ZN(n27942) );
  OAI21HSV2 U31499 ( .A1(n27940), .A2(n27941), .B(n27942), .ZN(n27943) );
  NAND2HSV0 U31500 ( .A1(n59601), .A2(n57560), .ZN(n27944) );
  CLKNAND2HSV0 U31501 ( .A1(n27944), .A2(n27943), .ZN(n27945) );
  OAI21HSV2 U31502 ( .A1(n27943), .A2(n27944), .B(n27945), .ZN(n27946) );
  NAND2HSV0 U31503 ( .A1(n59603), .A2(n25427), .ZN(n27947) );
  CLKNAND2HSV0 U31504 ( .A1(n27947), .A2(n27946), .ZN(n27948) );
  OAI21HSV2 U31505 ( .A1(n27946), .A2(n27947), .B(n27948), .ZN(n57192) );
  NOR4HSV2 U31506 ( .A1(n37991), .A2(n38005), .A3(n38006), .A4(n37865), .ZN(
        n27949) );
  IOA21HSV4 U31507 ( .A1(n37985), .A2(n27949), .B(n38106), .ZN(n59583) );
  CLKNAND2HSV0 U31508 ( .A1(n51798), .A2(n59984), .ZN(n27950) );
  CLKNAND2HSV0 U31509 ( .A1(n27950), .A2(n51562), .ZN(n27951) );
  OAI21HSV0 U31510 ( .A1(n51562), .A2(n27950), .B(n27951), .ZN(n27952) );
  XOR2HSV0 U31511 ( .A1(n51561), .A2(n27952), .Z(n27953) );
  NAND2HSV0 U31512 ( .A1(n51797), .A2(n51939), .ZN(n27954) );
  CLKNAND2HSV0 U31513 ( .A1(n27954), .A2(n27953), .ZN(n27955) );
  OAI21HSV0 U31514 ( .A1(n27953), .A2(n27954), .B(n27955), .ZN(n27956) );
  CLKNAND2HSV0 U31515 ( .A1(n59475), .A2(n52890), .ZN(n27957) );
  CLKNAND2HSV0 U31516 ( .A1(n27957), .A2(n27956), .ZN(n27958) );
  OAI21HSV0 U31517 ( .A1(n27956), .A2(n27957), .B(n27958), .ZN(n27959) );
  NAND2HSV0 U31518 ( .A1(n52414), .A2(\pe2/got [8]), .ZN(n27960) );
  CLKNAND2HSV0 U31519 ( .A1(n27960), .A2(n27959), .ZN(n27961) );
  OAI21HSV0 U31520 ( .A1(n27959), .A2(n27960), .B(n27961), .ZN(n27962) );
  OAI21HSV2 U31521 ( .A1(n27962), .A2(n27963), .B(n27964), .ZN(n27965) );
  NAND2HSV0 U31522 ( .A1(n59794), .A2(\pe2/got [10]), .ZN(n27966) );
  CLKNAND2HSV0 U31523 ( .A1(n27966), .A2(n27965), .ZN(n27967) );
  OAI21HSV0 U31524 ( .A1(n27965), .A2(n27966), .B(n27967), .ZN(\pe2/poht [22])
         );
  XOR2HSV0 U31525 ( .A1(n58653), .A2(n58652), .Z(n27968) );
  NAND2HSV0 U31526 ( .A1(n58611), .A2(n58709), .ZN(n27969) );
  CLKNAND2HSV0 U31527 ( .A1(n27969), .A2(n27968), .ZN(n27970) );
  OAI21HSV0 U31528 ( .A1(n27968), .A2(n27969), .B(n27970), .ZN(n27971) );
  CLKNAND2HSV0 U31529 ( .A1(n53109), .A2(\pe6/got [8]), .ZN(n27972) );
  CLKNAND2HSV0 U31530 ( .A1(n27972), .A2(n27971), .ZN(n27973) );
  OAI21HSV0 U31531 ( .A1(n27971), .A2(n27972), .B(n27973), .ZN(n27974) );
  NAND2HSV0 U31532 ( .A1(n59528), .A2(n58658), .ZN(n27975) );
  CLKNAND2HSV0 U31533 ( .A1(n27975), .A2(n27974), .ZN(n27976) );
  OAI21HSV0 U31534 ( .A1(n27974), .A2(n27975), .B(n27976), .ZN(n27977) );
  NAND2HSV0 U31535 ( .A1(n58657), .A2(n58812), .ZN(n27978) );
  CLKNAND2HSV0 U31536 ( .A1(n27978), .A2(n27977), .ZN(n27979) );
  OAI21HSV0 U31537 ( .A1(n27977), .A2(n27978), .B(n27979), .ZN(n27980) );
  CLKNAND2HSV0 U31538 ( .A1(n58656), .A2(n49742), .ZN(n27981) );
  CLKNAND2HSV0 U31539 ( .A1(n27981), .A2(n27980), .ZN(n27982) );
  OAI21HSV0 U31540 ( .A1(n27980), .A2(n27981), .B(n27982), .ZN(n27983) );
  CLKNAND2HSV0 U31541 ( .A1(n33039), .A2(n59024), .ZN(n27984) );
  CLKNAND2HSV0 U31542 ( .A1(n27984), .A2(n27983), .ZN(n27985) );
  OAI21HSV0 U31543 ( .A1(n27983), .A2(n27984), .B(n27985), .ZN(n27986) );
  NAND2HSV0 U31544 ( .A1(n48888), .A2(n58654), .ZN(n27987) );
  CLKNAND2HSV0 U31545 ( .A1(n27987), .A2(n27986), .ZN(n27988) );
  OAI21HSV0 U31546 ( .A1(n27986), .A2(n27987), .B(n27988), .ZN(n27989) );
  CLKNAND2HSV0 U31547 ( .A1(n27989), .A2(n27990), .ZN(n27991) );
  OAI21HSV0 U31548 ( .A1(n27989), .A2(n27990), .B(n27991), .ZN(\pe6/poht [18])
         );
  XOR2HSV0 U31549 ( .A1(n48884), .A2(n48883), .Z(n27992) );
  NAND2HSV0 U31550 ( .A1(n52670), .A2(n48742), .ZN(n27993) );
  CLKNAND2HSV0 U31551 ( .A1(n27993), .A2(n27992), .ZN(n27994) );
  OAI21HSV0 U31552 ( .A1(n27992), .A2(n27993), .B(n27994), .ZN(n27995) );
  NAND2HSV0 U31553 ( .A1(n52693), .A2(\pe5/got [27]), .ZN(n27996) );
  CLKNAND2HSV0 U31554 ( .A1(n27996), .A2(n27995), .ZN(n27997) );
  OAI21HSV0 U31555 ( .A1(n27995), .A2(n27996), .B(n27997), .ZN(n27998) );
  NAND2HSV0 U31556 ( .A1(n51272), .A2(n30779), .ZN(n27999) );
  CLKNAND2HSV0 U31557 ( .A1(n27999), .A2(n27998), .ZN(n28000) );
  OAI21HSV0 U31558 ( .A1(n27998), .A2(n27999), .B(n28000), .ZN(n28001) );
  NAND2HSV0 U31559 ( .A1(n59933), .A2(n30142), .ZN(n28002) );
  CLKNAND2HSV0 U31560 ( .A1(n28002), .A2(n28001), .ZN(n28003) );
  OAI21HSV0 U31561 ( .A1(n28001), .A2(n28002), .B(n28003), .ZN(n28004) );
  NAND2HSV0 U31562 ( .A1(n48885), .A2(n51411), .ZN(n28005) );
  CLKNAND2HSV0 U31563 ( .A1(n28005), .A2(n28004), .ZN(n28006) );
  OAI21HSV0 U31564 ( .A1(n28004), .A2(n28005), .B(n28006), .ZN(n28007) );
  CLKNAND2HSV0 U31565 ( .A1(n48741), .A2(n59580), .ZN(n28008) );
  CLKNAND2HSV0 U31566 ( .A1(n28008), .A2(n28007), .ZN(n28009) );
  OAI21HSV0 U31567 ( .A1(n28007), .A2(n28008), .B(n28009), .ZN(n28010) );
  CLKNAND2HSV0 U31568 ( .A1(n48886), .A2(n52767), .ZN(n28011) );
  CLKNAND2HSV0 U31569 ( .A1(n28011), .A2(n28010), .ZN(n28012) );
  OAI21HSV0 U31570 ( .A1(n28010), .A2(n28011), .B(n28012), .ZN(po5) );
  NAND2HSV0 U31571 ( .A1(n34879), .A2(n59388), .ZN(n28013) );
  OAI21HSV0 U31572 ( .A1(n34470), .A2(n48070), .B(n28013), .ZN(n28014) );
  OAI31HSV0 U31573 ( .A1(n34470), .A2(n28013), .A3(n48070), .B(n28014), .ZN(
        n34474) );
  NAND2HSV0 U31574 ( .A1(\pe6/bq[14] ), .A2(n32740), .ZN(n28015) );
  CLKNAND2HSV0 U31575 ( .A1(n28015), .A2(n32471), .ZN(n28016) );
  OAI21HSV0 U31576 ( .A1(n32471), .A2(n28015), .B(n28016), .ZN(n28017) );
  XOR2HSV0 U31577 ( .A1(n32475), .A2(n32476), .Z(n28018) );
  XOR2HSV0 U31578 ( .A1(n32474), .A2(n32473), .Z(n28019) );
  XOR2HSV0 U31579 ( .A1(n28018), .A2(n28019), .Z(n28020) );
  XOR2HSV0 U31580 ( .A1(n28020), .A2(n28017), .Z(n28021) );
  XOR2HSV0 U31581 ( .A1(n32470), .A2(n32472), .Z(n28022) );
  XOR2HSV0 U31582 ( .A1(n28021), .A2(n28022), .Z(n28023) );
  XOR2HSV0 U31583 ( .A1(n32479), .A2(n32480), .Z(n28024) );
  XOR2HSV0 U31584 ( .A1(n32478), .A2(n32477), .Z(n28025) );
  XOR2HSV0 U31585 ( .A1(n28024), .A2(n28025), .Z(n28026) );
  XOR2HSV0 U31586 ( .A1(\pe6/phq [19]), .A2(n32483), .Z(n28027) );
  XOR2HSV0 U31587 ( .A1(n32482), .A2(n32481), .Z(n28028) );
  XOR2HSV0 U31588 ( .A1(n28027), .A2(n28028), .Z(n28029) );
  CLKNHSV0 U31589 ( .I(n32490), .ZN(n28030) );
  OAI21HSV0 U31590 ( .A1(n32604), .A2(n32489), .B(n32488), .ZN(n28031) );
  CLKNAND2HSV0 U31591 ( .A1(n28031), .A2(n46636), .ZN(n28032) );
  OAI21HSV0 U31592 ( .A1(n28031), .A2(n46636), .B(n28032), .ZN(n28033) );
  OAI21HSV0 U31593 ( .A1(n32591), .A2(n35839), .B(n32485), .ZN(n28034) );
  CLKNAND2HSV0 U31594 ( .A1(n28034), .A2(n28033), .ZN(n28035) );
  OAI21HSV0 U31595 ( .A1(n28034), .A2(n28033), .B(n28035), .ZN(n28036) );
  MUX2NHSV0 U31596 ( .I0(n28030), .I1(n32490), .S(n28036), .ZN(n28037) );
  XOR2HSV0 U31597 ( .A1(n28037), .A2(n28029), .Z(n28038) );
  XOR2HSV0 U31598 ( .A1(n28023), .A2(n28026), .Z(n28039) );
  XOR2HSV0 U31599 ( .A1(n28038), .A2(n28039), .Z(n28040) );
  NAND2HSV0 U31600 ( .A1(n32596), .A2(n35612), .ZN(n28041) );
  NAND2HSV2 U31601 ( .A1(n28041), .A2(n28040), .ZN(n28042) );
  OAI21HSV2 U31602 ( .A1(n28040), .A2(n28041), .B(n28042), .ZN(n28043) );
  NAND2HSV0 U31603 ( .A1(n36106), .A2(n32286), .ZN(n28044) );
  NAND2HSV2 U31604 ( .A1(n28044), .A2(n28043), .ZN(n28045) );
  OAI21HSV2 U31605 ( .A1(n28043), .A2(n28044), .B(n28045), .ZN(n32492) );
  CLKNHSV0 U31606 ( .I(n33813), .ZN(n28046) );
  OAI22HSV0 U31607 ( .A1(n57509), .A2(n50248), .B1(n33250), .B2(n50129), .ZN(
        n28047) );
  OAI21HSV2 U31608 ( .A1(n33812), .A2(n33948), .B(n28047), .ZN(n28048) );
  MUX2NHSV1 U31609 ( .I0(n28046), .I1(n33813), .S(n28048), .ZN(n33814) );
  CLKNHSV0 U31610 ( .I(n49528), .ZN(n28049) );
  CLKNHSV0 U31611 ( .I(n49533), .ZN(n28050) );
  CLKNHSV0 U31612 ( .I(n52202), .ZN(n28051) );
  MUX2NHSV0 U31613 ( .I0(n28051), .I1(n52202), .S(n52455), .ZN(n28052) );
  MUX2NHSV0 U31614 ( .I0(n28050), .I1(n49533), .S(n28052), .ZN(n28053) );
  MUX2NHSV0 U31615 ( .I0(n28049), .I1(n49528), .S(n28053), .ZN(n28054) );
  AO22HSV0 U31616 ( .A1(n50956), .A2(n52448), .B1(n44750), .B2(n51805), .Z(
        n28055) );
  CLKNHSV0 U31617 ( .I(n51814), .ZN(n28056) );
  MUX2NHSV0 U31618 ( .I0(n51814), .I1(n28056), .S(n48936), .ZN(n28057) );
  AOI22HSV0 U31619 ( .A1(n52449), .A2(n52905), .B1(n52289), .B2(n51803), .ZN(
        n28058) );
  AOI21HSV0 U31620 ( .A1(n45293), .A2(n52947), .B(n28058), .ZN(n28059) );
  NAND2HSV0 U31621 ( .A1(n28059), .A2(n28057), .ZN(n28060) );
  OAI21HSV0 U31622 ( .A1(n28059), .A2(n28057), .B(n28060), .ZN(n28061) );
  OAI21HSV0 U31623 ( .A1(n45294), .A2(n52219), .B(n28055), .ZN(n28062) );
  CLKNAND2HSV0 U31624 ( .A1(n28062), .A2(n28061), .ZN(n28063) );
  OAI21HSV0 U31625 ( .A1(n28062), .A2(n28061), .B(n28063), .ZN(n28064) );
  XOR2HSV0 U31626 ( .A1(n28054), .A2(n28064), .Z(n45343) );
  XOR2HSV0 U31627 ( .A1(n41862), .A2(n41863), .Z(n28065) );
  XOR2HSV0 U31628 ( .A1(n41857), .A2(n41856), .Z(n28066) );
  XOR2HSV0 U31629 ( .A1(n28065), .A2(n28066), .Z(n28067) );
  XOR2HSV0 U31630 ( .A1(n41875), .A2(n41876), .Z(n28068) );
  XOR2HSV0 U31631 ( .A1(n41869), .A2(n41868), .Z(n28069) );
  XOR2HSV0 U31632 ( .A1(n28068), .A2(n28069), .Z(n28070) );
  XOR2HSV0 U31633 ( .A1(n41891), .A2(n41892), .Z(n28071) );
  XOR2HSV0 U31634 ( .A1(n41884), .A2(n41883), .Z(n28072) );
  XOR2HSV0 U31635 ( .A1(n28071), .A2(n28072), .Z(n28073) );
  XOR2HSV0 U31636 ( .A1(n28067), .A2(n28070), .Z(n28074) );
  XOR2HSV0 U31637 ( .A1(n28073), .A2(n28074), .Z(n28075) );
  NAND2HSV0 U31638 ( .A1(n59529), .A2(n55337), .ZN(n28076) );
  CLKNAND2HSV0 U31639 ( .A1(n28076), .A2(n28075), .ZN(n28077) );
  OAI21HSV0 U31640 ( .A1(n28075), .A2(n28076), .B(n28077), .ZN(n28078) );
  NAND2HSV0 U31641 ( .A1(n42275), .A2(n42155), .ZN(n28079) );
  CLKNAND2HSV0 U31642 ( .A1(n28079), .A2(n28078), .ZN(n28080) );
  OAI21HSV0 U31643 ( .A1(n28078), .A2(n28079), .B(n28080), .ZN(n28081) );
  NAND2HSV0 U31644 ( .A1(n41609), .A2(n54969), .ZN(n28082) );
  CLKNAND2HSV0 U31645 ( .A1(n28082), .A2(n28081), .ZN(n28083) );
  OAI21HSV0 U31646 ( .A1(n28081), .A2(n28082), .B(n28083), .ZN(n28084) );
  CLKNAND2HSV0 U31647 ( .A1(n53602), .A2(n41550), .ZN(n28085) );
  CLKNAND2HSV0 U31648 ( .A1(n28085), .A2(n28084), .ZN(n28086) );
  OAI21HSV0 U31649 ( .A1(n28084), .A2(n28085), .B(n28086), .ZN(n28087) );
  NAND2HSV0 U31650 ( .A1(n59919), .A2(n42162), .ZN(n28088) );
  CLKNAND2HSV0 U31651 ( .A1(n28088), .A2(n28087), .ZN(n28089) );
  OAI21HSV0 U31652 ( .A1(n28087), .A2(n28088), .B(n28089), .ZN(n28090) );
  NAND2HSV0 U31653 ( .A1(n42089), .A2(n41851), .ZN(n28091) );
  CLKNAND2HSV0 U31654 ( .A1(n28091), .A2(n28090), .ZN(n28092) );
  OAI21HSV0 U31655 ( .A1(n28090), .A2(n28091), .B(n28092), .ZN(n28093) );
  NAND2HSV0 U31656 ( .A1(n42359), .A2(n29773), .ZN(n28094) );
  CLKNAND2HSV0 U31657 ( .A1(n28094), .A2(n28093), .ZN(n28095) );
  OAI21HSV0 U31658 ( .A1(n28093), .A2(n28094), .B(n28095), .ZN(n28096) );
  OAI21HSV0 U31659 ( .A1(n41802), .A2(n41928), .B(n28096), .ZN(n28097) );
  OAI31HSV0 U31660 ( .A1(n41802), .A2(n28096), .A3(n41928), .B(n28097), .ZN(
        n28098) );
  NAND2HSV0 U31661 ( .A1(n41676), .A2(n41894), .ZN(n28099) );
  CLKNAND2HSV0 U31662 ( .A1(n28099), .A2(n28098), .ZN(n28100) );
  OAI21HSV0 U31663 ( .A1(n28098), .A2(n28099), .B(n28100), .ZN(n28101) );
  NAND2HSV0 U31664 ( .A1(n54724), .A2(n54264), .ZN(n28102) );
  CLKNAND2HSV0 U31665 ( .A1(n28102), .A2(n28101), .ZN(n28103) );
  OAI21HSV0 U31666 ( .A1(n28101), .A2(n28102), .B(n28103), .ZN(n41895) );
  INAND2HSV0 U31667 ( .A1(n33660), .B1(n52723), .ZN(n33401) );
  NAND2HSV0 U31668 ( .A1(n59420), .A2(\pe6/got [13]), .ZN(n59311) );
  NOR2HSV0 U31669 ( .A1(n38269), .A2(n38268), .ZN(n28104) );
  NAND2HSV2 U31670 ( .A1(n28104), .A2(n38444), .ZN(n38363) );
  XOR2HSV0 U31671 ( .A1(n56540), .A2(n56539), .Z(n28105) );
  XOR2HSV0 U31672 ( .A1(n56538), .A2(n28105), .Z(n28106) );
  NAND2HSV0 U31673 ( .A1(n59811), .A2(n56541), .ZN(n28107) );
  CLKNAND2HSV0 U31674 ( .A1(n28107), .A2(n28106), .ZN(n28108) );
  OAI21HSV0 U31675 ( .A1(n28106), .A2(n28107), .B(n28108), .ZN(n28109) );
  NAND2HSV0 U31676 ( .A1(n56624), .A2(n56781), .ZN(n28110) );
  CLKNAND2HSV0 U31677 ( .A1(n28110), .A2(n28109), .ZN(n28111) );
  OAI21HSV0 U31678 ( .A1(n28109), .A2(n28110), .B(n28111), .ZN(n28112) );
  NAND2HSV0 U31679 ( .A1(n45582), .A2(n56623), .ZN(n28113) );
  CLKNAND2HSV0 U31680 ( .A1(n28113), .A2(n28112), .ZN(n28114) );
  OAI21HSV0 U31681 ( .A1(n28112), .A2(n28113), .B(n28114), .ZN(n28115) );
  NAND2HSV0 U31682 ( .A1(n56562), .A2(n56560), .ZN(n28116) );
  CLKNAND2HSV0 U31683 ( .A1(n28116), .A2(n28115), .ZN(n28117) );
  OAI21HSV0 U31684 ( .A1(n28115), .A2(n28116), .B(n28117), .ZN(n28118) );
  NAND2HSV0 U31685 ( .A1(n56497), .A2(n56888), .ZN(n28119) );
  CLKNAND2HSV0 U31686 ( .A1(n28119), .A2(n28118), .ZN(n28120) );
  OAI21HSV2 U31687 ( .A1(n28118), .A2(n28119), .B(n28120), .ZN(n28121) );
  NAND2HSV0 U31688 ( .A1(n56622), .A2(n56855), .ZN(n28122) );
  NAND2HSV2 U31689 ( .A1(n28122), .A2(n28121), .ZN(n28123) );
  OAI21HSV2 U31690 ( .A1(n28121), .A2(n28122), .B(n28123), .ZN(n28124) );
  NAND2HSV0 U31691 ( .A1(n56783), .A2(n56559), .ZN(n28125) );
  NAND2HSV2 U31692 ( .A1(n28125), .A2(n28124), .ZN(n28126) );
  OAI21HSV2 U31693 ( .A1(n28124), .A2(n28125), .B(n28126), .ZN(n56542) );
  CLKNHSV0 U31694 ( .I(\pe3/ti_7t [30]), .ZN(n28127) );
  AOI21HSV0 U31695 ( .A1(n45932), .A2(n28127), .B(n45931), .ZN(n46558) );
  XOR2HSV0 U31696 ( .A1(n57306), .A2(n57305), .Z(n28128) );
  AOI21HSV0 U31697 ( .A1(n33918), .A2(n57820), .B(n28128), .ZN(n28129) );
  AO31HSV2 U31698 ( .A1(n33918), .A2(n57820), .A3(n28128), .B(n28129), .Z(
        n28130) );
  NAND2HSV0 U31699 ( .A1(n57675), .A2(n57424), .ZN(n28131) );
  CLKNAND2HSV0 U31700 ( .A1(n28131), .A2(n28130), .ZN(n28132) );
  OAI21HSV0 U31701 ( .A1(n28130), .A2(n28131), .B(n28132), .ZN(n28133) );
  NAND2HSV0 U31702 ( .A1(n57307), .A2(n57985), .ZN(n28134) );
  CLKNAND2HSV0 U31703 ( .A1(n28134), .A2(n28133), .ZN(n28135) );
  OAI21HSV0 U31704 ( .A1(n28133), .A2(n28134), .B(n28135), .ZN(n28136) );
  NAND2HSV0 U31705 ( .A1(\pe4/got [16]), .A2(n57984), .ZN(n28137) );
  CLKNAND2HSV0 U31706 ( .A1(n28137), .A2(n28136), .ZN(n28138) );
  OAI21HSV0 U31707 ( .A1(n28136), .A2(n28137), .B(n28138), .ZN(n28139) );
  CLKNAND2HSV0 U31708 ( .A1(n57427), .A2(n57457), .ZN(n28140) );
  CLKNAND2HSV0 U31709 ( .A1(n28140), .A2(n28139), .ZN(n28141) );
  OAI21HSV0 U31710 ( .A1(n28139), .A2(n28140), .B(n28141), .ZN(n28142) );
  CLKNAND2HSV0 U31711 ( .A1(\pe4/got [19]), .A2(n57308), .ZN(n28143) );
  CLKNAND2HSV0 U31712 ( .A1(n28143), .A2(n28142), .ZN(n28144) );
  OAI21HSV0 U31713 ( .A1(n28142), .A2(n28143), .B(n28144), .ZN(n28145) );
  CLKNAND2HSV0 U31714 ( .A1(n57554), .A2(n34042), .ZN(n28146) );
  CLKNAND2HSV0 U31715 ( .A1(n28146), .A2(n28145), .ZN(n28147) );
  OAI21HSV0 U31716 ( .A1(n28145), .A2(n28146), .B(n28147), .ZN(n28148) );
  NAND2HSV0 U31717 ( .A1(n59386), .A2(n34429), .ZN(n28149) );
  CLKNAND2HSV0 U31718 ( .A1(n28149), .A2(n28148), .ZN(n28150) );
  OAI21HSV0 U31719 ( .A1(n28148), .A2(n28149), .B(n28150), .ZN(n28151) );
  NAND2HSV0 U31720 ( .A1(n59601), .A2(n57819), .ZN(n28152) );
  CLKNAND2HSV0 U31721 ( .A1(n28152), .A2(n28151), .ZN(n28153) );
  OAI21HSV2 U31722 ( .A1(n28151), .A2(n28152), .B(n28153), .ZN(n28154) );
  NAND2HSV0 U31723 ( .A1(n57760), .A2(n57560), .ZN(n28155) );
  NAND2HSV2 U31724 ( .A1(n28155), .A2(n28154), .ZN(n28156) );
  OAI21HSV2 U31725 ( .A1(n28154), .A2(n28155), .B(n28156), .ZN(n28157) );
  CLKNAND2HSV0 U31726 ( .A1(n57309), .A2(n47904), .ZN(n28158) );
  NAND2HSV2 U31727 ( .A1(n28158), .A2(n28157), .ZN(n28159) );
  OAI21HSV2 U31728 ( .A1(n28157), .A2(n28158), .B(n28159), .ZN(n28160) );
  NAND2HSV0 U31729 ( .A1(n57574), .A2(n57310), .ZN(n28161) );
  CLKNAND2HSV0 U31730 ( .A1(n28161), .A2(n28160), .ZN(n28162) );
  OAI21HSV0 U31731 ( .A1(n28160), .A2(n28161), .B(n28162), .ZN(n57311) );
  CLKNHSV0 U31732 ( .I(\pe2/ti_7t [16]), .ZN(n28163) );
  AOI21HSV0 U31733 ( .A1(ctro2), .A2(n28163), .B(n38375), .ZN(n46121) );
  XOR2HSV0 U31734 ( .A1(n58475), .A2(n58474), .Z(n28164) );
  NAND2HSV0 U31735 ( .A1(n58611), .A2(\pe6/got [3]), .ZN(n28165) );
  CLKNAND2HSV0 U31736 ( .A1(n28165), .A2(n28164), .ZN(n28166) );
  OAI21HSV0 U31737 ( .A1(n28164), .A2(n28165), .B(n28166), .ZN(n28167) );
  NAND2HSV0 U31738 ( .A1(n58716), .A2(n46173), .ZN(n28168) );
  CLKNAND2HSV0 U31739 ( .A1(n28168), .A2(n28167), .ZN(n28169) );
  OAI21HSV0 U31740 ( .A1(n28167), .A2(n28168), .B(n28169), .ZN(n28170) );
  NAND2HSV0 U31741 ( .A1(n29753), .A2(n58661), .ZN(n28171) );
  CLKNAND2HSV0 U31742 ( .A1(n28171), .A2(n28170), .ZN(n28172) );
  OAI21HSV0 U31743 ( .A1(n28170), .A2(n28171), .B(n28172), .ZN(n28173) );
  NAND2HSV0 U31744 ( .A1(n59026), .A2(n58659), .ZN(n28174) );
  CLKNAND2HSV0 U31745 ( .A1(n28174), .A2(n28173), .ZN(n28175) );
  OAI21HSV0 U31746 ( .A1(n28173), .A2(n28174), .B(n28175), .ZN(n28176) );
  CLKNAND2HSV0 U31747 ( .A1(n46156), .A2(n58562), .ZN(n28177) );
  CLKNAND2HSV0 U31748 ( .A1(n28177), .A2(n28176), .ZN(n28178) );
  OAI21HSV0 U31749 ( .A1(n28176), .A2(n28177), .B(n28178), .ZN(n28179) );
  NAND2HSV0 U31750 ( .A1(n58526), .A2(n46145), .ZN(n28180) );
  CLKNAND2HSV0 U31751 ( .A1(n28180), .A2(n28179), .ZN(n28181) );
  OAI21HSV0 U31752 ( .A1(n28179), .A2(n28180), .B(n28181), .ZN(n28182) );
  NAND2HSV0 U31753 ( .A1(n58477), .A2(n48888), .ZN(n28183) );
  CLKNAND2HSV0 U31754 ( .A1(n28183), .A2(n28182), .ZN(n28184) );
  CLKNAND2HSV0 U31755 ( .A1(n28185), .A2(n28186), .ZN(n28187) );
  XOR2HSV0 U31756 ( .A1(n51009), .A2(n51008), .Z(n28188) );
  NAND2HSV0 U31757 ( .A1(n51728), .A2(n52050), .ZN(n28189) );
  CLKNAND2HSV0 U31758 ( .A1(n28189), .A2(n28188), .ZN(n28190) );
  OAI21HSV0 U31759 ( .A1(n28188), .A2(n28189), .B(n28190), .ZN(n28191) );
  XOR2HSV0 U31760 ( .A1(n51010), .A2(n28191), .Z(n28192) );
  NAND2HSV0 U31761 ( .A1(n51797), .A2(n59685), .ZN(n28193) );
  CLKNAND2HSV0 U31762 ( .A1(n28193), .A2(n28192), .ZN(n28194) );
  OAI21HSV0 U31763 ( .A1(n28192), .A2(n28193), .B(n28194), .ZN(n28195) );
  NAND2HSV0 U31764 ( .A1(n51120), .A2(n52922), .ZN(n28196) );
  CLKNAND2HSV0 U31765 ( .A1(n28196), .A2(n28195), .ZN(n28197) );
  OAI21HSV0 U31766 ( .A1(n28195), .A2(n28196), .B(n28197), .ZN(n28198) );
  NAND2HSV0 U31767 ( .A1(n52840), .A2(n45249), .ZN(n28200) );
  NAND2HSV0 U31768 ( .A1(n39008), .A2(n51961), .ZN(n28203) );
  CLKNAND2HSV0 U31769 ( .A1(n28203), .A2(n28202), .ZN(n28204) );
  OAI21HSV0 U31770 ( .A1(n28202), .A2(n28203), .B(n28204), .ZN(\pe2/poht [8])
         );
  XOR2HSV0 U31771 ( .A1(n48738), .A2(n48737), .Z(n28205) );
  AOI21HSV0 U31772 ( .A1(n48743), .A2(n52670), .B(n28205), .ZN(n28206) );
  AO31HSV2 U31773 ( .A1(n48743), .A2(n52670), .A3(n28205), .B(n28206), .Z(
        n28207) );
  NAND2HSV0 U31774 ( .A1(n51227), .A2(n48739), .ZN(n28208) );
  CLKNAND2HSV0 U31775 ( .A1(n28208), .A2(n28207), .ZN(n28209) );
  OAI21HSV0 U31776 ( .A1(n28207), .A2(n28208), .B(n28209), .ZN(n28210) );
  NAND2HSV0 U31777 ( .A1(n52835), .A2(n48742), .ZN(n28211) );
  CLKNAND2HSV0 U31778 ( .A1(n28211), .A2(n28210), .ZN(n28212) );
  OAI21HSV0 U31779 ( .A1(n28210), .A2(n28211), .B(n28212), .ZN(n28213) );
  NAND2HSV0 U31780 ( .A1(n59933), .A2(\pe5/got [27]), .ZN(n28214) );
  CLKNAND2HSV0 U31781 ( .A1(n28214), .A2(n28213), .ZN(n28215) );
  OAI21HSV0 U31782 ( .A1(n28213), .A2(n28214), .B(n28215), .ZN(n28216) );
  NAND2HSV0 U31783 ( .A1(n29777), .A2(n39430), .ZN(n28217) );
  CLKNAND2HSV0 U31784 ( .A1(n28217), .A2(n28216), .ZN(n28218) );
  OAI21HSV0 U31785 ( .A1(n28216), .A2(n28217), .B(n28218), .ZN(n28219) );
  NAND2HSV0 U31786 ( .A1(\pe5/got [29]), .A2(n59580), .ZN(n28220) );
  CLKNAND2HSV0 U31787 ( .A1(n48886), .A2(n48740), .ZN(n28223) );
  CLKNAND2HSV0 U31788 ( .A1(n28223), .A2(n28222), .ZN(n28224) );
  OAI21HSV0 U31789 ( .A1(n28222), .A2(n28223), .B(n28224), .ZN(\pe5/poht [2])
         );
  OAI22HSV0 U31790 ( .A1(n46663), .A2(n59094), .B1(n44403), .B2(n32858), .ZN(
        n28225) );
  OAI21HSV0 U31791 ( .A1(n58863), .A2(n36120), .B(n28225), .ZN(n36121) );
  XOR2HSV0 U31792 ( .A1(n33418), .A2(n33419), .Z(n28226) );
  CLKXOR2HSV4 U31793 ( .A1(n33417), .A2(n33416), .Z(n28227) );
  XOR2HSV4 U31794 ( .A1(n28226), .A2(n28227), .Z(n28228) );
  CLKXOR2HSV2 U31795 ( .A1(n33424), .A2(n33425), .Z(n28229) );
  XOR2HSV0 U31796 ( .A1(n33422), .A2(n33421), .Z(n28230) );
  CLKXOR2HSV2 U31797 ( .A1(n28229), .A2(n28230), .Z(n28231) );
  XOR2HSV4 U31798 ( .A1(n28228), .A2(n28231), .Z(n33434) );
  INOR2HSV1 U31799 ( .A1(\pe1/ti_7t [11]), .B1(n41217), .ZN(n40809) );
  AOI22HSV0 U31800 ( .A1(n52344), .A2(n36608), .B1(n52438), .B2(n39052), .ZN(
        n28232) );
  IAO21HSV0 U31801 ( .A1(n52437), .A2(n52436), .B(n28232), .ZN(n52439) );
  CLKNHSV0 U31802 ( .I(\pe2/phq [10]), .ZN(n28233) );
  NAND2HSV4 U31803 ( .A1(n48078), .A2(\pe2/pvq [10]), .ZN(n28234) );
  MUX2NHSV4 U31804 ( .I0(\pe2/phq [10]), .I1(n28233), .S(n28234), .ZN(n36339)
         );
  XOR2HSV0 U31805 ( .A1(n33979), .A2(n33978), .Z(n28235) );
  XOR2HSV0 U31806 ( .A1(n33977), .A2(n28235), .Z(n28236) );
  NAND2HSV0 U31807 ( .A1(n34410), .A2(n34458), .ZN(n28237) );
  NAND2HSV0 U31808 ( .A1(n28237), .A2(n28236), .ZN(n28238) );
  OAI21HSV2 U31809 ( .A1(n28236), .A2(n28237), .B(n28238), .ZN(n33980) );
  XOR2HSV0 U31810 ( .A1(n38254), .A2(n38252), .Z(n28239) );
  XOR2HSV0 U31811 ( .A1(n38251), .A2(n38253), .Z(n28240) );
  XOR2HSV0 U31812 ( .A1(n28239), .A2(n28240), .Z(n28241) );
  AOI21HSV0 U31813 ( .A1(n38781), .A2(n38702), .B(n28241), .ZN(n28242) );
  AO31HSV0 U31814 ( .A1(n38781), .A2(n38702), .A3(n28241), .B(n28242), .Z(
        n28243) );
  NAND2HSV0 U31815 ( .A1(n59982), .A2(n52934), .ZN(n28244) );
  CLKNAND2HSV0 U31816 ( .A1(n28244), .A2(n28243), .ZN(n28245) );
  OAI21HSV0 U31817 ( .A1(n28243), .A2(n28244), .B(n28245), .ZN(n28246) );
  NAND2HSV0 U31818 ( .A1(n39011), .A2(n39010), .ZN(n28247) );
  CLKNAND2HSV0 U31819 ( .A1(n28247), .A2(n28246), .ZN(n28248) );
  OAI21HSV0 U31820 ( .A1(n28246), .A2(n28247), .B(n28248), .ZN(n28249) );
  NAND2HSV0 U31821 ( .A1(n52367), .A2(n52167), .ZN(n28250) );
  CLKNAND2HSV0 U31822 ( .A1(n28250), .A2(n28249), .ZN(n28251) );
  OAI21HSV0 U31823 ( .A1(n28249), .A2(n28250), .B(n28251), .ZN(n28252) );
  NAND2HSV0 U31824 ( .A1(n45218), .A2(n38904), .ZN(n28253) );
  CLKNAND2HSV0 U31825 ( .A1(n28253), .A2(n28252), .ZN(n28254) );
  OAI21HSV0 U31826 ( .A1(n28252), .A2(n28253), .B(n28254), .ZN(n28255) );
  NAND2HSV0 U31827 ( .A1(\pe2/got [23]), .A2(n38780), .ZN(n28256) );
  CLKNAND2HSV0 U31828 ( .A1(n28256), .A2(n28255), .ZN(n28257) );
  OAI21HSV2 U31829 ( .A1(n28255), .A2(n28256), .B(n28257), .ZN(n38256) );
  XOR2HSV0 U31830 ( .A1(n51192), .A2(n51193), .Z(n28258) );
  XOR2HSV0 U31831 ( .A1(n51190), .A2(n51189), .Z(n28259) );
  XOR2HSV0 U31832 ( .A1(n28258), .A2(n28259), .Z(n28260) );
  XOR2HSV0 U31833 ( .A1(n51180), .A2(n51181), .Z(n28261) );
  XOR2HSV0 U31834 ( .A1(n51179), .A2(n51178), .Z(n28262) );
  XOR2HSV0 U31835 ( .A1(n28261), .A2(n28262), .Z(n28263) );
  XOR2HSV0 U31836 ( .A1(n51185), .A2(n51186), .Z(n28264) );
  XOR2HSV0 U31837 ( .A1(n51184), .A2(n51183), .Z(n28265) );
  XOR2HSV0 U31838 ( .A1(n28264), .A2(n28265), .Z(n28266) );
  XOR2HSV0 U31839 ( .A1(n51196), .A2(n51197), .Z(n28267) );
  XOR2HSV0 U31840 ( .A1(n51195), .A2(n51194), .Z(n28268) );
  XOR2HSV0 U31841 ( .A1(n28267), .A2(n28268), .Z(n28269) );
  CLKNHSV0 U31842 ( .I(n51174), .ZN(n28270) );
  OAI21HSV0 U31843 ( .A1(n51166), .A2(n51165), .B(n51175), .ZN(n28271) );
  OAI31HSV0 U31844 ( .A1(n51166), .A2(n51175), .A3(n51165), .B(n28271), .ZN(
        n28272) );
  MUX2NHSV0 U31845 ( .I0(n28270), .I1(n51174), .S(n28272), .ZN(n28273) );
  XOR2HSV0 U31846 ( .A1(n28273), .A2(n51168), .Z(n28274) );
  XOR2HSV0 U31847 ( .A1(n28269), .A2(n51169), .Z(n28275) );
  XOR2HSV0 U31848 ( .A1(n28274), .A2(n28275), .Z(n28276) );
  XOR2HSV0 U31849 ( .A1(n28276), .A2(n28266), .Z(n28277) );
  XOR2HSV0 U31850 ( .A1(n28260), .A2(n28263), .Z(n28278) );
  XOR2HSV0 U31851 ( .A1(n28277), .A2(n28278), .Z(n28279) );
  NAND2HSV0 U31852 ( .A1(n51362), .A2(n51162), .ZN(n28280) );
  CLKNAND2HSV0 U31853 ( .A1(n28280), .A2(n28279), .ZN(n28281) );
  OAI21HSV0 U31854 ( .A1(n28279), .A2(n28280), .B(n28281), .ZN(n28282) );
  NAND2HSV0 U31855 ( .A1(n51161), .A2(n29770), .ZN(n28283) );
  NAND2HSV0 U31856 ( .A1(n28283), .A2(n28282), .ZN(n28284) );
  OAI21HSV2 U31857 ( .A1(n28282), .A2(n28283), .B(n28284), .ZN(n28285) );
  NAND2HSV0 U31858 ( .A1(n51331), .A2(n52575), .ZN(n28286) );
  NAND2HSV2 U31859 ( .A1(n28286), .A2(n28285), .ZN(n28287) );
  OAI21HSV2 U31860 ( .A1(n28285), .A2(n28286), .B(n28287), .ZN(n28288) );
  NAND2HSV0 U31861 ( .A1(n52574), .A2(n51302), .ZN(n28289) );
  NAND2HSV0 U31862 ( .A1(n28289), .A2(n28288), .ZN(n28290) );
  OAI21HSV0 U31863 ( .A1(n28288), .A2(n28289), .B(n28290), .ZN(n51198) );
  INAND2HSV0 U31864 ( .A1(\pe2/ti_7t [20]), .B1(n38630), .ZN(n38878) );
  AOI21HSV4 U31865 ( .A1(n47943), .A2(n34841), .B(n34840), .ZN(n28291) );
  CLKNAND2HSV4 U31866 ( .A1(n34848), .A2(n28291), .ZN(n35026) );
  INOR2HSV0 U31867 ( .A1(\pe3/ti_7t [24]), .B1(n43604), .ZN(n45509) );
  XOR2HSV0 U31868 ( .A1(n57887), .A2(n57886), .Z(n28292) );
  NAND2HSV0 U31869 ( .A1(n59378), .A2(\pe4/got [3]), .ZN(n28293) );
  CLKNAND2HSV0 U31870 ( .A1(n28293), .A2(n28292), .ZN(n28294) );
  OAI21HSV0 U31871 ( .A1(n28292), .A2(n28293), .B(n28294), .ZN(n28295) );
  NAND2HSV0 U31872 ( .A1(n58206), .A2(n25284), .ZN(n28296) );
  CLKNAND2HSV0 U31873 ( .A1(n28296), .A2(n28295), .ZN(n28297) );
  OAI21HSV0 U31874 ( .A1(n28295), .A2(n28296), .B(n28297), .ZN(n28298) );
  NAND2HSV0 U31875 ( .A1(n57951), .A2(n57984), .ZN(n28299) );
  CLKNAND2HSV0 U31876 ( .A1(n28299), .A2(n28298), .ZN(n28300) );
  OAI21HSV0 U31877 ( .A1(n28298), .A2(n28299), .B(n28300), .ZN(n28301) );
  NAND2HSV0 U31878 ( .A1(n57427), .A2(\pe4/got [6]), .ZN(n28302) );
  CLKNAND2HSV0 U31879 ( .A1(n28302), .A2(n28301), .ZN(n28303) );
  OAI21HSV0 U31880 ( .A1(n28301), .A2(n28302), .B(n28303), .ZN(n28304) );
  NAND2HSV0 U31881 ( .A1(n58029), .A2(n58111), .ZN(n28305) );
  CLKNAND2HSV0 U31882 ( .A1(n28305), .A2(n28304), .ZN(n28306) );
  OAI21HSV0 U31883 ( .A1(n28304), .A2(n28305), .B(n28306), .ZN(n28307) );
  NAND2HSV0 U31884 ( .A1(n59935), .A2(n58102), .ZN(n28308) );
  CLKNAND2HSV0 U31885 ( .A1(n28308), .A2(n28307), .ZN(n28309) );
  OAI21HSV0 U31886 ( .A1(n28307), .A2(n28308), .B(n28309), .ZN(n28310) );
  CLKNAND2HSV0 U31887 ( .A1(n58112), .A2(n58041), .ZN(n28311) );
  CLKNAND2HSV0 U31888 ( .A1(n28311), .A2(n28310), .ZN(n28312) );
  OAI21HSV0 U31889 ( .A1(n28310), .A2(n28311), .B(n28312), .ZN(n28313) );
  NAND2HSV0 U31890 ( .A1(n58153), .A2(n58183), .ZN(n28314) );
  CLKNAND2HSV0 U31891 ( .A1(n28314), .A2(n28313), .ZN(n28315) );
  OAI21HSV0 U31892 ( .A1(n28313), .A2(n28314), .B(n28315), .ZN(n28316) );
  NAND2HSV0 U31893 ( .A1(n57960), .A2(n59663), .ZN(n28317) );
  CLKNAND2HSV0 U31894 ( .A1(n28317), .A2(n28316), .ZN(n28318) );
  OAI21HSV0 U31895 ( .A1(n28316), .A2(n28317), .B(n28318), .ZN(n28319) );
  CLKNAND2HSV0 U31896 ( .A1(n57889), .A2(n57888), .ZN(n28320) );
  CLKNAND2HSV0 U31897 ( .A1(n28320), .A2(n28319), .ZN(n28321) );
  OAI21HSV0 U31898 ( .A1(n28319), .A2(n28320), .B(n28321), .ZN(n28322) );
  CLKNAND2HSV0 U31899 ( .A1(\pe4/got [13]), .A2(n57755), .ZN(n28323) );
  CLKNAND2HSV0 U31900 ( .A1(n28323), .A2(n28322), .ZN(n28324) );
  OAI21HSV0 U31901 ( .A1(n28322), .A2(n28323), .B(n28324), .ZN(n57890) );
  NAND2HSV0 U31902 ( .A1(n51532), .A2(\pe2/aot [2]), .ZN(n28325) );
  AOI21HSV0 U31903 ( .A1(n51493), .A2(n53016), .B(n28325), .ZN(n28326) );
  AO31HSV2 U31904 ( .A1(n51493), .A2(n53016), .A3(n28325), .B(n28326), .Z(
        n28327) );
  NAND2HSV0 U31905 ( .A1(n52840), .A2(n52901), .ZN(n28328) );
  NAND2HSV0 U31906 ( .A1(n52895), .A2(n51961), .ZN(n28331) );
  CLKNAND2HSV0 U31907 ( .A1(n28331), .A2(n28330), .ZN(n28332) );
  OAI21HSV0 U31908 ( .A1(n28330), .A2(n28331), .B(n28332), .ZN(\pe2/poht [30])
         );
  XOR2HSV0 U31909 ( .A1(n58708), .A2(n58707), .Z(n28333) );
  XOR2HSV0 U31910 ( .A1(n58710), .A2(n28333), .Z(n28334) );
  AOI21HSV0 U31911 ( .A1(n59182), .A2(n35712), .B(n28334), .ZN(n28335) );
  AO31HSV2 U31912 ( .A1(n59182), .A2(n35712), .A3(n28334), .B(n28335), .Z(
        n28336) );
  NAND2HSV0 U31913 ( .A1(n58402), .A2(n58658), .ZN(n28337) );
  CLKNAND2HSV0 U31914 ( .A1(n28337), .A2(n28336), .ZN(n28338) );
  OAI21HSV0 U31915 ( .A1(n28336), .A2(n28337), .B(n28338), .ZN(n28339) );
  NAND2HSV0 U31916 ( .A1(n53172), .A2(n58812), .ZN(n28340) );
  CLKNAND2HSV0 U31917 ( .A1(n28340), .A2(n28339), .ZN(n28341) );
  OAI21HSV0 U31918 ( .A1(n28339), .A2(n28340), .B(n28341), .ZN(n28342) );
  CLKNAND2HSV0 U31919 ( .A1(n58657), .A2(n49742), .ZN(n28343) );
  CLKNAND2HSV0 U31920 ( .A1(n28343), .A2(n28342), .ZN(n28344) );
  OAI21HSV0 U31921 ( .A1(n28342), .A2(n28343), .B(n28344), .ZN(n28345) );
  NAND2HSV0 U31922 ( .A1(n58656), .A2(\pe6/got [12]), .ZN(n28346) );
  CLKNAND2HSV0 U31923 ( .A1(n28346), .A2(n28345), .ZN(n28347) );
  OAI21HSV0 U31924 ( .A1(n28345), .A2(n28346), .B(n28347), .ZN(n28348) );
  NAND2HSV0 U31925 ( .A1(n58712), .A2(n58711), .ZN(n28349) );
  CLKNAND2HSV0 U31926 ( .A1(n28349), .A2(n28348), .ZN(n28350) );
  OAI21HSV0 U31927 ( .A1(n28348), .A2(n28349), .B(n28350), .ZN(n28351) );
  NAND2HSV0 U31928 ( .A1(n58713), .A2(n48888), .ZN(n28352) );
  CLKNAND2HSV0 U31929 ( .A1(n28352), .A2(n28351), .ZN(n28353) );
  OAI21HSV2 U31930 ( .A1(n28351), .A2(n28352), .B(n28353), .ZN(n28354) );
  NAND2HSV0 U31931 ( .A1(n29772), .A2(\pe6/got [15]), .ZN(n28355) );
  CLKNAND2HSV0 U31932 ( .A1(n28354), .A2(n28355), .ZN(n28356) );
  OAI21HSV0 U31933 ( .A1(n28354), .A2(n28355), .B(n28356), .ZN(\pe6/poht [17])
         );
  CLKNAND2HSV0 U31934 ( .A1(n28357), .A2(n51119), .ZN(n28358) );
  OAI21HSV0 U31935 ( .A1(n51119), .A2(n28357), .B(n28358), .ZN(n28359) );
  NAND2HSV0 U31936 ( .A1(n52726), .A2(n56953), .ZN(n28360) );
  NAND2HSV0 U31937 ( .A1(n28360), .A2(n28359), .ZN(n28361) );
  OAI21HSV0 U31938 ( .A1(n28359), .A2(n28360), .B(n28361), .ZN(pov3[29]) );
  NAND2HSV0 U31939 ( .A1(n52856), .A2(n53094), .ZN(n28362) );
  NAND2HSV0 U31940 ( .A1(n28362), .A2(n47938), .ZN(n28363) );
  NAND2HSV0 U31941 ( .A1(n28365), .A2(n28364), .ZN(n28366) );
  OAI21HSV0 U31942 ( .A1(n28364), .A2(n28365), .B(n28366), .ZN(n60092) );
  XOR2HSV0 U31943 ( .A1(n52666), .A2(n52665), .Z(n28367) );
  NAND2HSV0 U31944 ( .A1(n52565), .A2(n45816), .ZN(n28368) );
  CLKNAND2HSV0 U31945 ( .A1(n28368), .A2(n28367), .ZN(n28369) );
  OAI21HSV0 U31946 ( .A1(n28367), .A2(n28368), .B(n28369), .ZN(n28370) );
  NAND2HSV0 U31947 ( .A1(n52693), .A2(n51228), .ZN(n28371) );
  CLKNAND2HSV0 U31948 ( .A1(n28371), .A2(n28370), .ZN(n28372) );
  OAI21HSV0 U31949 ( .A1(n28370), .A2(n28371), .B(n28372), .ZN(n28373) );
  CLKNAND2HSV0 U31950 ( .A1(n52835), .A2(\pe5/got [22]), .ZN(n28374) );
  CLKNAND2HSV0 U31951 ( .A1(n28374), .A2(n28373), .ZN(n28375) );
  OAI21HSV0 U31952 ( .A1(n28373), .A2(n28374), .B(n28375), .ZN(n28376) );
  CLKNAND2HSV0 U31953 ( .A1(n52563), .A2(n47200), .ZN(n28377) );
  CLKNAND2HSV0 U31954 ( .A1(n28377), .A2(n28376), .ZN(n28378) );
  OAI21HSV0 U31955 ( .A1(n28376), .A2(n28377), .B(n28378), .ZN(n28379) );
  CLKNAND2HSV0 U31956 ( .A1(n29779), .A2(n59637), .ZN(n28380) );
  CLKNAND2HSV0 U31957 ( .A1(n28380), .A2(n28379), .ZN(n28381) );
  OAI21HSV0 U31958 ( .A1(n28379), .A2(n28380), .B(n28381), .ZN(n28382) );
  NAND2HSV0 U31959 ( .A1(n52667), .A2(n37630), .ZN(n28383) );
  CLKNAND2HSV0 U31960 ( .A1(n28383), .A2(n28382), .ZN(n28384) );
  OAI21HSV0 U31961 ( .A1(n28382), .A2(n28383), .B(n28384), .ZN(n28385) );
  NAND2HSV0 U31962 ( .A1(n52562), .A2(\pe5/got [26]), .ZN(n28386) );
  CLKNAND2HSV0 U31963 ( .A1(n28386), .A2(n28385), .ZN(n28387) );
  OAI21HSV0 U31964 ( .A1(n28385), .A2(n28386), .B(n28387), .ZN(\pe5/poht [6])
         );
  CLKNHSV0 U31965 ( .I(n57235), .ZN(n28388) );
  NAND2HSV0 U31966 ( .A1(\pe4/pvq [30]), .A2(n59486), .ZN(n28389) );
  NAND2HSV0 U31967 ( .A1(n28389), .A2(\pe4/phq [30]), .ZN(n28390) );
  OAI21HSV2 U31968 ( .A1(\pe4/phq [30]), .A2(n28389), .B(n28390), .ZN(n28391)
         );
  MUX2NHSV1 U31969 ( .I0(n57235), .I1(n28388), .S(n28391), .ZN(n35497) );
  CLKNHSV0 U31970 ( .I(n33950), .ZN(n28392) );
  NAND2HSV0 U31971 ( .A1(\pe4/pvq [12]), .A2(n34054), .ZN(n28393) );
  NAND2HSV0 U31972 ( .A1(n28393), .A2(\pe4/phq [12]), .ZN(n28394) );
  OAI21HSV2 U31973 ( .A1(\pe4/phq [12]), .A2(n28393), .B(n28394), .ZN(n28395)
         );
  MUX2NHSV0 U31974 ( .I0(n33950), .I1(n28392), .S(n28395), .ZN(n33553) );
  XOR2HSV0 U31975 ( .A1(n34364), .A2(n34366), .Z(n28396) );
  XOR2HSV0 U31976 ( .A1(n34365), .A2(n28396), .Z(n28397) );
  CLKNAND2HSV0 U31977 ( .A1(n35227), .A2(n57888), .ZN(n28398) );
  CLKNAND2HSV0 U31978 ( .A1(n28398), .A2(n28397), .ZN(n28399) );
  OAI21HSV2 U31979 ( .A1(n28397), .A2(n28398), .B(n28399), .ZN(n28400) );
  CLKXOR2HSV2 U31980 ( .A1(n28400), .A2(n34393), .Z(n28401) );
  XOR2HSV0 U31981 ( .A1(n34395), .A2(n34394), .Z(n28402) );
  CLKXOR2HSV2 U31982 ( .A1(n28401), .A2(n28402), .Z(n28403) );
  AOI21HSV0 U31983 ( .A1(n59630), .A2(n57285), .B(n28403), .ZN(n28404) );
  AO31HSV0 U31984 ( .A1(n59630), .A2(n57285), .A3(n28403), .B(n28404), .Z(
        n28405) );
  NAND2HSV0 U31985 ( .A1(n59382), .A2(n47657), .ZN(n28406) );
  NAND2HSV2 U31986 ( .A1(n28406), .A2(n28405), .ZN(n28407) );
  OAI21HSV0 U31987 ( .A1(n28405), .A2(n28406), .B(n28407), .ZN(n28408) );
  NAND2HSV0 U31988 ( .A1(n57307), .A2(n34868), .ZN(n28409) );
  NAND2HSV0 U31989 ( .A1(n28409), .A2(n28408), .ZN(n28410) );
  OAI21HSV0 U31990 ( .A1(n28408), .A2(n28409), .B(n28410), .ZN(n28411) );
  NAND2HSV0 U31991 ( .A1(n57526), .A2(n59604), .ZN(n28412) );
  NAND2HSV0 U31992 ( .A1(n28412), .A2(n28411), .ZN(n28413) );
  OAI21HSV0 U31993 ( .A1(n28411), .A2(n28412), .B(n28413), .ZN(n34397) );
  CLKNHSV0 U31994 ( .I(n35927), .ZN(n28414) );
  OAI21HSV0 U31995 ( .A1(n35837), .A2(n32245), .B(n35928), .ZN(n28415) );
  OAI21HSV0 U31996 ( .A1(n36160), .A2(n28414), .B(n28415), .ZN(n28416) );
  OAI22HSV0 U31997 ( .A1(n32714), .A2(n48042), .B1(n32086), .B2(n48041), .ZN(
        n28417) );
  OAI21HSV0 U31998 ( .A1(n36127), .A2(n35926), .B(n28417), .ZN(n28418) );
  NAND2HSV0 U31999 ( .A1(n28418), .A2(n28416), .ZN(n28419) );
  OAI21HSV0 U32000 ( .A1(n28418), .A2(n28416), .B(n28419), .ZN(n35931) );
  NAND2HSV0 U32001 ( .A1(n53014), .A2(\pe2/pvq [28]), .ZN(n28420) );
  NAND2HSV0 U32002 ( .A1(n28420), .A2(\pe2/phq [28]), .ZN(n28421) );
  OAI21HSV2 U32003 ( .A1(\pe2/phq [28]), .A2(n28420), .B(n28421), .ZN(n44727)
         );
  CLKNHSV0 U32004 ( .I(\pe4/phq [5]), .ZN(n28422) );
  NAND2HSV4 U32005 ( .A1(\pe4/aot [28]), .A2(n35075), .ZN(n28423) );
  NAND3HSV2 U32006 ( .A1(n45590), .A2(n45591), .A3(n45592), .ZN(n28424) );
  OAI22HSV0 U32007 ( .A1(n33113), .A2(n34631), .B1(n34117), .B2(n33355), .ZN(
        n28425) );
  OAI21HSV2 U32008 ( .A1(n33203), .A2(n33946), .B(n28425), .ZN(n33117) );
  IOA21HSV4 U32009 ( .A1(n35026), .A2(n35025), .B(n34981), .ZN(n35016) );
  CLKNHSV0 U32010 ( .I(n41260), .ZN(n28426) );
  NAND2HSV0 U32011 ( .A1(\pe1/bq[23] ), .A2(n59385), .ZN(n28427) );
  AOI22HSV0 U32012 ( .A1(n40827), .A2(n41738), .B1(n40828), .B2(n28427), .ZN(
        n28428) );
  MUX2NHSV0 U32013 ( .I0(n41260), .I1(n28426), .S(n28428), .ZN(n28429) );
  NAND2HSV0 U32014 ( .A1(n40875), .A2(n41248), .ZN(n28430) );
  NAND2HSV0 U32015 ( .A1(n28430), .A2(n28429), .ZN(n28431) );
  OAI21HSV2 U32016 ( .A1(n28429), .A2(n28430), .B(n28431), .ZN(n40841) );
  INOR2HSV0 U32017 ( .A1(\pe1/ti_7t [12]), .B1(n41134), .ZN(n40767) );
  NAND2HSV0 U32018 ( .A1(n57190), .A2(n34865), .ZN(n28432) );
  NAND2HSV2 U32019 ( .A1(n28432), .A2(n34813), .ZN(n28433) );
  OAI21HSV2 U32020 ( .A1(n34813), .A2(n28432), .B(n28433), .ZN(n28434) );
  NAND2HSV0 U32021 ( .A1(n34864), .A2(n29758), .ZN(n28435) );
  NAND2HSV2 U32022 ( .A1(n28435), .A2(n28434), .ZN(n28436) );
  OAI21HSV2 U32023 ( .A1(n28434), .A2(n28435), .B(n28436), .ZN(n34815) );
  INHSV2 U32024 ( .I(n40419), .ZN(n28437) );
  NAND2HSV0 U32025 ( .A1(n42223), .A2(n40491), .ZN(n28438) );
  MUX2NHSV2 U32026 ( .I0(n40419), .I1(n28437), .S(n28438), .ZN(n40420) );
  CLKNHSV0 U32027 ( .I(n51611), .ZN(n28439) );
  CLKNAND2HSV0 U32028 ( .A1(n53019), .A2(\pe2/bq[12] ), .ZN(n28440) );
  NAND2HSV0 U32029 ( .A1(n28440), .A2(n51738), .ZN(n28441) );
  OAI21HSV0 U32030 ( .A1(n51738), .A2(n28440), .B(n28441), .ZN(n28442) );
  NAND2HSV0 U32031 ( .A1(n51759), .A2(\pe2/bq[4] ), .ZN(n28443) );
  NAND2HSV0 U32032 ( .A1(n28443), .A2(n28442), .ZN(n28444) );
  OAI21HSV0 U32033 ( .A1(n28442), .A2(n28443), .B(n28444), .ZN(n28445) );
  MUX2NHSV0 U32034 ( .I0(n28439), .I1(n51611), .S(n28445), .ZN(n51648) );
  CLKNHSV0 U32035 ( .I(n29847), .ZN(n28446) );
  CLKNHSV0 U32036 ( .I(n29876), .ZN(n28447) );
  CLKNHSV0 U32037 ( .I(n29871), .ZN(n28448) );
  MUX2NHSV0 U32038 ( .I0(n28448), .I1(n29871), .S(n29872), .ZN(n28449) );
  NOR2HSV0 U32039 ( .A1(n40719), .A2(n40505), .ZN(n28451) );
  CLKNHSV0 U32040 ( .I(n40502), .ZN(n28452) );
  MUX2NHSV0 U32041 ( .I0(n28452), .I1(n40502), .S(n40503), .ZN(n28453) );
  AOI21HSV2 U32042 ( .A1(n40822), .A2(n41422), .B(n28453), .ZN(n28454) );
  AOI21HSV2 U32043 ( .A1(n41422), .A2(n28451), .B(n28454), .ZN(n28455) );
  AOI21HSV2 U32044 ( .A1(n28455), .A2(n40527), .B(n40668), .ZN(n28456) );
  OAI21HSV2 U32045 ( .A1(n28455), .A2(n40527), .B(n28456), .ZN(n28457) );
  CLKNAND2HSV2 U32046 ( .A1(n40541), .A2(n28457), .ZN(n40641) );
  OR2HSV1 U32047 ( .A1(n33094), .A2(\pe4/ti_7t [6]), .Z(n33226) );
  NOR2HSV0 U32048 ( .A1(n33660), .A2(n33929), .ZN(n28458) );
  NAND4HSV2 U32049 ( .A1(n33661), .A2(n33663), .A3(n33662), .A4(n28458), .ZN(
        n33664) );
  INHSV2 U32050 ( .I(n38616), .ZN(n28459) );
  CLKNHSV0 U32051 ( .I(n38615), .ZN(n28460) );
  MUX2NHSV0 U32052 ( .I0(n28460), .I1(n38615), .S(n28461), .ZN(n28462) );
  INOR2HSV0 U32053 ( .A1(\pe2/ti_7t [9]), .B1(n38183), .ZN(n37923) );
  XOR2HSV0 U32054 ( .A1(n58182), .A2(n58181), .Z(n28463) );
  XOR2HSV0 U32055 ( .A1(n58180), .A2(n28463), .Z(n28464) );
  AOI21HSV0 U32056 ( .A1(n58314), .A2(n58154), .B(n28464), .ZN(n28465) );
  AO31HSV2 U32057 ( .A1(n58314), .A2(n58154), .A3(n28464), .B(n28465), .Z(
        n28466) );
  NAND2HSV0 U32058 ( .A1(n58183), .A2(n58258), .ZN(n28467) );
  CLKNAND2HSV0 U32059 ( .A1(n28467), .A2(n28466), .ZN(n28468) );
  OAI21HSV0 U32060 ( .A1(n28466), .A2(n28467), .B(n28468), .ZN(n28469) );
  NAND2HSV0 U32061 ( .A1(\pe4/got [3]), .A2(n59672), .ZN(n28470) );
  CLKNAND2HSV0 U32062 ( .A1(n28470), .A2(n28469), .ZN(n28471) );
  OAI21HSV0 U32063 ( .A1(n28469), .A2(n28470), .B(n28471), .ZN(n28472) );
  NAND2HSV0 U32064 ( .A1(n58220), .A2(n58246), .ZN(n28473) );
  CLKNAND2HSV0 U32065 ( .A1(n28473), .A2(n28472), .ZN(n28474) );
  OAI21HSV0 U32066 ( .A1(n28472), .A2(n28473), .B(n28474), .ZN(n28475) );
  NAND2HSV0 U32067 ( .A1(n58185), .A2(n58184), .ZN(n28476) );
  CLKNAND2HSV0 U32068 ( .A1(n28476), .A2(n28475), .ZN(n28477) );
  OAI21HSV0 U32069 ( .A1(n28475), .A2(n28476), .B(n28477), .ZN(n28478) );
  CLKNAND2HSV0 U32070 ( .A1(n58216), .A2(n59837), .ZN(n28479) );
  CLKNAND2HSV0 U32071 ( .A1(n28479), .A2(n28478), .ZN(n28480) );
  OAI21HSV0 U32072 ( .A1(n28478), .A2(n28479), .B(n28480), .ZN(n28481) );
  NAND2HSV0 U32073 ( .A1(n58111), .A2(n58141), .ZN(n28482) );
  CLKNAND2HSV0 U32074 ( .A1(n28482), .A2(n28481), .ZN(n28483) );
  OAI21HSV2 U32075 ( .A1(n28481), .A2(n28482), .B(n28483), .ZN(n28484) );
  NAND2HSV0 U32076 ( .A1(n57818), .A2(n58272), .ZN(n28485) );
  NAND2HSV2 U32077 ( .A1(n28485), .A2(n28484), .ZN(n28486) );
  OAI21HSV2 U32078 ( .A1(n28484), .A2(n28485), .B(n28486), .ZN(n28487) );
  NAND2HSV0 U32079 ( .A1(n57646), .A2(n58186), .ZN(n28488) );
  CLKNAND2HSV0 U32080 ( .A1(n28488), .A2(n28487), .ZN(n28489) );
  OAI21HSV2 U32081 ( .A1(n28487), .A2(n28488), .B(n28489), .ZN(n58187) );
  CLKNHSV0 U32082 ( .I(n47971), .ZN(n28490) );
  NAND2HSV0 U32083 ( .A1(n47970), .A2(n28490), .ZN(n28491) );
  OAI211HSV0 U32084 ( .A1(n28490), .A2(n47970), .B(n28491), .C(n44369), .ZN(
        n28492) );
  NAND2HSV0 U32085 ( .A1(n28492), .A2(poh6[17]), .ZN(n28493) );
  OAI21HSV2 U32086 ( .A1(poh6[17]), .A2(n28492), .B(n28493), .ZN(po[18]) );
  AOI21HSV0 U32087 ( .A1(n58658), .A2(n58611), .B(n46816), .ZN(n28494) );
  AO31HSV2 U32088 ( .A1(n58658), .A2(n58611), .A3(n46816), .B(n28494), .Z(
        n28495) );
  NAND2HSV0 U32089 ( .A1(n53109), .A2(n58812), .ZN(n28496) );
  CLKNAND2HSV0 U32090 ( .A1(n28496), .A2(n28495), .ZN(n28497) );
  OAI21HSV0 U32091 ( .A1(n28495), .A2(n28496), .B(n28497), .ZN(n28498) );
  NAND2HSV0 U32092 ( .A1(n53172), .A2(n58572), .ZN(n28499) );
  CLKNAND2HSV0 U32093 ( .A1(n28499), .A2(n28498), .ZN(n28500) );
  OAI21HSV0 U32094 ( .A1(n28498), .A2(n28499), .B(n28500), .ZN(n28501) );
  NAND2HSV0 U32095 ( .A1(n58657), .A2(\pe6/got [12]), .ZN(n28502) );
  CLKNAND2HSV0 U32096 ( .A1(n28502), .A2(n28501), .ZN(n28503) );
  OAI21HSV0 U32097 ( .A1(n28501), .A2(n28502), .B(n28503), .ZN(n28504) );
  NAND2HSV0 U32098 ( .A1(n58576), .A2(n58811), .ZN(n28505) );
  CLKNAND2HSV0 U32099 ( .A1(n28505), .A2(n28504), .ZN(n28506) );
  OAI21HSV0 U32100 ( .A1(n28504), .A2(n28505), .B(n28506), .ZN(n28507) );
  CLKNAND2HSV0 U32101 ( .A1(n49741), .A2(n59169), .ZN(n28508) );
  CLKNAND2HSV0 U32102 ( .A1(n28508), .A2(n28507), .ZN(n28509) );
  OAI21HSV0 U32103 ( .A1(n28507), .A2(n28508), .B(n28509), .ZN(n28510) );
  NAND2HSV0 U32104 ( .A1(n59167), .A2(\pe6/got [15]), .ZN(n28511) );
  CLKNAND2HSV0 U32105 ( .A1(n28511), .A2(n28510), .ZN(n28512) );
  OAI21HSV0 U32106 ( .A1(n28513), .A2(n28514), .B(n28515), .ZN(\pe6/poht [16])
         );
  NAND2HSV0 U32107 ( .A1(n36924), .A2(n59359), .ZN(n28516) );
  NAND2HSV0 U32108 ( .A1(n28516), .A2(n51011), .ZN(n28517) );
  OAI21HSV0 U32109 ( .A1(n51011), .A2(n28516), .B(n28517), .ZN(n28518) );
  NAND2HSV0 U32110 ( .A1(n52726), .A2(n55946), .ZN(n28519) );
  NAND2HSV0 U32111 ( .A1(n28519), .A2(n28518), .ZN(n28520) );
  OAI21HSV0 U32112 ( .A1(n28518), .A2(n28519), .B(n28520), .ZN(n60085) );
  XOR2HSV0 U32113 ( .A1(n47138), .A2(n47137), .Z(n28521) );
  AOI21HSV0 U32114 ( .A1(n47056), .A2(n47268), .B(n28521), .ZN(n28522) );
  AO31HSV0 U32115 ( .A1(n47056), .A2(n47268), .A3(n28521), .B(n28522), .Z(
        n28523) );
  NAND2HSV0 U32116 ( .A1(n51227), .A2(n45816), .ZN(n28524) );
  CLKNAND2HSV0 U32117 ( .A1(n28524), .A2(n28523), .ZN(n28525) );
  OAI21HSV0 U32118 ( .A1(n28523), .A2(n28524), .B(n28525), .ZN(n28526) );
  NAND2HSV0 U32119 ( .A1(n29779), .A2(\pe5/got [23]), .ZN(n28527) );
  NAND2HSV0 U32120 ( .A1(n37631), .A2(n59580), .ZN(n28529) );
  CLKNAND2HSV0 U32121 ( .A1(n28529), .A2(n28528), .ZN(n28530) );
  OAI21HSV0 U32122 ( .A1(n28528), .A2(n28529), .B(n28530), .ZN(n28531) );
  NAND2HSV0 U32123 ( .A1(n37630), .A2(n48886), .ZN(n28532) );
  CLKNAND2HSV0 U32124 ( .A1(n28532), .A2(n28531), .ZN(n28533) );
  OAI21HSV0 U32125 ( .A1(n28531), .A2(n28532), .B(n28533), .ZN(\pe5/poht [7])
         );
  XOR2HSV0 U32126 ( .A1(n51794), .A2(n51793), .Z(n28534) );
  CLKNAND2HSV0 U32127 ( .A1(n28535), .A2(n28534), .ZN(n28536) );
  OAI21HSV0 U32128 ( .A1(n28534), .A2(n28535), .B(n28536), .ZN(n28537) );
  NAND2HSV0 U32129 ( .A1(n25831), .A2(n52051), .ZN(n28538) );
  CLKNAND2HSV0 U32130 ( .A1(n28538), .A2(n28537), .ZN(n28539) );
  OAI21HSV0 U32131 ( .A1(n28537), .A2(n28538), .B(n28539), .ZN(n28540) );
  OAI21HSV2 U32132 ( .A1(n28543), .A2(n28544), .B(n28545), .ZN(n28546) );
  NAND2HSV0 U32133 ( .A1(n44712), .A2(n52558), .ZN(n28547) );
  CLKNAND2HSV0 U32134 ( .A1(n28547), .A2(n28546), .ZN(n28548) );
  OAI21HSV0 U32135 ( .A1(n28546), .A2(n28547), .B(n28548), .ZN(\pe2/poht [14])
         );
  NAND2HSV0 U32136 ( .A1(n59766), .A2(n47997), .ZN(n28549) );
  NAND2HSV0 U32137 ( .A1(n28549), .A2(n47998), .ZN(n28550) );
  OAI21HSV0 U32138 ( .A1(n47998), .A2(n28549), .B(n28550), .ZN(n60098) );
  OAI22HSV0 U32139 ( .A1(n32878), .A2(n46853), .B1(n59105), .B2(n32589), .ZN(
        n28551) );
  OAI21HSV0 U32140 ( .A1(n35739), .A2(n32590), .B(n28551), .ZN(n28552) );
  CLKNAND2HSV0 U32141 ( .A1(n28552), .A2(n32591), .ZN(n28553) );
  OAI21HSV0 U32142 ( .A1(n28552), .A2(n32591), .B(n28553), .ZN(n32592) );
  XOR2HSV0 U32143 ( .A1(n35774), .A2(n35773), .Z(n28554) );
  AOI21HSV0 U32144 ( .A1(n58715), .A2(n58815), .B(n28554), .ZN(n28555) );
  AO31HSV2 U32145 ( .A1(n58715), .A2(n58815), .A3(n28554), .B(n28555), .Z(
        n28556) );
  NAND2HSV0 U32146 ( .A1(n35722), .A2(n35922), .ZN(n28557) );
  CLKNAND2HSV0 U32147 ( .A1(n28557), .A2(n28556), .ZN(n28558) );
  OAI21HSV0 U32148 ( .A1(n28556), .A2(n28557), .B(n28558), .ZN(n28559) );
  CLKNAND2HSV0 U32149 ( .A1(n46818), .A2(n59034), .ZN(n28560) );
  CLKNAND2HSV0 U32150 ( .A1(n28560), .A2(n28559), .ZN(n28561) );
  OAI21HSV0 U32151 ( .A1(n28559), .A2(n28560), .B(n28561), .ZN(n28562) );
  NAND2HSV0 U32152 ( .A1(n36105), .A2(n59328), .ZN(n28563) );
  CLKNAND2HSV0 U32153 ( .A1(n28563), .A2(n28562), .ZN(n28564) );
  OAI21HSV0 U32154 ( .A1(n28562), .A2(n28563), .B(n28564), .ZN(n28565) );
  NAND2HSV0 U32155 ( .A1(n59032), .A2(n59175), .ZN(n28566) );
  CLKNAND2HSV0 U32156 ( .A1(n28566), .A2(n28565), .ZN(n28567) );
  OAI21HSV0 U32157 ( .A1(n28565), .A2(n28566), .B(n28567), .ZN(n28568) );
  NAND2HSV0 U32158 ( .A1(n59174), .A2(n35898), .ZN(n28569) );
  CLKNAND2HSV0 U32159 ( .A1(n28569), .A2(n28568), .ZN(n28570) );
  OAI21HSV0 U32160 ( .A1(n28568), .A2(n28569), .B(n28570), .ZN(n28571) );
  NAND2HSV0 U32161 ( .A1(n32970), .A2(n35775), .ZN(n28572) );
  CLKNAND2HSV0 U32162 ( .A1(n28572), .A2(n28571), .ZN(n28573) );
  OAI21HSV2 U32163 ( .A1(n28571), .A2(n28572), .B(n28573), .ZN(n28574) );
  NAND2HSV0 U32164 ( .A1(n31710), .A2(n35721), .ZN(n28575) );
  CLKNAND2HSV0 U32165 ( .A1(n28575), .A2(n28574), .ZN(n28576) );
  OAI21HSV0 U32166 ( .A1(n28574), .A2(n28575), .B(n28576), .ZN(n35776) );
  XOR2HSV0 U32167 ( .A1(n33974), .A2(n33975), .Z(n28577) );
  XOR2HSV0 U32168 ( .A1(n33957), .A2(n33956), .Z(n28578) );
  XOR2HSV0 U32169 ( .A1(n28577), .A2(n28578), .Z(n28579) );
  AOI21HSV0 U32170 ( .A1(n33976), .A2(n57753), .B(n28579), .ZN(n28580) );
  AO31HSV0 U32171 ( .A1(n33976), .A2(n57753), .A3(n28579), .B(n28580), .Z(
        n28581) );
  XOR2HSV0 U32172 ( .A1(n33955), .A2(n28581), .Z(n28582) );
  NAND2HSV0 U32173 ( .A1(n35340), .A2(n59602), .ZN(n28583) );
  CLKNAND2HSV0 U32174 ( .A1(n28583), .A2(n28582), .ZN(n28584) );
  OAI21HSV0 U32175 ( .A1(n28582), .A2(n28583), .B(n28584), .ZN(n28585) );
  NAND2HSV0 U32176 ( .A1(\pe4/got [20]), .A2(n47733), .ZN(n28586) );
  NAND2HSV2 U32177 ( .A1(n28586), .A2(n28585), .ZN(n28587) );
  OAI21HSV2 U32178 ( .A1(n28585), .A2(n28586), .B(n28587), .ZN(n28588) );
  NAND2HSV0 U32179 ( .A1(n57526), .A2(n59370), .ZN(n28589) );
  NAND2HSV2 U32180 ( .A1(n28589), .A2(n28588), .ZN(n28590) );
  OAI21HSV2 U32181 ( .A1(n28588), .A2(n28589), .B(n28590), .ZN(n28591) );
  NAND2HSV0 U32182 ( .A1(n34351), .A2(n57530), .ZN(n28592) );
  NAND2HSV2 U32183 ( .A1(n28592), .A2(n28591), .ZN(n28593) );
  OAI21HSV2 U32184 ( .A1(n28591), .A2(n28592), .B(n28593), .ZN(n28594) );
  NAND2HSV0 U32185 ( .A1(n59369), .A2(n34595), .ZN(n28595) );
  NAND2HSV0 U32186 ( .A1(n28595), .A2(n28594), .ZN(n28596) );
  OAI21HSV0 U32187 ( .A1(n28594), .A2(n28595), .B(n28596), .ZN(n33978) );
  NAND2HSV0 U32188 ( .A1(n51919), .A2(n53005), .ZN(n28598) );
  NOR2HSV0 U32189 ( .A1(n51704), .A2(n51703), .ZN(n28599) );
  AOI21HSV2 U32190 ( .A1(n28598), .A2(n51984), .B(n28599), .ZN(n51706) );
  INOR2HSV0 U32191 ( .A1(\pe1/ti_7t [28]), .B1(n44649), .ZN(n45781) );
  XOR2HSV0 U32192 ( .A1(n52598), .A2(n52599), .Z(n28600) );
  XOR2HSV0 U32193 ( .A1(n52589), .A2(n52588), .Z(n28601) );
  XOR2HSV0 U32194 ( .A1(n28600), .A2(n28601), .Z(n28602) );
  XOR2HSV0 U32195 ( .A1(n52614), .A2(n52615), .Z(n28603) );
  XOR2HSV0 U32196 ( .A1(n52606), .A2(n52605), .Z(n28604) );
  XOR2HSV0 U32197 ( .A1(n28603), .A2(n28604), .Z(n28605) );
  XOR2HSV0 U32198 ( .A1(n52628), .A2(n52629), .Z(n28606) );
  XOR2HSV0 U32199 ( .A1(n52617), .A2(n52616), .Z(n28607) );
  XOR2HSV0 U32200 ( .A1(n28606), .A2(n28607), .Z(n28608) );
  XOR2HSV0 U32201 ( .A1(n28608), .A2(n52637), .Z(n28609) );
  XOR2HSV0 U32202 ( .A1(n28605), .A2(n52638), .Z(n28610) );
  XOR2HSV0 U32203 ( .A1(n28609), .A2(n28610), .Z(n28611) );
  XOR2HSV0 U32204 ( .A1(n28602), .A2(n28611), .Z(n28612) );
  NAND2HSV0 U32205 ( .A1(n39654), .A2(n51362), .ZN(n28613) );
  CLKNAND2HSV0 U32206 ( .A1(n28613), .A2(n28612), .ZN(n28614) );
  OAI21HSV0 U32207 ( .A1(n28612), .A2(n28613), .B(n28614), .ZN(n28615) );
  CLKNAND2HSV0 U32208 ( .A1(n51161), .A2(n47338), .ZN(n28616) );
  CLKNAND2HSV0 U32209 ( .A1(n28616), .A2(n28615), .ZN(n28617) );
  OAI21HSV0 U32210 ( .A1(n28615), .A2(n28616), .B(n28617), .ZN(n28618) );
  NAND2HSV0 U32211 ( .A1(n52580), .A2(n52579), .ZN(n28619) );
  CLKNAND2HSV0 U32212 ( .A1(n28619), .A2(n28618), .ZN(n28620) );
  OAI21HSV0 U32213 ( .A1(n28618), .A2(n28619), .B(n28620), .ZN(n28621) );
  NAND2HSV0 U32214 ( .A1(n52577), .A2(n52578), .ZN(n28622) );
  CLKNAND2HSV0 U32215 ( .A1(n28622), .A2(n28621), .ZN(n28623) );
  OAI21HSV0 U32216 ( .A1(n28621), .A2(n28622), .B(n28623), .ZN(n28624) );
  NAND2HSV0 U32217 ( .A1(n52576), .A2(n29770), .ZN(n28625) );
  CLKNAND2HSV0 U32218 ( .A1(n28625), .A2(n28624), .ZN(n28626) );
  OAI21HSV2 U32219 ( .A1(n28624), .A2(n28625), .B(n28626), .ZN(n28627) );
  NAND2HSV0 U32220 ( .A1(n51200), .A2(n52575), .ZN(n28628) );
  NAND2HSV2 U32221 ( .A1(n28628), .A2(n28627), .ZN(n28629) );
  OAI21HSV2 U32222 ( .A1(n28627), .A2(n28628), .B(n28629), .ZN(n28630) );
  NAND2HSV0 U32223 ( .A1(n52574), .A2(n52573), .ZN(n28631) );
  CLKNAND2HSV0 U32224 ( .A1(n28631), .A2(n28630), .ZN(n28632) );
  OAI21HSV0 U32225 ( .A1(n28630), .A2(n28631), .B(n28632), .ZN(n52639) );
  XOR2HSV0 U32226 ( .A1(n40799), .A2(n40800), .Z(n28633) );
  XOR2HSV0 U32227 ( .A1(n40795), .A2(n40794), .Z(n28634) );
  XOR2HSV0 U32228 ( .A1(n28633), .A2(n28634), .Z(n28635) );
  CLKNHSV0 U32229 ( .I(n40827), .ZN(n28636) );
  AO22HSV2 U32230 ( .A1(n40898), .A2(\pe1/bq[23] ), .B1(\pe1/bq[18] ), .B2(
        n25226), .Z(n28637) );
  CLKNAND2HSV0 U32231 ( .A1(n42099), .A2(n40897), .ZN(n28638) );
  CLKNAND2HSV0 U32232 ( .A1(n28638), .A2(n53671), .ZN(n28639) );
  OAI21HSV0 U32233 ( .A1(n53671), .A2(n28638), .B(n28639), .ZN(n28640) );
  OAI21HSV0 U32234 ( .A1(n42214), .A2(n41363), .B(n28637), .ZN(n28641) );
  CLKNAND2HSV0 U32235 ( .A1(n28641), .A2(n28640), .ZN(n28642) );
  OAI21HSV0 U32236 ( .A1(n28641), .A2(n28640), .B(n28642), .ZN(n28643) );
  NAND2HSV0 U32237 ( .A1(n41676), .A2(n41248), .ZN(n28644) );
  CLKNAND2HSV0 U32238 ( .A1(n28644), .A2(n28643), .ZN(n28645) );
  OAI21HSV0 U32239 ( .A1(n28643), .A2(n28644), .B(n28645), .ZN(n28646) );
  XOR2HSV0 U32240 ( .A1(n40791), .A2(n40790), .Z(n28647) );
  XOR2HSV0 U32241 ( .A1(n28646), .A2(n28647), .Z(n28648) );
  MUX2NHSV0 U32242 ( .I0(n28636), .I1(n40827), .S(n28648), .ZN(n28649) );
  XOR2HSV0 U32243 ( .A1(n40796), .A2(n28635), .Z(n28650) );
  XOR2HSV0 U32244 ( .A1(n28649), .A2(n28650), .Z(n28651) );
  CLKNAND2HSV0 U32245 ( .A1(n40886), .A2(n41549), .ZN(n28652) );
  CLKNAND2HSV0 U32246 ( .A1(n28652), .A2(n28651), .ZN(n28653) );
  OAI21HSV0 U32247 ( .A1(n28651), .A2(n28652), .B(n28653), .ZN(n28654) );
  NAND2HSV0 U32248 ( .A1(n41387), .A2(n40910), .ZN(n28655) );
  CLKNAND2HSV0 U32249 ( .A1(n28655), .A2(n28654), .ZN(n28656) );
  OAI21HSV0 U32250 ( .A1(n28654), .A2(n28655), .B(n28656), .ZN(n28657) );
  NAND2HSV0 U32251 ( .A1(n41144), .A2(\pe1/got [23]), .ZN(n28658) );
  CLKNAND2HSV0 U32252 ( .A1(n28658), .A2(n28657), .ZN(n28659) );
  OAI21HSV0 U32253 ( .A1(n28657), .A2(n28658), .B(n28659), .ZN(n28660) );
  CLKNAND2HSV0 U32254 ( .A1(n40913), .A2(n40917), .ZN(n28661) );
  CLKNAND2HSV0 U32255 ( .A1(n28661), .A2(n28660), .ZN(n28662) );
  OAI21HSV0 U32256 ( .A1(n28660), .A2(n28661), .B(n28662), .ZN(n28663) );
  NAND2HSV0 U32257 ( .A1(n41201), .A2(n42431), .ZN(n28664) );
  CLKNAND2HSV0 U32258 ( .A1(n28664), .A2(n28663), .ZN(n28665) );
  OAI21HSV0 U32259 ( .A1(n28663), .A2(n28664), .B(n28665), .ZN(n28666) );
  NAND2HSV0 U32260 ( .A1(n41689), .A2(n41929), .ZN(n28667) );
  CLKNAND2HSV0 U32261 ( .A1(n28667), .A2(n28666), .ZN(n28668) );
  OAI21HSV2 U32262 ( .A1(n28666), .A2(n28667), .B(n28668), .ZN(n40814) );
  NAND3HSV4 U32263 ( .A1(n36260), .A2(n36259), .A3(n36258), .ZN(n36363) );
  CLKNHSV0 U32264 ( .I(n46566), .ZN(n28669) );
  XOR2HSV0 U32265 ( .A1(n57815), .A2(n57814), .Z(n28670) );
  XOR2HSV0 U32266 ( .A1(n57813), .A2(n28670), .Z(n28671) );
  CLKNAND2HSV0 U32267 ( .A1(n28672), .A2(n28671), .ZN(n28673) );
  OAI21HSV0 U32268 ( .A1(n28671), .A2(n28672), .B(n28673), .ZN(n28674) );
  NAND2HSV0 U32269 ( .A1(n59378), .A2(n58206), .ZN(n28675) );
  CLKNAND2HSV0 U32270 ( .A1(n28675), .A2(n28674), .ZN(n28676) );
  OAI21HSV0 U32271 ( .A1(n28674), .A2(n28675), .B(n28676), .ZN(n28677) );
  NAND2HSV0 U32272 ( .A1(n58246), .A2(n25284), .ZN(n28678) );
  CLKNAND2HSV0 U32273 ( .A1(n28678), .A2(n28677), .ZN(n28679) );
  OAI21HSV0 U32274 ( .A1(n28677), .A2(n28678), .B(n28679), .ZN(n28680) );
  NAND2HSV0 U32275 ( .A1(n58184), .A2(n57984), .ZN(n28681) );
  CLKNAND2HSV0 U32276 ( .A1(n28681), .A2(n28680), .ZN(n28682) );
  OAI21HSV0 U32277 ( .A1(n28680), .A2(n28681), .B(n28682), .ZN(n28683) );
  CLKNAND2HSV0 U32278 ( .A1(n58036), .A2(n57817), .ZN(n28684) );
  CLKNAND2HSV0 U32279 ( .A1(n28684), .A2(n28683), .ZN(n28685) );
  OAI21HSV0 U32280 ( .A1(n28683), .A2(n28684), .B(n28685), .ZN(n28686) );
  CLKNAND2HSV0 U32281 ( .A1(n57818), .A2(n34733), .ZN(n28687) );
  CLKNAND2HSV0 U32282 ( .A1(n28687), .A2(n28686), .ZN(n28688) );
  OAI21HSV0 U32283 ( .A1(n28686), .A2(n28687), .B(n28688), .ZN(n28689) );
  NAND2HSV0 U32284 ( .A1(n59935), .A2(n57177), .ZN(n28690) );
  CLKNAND2HSV0 U32285 ( .A1(n28690), .A2(n28689), .ZN(n28691) );
  OAI21HSV0 U32286 ( .A1(n28689), .A2(n28690), .B(n28691), .ZN(n28692) );
  NAND2HSV0 U32287 ( .A1(n58154), .A2(n59663), .ZN(n28693) );
  CLKNAND2HSV0 U32288 ( .A1(n28693), .A2(n28692), .ZN(n28694) );
  OAI21HSV0 U32289 ( .A1(n28692), .A2(n28693), .B(n28694), .ZN(n28695) );
  CLKNAND2HSV0 U32290 ( .A1(n58110), .A2(n57819), .ZN(n28696) );
  CLKNAND2HSV0 U32291 ( .A1(n28696), .A2(n28695), .ZN(n28697) );
  OAI21HSV2 U32292 ( .A1(n28695), .A2(n28696), .B(n28697), .ZN(n28698) );
  NAND2HSV0 U32293 ( .A1(n57960), .A2(n58153), .ZN(n28699) );
  CLKNAND2HSV0 U32294 ( .A1(n28699), .A2(n28698), .ZN(n28700) );
  OAI21HSV2 U32295 ( .A1(n28698), .A2(n28699), .B(n28700), .ZN(n28701) );
  NAND2HSV0 U32296 ( .A1(n57889), .A2(n57820), .ZN(n28702) );
  CLKNAND2HSV0 U32297 ( .A1(n28702), .A2(n28701), .ZN(n28703) );
  OAI21HSV2 U32298 ( .A1(n28701), .A2(n28702), .B(n28703), .ZN(n28704) );
  CLKNAND2HSV0 U32299 ( .A1(n58052), .A2(n57310), .ZN(n28705) );
  CLKNAND2HSV0 U32300 ( .A1(n28705), .A2(n28704), .ZN(n28706) );
  OAI21HSV0 U32301 ( .A1(n28704), .A2(n28705), .B(n28706), .ZN(n57821) );
  XOR2HSV0 U32302 ( .A1(n49311), .A2(n49308), .Z(n28707) );
  XOR2HSV0 U32303 ( .A1(n49307), .A2(n49309), .Z(n28708) );
  XOR2HSV0 U32304 ( .A1(n28707), .A2(n28708), .Z(n28709) );
  XOR2HSV0 U32305 ( .A1(n49310), .A2(n28709), .Z(n28710) );
  NAND2HSV0 U32306 ( .A1(n56855), .A2(n45636), .ZN(n28711) );
  CLKNAND2HSV0 U32307 ( .A1(n28711), .A2(n28710), .ZN(n28712) );
  OAI21HSV0 U32308 ( .A1(n28710), .A2(n28711), .B(n28712), .ZN(n28713) );
  NAND2HSV0 U32309 ( .A1(n55912), .A2(n56266), .ZN(n28714) );
  CLKNAND2HSV0 U32310 ( .A1(n28714), .A2(n28713), .ZN(n28715) );
  OAI21HSV0 U32311 ( .A1(n28713), .A2(n28714), .B(n28715), .ZN(n28716) );
  NAND2HSV0 U32312 ( .A1(n56559), .A2(n53228), .ZN(n28717) );
  CLKNAND2HSV0 U32313 ( .A1(n28717), .A2(n28716), .ZN(n28718) );
  OAI21HSV0 U32314 ( .A1(n28716), .A2(n28717), .B(n28718), .ZN(n28719) );
  NAND2HSV0 U32315 ( .A1(n56495), .A2(n56662), .ZN(n28720) );
  CLKNAND2HSV0 U32316 ( .A1(n28720), .A2(n28719), .ZN(n28721) );
  OAI21HSV0 U32317 ( .A1(n28719), .A2(n28720), .B(n28721), .ZN(n28722) );
  NAND2HSV0 U32318 ( .A1(n56066), .A2(n56342), .ZN(n28723) );
  CLKNAND2HSV0 U32319 ( .A1(n28723), .A2(n28722), .ZN(n28724) );
  OAI21HSV0 U32320 ( .A1(n28722), .A2(n28723), .B(n28724), .ZN(n28725) );
  NAND2HSV0 U32321 ( .A1(n56618), .A2(n56737), .ZN(n28726) );
  CLKNAND2HSV0 U32322 ( .A1(n28726), .A2(n28725), .ZN(n28727) );
  OAI21HSV0 U32323 ( .A1(n28725), .A2(n28726), .B(n28727), .ZN(n28728) );
  NAND2HSV0 U32324 ( .A1(n56421), .A2(n56622), .ZN(n28729) );
  CLKNAND2HSV0 U32325 ( .A1(n28729), .A2(n28728), .ZN(n28730) );
  OAI21HSV2 U32326 ( .A1(n28728), .A2(n28729), .B(n28730), .ZN(n28731) );
  NAND2HSV0 U32327 ( .A1(\pe3/got [14]), .A2(n50757), .ZN(n28732) );
  CLKNAND2HSV0 U32328 ( .A1(n28732), .A2(n28731), .ZN(n28733) );
  OAI21HSV0 U32329 ( .A1(n28731), .A2(n28732), .B(n28733), .ZN(n49312) );
  NOR2HSV0 U32330 ( .A1(n51439), .A2(n51438), .ZN(n28734) );
  NOR2HSV2 U32331 ( .A1(n51440), .A2(n28734), .ZN(n28735) );
  AOI211HSV1 U32332 ( .A1(n51440), .A2(n28734), .B(n32047), .C(n28735), .ZN(
        n28736) );
  XOR2HSV0 U32333 ( .A1(poh6[8]), .A2(n28736), .Z(po[9]) );
  OAI21HSV0 U32334 ( .A1(n46560), .A2(n46559), .B(n46558), .ZN(n28737) );
  CLKNAND2HSV0 U32335 ( .A1(n28737), .A2(n46562), .ZN(n28738) );
  OAI21HSV0 U32336 ( .A1(n28737), .A2(n46562), .B(n28738), .ZN(n60022) );
  XOR2HSV0 U32337 ( .A1(n46149), .A2(n46148), .Z(n28739) );
  NAND2HSV0 U32338 ( .A1(n58480), .A2(n58816), .ZN(n28740) );
  CLKNAND2HSV0 U32339 ( .A1(n28740), .A2(n28739), .ZN(n28741) );
  OAI21HSV0 U32340 ( .A1(n28739), .A2(n28740), .B(n28741), .ZN(n28742) );
  NAND2HSV0 U32341 ( .A1(n58716), .A2(n58423), .ZN(n28743) );
  CLKNAND2HSV0 U32342 ( .A1(n28743), .A2(n28742), .ZN(n28744) );
  OAI21HSV0 U32343 ( .A1(n28742), .A2(n28743), .B(n28744), .ZN(n28745) );
  CLKNAND2HSV0 U32344 ( .A1(n28746), .A2(n28745), .ZN(n28747) );
  OAI21HSV0 U32345 ( .A1(n28745), .A2(n28746), .B(n28747), .ZN(n28748) );
  NAND2HSV0 U32346 ( .A1(n58809), .A2(n58400), .ZN(n28749) );
  CLKNAND2HSV0 U32347 ( .A1(n28749), .A2(n28748), .ZN(n28750) );
  OAI21HSV0 U32348 ( .A1(n28748), .A2(n28749), .B(n28750), .ZN(n28751) );
  CLKNAND2HSV0 U32349 ( .A1(n58576), .A2(n58399), .ZN(n28752) );
  CLKNAND2HSV0 U32350 ( .A1(n28752), .A2(n28751), .ZN(n28753) );
  OAI21HSV0 U32351 ( .A1(n28751), .A2(n28752), .B(n28753), .ZN(n28754) );
  CLKNAND2HSV0 U32352 ( .A1(n36109), .A2(n58575), .ZN(n28755) );
  CLKNAND2HSV0 U32353 ( .A1(n28755), .A2(n28754), .ZN(n28756) );
  OAI21HSV0 U32354 ( .A1(n28754), .A2(n28755), .B(n28756), .ZN(n28757) );
  CLKNAND2HSV0 U32355 ( .A1(n28758), .A2(n28757), .ZN(n28759) );
  OAI21HSV0 U32356 ( .A1(n28757), .A2(n28758), .B(n28759), .ZN(n28760) );
  OAI21HSV0 U32357 ( .A1(n28760), .A2(n28761), .B(n28762), .ZN(\pe6/poht [23])
         );
  XOR2HSV0 U32358 ( .A1(n51226), .A2(n51225), .Z(n28763) );
  AOI21HSV0 U32359 ( .A1(n51156), .A2(n52565), .B(n28763), .ZN(n28764) );
  AO31HSV2 U32360 ( .A1(n51156), .A2(n52565), .A3(n28763), .B(n28764), .Z(
        n28765) );
  NAND2HSV0 U32361 ( .A1(n51227), .A2(n52566), .ZN(n28766) );
  CLKNAND2HSV0 U32362 ( .A1(n28766), .A2(n28765), .ZN(n28767) );
  OAI21HSV0 U32363 ( .A1(n28765), .A2(n28766), .B(n28767), .ZN(n28768) );
  NAND2HSV0 U32364 ( .A1(n51014), .A2(n37556), .ZN(n28769) );
  CLKNAND2HSV0 U32365 ( .A1(n28769), .A2(n28768), .ZN(n28770) );
  OAI21HSV0 U32366 ( .A1(n28768), .A2(n28769), .B(n28770), .ZN(n28771) );
  NAND2HSV0 U32367 ( .A1(n51155), .A2(n45816), .ZN(n28772) );
  CLKNAND2HSV0 U32368 ( .A1(n28772), .A2(n28771), .ZN(n28773) );
  OAI21HSV0 U32369 ( .A1(n28771), .A2(n28772), .B(n28773), .ZN(n28774) );
  NAND2HSV0 U32370 ( .A1(n29777), .A2(n51228), .ZN(n28775) );
  CLKNAND2HSV0 U32371 ( .A1(n28775), .A2(n28774), .ZN(n28776) );
  OAI21HSV0 U32372 ( .A1(n28774), .A2(n28775), .B(n28776), .ZN(n28777) );
  NAND2HSV0 U32373 ( .A1(n52668), .A2(n47267), .ZN(n28778) );
  CLKNAND2HSV0 U32374 ( .A1(n28778), .A2(n28777), .ZN(n28779) );
  OAI21HSV2 U32375 ( .A1(n28777), .A2(n28778), .B(n28779), .ZN(n28780) );
  NAND2HSV0 U32376 ( .A1(n29771), .A2(n59948), .ZN(n28781) );
  CLKNAND2HSV0 U32377 ( .A1(n28781), .A2(n28780), .ZN(n28782) );
  OAI21HSV0 U32378 ( .A1(n28780), .A2(n28781), .B(n28782), .ZN(\pe5/poht [9])
         );
  XOR2HSV0 U32379 ( .A1(n50925), .A2(n50924), .Z(n28783) );
  XOR2HSV0 U32380 ( .A1(n50927), .A2(n28783), .Z(n28784) );
  CLKNAND2HSV0 U32381 ( .A1(n28785), .A2(n28784), .ZN(n28786) );
  OAI21HSV0 U32382 ( .A1(n28784), .A2(n28785), .B(n28786), .ZN(n28787) );
  NAND2HSV0 U32383 ( .A1(n52048), .A2(n52855), .ZN(n28788) );
  CLKNAND2HSV0 U32384 ( .A1(n28788), .A2(n28787), .ZN(n28789) );
  OAI21HSV0 U32385 ( .A1(n28787), .A2(n28788), .B(n28789), .ZN(n28790) );
  NAND2HSV0 U32386 ( .A1(n52047), .A2(n51686), .ZN(n28791) );
  CLKNAND2HSV0 U32387 ( .A1(n28791), .A2(n28790), .ZN(n28792) );
  NAND2HSV0 U32388 ( .A1(n52890), .A2(n52558), .ZN(n28797) );
  INAND3HSV0 U32389 ( .A1(n47978), .B1(n25850), .B2(n47980), .ZN(n28799) );
  NAND2HSV0 U32390 ( .A1(n28799), .A2(n47982), .ZN(n28800) );
  OAI21HSV0 U32391 ( .A1(n47982), .A2(n28799), .B(n28800), .ZN(n60096) );
  NAND2HSV0 U32392 ( .A1(n53014), .A2(\pe2/pvq [26]), .ZN(n28801) );
  NAND2HSV0 U32393 ( .A1(n28801), .A2(\pe2/phq [26]), .ZN(n28802) );
  OAI21HSV2 U32394 ( .A1(\pe2/phq [26]), .A2(n28801), .B(n28802), .ZN(n44052)
         );
  NAND2HSV0 U32395 ( .A1(n34240), .A2(n33533), .ZN(n28803) );
  AOI21HSV0 U32396 ( .A1(n33615), .A2(n33631), .B(n28803), .ZN(n28804) );
  AO31HSV0 U32397 ( .A1(n33615), .A2(n33631), .A3(n28803), .B(n28804), .Z(
        n33488) );
  NAND2HSV0 U32398 ( .A1(n33474), .A2(n33103), .ZN(n28805) );
  AOI21HSV0 U32399 ( .A1(n33248), .A2(n59523), .B(n28805), .ZN(n28806) );
  AO31HSV2 U32400 ( .A1(n33248), .A2(n59523), .A3(n28805), .B(n28806), .Z(
        n33207) );
  XOR2HSV0 U32401 ( .A1(n39663), .A2(n39662), .Z(n28807) );
  XOR2HSV0 U32402 ( .A1(n39661), .A2(n28807), .Z(n28808) );
  AOI21HSV0 U32403 ( .A1(n46974), .A2(n48748), .B(n28808), .ZN(n28809) );
  AO31HSV2 U32404 ( .A1(n46974), .A2(n48748), .A3(n28808), .B(n28809), .Z(
        n28810) );
  CLKNAND2HSV0 U32405 ( .A1(n50495), .A2(n31147), .ZN(n28811) );
  CLKNAND2HSV0 U32406 ( .A1(n28811), .A2(n28810), .ZN(n28812) );
  OAI21HSV0 U32407 ( .A1(n28810), .A2(n28811), .B(n28812), .ZN(n28813) );
  CLKNAND2HSV0 U32408 ( .A1(n47056), .A2(n39257), .ZN(n28814) );
  CLKNAND2HSV0 U32409 ( .A1(n28814), .A2(n28813), .ZN(n28815) );
  OAI21HSV0 U32410 ( .A1(n28813), .A2(n28814), .B(n28815), .ZN(n28816) );
  NAND2HSV0 U32411 ( .A1(n45816), .A2(n44694), .ZN(n28817) );
  CLKNAND2HSV0 U32412 ( .A1(n28817), .A2(n28816), .ZN(n28818) );
  OAI21HSV0 U32413 ( .A1(n28816), .A2(n28817), .B(n28818), .ZN(n28819) );
  NAND2HSV0 U32414 ( .A1(n37656), .A2(n45417), .ZN(n28820) );
  CLKNAND2HSV0 U32415 ( .A1(n28820), .A2(n28819), .ZN(n28821) );
  OAI21HSV0 U32416 ( .A1(n28819), .A2(n28820), .B(n28821), .ZN(n28822) );
  NAND2HSV0 U32417 ( .A1(n59517), .A2(n48744), .ZN(n28823) );
  CLKNAND2HSV0 U32418 ( .A1(n28823), .A2(n28822), .ZN(n28824) );
  OAI21HSV0 U32419 ( .A1(n28822), .A2(n28823), .B(n28824), .ZN(n28825) );
  CLKNAND2HSV0 U32420 ( .A1(n59882), .A2(n59948), .ZN(n28826) );
  CLKNAND2HSV0 U32421 ( .A1(n28826), .A2(n28825), .ZN(n28827) );
  OAI21HSV0 U32422 ( .A1(n28825), .A2(n28826), .B(n28827), .ZN(n28828) );
  CLKNAND2HSV0 U32423 ( .A1(n48743), .A2(n48746), .ZN(n28829) );
  CLKNAND2HSV0 U32424 ( .A1(n28829), .A2(n28828), .ZN(n28830) );
  OAI21HSV0 U32425 ( .A1(n28828), .A2(n28829), .B(n28830), .ZN(n28831) );
  NAND2HSV0 U32426 ( .A1(n37630), .A2(n40116), .ZN(n28832) );
  CLKNAND2HSV0 U32427 ( .A1(n28832), .A2(n28831), .ZN(n28833) );
  OAI21HSV0 U32428 ( .A1(n28831), .A2(n28832), .B(n28833), .ZN(n39665) );
  OAI22HSV0 U32429 ( .A1(n41425), .A2(n44705), .B1(n41650), .B2(n53553), .ZN(
        n28834) );
  OAI21HSV2 U32430 ( .A1(n41350), .A2(n41251), .B(n28834), .ZN(n41255) );
  NAND2HSV0 U32431 ( .A1(n48243), .A2(\pe5/bq[11] ), .ZN(n28835) );
  AOI21HSV0 U32432 ( .A1(n50444), .A2(n40210), .B(n28835), .ZN(n28836) );
  AO31HSV0 U32433 ( .A1(n50444), .A2(n40210), .A3(n28835), .B(n28836), .Z(
        n40211) );
  XOR2HSV0 U32434 ( .A1(n38488), .A2(n38487), .Z(n28837) );
  NAND2HSV0 U32435 ( .A1(\pe2/got [16]), .A2(n43950), .ZN(n28838) );
  NAND2HSV2 U32436 ( .A1(n28838), .A2(n28837), .ZN(n28839) );
  OAI21HSV0 U32437 ( .A1(n28837), .A2(n28838), .B(n28839), .ZN(n28840) );
  XOR2HSV0 U32438 ( .A1(n38496), .A2(n38497), .Z(n28841) );
  XOR2HSV0 U32439 ( .A1(n38491), .A2(n38490), .Z(n28842) );
  XOR2HSV0 U32440 ( .A1(n28841), .A2(n28842), .Z(n28843) );
  XOR2HSV0 U32441 ( .A1(n38500), .A2(n38501), .Z(n28844) );
  XOR2HSV0 U32442 ( .A1(n38507), .A2(n38506), .Z(n28845) );
  XOR2HSV0 U32443 ( .A1(n28844), .A2(n28845), .Z(n28846) );
  XOR2HSV0 U32444 ( .A1(n28840), .A2(n28843), .Z(n28847) );
  XOR2HSV0 U32445 ( .A1(n28846), .A2(n28847), .Z(n28848) );
  CLKNAND2HSV0 U32446 ( .A1(n38781), .A2(n38539), .ZN(n28849) );
  NAND2HSV2 U32447 ( .A1(n28849), .A2(n28848), .ZN(n28850) );
  OAI21HSV2 U32448 ( .A1(n28848), .A2(n28849), .B(n28850), .ZN(n28851) );
  OAI21HSV0 U32449 ( .A1(n38489), .A2(n53064), .B(n28851), .ZN(n28852) );
  OAI31HSV0 U32450 ( .A1(n38489), .A2(n28851), .A3(n53064), .B(n28852), .ZN(
        n28853) );
  NAND2HSV0 U32451 ( .A1(n44715), .A2(\pe2/got [19]), .ZN(n28854) );
  NAND2HSV0 U32452 ( .A1(n28854), .A2(n28853), .ZN(n28855) );
  OAI21HSV0 U32453 ( .A1(n28853), .A2(n28854), .B(n28855), .ZN(n28856) );
  NAND2HSV0 U32454 ( .A1(n38702), .A2(n39010), .ZN(n28857) );
  CLKNAND2HSV0 U32455 ( .A1(n28857), .A2(n28856), .ZN(n28858) );
  OAI21HSV2 U32456 ( .A1(n28856), .A2(n28857), .B(n28858), .ZN(n28859) );
  NAND2HSV0 U32457 ( .A1(n52167), .A2(n52053), .ZN(n28860) );
  CLKNAND2HSV0 U32458 ( .A1(n28860), .A2(n28859), .ZN(n28861) );
  OAI21HSV0 U32459 ( .A1(n28859), .A2(n28860), .B(n28861), .ZN(n38508) );
  AOI22HSV0 U32460 ( .A1(n59189), .A2(\pe6/bq[11] ), .B1(n50829), .B2(n58857), 
        .ZN(n28862) );
  IAO21HSV0 U32461 ( .A1(n50828), .A2(n53128), .B(n28862), .ZN(n50830) );
  OAI22HSV0 U32462 ( .A1(n40445), .A2(n45814), .B1(n53833), .B2(n48060), .ZN(
        n28863) );
  OAI21HSV0 U32463 ( .A1(n41075), .A2(n41630), .B(n28863), .ZN(n28864) );
  OAI22HSV0 U32464 ( .A1(n41076), .A2(n54973), .B1(n46629), .B2(n44703), .ZN(
        n28865) );
  OAI21HSV0 U32465 ( .A1(n41077), .A2(n54074), .B(n28865), .ZN(n28866) );
  CLKNAND2HSV0 U32466 ( .A1(n28866), .A2(n28864), .ZN(n28867) );
  OAI21HSV0 U32467 ( .A1(n28866), .A2(n28864), .B(n28867), .ZN(n28868) );
  NAND2HSV0 U32468 ( .A1(n41284), .A2(n41160), .ZN(n28869) );
  CLKNAND2HSV0 U32469 ( .A1(n28869), .A2(n28868), .ZN(n28870) );
  OAI21HSV2 U32470 ( .A1(n28868), .A2(n28869), .B(n28870), .ZN(n41078) );
  NAND2HSV0 U32471 ( .A1(n59165), .A2(n35898), .ZN(n28871) );
  NAND2HSV0 U32472 ( .A1(n35812), .A2(n59032), .ZN(n28872) );
  NAND2HSV0 U32473 ( .A1(n28872), .A2(n28871), .ZN(n28873) );
  OAI21HSV2 U32474 ( .A1(n28871), .A2(n28872), .B(n28873), .ZN(n32776) );
  INOR2HSV1 U32475 ( .A1(\pe1/ti_7t [9]), .B1(n41134), .ZN(n40671) );
  NAND2HSV0 U32476 ( .A1(n46672), .A2(\pe6/aot [17]), .ZN(n28874) );
  AOI21HSV0 U32477 ( .A1(n32740), .A2(n59045), .B(n28874), .ZN(n28875) );
  AO31HSV2 U32478 ( .A1(n59276), .A2(n59045), .A3(n28874), .B(n28875), .Z(
        n32374) );
  CLKNHSV0 U32479 ( .I(\pe4/phq [1]), .ZN(n28876) );
  INAND2HSV0 U32480 ( .A1(\pe1/ti_7t [13]), .B1(n41712), .ZN(n41229) );
  NOR2HSV0 U32481 ( .A1(n34221), .A2(n46581), .ZN(n28877) );
  XOR2HSV0 U32482 ( .A1(n56244), .A2(n56245), .Z(n28878) );
  XOR2HSV0 U32483 ( .A1(n56246), .A2(n56243), .Z(n28879) );
  XOR2HSV0 U32484 ( .A1(n28878), .A2(n28879), .Z(n28880) );
  NAND2HSV0 U32485 ( .A1(n59811), .A2(\pe3/got [8]), .ZN(n28881) );
  CLKNAND2HSV0 U32486 ( .A1(n28881), .A2(n28880), .ZN(n28882) );
  OAI21HSV0 U32487 ( .A1(n28880), .A2(n28881), .B(n28882), .ZN(n28883) );
  NAND2HSV0 U32488 ( .A1(n56624), .A2(n56495), .ZN(n28884) );
  CLKNAND2HSV0 U32489 ( .A1(n28884), .A2(n28883), .ZN(n28885) );
  OAI21HSV0 U32490 ( .A1(n28883), .A2(n28884), .B(n28885), .ZN(n28886) );
  NAND2HSV0 U32491 ( .A1(n56662), .A2(n56247), .ZN(n28887) );
  CLKNAND2HSV0 U32492 ( .A1(n28887), .A2(n28886), .ZN(n28888) );
  OAI21HSV0 U32493 ( .A1(n28886), .A2(n28887), .B(n28888), .ZN(n28889) );
  NAND2HSV0 U32494 ( .A1(n56562), .A2(n56176), .ZN(n28890) );
  CLKNAND2HSV0 U32495 ( .A1(n28890), .A2(n28889), .ZN(n28891) );
  OAI21HSV0 U32496 ( .A1(n28889), .A2(n28890), .B(n28891), .ZN(n28892) );
  NAND2HSV0 U32497 ( .A1(\pe3/got [13]), .A2(n56497), .ZN(n28893) );
  CLKNAND2HSV0 U32498 ( .A1(n28893), .A2(n28892), .ZN(n28894) );
  OAI21HSV2 U32499 ( .A1(n28892), .A2(n28893), .B(n28894), .ZN(n28895) );
  NAND2HSV0 U32500 ( .A1(n56622), .A2(n56493), .ZN(n28896) );
  NAND2HSV2 U32501 ( .A1(n28896), .A2(n28895), .ZN(n28897) );
  OAI21HSV2 U32502 ( .A1(n28895), .A2(n28896), .B(n28897), .ZN(n28898) );
  NAND2HSV0 U32503 ( .A1(n56175), .A2(n56174), .ZN(n28899) );
  NAND2HSV2 U32504 ( .A1(n28899), .A2(n28898), .ZN(n28900) );
  OAI21HSV2 U32505 ( .A1(n28898), .A2(n28899), .B(n28900), .ZN(n56248) );
  CLKNHSV0 U32506 ( .I(n50917), .ZN(n28901) );
  NAND2HSV0 U32507 ( .A1(n52905), .A2(n59792), .ZN(n28902) );
  NAND2HSV0 U32508 ( .A1(n51486), .A2(n53226), .ZN(n28903) );
  NAND2HSV0 U32509 ( .A1(n28903), .A2(n28902), .ZN(n28904) );
  OAI21HSV2 U32510 ( .A1(n28902), .A2(n28903), .B(n28904), .ZN(n28905) );
  MUX2NHSV1 U32511 ( .I0(n28901), .I1(n50917), .S(n28905), .ZN(n48623) );
  CLKNHSV0 U32512 ( .I(n54631), .ZN(n55589) );
  INOR2HSV0 U32513 ( .A1(n38878), .B1(n44307), .ZN(n52824) );
  NAND2HSV0 U32514 ( .A1(n25866), .A2(n32329), .ZN(n28906) );
  NAND2HSV0 U32515 ( .A1(n28906), .A2(poh6[10]), .ZN(n28907) );
  OAI21HSV2 U32516 ( .A1(poh6[10]), .A2(n28906), .B(n28907), .ZN(po[11]) );
  NOR2HSV0 U32517 ( .A1(n48010), .A2(n48011), .ZN(n28908) );
  NAND2HSV0 U32518 ( .A1(n28908), .A2(n48012), .ZN(n28909) );
  OAI211HSV0 U32519 ( .A1(n48012), .A2(n28908), .B(n28909), .C(n48013), .ZN(
        n28910) );
  NAND2HSV0 U32520 ( .A1(n28910), .A2(poh6[5]), .ZN(n28911) );
  OAI21HSV2 U32521 ( .A1(poh6[5]), .A2(n28910), .B(n28911), .ZN(po[6]) );
  CLKNHSV0 U32522 ( .I(n58382), .ZN(n28912) );
  CLKNHSV0 U32523 ( .I(n58381), .ZN(n28913) );
  XOR2HSV0 U32524 ( .A1(n58379), .A2(n58380), .Z(n28914) );
  XOR2HSV0 U32525 ( .A1(n58377), .A2(n58376), .Z(n28915) );
  XOR2HSV0 U32526 ( .A1(n28914), .A2(n28915), .Z(n28916) );
  MUX2NHSV0 U32527 ( .I0(n28913), .I1(n58381), .S(n28916), .ZN(n28917) );
  MUX2NHSV0 U32528 ( .I0(n28912), .I1(n58382), .S(n28917), .ZN(n28918) );
  NAND2HSV0 U32529 ( .A1(n53172), .A2(n58403), .ZN(n28919) );
  CLKNAND2HSV0 U32530 ( .A1(n28919), .A2(n28918), .ZN(n28920) );
  OAI21HSV0 U32531 ( .A1(n28918), .A2(n28919), .B(n28920), .ZN(n28921) );
  NAND2HSV0 U32532 ( .A1(n58809), .A2(n58724), .ZN(n28922) );
  CLKNAND2HSV0 U32533 ( .A1(n28922), .A2(n28921), .ZN(n28923) );
  OAI21HSV0 U32534 ( .A1(n28921), .A2(n28922), .B(n28923), .ZN(n28924) );
  CLKNAND2HSV0 U32535 ( .A1(n49181), .A2(n58423), .ZN(n28925) );
  CLKNAND2HSV0 U32536 ( .A1(n28925), .A2(n28924), .ZN(n28926) );
  OAI21HSV0 U32537 ( .A1(n28924), .A2(n28925), .B(n28926), .ZN(n28927) );
  NAND2HSV0 U32538 ( .A1(n58401), .A2(n58575), .ZN(n28928) );
  CLKNAND2HSV0 U32539 ( .A1(n28928), .A2(n28927), .ZN(n28929) );
  OAI21HSV0 U32540 ( .A1(n28927), .A2(n28928), .B(n28929), .ZN(n28930) );
  NAND2HSV0 U32541 ( .A1(n48888), .A2(n58384), .ZN(n28931) );
  CLKNAND2HSV0 U32542 ( .A1(n28931), .A2(n28930), .ZN(n28932) );
  OAI21HSV2 U32543 ( .A1(n28930), .A2(n28931), .B(n28932), .ZN(n28933) );
  NAND2HSV0 U32544 ( .A1(n58398), .A2(n59023), .ZN(n28934) );
  CLKNAND2HSV0 U32545 ( .A1(n28934), .A2(n28933), .ZN(n28935) );
  OAI21HSV0 U32546 ( .A1(n28933), .A2(n28934), .B(n28935), .ZN(\pe6/poht [26])
         );
  NAND2HSV0 U32547 ( .A1(n51399), .A2(n48841), .ZN(n28936) );
  CLKNAND2HSV0 U32548 ( .A1(n28936), .A2(n47425), .ZN(n28937) );
  OAI21HSV0 U32549 ( .A1(n47425), .A2(n28936), .B(n28937), .ZN(n28938) );
  NAND2HSV0 U32550 ( .A1(n53290), .A2(n51200), .ZN(n28939) );
  CLKNAND2HSV0 U32551 ( .A1(n28939), .A2(n28938), .ZN(n28940) );
  OAI21HSV0 U32552 ( .A1(n28938), .A2(n28939), .B(n28940), .ZN(n28941) );
  CLKNAND2HSV0 U32553 ( .A1(n51335), .A2(n59905), .ZN(n28942) );
  CLKNAND2HSV0 U32554 ( .A1(n28942), .A2(n28941), .ZN(n28943) );
  OAI21HSV0 U32555 ( .A1(n28941), .A2(n28942), .B(n28943), .ZN(n28944) );
  CLKNAND2HSV0 U32556 ( .A1(n51014), .A2(\pe5/got [8]), .ZN(n28945) );
  CLKNAND2HSV0 U32557 ( .A1(n28945), .A2(n28944), .ZN(n28946) );
  OAI21HSV0 U32558 ( .A1(n28944), .A2(n28945), .B(n28946), .ZN(n28947) );
  NAND2HSV0 U32559 ( .A1(n52669), .A2(n51358), .ZN(n28948) );
  CLKNAND2HSV0 U32560 ( .A1(n28948), .A2(n28947), .ZN(n28949) );
  OAI21HSV0 U32561 ( .A1(n28947), .A2(n28948), .B(n28949), .ZN(n28950) );
  NAND2HSV0 U32562 ( .A1(n53289), .A2(n51411), .ZN(n28951) );
  CLKNAND2HSV0 U32563 ( .A1(n28951), .A2(n28950), .ZN(n28952) );
  OAI21HSV0 U32564 ( .A1(n28950), .A2(n28951), .B(n28952), .ZN(n28953) );
  NAND2HSV0 U32565 ( .A1(n59643), .A2(n59580), .ZN(n28954) );
  CLKNAND2HSV0 U32566 ( .A1(n28954), .A2(n28953), .ZN(n28955) );
  OAI21HSV0 U32567 ( .A1(n28953), .A2(n28954), .B(n28955), .ZN(n28956) );
  NAND2HSV0 U32568 ( .A1(\pe5/got [12]), .A2(n29771), .ZN(n28957) );
  CLKNAND2HSV0 U32569 ( .A1(n28957), .A2(n28956), .ZN(n28958) );
  OAI21HSV0 U32570 ( .A1(n28956), .A2(n28957), .B(n28958), .ZN(\pe5/poht [20])
         );
  NAND2HSV0 U32571 ( .A1(n48482), .A2(\pe3/got [23]), .ZN(n28960) );
  CLKNAND2HSV0 U32572 ( .A1(n28960), .A2(n46544), .ZN(n28961) );
  OAI21HSV0 U32573 ( .A1(n46544), .A2(n28960), .B(n28961), .ZN(n28962) );
  NAND2HSV0 U32574 ( .A1(n56863), .A2(n55701), .ZN(n28963) );
  CLKNAND2HSV0 U32575 ( .A1(n28963), .A2(n28962), .ZN(n28964) );
  OAI21HSV0 U32576 ( .A1(n28962), .A2(n28963), .B(n28964), .ZN(n28965) );
  NAND2HSV0 U32577 ( .A1(n46441), .A2(n48481), .ZN(n28966) );
  CLKNAND2HSV0 U32578 ( .A1(n28966), .A2(n28965), .ZN(n28967) );
  OAI21HSV0 U32579 ( .A1(n28965), .A2(n28966), .B(n28967), .ZN(n28968) );
  NAND2HSV0 U32580 ( .A1(n45947), .A2(n55944), .ZN(n28969) );
  CLKNAND2HSV0 U32581 ( .A1(n28969), .A2(n28968), .ZN(n28970) );
  OAI21HSV0 U32582 ( .A1(n28968), .A2(n28969), .B(n28970), .ZN(n28971) );
  CLKNAND2HSV0 U32583 ( .A1(n28972), .A2(n28971), .ZN(n28973) );
  OAI21HSV0 U32584 ( .A1(n28971), .A2(n28972), .B(n28973), .ZN(n28974) );
  OAI21HSV0 U32585 ( .A1(n36799), .A2(n28959), .B(n28974), .ZN(n28975) );
  NAND2HSV0 U32586 ( .A1(n59963), .A2(n56260), .ZN(n28977) );
  CLKNAND2HSV0 U32587 ( .A1(n28977), .A2(n28976), .ZN(n28978) );
  OAI21HSV0 U32588 ( .A1(n28976), .A2(n28977), .B(n28978), .ZN(n28979) );
  NAND2HSV0 U32589 ( .A1(n59347), .A2(n56948), .ZN(n28980) );
  CLKNAND2HSV0 U32590 ( .A1(n28980), .A2(n28979), .ZN(n28981) );
  OAI21HSV0 U32591 ( .A1(n28979), .A2(n28980), .B(n28981), .ZN(\pe3/poht [2])
         );
  CLKNHSV0 U32592 ( .I(n52714), .ZN(n28982) );
  MUX2NHSV0 U32593 ( .I0(n28982), .I1(n52714), .S(n52713), .ZN(n28983) );
  NAND3HSV0 U32594 ( .A1(n52715), .A2(n52716), .A3(n52717), .ZN(n28984) );
  NAND2HSV0 U32595 ( .A1(n28984), .A2(n28983), .ZN(n28985) );
  OAI21HSV0 U32596 ( .A1(n28983), .A2(n28984), .B(n28985), .ZN(n60075) );
  CLKNHSV0 U32597 ( .I(n52775), .ZN(n28986) );
  OAI211HSV0 U32598 ( .A1(n52772), .A2(n52773), .B(n52774), .C(n52771), .ZN(
        n28987) );
  MUX2NHSV1 U32599 ( .I0(n28986), .I1(n52775), .S(n28987), .ZN(pov2[15]) );
  NAND2HSV2 U32600 ( .A1(n48019), .A2(\pe3/pvq [30]), .ZN(n28988) );
  NAND2HSV2 U32601 ( .A1(n28988), .A2(\pe3/phq [30]), .ZN(n28989) );
  OAI21HSV2 U32602 ( .A1(\pe3/phq [30]), .A2(n28988), .B(n28989), .ZN(n45685)
         );
  OAI22HSV0 U32603 ( .A1(n41460), .A2(n53723), .B1(n53447), .B2(n53691), .ZN(
        n28990) );
  OAI21HSV2 U32604 ( .A1(n41776), .A2(n42217), .B(n28990), .ZN(n41463) );
  OAI22HSV0 U32605 ( .A1(n36389), .A2(n38655), .B1(n48934), .B2(n36434), .ZN(
        n28991) );
  OAI21HSV2 U32606 ( .A1(n45192), .A2(n37896), .B(n28991), .ZN(n37898) );
  INHSV2 U32607 ( .I(n35427), .ZN(n28992) );
  CLKXOR2HSV4 U32608 ( .A1(n35426), .A2(n35425), .Z(n28993) );
  MUX2NHSV2 U32609 ( .I0(n28992), .I1(n35427), .S(n28993), .ZN(n35430) );
  NOR2HSV0 U32610 ( .A1(n41425), .A2(n54843), .ZN(n28994) );
  OAI22HSV0 U32611 ( .A1(n41888), .A2(n28994), .B1(n41890), .B2(n41889), .ZN(
        n28995) );
  OAI22HSV0 U32612 ( .A1(n46142), .A2(n41512), .B1(n41885), .B2(n41963), .ZN(
        n28996) );
  OAI21HSV0 U32613 ( .A1(n41886), .A2(n41887), .B(n28996), .ZN(n28997) );
  NAND2HSV0 U32614 ( .A1(n28997), .A2(n28995), .ZN(n28998) );
  OAI21HSV0 U32615 ( .A1(n28997), .A2(n28995), .B(n28998), .ZN(n41892) );
  NAND2HSV0 U32616 ( .A1(n39615), .A2(\pe5/aot [23]), .ZN(n28999) );
  AOI21HSV0 U32617 ( .A1(\pe5/bq[13] ), .A2(n48171), .B(n28999), .ZN(n29000)
         );
  AO31HSV2 U32618 ( .A1(\pe5/bq[13] ), .A2(n48171), .A3(n28999), .B(n29000), 
        .Z(n40215) );
  CLKNHSV0 U32619 ( .I(n52443), .ZN(n29001) );
  AOI22HSV0 U32620 ( .A1(n51547), .A2(n52444), .B1(\pe2/aot [7]), .B2(n52950), 
        .ZN(n29002) );
  AOI21HSV2 U32621 ( .A1(n52445), .A2(n29001), .B(n29002), .ZN(n52453) );
  NOR2HSV0 U32622 ( .A1(n45844), .A2(n59869), .ZN(n29003) );
  OAI22HSV0 U32623 ( .A1(n52627), .A2(n46920), .B1(n47303), .B2(n29003), .ZN(
        n45845) );
  CLKNHSV0 U32624 ( .I(n57016), .ZN(n29004) );
  AOI22HSV0 U32625 ( .A1(\pe4/aot [1]), .A2(n34598), .B1(n57850), .B2(n59683), 
        .ZN(n29005) );
  IAO21HSV0 U32626 ( .A1(n50360), .A2(n57988), .B(n29005), .ZN(n29006) );
  MUX2NHSV0 U32627 ( .I0(n57016), .I1(n29004), .S(n29006), .ZN(n50361) );
  AO22HSV0 U32628 ( .A1(n59217), .A2(n59250), .B1(n58464), .B2(n59247), .Z(
        n29007) );
  AOI21HSV0 U32629 ( .A1(\pe6/aot [13]), .A2(\pe6/bq[18] ), .B(n59106), .ZN(
        n29008) );
  AOI21HSV0 U32630 ( .A1(n59198), .A2(n59107), .B(n29008), .ZN(n29009) );
  OAI21HSV2 U32631 ( .A1(n59109), .A2(n59108), .B(n29007), .ZN(n29010) );
  NAND2HSV2 U32632 ( .A1(n29010), .A2(n29009), .ZN(n29011) );
  OAI21HSV2 U32633 ( .A1(n29010), .A2(n29009), .B(n29011), .ZN(n59113) );
  AOI22HSV0 U32634 ( .A1(n58731), .A2(n46662), .B1(n59088), .B2(\pe6/bq[14] ), 
        .ZN(n29012) );
  IAO21HSV2 U32635 ( .A1(n46661), .A2(n49852), .B(n29012), .ZN(n46665) );
  CLKNHSV0 U32636 ( .I(n33450), .ZN(n29013) );
  OAI21HSV2 U32637 ( .A1(n33909), .A2(n29013), .B(n45803), .ZN(n33569) );
  INAND2HSV0 U32638 ( .A1(n38728), .B1(n38729), .ZN(n38730) );
  NAND2HSV0 U32639 ( .A1(n53411), .A2(n40898), .ZN(n29014) );
  OAI21HSV0 U32640 ( .A1(n40412), .A2(n41622), .B(n41162), .ZN(n29015) );
  OAI21HSV0 U32641 ( .A1(n29014), .A2(n40413), .B(n29015), .ZN(n40414) );
  NAND2HSV2 U32642 ( .A1(n29016), .A2(n48311), .ZN(n29017) );
  OAI21HSV4 U32643 ( .A1(n48311), .A2(n29016), .B(n29017), .ZN(n45783) );
  NOR2HSV2 U32644 ( .A1(n34207), .A2(n34208), .ZN(n29018) );
  INAND3HSV2 U32645 ( .A1(n34317), .B1(n34319), .B2(n34320), .ZN(n52820) );
  NAND2HSV0 U32646 ( .A1(n47940), .A2(n48001), .ZN(n29019) );
  NAND2HSV0 U32647 ( .A1(n29019), .A2(poh6[26]), .ZN(n29020) );
  OAI21HSV2 U32648 ( .A1(poh6[26]), .A2(n29019), .B(n29020), .ZN(po[27]) );
  CLKNHSV0 U32649 ( .I(n32838), .ZN(n29021) );
  AOI21HSV4 U32650 ( .A1(n29021), .A2(n32416), .B(n32417), .ZN(n32648) );
  XOR2HSV0 U32651 ( .A1(n58804), .A2(n58803), .Z(n29023) );
  XOR2HSV0 U32652 ( .A1(n58806), .A2(n29023), .Z(n29024) );
  NAND2HSV0 U32653 ( .A1(n58717), .A2(n59178), .ZN(n29025) );
  CLKNAND2HSV0 U32654 ( .A1(n29025), .A2(n29024), .ZN(n29026) );
  OAI21HSV0 U32655 ( .A1(n29024), .A2(n29025), .B(n29026), .ZN(n29027) );
  NAND2HSV0 U32656 ( .A1(n58716), .A2(n58715), .ZN(n29028) );
  CLKNAND2HSV0 U32657 ( .A1(n29028), .A2(n29027), .ZN(n29029) );
  OAI21HSV0 U32658 ( .A1(n29027), .A2(n29028), .B(n29029), .ZN(n29030) );
  NAND2HSV0 U32659 ( .A1(n29753), .A2(n58807), .ZN(n29031) );
  CLKNAND2HSV0 U32660 ( .A1(n29031), .A2(n29030), .ZN(n29032) );
  OAI21HSV0 U32661 ( .A1(n29030), .A2(n29031), .B(n29032), .ZN(n29033) );
  NAND2HSV0 U32662 ( .A1(n59172), .A2(n59029), .ZN(n29034) );
  CLKNAND2HSV0 U32663 ( .A1(n29034), .A2(n29033), .ZN(n29035) );
  OAI21HSV0 U32664 ( .A1(n29033), .A2(n29034), .B(n29035), .ZN(n29036) );
  NAND2HSV0 U32665 ( .A1(n59170), .A2(n59328), .ZN(n29037) );
  CLKNAND2HSV0 U32666 ( .A1(n29037), .A2(n29036), .ZN(n29038) );
  OAI21HSV0 U32667 ( .A1(n29036), .A2(n29037), .B(n29038), .ZN(n29039) );
  NAND2HSV0 U32668 ( .A1(n58714), .A2(n59169), .ZN(n29040) );
  CLKNAND2HSV0 U32669 ( .A1(n29040), .A2(n29039), .ZN(n29041) );
  OAI21HSV0 U32670 ( .A1(n29039), .A2(n29040), .B(n29041), .ZN(n29042) );
  OAI21HSV2 U32671 ( .A1(n29042), .A2(n29043), .B(n29044), .ZN(n29045) );
  CLKNAND2HSV0 U32672 ( .A1(n59165), .A2(n29772), .ZN(n29046) );
  CLKNAND2HSV0 U32673 ( .A1(n29046), .A2(n29045), .ZN(n29047) );
  OAI21HSV0 U32674 ( .A1(n29045), .A2(n29046), .B(n29047), .ZN(\pe6/poht [8])
         );
  NAND2HSV0 U32675 ( .A1(n34843), .A2(n57755), .ZN(n29048) );
  NAND2HSV0 U32676 ( .A1(n29048), .A2(n46582), .ZN(n29049) );
  OAI21HSV0 U32677 ( .A1(n46582), .A2(n29048), .B(n29049), .ZN(n29050) );
  NAND2HSV0 U32678 ( .A1(n47772), .A2(n58193), .ZN(n29051) );
  CLKNAND2HSV0 U32679 ( .A1(n29051), .A2(n29050), .ZN(n29052) );
  OAI21HSV0 U32680 ( .A1(n29050), .A2(n29051), .B(n29052), .ZN(n60078) );
  CLKNHSV0 U32681 ( .I(n41236), .ZN(n29053) );
  CLKNHSV0 U32682 ( .I(n41233), .ZN(n29055) );
  CLKNHSV0 U32683 ( .I(n41231), .ZN(n29056) );
  OAI211HSV0 U32684 ( .A1(n59576), .A2(n41230), .B(n53512), .C(n41229), .ZN(
        n29058) );
  MUX2NHSV0 U32685 ( .I0(n41232), .I1(n29057), .S(n29058), .ZN(n29059) );
  MUX2NHSV0 U32686 ( .I0(n29056), .I1(n41231), .S(n29059), .ZN(n29060) );
  MUX2NHSV2 U32687 ( .I0(n41237), .I1(n29054), .S(n29061), .ZN(n60107) );
  XOR2HSV0 U32688 ( .A1(n51304), .A2(n51303), .Z(n29062) );
  NAND2HSV0 U32689 ( .A1(n52670), .A2(n51334), .ZN(n29063) );
  CLKNAND2HSV0 U32690 ( .A1(n29063), .A2(n29062), .ZN(n29064) );
  OAI21HSV0 U32691 ( .A1(n29062), .A2(n29063), .B(n29064), .ZN(n29065) );
  NAND2HSV0 U32692 ( .A1(n51335), .A2(\pe5/got [6]), .ZN(n29066) );
  CLKNAND2HSV0 U32693 ( .A1(n29066), .A2(n29065), .ZN(n29067) );
  OAI21HSV0 U32694 ( .A1(n29065), .A2(n29066), .B(n29067), .ZN(n29068) );
  NAND2HSV0 U32695 ( .A1(n51272), .A2(n51017), .ZN(n29069) );
  CLKNAND2HSV0 U32696 ( .A1(n29069), .A2(n29068), .ZN(n29070) );
  OAI21HSV0 U32697 ( .A1(n29068), .A2(n29069), .B(n29070), .ZN(n29071) );
  NAND2HSV0 U32698 ( .A1(n52563), .A2(\pe5/got [8]), .ZN(n29072) );
  CLKNAND2HSV0 U32699 ( .A1(n29072), .A2(n29071), .ZN(n29073) );
  OAI21HSV0 U32700 ( .A1(n29071), .A2(n29072), .B(n29073), .ZN(n29074) );
  NAND2HSV0 U32701 ( .A1(n52641), .A2(n51411), .ZN(n29075) );
  CLKNAND2HSV0 U32702 ( .A1(n29075), .A2(n29074), .ZN(n29076) );
  OAI21HSV0 U32703 ( .A1(n29074), .A2(n29075), .B(n29076), .ZN(n29077) );
  CLKNAND2HSV0 U32704 ( .A1(n53198), .A2(n53289), .ZN(n29078) );
  CLKNAND2HSV0 U32705 ( .A1(n29078), .A2(n29077), .ZN(n29079) );
  OAI21HSV0 U32706 ( .A1(n29077), .A2(n29078), .B(n29079), .ZN(n29080) );
  NAND2HSV0 U32707 ( .A1(n29771), .A2(n51305), .ZN(n29081) );
  CLKNAND2HSV0 U32708 ( .A1(n29081), .A2(n29080), .ZN(n29082) );
  OAI21HSV0 U32709 ( .A1(n29080), .A2(n29081), .B(n29082), .ZN(\pe5/poht [21])
         );
  XOR2HSV0 U32710 ( .A1(n49313), .A2(n49312), .Z(n29083) );
  AOI21HSV0 U32711 ( .A1(n49252), .A2(n55946), .B(n29083), .ZN(n29084) );
  AO31HSV0 U32712 ( .A1(n49252), .A2(n55946), .A3(n29083), .B(n29084), .Z(
        n29085) );
  NAND2HSV0 U32713 ( .A1(n56340), .A2(n56335), .ZN(n29086) );
  CLKNAND2HSV0 U32714 ( .A1(n29086), .A2(n29085), .ZN(n29087) );
  OAI21HSV0 U32715 ( .A1(n29085), .A2(n29086), .B(n29087), .ZN(n29088) );
  NAND2HSV0 U32716 ( .A1(\pe3/got [18]), .A2(n25989), .ZN(n29089) );
  CLKNAND2HSV0 U32717 ( .A1(n29089), .A2(n29088), .ZN(n29090) );
  OAI21HSV0 U32718 ( .A1(n29088), .A2(n29089), .B(n29090), .ZN(n29091) );
  NAND2HSV0 U32719 ( .A1(n56907), .A2(n56489), .ZN(n29092) );
  CLKNAND2HSV0 U32720 ( .A1(n29092), .A2(n29091), .ZN(n29093) );
  OAI21HSV0 U32721 ( .A1(n29091), .A2(n29092), .B(n29093), .ZN(n29094) );
  NAND2HSV0 U32722 ( .A1(n56172), .A2(n45581), .ZN(n29095) );
  CLKNAND2HSV0 U32723 ( .A1(n29095), .A2(n29094), .ZN(n29096) );
  OAI21HSV0 U32724 ( .A1(n29094), .A2(n29095), .B(n29096), .ZN(n29097) );
  NAND2HSV0 U32725 ( .A1(\pe3/got [22]), .A2(n56948), .ZN(n29101) );
  CLKNAND2HSV0 U32726 ( .A1(n29101), .A2(n29100), .ZN(n29102) );
  OAI21HSV0 U32727 ( .A1(n29100), .A2(n29101), .B(n29102), .ZN(\pe3/poht [10])
         );
  CLKNHSV0 U32728 ( .I(n47990), .ZN(n29103) );
  MUX2NHSV0 U32729 ( .I0(n29103), .I1(n47990), .S(n47989), .ZN(n60058) );
  CLKNHSV0 U32730 ( .I(n52792), .ZN(n29104) );
  NOR3HSV0 U32731 ( .A1(n26565), .A2(n52791), .A3(n42603), .ZN(n29105) );
  MUX2NHSV0 U32732 ( .I0(n52792), .I1(n29104), .S(n29105), .ZN(pov3[17]) );
  CLKNHSV0 U32733 ( .I(n52749), .ZN(n29106) );
  NAND2HSV0 U32734 ( .A1(n52747), .A2(n52748), .ZN(n29107) );
  AOI21HSV0 U32735 ( .A1(n52746), .A2(n52745), .B(n29107), .ZN(n29108) );
  MUX2NHSV0 U32736 ( .I0(n52749), .I1(n29106), .S(n29108), .ZN(n60043) );
  INOR2HSV0 U32737 ( .A1(n52776), .B1(n52777), .ZN(n29109) );
  CLKNAND2HSV0 U32738 ( .A1(n29109), .A2(n26790), .ZN(n29110) );
  OAI21HSV0 U32739 ( .A1(n29109), .A2(n26790), .B(n29110), .ZN(n60050) );
  OAI22HSV0 U32740 ( .A1(n36124), .A2(n58483), .B1(n36123), .B2(n59193), .ZN(
        n29111) );
  OAI21HSV2 U32741 ( .A1(n36125), .A2(n36126), .B(n29111), .ZN(n36129) );
  OAI22HSV0 U32742 ( .A1(n42264), .A2(n42361), .B1(n54829), .B2(n41461), .ZN(
        n29112) );
  OAI21HSV0 U32743 ( .A1(n41739), .A2(n42211), .B(n29112), .ZN(n41462) );
  OAI22HSV0 U32744 ( .A1(n49518), .A2(n38655), .B1(n48934), .B2(n44854), .ZN(
        n29113) );
  OAI21HSV0 U32745 ( .A1(n38123), .A2(n38295), .B(n29113), .ZN(n38124) );
  NOR2HSV0 U32746 ( .A1(n58013), .A2(n33250), .ZN(n29114) );
  OAI22HSV0 U32747 ( .A1(n58287), .A2(n50339), .B1(n50340), .B2(n29114), .ZN(
        n50344) );
  INOR2HSV0 U32748 ( .A1(\pe2/ti_7t [23]), .B1(n36473), .ZN(n43920) );
  AOI22HSV0 U32749 ( .A1(n44435), .A2(\pe6/aot [10]), .B1(n46658), .B2(
        \pe6/aot [1]), .ZN(n29115) );
  IAO21HSV0 U32750 ( .A1(n46657), .A2(n49841), .B(n29115), .ZN(n46659) );
  AOI22HSV0 U32751 ( .A1(n48530), .A2(\pe3/bq[4] ), .B1(n59809), .B2(n56971), 
        .ZN(n29116) );
  IAO21HSV0 U32752 ( .A1(n55859), .A2(n56097), .B(n29116), .ZN(n55860) );
  AOI21HSV0 U32753 ( .A1(n59088), .A2(n58619), .B(n49833), .ZN(n29117) );
  AOI21HSV0 U32754 ( .A1(n49762), .A2(n49683), .B(n29117), .ZN(n49338) );
  AOI22HSV0 U32755 ( .A1(n54078), .A2(n41623), .B1(n41760), .B2(n59985), .ZN(
        n29118) );
  AOI21HSV0 U32756 ( .A1(n41763), .A2(n40788), .B(n29118), .ZN(n40791) );
  OAI21HSV0 U32757 ( .A1(n35817), .A2(n59105), .B(n49682), .ZN(n29119) );
  CLKNAND2HSV0 U32758 ( .A1(n32596), .A2(n59236), .ZN(n29120) );
  NAND2HSV2 U32759 ( .A1(n29120), .A2(\pe6/phq [18]), .ZN(n29121) );
  OAI21HSV2 U32760 ( .A1(\pe6/phq [18]), .A2(n29120), .B(n29121), .ZN(n29122)
         );
  OAI21HSV0 U32761 ( .A1(n32372), .A2(n35929), .B(n29119), .ZN(n29123) );
  NAND2HSV0 U32762 ( .A1(n29123), .A2(n29122), .ZN(n29124) );
  OAI21HSV2 U32763 ( .A1(n29123), .A2(n29122), .B(n29124), .ZN(n32378) );
  NOR2HSV0 U32764 ( .A1(n49423), .A2(n56704), .ZN(n29125) );
  OAI22HSV0 U32765 ( .A1(n56940), .A2(n56116), .B1(n56578), .B2(n29125), .ZN(
        n53251) );
  CLKNHSV0 U32766 ( .I(n53322), .ZN(n29126) );
  NAND2HSV0 U32767 ( .A1(n53323), .A2(n50526), .ZN(n29127) );
  NAND2HSV0 U32768 ( .A1(n29127), .A2(n53321), .ZN(n29128) );
  OAI21HSV0 U32769 ( .A1(n53321), .A2(n29127), .B(n29128), .ZN(n29129) );
  NAND2HSV0 U32770 ( .A1(\pe5/aot [3]), .A2(\pe5/bq[14] ), .ZN(n29130) );
  NAND2HSV0 U32771 ( .A1(n29130), .A2(n29129), .ZN(n29131) );
  OAI21HSV0 U32772 ( .A1(n29129), .A2(n29130), .B(n29131), .ZN(n29132) );
  MUX2NHSV0 U32773 ( .I0(n29126), .I1(n53322), .S(n29132), .ZN(n53324) );
  CLKNHSV0 U32774 ( .I(\pe5/ti_7t [5]), .ZN(n29133) );
  XOR2HSV0 U32775 ( .A1(n47883), .A2(n47882), .Z(n29134) );
  XOR2HSV0 U32776 ( .A1(n47884), .A2(n29134), .Z(n29135) );
  NAND2HSV0 U32777 ( .A1(n58300), .A2(n59672), .ZN(n29136) );
  CLKNAND2HSV0 U32778 ( .A1(n29136), .A2(n29135), .ZN(n29137) );
  OAI21HSV0 U32779 ( .A1(n29135), .A2(n29136), .B(n29137), .ZN(n29138) );
  NAND2HSV0 U32780 ( .A1(n58220), .A2(\pe4/got [3]), .ZN(n29139) );
  CLKNAND2HSV0 U32781 ( .A1(n29139), .A2(n29138), .ZN(n29140) );
  OAI21HSV0 U32782 ( .A1(n29138), .A2(n29139), .B(n29140), .ZN(n29141) );
  NAND2HSV0 U32783 ( .A1(n58185), .A2(n58258), .ZN(n29142) );
  CLKNAND2HSV0 U32784 ( .A1(n29142), .A2(n29141), .ZN(n29143) );
  OAI21HSV0 U32785 ( .A1(n29141), .A2(n29142), .B(n29143), .ZN(n29144) );
  NAND2HSV0 U32786 ( .A1(n58218), .A2(n58246), .ZN(n29145) );
  CLKNAND2HSV0 U32787 ( .A1(n29145), .A2(n29144), .ZN(n29146) );
  OAI21HSV0 U32788 ( .A1(n29144), .A2(n29145), .B(n29146), .ZN(n29147) );
  CLKNAND2HSV0 U32789 ( .A1(n29148), .A2(n29147), .ZN(n29149) );
  NAND2HSV0 U32790 ( .A1(n58216), .A2(n59348), .ZN(n29151) );
  NAND2HSV0 U32791 ( .A1(n29151), .A2(n29150), .ZN(n29152) );
  OAI21HSV0 U32792 ( .A1(n29150), .A2(n29151), .B(n29152), .ZN(n29153) );
  NAND2HSV0 U32793 ( .A1(n57177), .A2(n26692), .ZN(n29154) );
  CLKNAND2HSV0 U32794 ( .A1(n29154), .A2(n29153), .ZN(n29155) );
  OAI21HSV2 U32795 ( .A1(n29153), .A2(n29154), .B(n29155), .ZN(n47886) );
  INOR2HSV2 U32796 ( .A1(n36650), .B1(n37835), .ZN(n36662) );
  CLKNHSV0 U32797 ( .I(n41231), .ZN(n29156) );
  CLKNHSV0 U32798 ( .I(n41232), .ZN(n29157) );
  MUX2NHSV1 U32799 ( .I0(n29157), .I1(n41232), .S(n29158), .ZN(n29159) );
  MUX2NHSV1 U32800 ( .I0(n29156), .I1(n41231), .S(n29159), .ZN(n41213) );
  CLKNHSV0 U32801 ( .I(n47942), .ZN(n29160) );
  NAND2HSV2 U32802 ( .A1(n47941), .A2(n29160), .ZN(n29161) );
  OAI211HSV1 U32803 ( .A1(n29160), .A2(n47941), .B(n29161), .C(n48013), .ZN(
        n29162) );
  NAND2HSV0 U32804 ( .A1(n29162), .A2(poh6[25]), .ZN(n29163) );
  OAI21HSV2 U32805 ( .A1(poh6[25]), .A2(n29162), .B(n29163), .ZN(po[26]) );
  CLKNHSV0 U32806 ( .I(n32685), .ZN(n29164) );
  AOI21HSV2 U32807 ( .A1(n29742), .A2(n52780), .B(n29164), .ZN(n32521) );
  NAND3HSV0 U32808 ( .A1(n34427), .A2(n57204), .A3(n34426), .ZN(n29165) );
  NAND2HSV0 U32809 ( .A1(n29165), .A2(n34419), .ZN(n34721) );
  CLKNHSV0 U32810 ( .I(n55514), .ZN(n29166) );
  XOR2HSV0 U32811 ( .A1(n55511), .A2(n55510), .Z(n29167) );
  NAND2HSV0 U32812 ( .A1(n59751), .A2(n54455), .ZN(n29168) );
  CLKNAND2HSV0 U32813 ( .A1(n29168), .A2(n29167), .ZN(n29169) );
  OAI21HSV0 U32814 ( .A1(n29167), .A2(n29168), .B(n29169), .ZN(n29170) );
  NAND2HSV0 U32815 ( .A1(n59736), .A2(n55340), .ZN(n29171) );
  CLKNAND2HSV0 U32816 ( .A1(n29171), .A2(n29170), .ZN(n29172) );
  OAI21HSV0 U32817 ( .A1(n29170), .A2(n29171), .B(n29172), .ZN(n29173) );
  CLKNAND2HSV0 U32818 ( .A1(\pe1/got [4]), .A2(n55490), .ZN(n29174) );
  CLKNAND2HSV0 U32819 ( .A1(n29174), .A2(n29173), .ZN(n29175) );
  OAI21HSV0 U32820 ( .A1(n29173), .A2(n29174), .B(n29175), .ZN(n29176) );
  OAI21HSV0 U32821 ( .A1(n55512), .A2(n29166), .B(n29176), .ZN(n29177) );
  OAI31HSV0 U32822 ( .A1(n55512), .A2(n29176), .A3(n29166), .B(n29177), .ZN(
        n29178) );
  NAND2HSV0 U32823 ( .A1(n55489), .A2(n55475), .ZN(n29179) );
  CLKNAND2HSV0 U32824 ( .A1(n29179), .A2(n29178), .ZN(n29180) );
  OAI21HSV0 U32825 ( .A1(n29178), .A2(n29179), .B(n29180), .ZN(n29181) );
  NAND2HSV0 U32826 ( .A1(n55488), .A2(n55448), .ZN(n29182) );
  CLKNAND2HSV0 U32827 ( .A1(n29182), .A2(n29181), .ZN(n29183) );
  OAI21HSV0 U32828 ( .A1(n29181), .A2(n29182), .B(n29183), .ZN(n29184) );
  CLKNAND2HSV0 U32829 ( .A1(n29185), .A2(n29184), .ZN(n29186) );
  OAI21HSV2 U32830 ( .A1(n29184), .A2(n29185), .B(n29186), .ZN(n29187) );
  NAND2HSV0 U32831 ( .A1(n55339), .A2(n59520), .ZN(n29188) );
  CLKNAND2HSV0 U32832 ( .A1(n29188), .A2(n29187), .ZN(n29189) );
  OAI21HSV0 U32833 ( .A1(n29187), .A2(n29188), .B(n29189), .ZN(\pe1/poht [24])
         );
  NAND2HSV0 U32834 ( .A1(n59022), .A2(n59167), .ZN(n29190) );
  CLKNAND2HSV0 U32835 ( .A1(n59025), .A2(n59514), .ZN(n29191) );
  NAND2HSV0 U32836 ( .A1(n32970), .A2(n53172), .ZN(n29192) );
  CLKNHSV0 U32837 ( .I(n49735), .ZN(n29193) );
  NAND2HSV0 U32838 ( .A1(n59028), .A2(n59175), .ZN(n29194) );
  MUX2NHSV0 U32839 ( .I0(n49735), .I1(n29193), .S(n29194), .ZN(n29195) );
  NAND2HSV0 U32840 ( .A1(n59027), .A2(n58934), .ZN(n29196) );
  XOR2HSV0 U32841 ( .A1(n29195), .A2(n29196), .Z(n29197) );
  XOR2HSV0 U32842 ( .A1(n29192), .A2(n29197), .Z(n29198) );
  NAND2HSV0 U32843 ( .A1(n59173), .A2(n58385), .ZN(n29199) );
  XOR2HSV0 U32844 ( .A1(n29198), .A2(n29199), .Z(n29200) );
  XOR2HSV0 U32845 ( .A1(n29191), .A2(n29200), .Z(n29201) );
  NAND2HSV0 U32846 ( .A1(n59024), .A2(n49665), .ZN(n29202) );
  XOR2HSV0 U32847 ( .A1(n29201), .A2(n29202), .Z(n29203) );
  XOR2HSV0 U32848 ( .A1(n29204), .A2(n29205), .Z(\pe6/poht [3]) );
  CLKNHSV0 U32849 ( .I(n37414), .ZN(n29206) );
  MUX2NHSV0 U32850 ( .I0(n29206), .I1(n37414), .S(n42682), .ZN(n60046) );
  AOI21HSV4 U32851 ( .A1(n41592), .A2(n40654), .B(n29208), .ZN(n29209) );
  XOR2HSV0 U32852 ( .A1(n51333), .A2(n51332), .Z(n29210) );
  NAND2HSV0 U32853 ( .A1(n52565), .A2(n51418), .ZN(n29211) );
  CLKNAND2HSV0 U32854 ( .A1(n29211), .A2(n29210), .ZN(n29212) );
  OAI21HSV0 U32855 ( .A1(n29210), .A2(n29211), .B(n29212), .ZN(n29213) );
  CLKNAND2HSV0 U32856 ( .A1(n51404), .A2(n51334), .ZN(n29214) );
  CLKNAND2HSV0 U32857 ( .A1(n29214), .A2(n29213), .ZN(n29215) );
  OAI21HSV0 U32858 ( .A1(n29213), .A2(n29214), .B(n29215), .ZN(n29216) );
  NAND2HSV0 U32859 ( .A1(n52564), .A2(n51200), .ZN(n29217) );
  CLKNAND2HSV0 U32860 ( .A1(n29217), .A2(n29216), .ZN(n29218) );
  OAI21HSV0 U32861 ( .A1(n29216), .A2(n29217), .B(n29218), .ZN(n29219) );
  NAND2HSV0 U32862 ( .A1(n52669), .A2(n59905), .ZN(n29220) );
  CLKNAND2HSV0 U32863 ( .A1(n29220), .A2(n29219), .ZN(n29221) );
  OAI21HSV0 U32864 ( .A1(n29219), .A2(n29220), .B(n29221), .ZN(n29222) );
  NAND2HSV0 U32865 ( .A1(n29777), .A2(n50698), .ZN(n29223) );
  CLKNAND2HSV0 U32866 ( .A1(n29223), .A2(n29222), .ZN(n29224) );
  OAI21HSV0 U32867 ( .A1(n29222), .A2(n29223), .B(n29224), .ZN(n29225) );
  CLKNAND2HSV0 U32868 ( .A1(n52668), .A2(n59891), .ZN(n29226) );
  CLKNAND2HSV0 U32869 ( .A1(n29226), .A2(n29225), .ZN(n29227) );
  OAI21HSV2 U32870 ( .A1(n29225), .A2(n29226), .B(n29227), .ZN(n29228) );
  NAND2HSV0 U32871 ( .A1(n53210), .A2(n53289), .ZN(n29229) );
  CLKNAND2HSV0 U32872 ( .A1(n29229), .A2(n29228), .ZN(n29230) );
  OAI21HSV0 U32873 ( .A1(n29228), .A2(n29229), .B(n29230), .ZN(\pe5/poht [22])
         );
  XOR2HSV0 U32874 ( .A1(n47495), .A2(n47494), .Z(n29231) );
  NAND2HSV0 U32875 ( .A1(n56863), .A2(n56174), .ZN(n29232) );
  CLKNAND2HSV0 U32876 ( .A1(n29232), .A2(n29231), .ZN(n29233) );
  OAI21HSV0 U32877 ( .A1(n29231), .A2(n29232), .B(n29233), .ZN(n29234) );
  NAND2HSV0 U32878 ( .A1(n56173), .A2(n56065), .ZN(n29235) );
  CLKNAND2HSV0 U32879 ( .A1(n29235), .A2(n29234), .ZN(n29236) );
  OAI21HSV0 U32880 ( .A1(n29234), .A2(n29235), .B(n29236), .ZN(n29237) );
  NAND2HSV0 U32881 ( .A1(n25989), .A2(n56335), .ZN(n29238) );
  CLKNAND2HSV0 U32882 ( .A1(n29238), .A2(n29237), .ZN(n29239) );
  OAI21HSV0 U32883 ( .A1(n29237), .A2(n29238), .B(n29239), .ZN(n29240) );
  NAND2HSV0 U32884 ( .A1(n48480), .A2(\pe3/got [18]), .ZN(n29241) );
  CLKNAND2HSV0 U32885 ( .A1(n29241), .A2(n29240), .ZN(n29242) );
  OAI21HSV0 U32886 ( .A1(n29240), .A2(n29241), .B(n29242), .ZN(n29243) );
  NAND2HSV0 U32887 ( .A1(n56172), .A2(n59965), .ZN(n29244) );
  CLKNAND2HSV0 U32888 ( .A1(n29244), .A2(n29243), .ZN(n29245) );
  OAI21HSV0 U32889 ( .A1(n29243), .A2(n29244), .B(n29245), .ZN(n29246) );
  NAND2HSV0 U32890 ( .A1(n29247), .A2(n29246), .ZN(n29248) );
  NAND2HSV0 U32891 ( .A1(n56965), .A2(n56171), .ZN(n29250) );
  CLKNAND2HSV0 U32892 ( .A1(n29250), .A2(n29249), .ZN(n29251) );
  OAI21HSV0 U32893 ( .A1(n29249), .A2(n29250), .B(n29251), .ZN(\pe3/poht [11])
         );
  XOR2HSV0 U32894 ( .A1(n47900), .A2(n47899), .Z(n29252) );
  NAND2HSV0 U32895 ( .A1(n51878), .A2(n52901), .ZN(n29253) );
  CLKNAND2HSV0 U32896 ( .A1(n29253), .A2(n29252), .ZN(n29254) );
  OAI21HSV0 U32897 ( .A1(n29252), .A2(n29253), .B(n29254), .ZN(n29255) );
  NAND2HSV0 U32898 ( .A1(n51797), .A2(n52895), .ZN(n29256) );
  CLKNAND2HSV0 U32899 ( .A1(n29256), .A2(n29255), .ZN(n29257) );
  OAI21HSV0 U32900 ( .A1(n29255), .A2(n29256), .B(n29257), .ZN(n29258) );
  CLKNAND2HSV0 U32901 ( .A1(n29259), .A2(n29258), .ZN(n29260) );
  OAI21HSV0 U32902 ( .A1(n29258), .A2(n29259), .B(n29260), .ZN(n29261) );
  NAND2HSV0 U32903 ( .A1(n52414), .A2(n52855), .ZN(n29262) );
  CLKNAND2HSV0 U32904 ( .A1(n29262), .A2(n29261), .ZN(n29263) );
  OAI21HSV0 U32905 ( .A1(n29261), .A2(n29262), .B(n29263), .ZN(n29264) );
  CLKNAND2HSV0 U32906 ( .A1(n52840), .A2(n59778), .ZN(n29265) );
  CLKNAND2HSV0 U32907 ( .A1(n29265), .A2(n29264), .ZN(n29266) );
  NAND2HSV0 U32908 ( .A1(n59794), .A2(n59777), .ZN(n29268) );
  CLKNAND2HSV0 U32909 ( .A1(n29268), .A2(n29267), .ZN(n29269) );
  OAI21HSV0 U32910 ( .A1(n29267), .A2(n29268), .B(n29269), .ZN(\pe2/poht [26])
         );
  CLKNHSV0 U32911 ( .I(n52754), .ZN(n29270) );
  MUX2NHSV0 U32912 ( .I0(n52754), .I1(n29270), .S(n52753), .ZN(n29271) );
  CLKNAND2HSV0 U32913 ( .A1(n52834), .A2(n59871), .ZN(n29272) );
  CLKNAND2HSV0 U32914 ( .A1(n29272), .A2(n29271), .ZN(n29273) );
  OAI21HSV0 U32915 ( .A1(n29271), .A2(n29272), .B(n29273), .ZN(pov5[12]) );
  CLKNHSV0 U32916 ( .I(n52699), .ZN(n29274) );
  AOI21HSV0 U32917 ( .A1(n52697), .A2(n52698), .B(n33184), .ZN(n29275) );
  MUX2NHSV0 U32918 ( .I0(n29274), .I1(n52699), .S(n29275), .ZN(n60034) );
  CLKNHSV0 U32919 ( .I(n52730), .ZN(n29276) );
  MUX2NHSV0 U32920 ( .I0(n29276), .I1(n52730), .S(n52729), .ZN(n29277) );
  XOR2HSV0 U32921 ( .A1(n29277), .A2(n52731), .Z(n60080) );
  CLKNHSV0 U32922 ( .I(n48620), .ZN(n29278) );
  MUX2NHSV0 U32923 ( .I0(n29278), .I1(n48620), .S(n48619), .ZN(n29279) );
  INHSV2 U32924 ( .I(n46122), .ZN(n29280) );
  INAND3HSV0 U32925 ( .A1(n46120), .B1(n38606), .B2(n46121), .ZN(n29281) );
  MUX2NHSV1 U32926 ( .I0(n29280), .I1(n46122), .S(n29281), .ZN(pov2[17]) );
  XOR2HSV0 U32927 ( .A1(n40369), .A2(n51113), .Z(n29282) );
  NAND2HSV0 U32928 ( .A1(n59675), .A2(n51114), .ZN(n29283) );
  NAND2HSV0 U32929 ( .A1(n29283), .A2(n29282), .ZN(n29284) );
  OAI21HSV2 U32930 ( .A1(n29282), .A2(n29283), .B(n29284), .ZN(n60109) );
  INOR2HSV0 U32931 ( .A1(n34453), .B1(n34452), .ZN(n34455) );
  CLKNHSV0 U32932 ( .I(\pe4/phq [8]), .ZN(n29285) );
  NAND2HSV0 U32933 ( .A1(n33808), .A2(\pe4/pvq [8]), .ZN(n29286) );
  MUX2NHSV1 U32934 ( .I0(\pe4/phq [8]), .I1(n29285), .S(n29286), .ZN(n33139)
         );
  OAI22HSV0 U32935 ( .A1(n37940), .A2(n47608), .B1(n48934), .B2(n38687), .ZN(
        n29287) );
  OAI21HSV0 U32936 ( .A1(n38548), .A2(n38300), .B(n29287), .ZN(n29288) );
  NAND2HSV0 U32937 ( .A1(n29288), .A2(n38494), .ZN(n29289) );
  OAI21HSV0 U32938 ( .A1(n29288), .A2(n38494), .B(n29289), .ZN(n38301) );
  XOR2HSV0 U32939 ( .A1(n33906), .A2(n33908), .Z(n29290) );
  XOR2HSV0 U32940 ( .A1(n33907), .A2(n29290), .Z(n29291) );
  CLKNAND2HSV0 U32941 ( .A1(n47733), .A2(n59372), .ZN(n29292) );
  NAND2HSV2 U32942 ( .A1(n29292), .A2(n29291), .ZN(n29293) );
  OAI21HSV2 U32943 ( .A1(n29291), .A2(n29292), .B(n29293), .ZN(n29294) );
  NAND2HSV0 U32944 ( .A1(n34396), .A2(n59602), .ZN(n29295) );
  NAND2HSV2 U32945 ( .A1(n29295), .A2(n29294), .ZN(n29296) );
  OAI21HSV2 U32946 ( .A1(n29294), .A2(n29295), .B(n29296), .ZN(n29297) );
  NAND2HSV0 U32947 ( .A1(n35036), .A2(\pe4/got [20]), .ZN(n29298) );
  NAND2HSV2 U32948 ( .A1(n29298), .A2(n29297), .ZN(n29299) );
  OAI21HSV2 U32949 ( .A1(n29297), .A2(n29298), .B(n29299), .ZN(n29300) );
  NAND2HSV0 U32950 ( .A1(n59681), .A2(n59370), .ZN(n29301) );
  NAND2HSV0 U32951 ( .A1(n29301), .A2(n29300), .ZN(n29302) );
  OAI21HSV0 U32952 ( .A1(n29300), .A2(n29301), .B(n29302), .ZN(n33911) );
  NAND2HSV0 U32953 ( .A1(n38134), .A2(\pe2/bq[21] ), .ZN(n29303) );
  AOI21HSV0 U32954 ( .A1(n38303), .A2(n51639), .B(n29303), .ZN(n29304) );
  AO31HSV0 U32955 ( .A1(n38303), .A2(n51639), .A3(n29303), .B(n29304), .Z(
        n29305) );
  NAND2HSV0 U32956 ( .A1(n36608), .A2(n59758), .ZN(n29306) );
  NAND2HSV2 U32957 ( .A1(n29306), .A2(n29305), .ZN(n29307) );
  OAI21HSV2 U32958 ( .A1(n29305), .A2(n29306), .B(n29307), .ZN(n29308) );
  NAND2HSV0 U32959 ( .A1(n38393), .A2(n39052), .ZN(n29309) );
  NAND2HSV2 U32960 ( .A1(n29309), .A2(n29308), .ZN(n29310) );
  OAI21HSV2 U32961 ( .A1(n29308), .A2(n29309), .B(n29310), .ZN(n38142) );
  NAND2HSV0 U32962 ( .A1(n32971), .A2(n35813), .ZN(n29311) );
  NAND2HSV2 U32963 ( .A1(\pe6/got [19]), .A2(n36185), .ZN(n29312) );
  CLKNAND2HSV0 U32964 ( .A1(n29312), .A2(n29311), .ZN(n29313) );
  OAI21HSV0 U32965 ( .A1(n29311), .A2(n29312), .B(n29313), .ZN(n32834) );
  OAI22HSV0 U32966 ( .A1(n31044), .A2(n48031), .B1(n48219), .B2(n47162), .ZN(
        n29314) );
  NAND2HSV0 U32967 ( .A1(\pe5/pvq [30]), .A2(n48029), .ZN(n29315) );
  CLKNAND2HSV0 U32968 ( .A1(n29315), .A2(\pe5/phq [30]), .ZN(n29316) );
  OAI21HSV0 U32969 ( .A1(\pe5/phq [30]), .A2(n29315), .B(n29316), .ZN(n29317)
         );
  OAI21HSV2 U32970 ( .A1(n40227), .A2(n47325), .B(n29314), .ZN(n29318) );
  NAND2HSV0 U32971 ( .A1(n29318), .A2(n29317), .ZN(n29319) );
  OAI21HSV0 U32972 ( .A1(n29318), .A2(n29317), .B(n29319), .ZN(n40228) );
  AOI22HSV0 U32973 ( .A1(\pe4/bq[20] ), .A2(n59683), .B1(n57234), .B2(n57846), 
        .ZN(n29320) );
  IAO21HSV0 U32974 ( .A1(n57349), .A2(n57731), .B(n29320), .ZN(n57350) );
  NOR2HSV0 U32975 ( .A1(n43724), .A2(n43235), .ZN(n29321) );
  NAND2HSV0 U32976 ( .A1(n29321), .A2(n49253), .ZN(n43728) );
  AOI22HSV0 U32977 ( .A1(n59866), .A2(n52594), .B1(n47305), .B2(n50588), .ZN(
        n29322) );
  AOI21HSV0 U32978 ( .A1(n47238), .A2(n48675), .B(n29322), .ZN(n47239) );
  AOI22HSV0 U32979 ( .A1(n56972), .A2(n48522), .B1(n55976), .B2(n56864), .ZN(
        n29323) );
  IAO21HSV2 U32980 ( .A1(n48521), .A2(n49420), .B(n29323), .ZN(n48524) );
  NAND2HSV0 U32981 ( .A1(n56094), .A2(n55864), .ZN(n29324) );
  NOR2HSV0 U32982 ( .A1(n55724), .A2(n56650), .ZN(n29325) );
  AOI21HSV2 U32983 ( .A1(n29324), .A2(n55725), .B(n29325), .ZN(n55726) );
  CLKNHSV0 U32984 ( .I(n56116), .ZN(n29326) );
  IOA21HSV2 U32985 ( .A1(n56113), .A2(\pe3/bq[9] ), .B(n56115), .ZN(n29327) );
  OAI21HSV2 U32986 ( .A1(n56114), .A2(n56426), .B(n29327), .ZN(n29328) );
  MUX2NHSV1 U32987 ( .I0(n29326), .I1(n56116), .S(n29328), .ZN(n56120) );
  AOI22HSV0 U32988 ( .A1(n46614), .A2(n56970), .B1(n56575), .B2(n56106), .ZN(
        n29329) );
  IAO21HSV0 U32989 ( .A1(n46347), .A2(n47434), .B(n29329), .ZN(n46360) );
  CLKNHSV0 U32990 ( .I(n44163), .ZN(n29330) );
  CLKNHSV0 U32991 ( .I(\pe2/phq [8]), .ZN(n29331) );
  NAND2HSV2 U32992 ( .A1(\pe2/pvq [8]), .A2(n45811), .ZN(n29332) );
  MUX2NHSV2 U32993 ( .I0(n29331), .I1(\pe2/phq [8]), .S(n29332), .ZN(n29333)
         );
  NAND2HSV0 U32994 ( .A1(n36603), .A2(n38064), .ZN(n29334) );
  CLKXOR2HSV2 U32995 ( .A1(n29333), .A2(n29334), .Z(n36544) );
  NAND2HSV0 U32996 ( .A1(n53718), .A2(n44569), .ZN(n29335) );
  NAND2HSV0 U32997 ( .A1(n40898), .A2(n41771), .ZN(n29336) );
  CLKNAND2HSV0 U32998 ( .A1(n29336), .A2(n29335), .ZN(n29337) );
  OAI21HSV0 U32999 ( .A1(n29335), .A2(n29336), .B(n29337), .ZN(n29338) );
  NAND2HSV0 U33000 ( .A1(n41298), .A2(n40741), .ZN(n29339) );
  CLKNAND2HSV0 U33001 ( .A1(n29339), .A2(n29338), .ZN(n29340) );
  OAI21HSV2 U33002 ( .A1(n29338), .A2(n29339), .B(n29340), .ZN(n40695) );
  CLKNAND2HSV0 U33003 ( .A1(n44702), .A2(n33022), .ZN(n29341) );
  OAI21HSV0 U33004 ( .A1(n35864), .A2(n46192), .B(n29341), .ZN(n29342) );
  OAI31HSV0 U33005 ( .A1(n35864), .A2(n29341), .A3(n46192), .B(n29342), .ZN(
        n32375) );
  AOI22HSV0 U33006 ( .A1(n54999), .A2(n55433), .B1(n59993), .B2(n54179), .ZN(
        n29343) );
  IAO21HSV2 U33007 ( .A1(n54998), .A2(n55118), .B(n29343), .ZN(n55000) );
  OAI21HSV0 U33008 ( .A1(n56914), .A2(n47447), .B(n56572), .ZN(n29344) );
  OAI21HSV0 U33009 ( .A1(n56574), .A2(n56573), .B(n29344), .ZN(n56580) );
  CLKNHSV0 U33010 ( .I(n40350), .ZN(n29345) );
  NAND2HSV2 U33011 ( .A1(n40349), .A2(n40348), .ZN(n29346) );
  MUX2NHSV0 U33012 ( .I0(n40350), .I1(n29345), .S(n29346), .ZN(n40351) );
  XOR2HSV0 U33013 ( .A1(n47767), .A2(n47769), .Z(n29347) );
  XOR2HSV0 U33014 ( .A1(n47768), .A2(n29347), .Z(n29348) );
  NAND2HSV0 U33015 ( .A1(\pe4/got [25]), .A2(n47904), .ZN(n29349) );
  CLKNAND2HSV0 U33016 ( .A1(n29349), .A2(n29348), .ZN(n29350) );
  OAI21HSV0 U33017 ( .A1(n29348), .A2(n29349), .B(n29350), .ZN(n29351) );
  NAND2HSV0 U33018 ( .A1(n47771), .A2(n57310), .ZN(n29352) );
  CLKNAND2HSV0 U33019 ( .A1(n29351), .A2(n29352), .ZN(n29353) );
  OAI21HSV0 U33020 ( .A1(n29351), .A2(n29352), .B(n29353), .ZN(n29354) );
  NAND2HSV0 U33021 ( .A1(n59837), .A2(n59350), .ZN(n29355) );
  CLKNAND2HSV0 U33022 ( .A1(n29355), .A2(n29354), .ZN(n29356) );
  NAND2HSV0 U33023 ( .A1(n58449), .A2(n58360), .ZN(n29360) );
  OAI21HSV0 U33024 ( .A1(n58537), .A2(n48887), .B(n29360), .ZN(n29361) );
  OAI31HSV0 U33025 ( .A1(n58537), .A2(n29360), .A3(n48887), .B(n29361), .ZN(
        n29362) );
  AOI21HSV0 U33026 ( .A1(n58460), .A2(n58734), .B(n29362), .ZN(n29363) );
  AO31HSV0 U33027 ( .A1(n58460), .A2(n58734), .A3(n29362), .B(n29363), .Z(
        n29364) );
  NAND2HSV0 U33028 ( .A1(n58405), .A2(n58459), .ZN(n29365) );
  CLKNAND2HSV0 U33029 ( .A1(n29365), .A2(n29364), .ZN(n29366) );
  OAI21HSV2 U33030 ( .A1(n29364), .A2(n29365), .B(n29366), .ZN(n29367) );
  NAND2HSV0 U33031 ( .A1(n58619), .A2(n58464), .ZN(n29368) );
  NAND2HSV0 U33032 ( .A1(n59062), .A2(\pe6/aot [6]), .ZN(n29369) );
  CLKNAND2HSV0 U33033 ( .A1(n29369), .A2(n29368), .ZN(n29370) );
  OAI21HSV0 U33034 ( .A1(n29368), .A2(n29369), .B(n29370), .ZN(n29371) );
  NAND2HSV0 U33035 ( .A1(n58496), .A2(\pe6/aot [7]), .ZN(n29372) );
  CLKNAND2HSV0 U33036 ( .A1(n29372), .A2(n29371), .ZN(n29373) );
  OAI21HSV0 U33037 ( .A1(n29371), .A2(n29372), .B(n29373), .ZN(n29374) );
  NAND2HSV0 U33038 ( .A1(\pe6/aot [1]), .A2(\pe6/bq[9] ), .ZN(n29375) );
  CLKNAND2HSV0 U33039 ( .A1(n29375), .A2(n29374), .ZN(n29376) );
  OAI21HSV0 U33040 ( .A1(n29374), .A2(n29375), .B(n29376), .ZN(n29377) );
  CLKNAND2HSV0 U33041 ( .A1(n49847), .A2(n58452), .ZN(n29378) );
  CLKNAND2HSV0 U33042 ( .A1(n29378), .A2(n29377), .ZN(n29379) );
  OAI21HSV0 U33043 ( .A1(n29377), .A2(n29378), .B(n29379), .ZN(n29380) );
  XOR2HSV0 U33044 ( .A1(n29367), .A2(n29380), .Z(n46148) );
  NAND2HSV0 U33045 ( .A1(n58197), .A2(n58230), .ZN(n29381) );
  AOI21HSV0 U33046 ( .A1(n58306), .A2(n58196), .B(n29381), .ZN(n29382) );
  AO31HSV2 U33047 ( .A1(n58306), .A2(n58196), .A3(n29381), .B(n29382), .Z(
        n29383) );
  NAND2HSV0 U33048 ( .A1(\pe4/aot [2]), .A2(n58195), .ZN(n29384) );
  OAI21HSV0 U33049 ( .A1(n48032), .A2(n58194), .B(n29384), .ZN(n29385) );
  OAI31HSV0 U33050 ( .A1(n48032), .A2(n29384), .A3(n58194), .B(n29385), .ZN(
        n29386) );
  NAND2HSV0 U33051 ( .A1(n58198), .A2(\pe4/bq[1] ), .ZN(n29387) );
  NAND2HSV0 U33052 ( .A1(\pe4/bq[2] ), .A2(n59352), .ZN(n29388) );
  CLKNAND2HSV0 U33053 ( .A1(n29388), .A2(n29387), .ZN(n29389) );
  OAI21HSV0 U33054 ( .A1(n29387), .A2(n29388), .B(n29389), .ZN(n29390) );
  NAND2HSV0 U33055 ( .A1(n58199), .A2(n58156), .ZN(n29391) );
  CLKNAND2HSV0 U33056 ( .A1(n29391), .A2(n29390), .ZN(n29392) );
  OAI21HSV0 U33057 ( .A1(n29390), .A2(n29391), .B(n29392), .ZN(n29393) );
  XOR2HSV0 U33058 ( .A1(n29383), .A2(n29386), .Z(n29394) );
  XOR2HSV0 U33059 ( .A1(n29393), .A2(n29394), .Z(n58200) );
  INOR2HSV0 U33060 ( .A1(\pe1/ti_7t [29]), .B1(n42335), .ZN(n44524) );
  NAND2HSV0 U33061 ( .A1(n32156), .A2(n33079), .ZN(n29395) );
  NAND2HSV0 U33062 ( .A1(n29395), .A2(poh6[13]), .ZN(n29396) );
  OAI21HSV2 U33063 ( .A1(poh6[13]), .A2(n29395), .B(n29396), .ZN(po[14]) );
  CLKNHSV0 U33064 ( .I(n48001), .ZN(n29397) );
  OAI21HSV0 U33065 ( .A1(n48000), .A2(n29397), .B(poh6[7]), .ZN(n29398) );
  OAI31HSV0 U33066 ( .A1(n48000), .A2(poh6[7]), .A3(n29397), .B(n29398), .ZN(
        po[8]) );
  INHSV2 U33067 ( .I(n48003), .ZN(n29399) );
  OAI21HSV0 U33068 ( .A1(n48002), .A2(n29399), .B(n48013), .ZN(n29400) );
  AOI21HSV2 U33069 ( .A1(n29399), .A2(n48004), .B(n29400), .ZN(n29401) );
  XOR2HSV0 U33070 ( .A1(n29401), .A2(poh6[6]), .Z(po[7]) );
  INAND2HSV0 U33071 ( .A1(\pe1/ti_7t [23]), .B1(n41712), .ZN(n42352) );
  NAND2HSV0 U33072 ( .A1(n46125), .A2(n46126), .ZN(n29402) );
  OAI21HSV0 U33073 ( .A1(\pe3/pq ), .A2(n46125), .B(n29402), .ZN(\pe3/ti_1t )
         );
  AOI21HSV0 U33074 ( .A1(n59489), .A2(n53367), .B(n53368), .ZN(n29403) );
  AO31HSV0 U33075 ( .A1(n59489), .A2(n53367), .A3(n53368), .B(n29403), .Z(
        n60103) );
  IOA21HSV4 U33076 ( .A1(n47996), .A2(n31900), .B(n31901), .ZN(n59596) );
  XOR2HSV0 U33077 ( .A1(n45922), .A2(n45921), .Z(n29404) );
  AOI21HSV0 U33078 ( .A1(n59355), .A2(n47268), .B(n29404), .ZN(n29405) );
  AO31HSV0 U33079 ( .A1(n59355), .A2(n47268), .A3(n29404), .B(n29405), .Z(
        n29406) );
  CLKNAND2HSV0 U33080 ( .A1(n51404), .A2(n52577), .ZN(n29407) );
  CLKNAND2HSV0 U33081 ( .A1(n29407), .A2(n29406), .ZN(n29408) );
  OAI21HSV0 U33082 ( .A1(n29406), .A2(n29407), .B(n29408), .ZN(n29409) );
  CLKNAND2HSV0 U33083 ( .A1(n53288), .A2(\pe5/got [5]), .ZN(n29410) );
  CLKNAND2HSV0 U33084 ( .A1(n29410), .A2(n29409), .ZN(n29411) );
  OAI21HSV0 U33085 ( .A1(n29409), .A2(n29410), .B(n29411), .ZN(n29412) );
  NAND2HSV0 U33086 ( .A1(n52669), .A2(n51200), .ZN(n29413) );
  CLKNAND2HSV0 U33087 ( .A1(n29413), .A2(n29412), .ZN(n29414) );
  OAI21HSV0 U33088 ( .A1(n29412), .A2(n29413), .B(n29414), .ZN(n29415) );
  CLKNAND2HSV0 U33089 ( .A1(n29775), .A2(n59905), .ZN(n29416) );
  CLKNAND2HSV0 U33090 ( .A1(n29416), .A2(n29415), .ZN(n29417) );
  OAI21HSV0 U33091 ( .A1(n29415), .A2(n29416), .B(n29417), .ZN(n29418) );
  NAND2HSV0 U33092 ( .A1(n50698), .A2(n53198), .ZN(n29419) );
  CLKNAND2HSV0 U33093 ( .A1(n29419), .A2(n29418), .ZN(n29420) );
  OAI21HSV2 U33094 ( .A1(n29418), .A2(n29419), .B(n29420), .ZN(n29421) );
  CLKNAND2HSV0 U33095 ( .A1(n59891), .A2(n52562), .ZN(n29422) );
  CLKNAND2HSV0 U33096 ( .A1(n29422), .A2(n29421), .ZN(n29423) );
  OAI21HSV0 U33097 ( .A1(n29421), .A2(n29422), .B(n29423), .ZN(\pe5/poht [23])
         );
  XOR2HSV0 U33098 ( .A1(n56416), .A2(n56415), .Z(n29424) );
  NAND2HSV0 U33099 ( .A1(n55822), .A2(n56421), .ZN(n29425) );
  CLKNAND2HSV0 U33100 ( .A1(n29425), .A2(n29424), .ZN(n29426) );
  OAI21HSV0 U33101 ( .A1(n29424), .A2(n29425), .B(n29426), .ZN(n29427) );
  NAND2HSV0 U33102 ( .A1(n55946), .A2(n56493), .ZN(n29428) );
  CLKNAND2HSV0 U33103 ( .A1(n29428), .A2(n29427), .ZN(n29429) );
  OAI21HSV0 U33104 ( .A1(n29427), .A2(n29428), .B(n29429), .ZN(n29430) );
  CLKNAND2HSV0 U33105 ( .A1(n56340), .A2(n56419), .ZN(n29431) );
  CLKNAND2HSV0 U33106 ( .A1(n29431), .A2(n29430), .ZN(n29432) );
  OAI21HSV0 U33107 ( .A1(n29430), .A2(n29431), .B(n29432), .ZN(n29433) );
  CLKNAND2HSV0 U33108 ( .A1(n29434), .A2(n29433), .ZN(n29435) );
  OAI21HSV0 U33109 ( .A1(n29433), .A2(n29434), .B(n29435), .ZN(n29436) );
  NAND2HSV0 U33110 ( .A1(n56339), .A2(n56335), .ZN(n29437) );
  CLKNAND2HSV0 U33111 ( .A1(n29437), .A2(n29436), .ZN(n29438) );
  OAI21HSV0 U33112 ( .A1(n29436), .A2(n29437), .B(n29438), .ZN(n29439) );
  NAND2HSV0 U33113 ( .A1(n56935), .A2(\pe3/got [18]), .ZN(n29440) );
  CLKNAND2HSV0 U33114 ( .A1(n29440), .A2(n29439), .ZN(n29441) );
  OAI21HSV0 U33115 ( .A1(n29439), .A2(n29440), .B(n29441), .ZN(n29442) );
  NAND3HSV0 U33116 ( .A1(n56418), .A2(n56489), .A3(n56417), .ZN(n29444) );
  CLKNHSV0 U33117 ( .I(n52898), .ZN(n29446) );
  CLKNHSV0 U33118 ( .I(n52897), .ZN(n29447) );
  OAI21HSV0 U33119 ( .A1(n49618), .A2(n47893), .B(n52899), .ZN(n29448) );
  OAI31HSV0 U33120 ( .A1(n49618), .A2(n52899), .A3(n47893), .B(n29448), .ZN(
        n29449) );
  MUX2NHSV0 U33121 ( .I0(n29447), .I1(n52897), .S(n29449), .ZN(n29450) );
  MUX2NHSV0 U33122 ( .I0(n52898), .I1(n29446), .S(n29450), .ZN(n29451) );
  NAND2HSV0 U33123 ( .A1(n52896), .A2(n59475), .ZN(n29452) );
  CLKNAND2HSV0 U33124 ( .A1(n29452), .A2(n29451), .ZN(n29453) );
  OAI21HSV0 U33125 ( .A1(n29451), .A2(n29452), .B(n29453), .ZN(n29454) );
  NAND2HSV0 U33126 ( .A1(n52895), .A2(n53093), .ZN(n29455) );
  CLKNAND2HSV0 U33127 ( .A1(n29455), .A2(n29454), .ZN(n29456) );
  CLKNAND2HSV0 U33128 ( .A1(n25709), .A2(n52900), .ZN(n29458) );
  NAND2HSV2 U33129 ( .A1(n29458), .A2(n29457), .ZN(n29459) );
  OAI21HSV2 U33130 ( .A1(n29457), .A2(n29458), .B(n29459), .ZN(n29460) );
  NAND2HSV0 U33131 ( .A1(n51896), .A2(n59794), .ZN(n29461) );
  CLKNAND2HSV0 U33132 ( .A1(n29461), .A2(n29460), .ZN(n29462) );
  OAI21HSV0 U33133 ( .A1(n29460), .A2(n29461), .B(n29462), .ZN(\pe2/poht [28])
         );
  NAND3HSV0 U33134 ( .A1(n52787), .A2(n52786), .A3(n52785), .ZN(n29463) );
  NAND2HSV0 U33135 ( .A1(n29463), .A2(n52788), .ZN(n29464) );
  OAI21HSV0 U33136 ( .A1(n52788), .A2(n29463), .B(n29464), .ZN(n60070) );
  INOR2HSV0 U33137 ( .A1(n52758), .B1(n52757), .ZN(n29465) );
  CLKNHSV0 U33138 ( .I(n52756), .ZN(n29466) );
  CLKNAND2HSV0 U33139 ( .A1(n59833), .A2(n52755), .ZN(n29467) );
  MUX2NHSV1 U33140 ( .I0(n29466), .I1(n25859), .S(n29467), .ZN(n29468) );
  OAI21HSV0 U33141 ( .A1(n52759), .A2(n29465), .B(n29718), .ZN(n29469) );
  CLKNAND2HSV0 U33142 ( .A1(n29469), .A2(n29468), .ZN(n29470) );
  OAI21HSV0 U33143 ( .A1(n29469), .A2(n29468), .B(n29470), .ZN(n60023) );
  INOR2HSV0 U33144 ( .A1(n52750), .B1(n52751), .ZN(n29471) );
  CLKNAND2HSV0 U33145 ( .A1(n29471), .A2(n52752), .ZN(n29472) );
  OAI21HSV0 U33146 ( .A1(n29471), .A2(n52752), .B(n29472), .ZN(n60059) );
  INHSV2 U33147 ( .I(n47949), .ZN(n29473) );
  MUX2NHSV1 U33148 ( .I0(n47949), .I1(n29473), .S(n29474), .ZN(pov3[22]) );
  INHSV2 U33149 ( .I(n53386), .ZN(n29475) );
  CLKNHSV0 U33150 ( .I(n53384), .ZN(n29476) );
  MUX2NHSV0 U33151 ( .I0(n29476), .I1(n53384), .S(n53385), .ZN(n29477) );
  MUX2NHSV1 U33152 ( .I0(n29475), .I1(n53386), .S(n29477), .ZN(n60097) );
  CLKNHSV0 U33153 ( .I(n52815), .ZN(n29478) );
  OAI211HSV0 U33154 ( .A1(n52813), .A2(n52814), .B(n52812), .C(n52811), .ZN(
        n29479) );
  MUX2NHSV0 U33155 ( .I0(n52815), .I1(n29478), .S(n29479), .ZN(n60047) );
  CLKNAND2HSV0 U33156 ( .A1(n41144), .A2(n51114), .ZN(n29480) );
  NAND2HSV0 U33157 ( .A1(n29480), .A2(n46610), .ZN(n29481) );
  OAI21HSV0 U33158 ( .A1(n46610), .A2(n29480), .B(n29481), .ZN(pov1[6]) );
  AOI22HSV0 U33159 ( .A1(n38803), .A2(n52104), .B1(n51825), .B2(n52941), .ZN(
        n29482) );
  AOI21HSV0 U33160 ( .A1(n45191), .A2(n44729), .B(n29482), .ZN(n44730) );
  CLKNHSV0 U33161 ( .I(n41757), .ZN(n29483) );
  OAI21HSV0 U33162 ( .A1(n53672), .A2(n53410), .B(n29483), .ZN(n41758) );
  OAI22HSV0 U33163 ( .A1(n53447), .A2(n45814), .B1(n46629), .B2(n41512), .ZN(
        n29484) );
  OAI21HSV0 U33164 ( .A1(n41777), .A2(n41634), .B(n29484), .ZN(n41513) );
  AOI22HSV0 U33165 ( .A1(n57459), .A2(n58283), .B1(n59605), .B2(n58116), .ZN(
        n29485) );
  IAO21HSV0 U33166 ( .A1(n50342), .A2(n50341), .B(n29485), .ZN(n50343) );
  AOI22HSV0 U33167 ( .A1(n59098), .A2(\pe6/aot [11]), .B1(n59100), .B2(n59099), 
        .ZN(n29486) );
  IAO21HSV0 U33168 ( .A1(n59097), .A2(n59187), .B(n29486), .ZN(n59101) );
  AOI22HSV0 U33169 ( .A1(\pe3/bq[19] ), .A2(n56911), .B1(\pe3/aot [22]), .B2(
        n56529), .ZN(n29487) );
  IAO21HSV0 U33170 ( .A1(n55638), .A2(n56837), .B(n29487), .ZN(n55639) );
  AOI22HSV0 U33171 ( .A1(n49836), .A2(n58962), .B1(n45812), .B2(n58353), .ZN(
        n29488) );
  IAO21HSV0 U33172 ( .A1(n49682), .A2(n58544), .B(n29488), .ZN(n49684) );
  AOI22HSV0 U33173 ( .A1(n56106), .A2(\pe3/aot [8]), .B1(n59808), .B2(n42971), 
        .ZN(n29489) );
  IAO21HSV0 U33174 ( .A1(n55848), .A2(n55991), .B(n29489), .ZN(n55853) );
  AO22HSV0 U33175 ( .A1(n48802), .A2(n59945), .B1(n52619), .B2(n48242), .Z(
        n29490) );
  AOI22HSV0 U33176 ( .A1(n50500), .A2(\pe5/aot [18]), .B1(\pe5/aot [3]), .B2(
        n48804), .ZN(n29491) );
  IAO21HSV0 U33177 ( .A1(n48803), .A2(n50584), .B(n29491), .ZN(n29492) );
  OAI21HSV0 U33178 ( .A1(n48801), .A2(n53321), .B(n29490), .ZN(n29493) );
  CLKNAND2HSV0 U33179 ( .A1(n29493), .A2(n29492), .ZN(n29494) );
  OAI21HSV0 U33180 ( .A1(n29493), .A2(n29492), .B(n29494), .ZN(n48805) );
  OAI21HSV0 U33181 ( .A1(n41650), .A2(n41622), .B(n40984), .ZN(n29495) );
  OAI21HSV0 U33182 ( .A1(n40789), .A2(n41352), .B(n29495), .ZN(n40790) );
  OAI22HSV0 U33183 ( .A1(n35816), .A2(n44397), .B1(n36132), .B2(n32373), .ZN(
        n29496) );
  OAI21HSV0 U33184 ( .A1(n32739), .A2(n32744), .B(n29496), .ZN(n29497) );
  CLKNAND2HSV0 U33185 ( .A1(n29497), .A2(n35839), .ZN(n29498) );
  OAI21HSV0 U33186 ( .A1(n29497), .A2(n35839), .B(n29498), .ZN(n32377) );
  INAND2HSV0 U33187 ( .A1(n34579), .B1(n34577), .ZN(n34582) );
  CLKNAND2HSV0 U33188 ( .A1(n54999), .A2(n59495), .ZN(n29499) );
  CLKNAND2HSV0 U33189 ( .A1(n48380), .A2(n54904), .ZN(n29500) );
  CLKNAND2HSV0 U33190 ( .A1(n29500), .A2(n29499), .ZN(n29501) );
  OAI21HSV0 U33191 ( .A1(n29499), .A2(n29500), .B(n29501), .ZN(n54644) );
  CLKNAND2HSV0 U33192 ( .A1(n59034), .A2(n59180), .ZN(n46725) );
  INOR2HSV0 U33193 ( .A1(n40141), .B1(n40142), .ZN(n40145) );
  INAND2HSV0 U33194 ( .A1(n30206), .B1(\pe5/ti_7t [3]), .ZN(n29859) );
  INAND2HSV0 U33195 ( .A1(\pe1/ti_7t [19]), .B1(n41242), .ZN(n41697) );
  INOR2HSV0 U33196 ( .A1(\pe2/ti_7t [11]), .B1(n44315), .ZN(n52746) );
  CLKNHSV0 U33197 ( .I(n48013), .ZN(n29502) );
  OAI21HSV0 U33198 ( .A1(n48009), .A2(n29502), .B(poh6[4]), .ZN(n29503) );
  OAI31HSV0 U33199 ( .A1(n48009), .A2(poh6[4]), .A3(n29502), .B(n29503), .ZN(
        po[5]) );
  CLKNHSV0 U33200 ( .I(n48018), .ZN(n29504) );
  OAI21HSV0 U33201 ( .A1(n48017), .A2(n29504), .B(poh6[1]), .ZN(n29505) );
  OAI31HSV0 U33202 ( .A1(n48017), .A2(poh6[1]), .A3(n29504), .B(n29505), .ZN(
        po[2]) );
  CLKNAND2HSV0 U33203 ( .A1(n59965), .A2(n55822), .ZN(n29506) );
  CLKNAND2HSV0 U33204 ( .A1(n29506), .A2(n49491), .ZN(n29507) );
  OAI21HSV0 U33205 ( .A1(n49491), .A2(n29506), .B(n29507), .ZN(n29508) );
  CLKNAND2HSV0 U33206 ( .A1(n55946), .A2(n49404), .ZN(n29509) );
  CLKNAND2HSV0 U33207 ( .A1(n29509), .A2(n29508), .ZN(n29510) );
  OAI21HSV0 U33208 ( .A1(n29508), .A2(n29509), .B(n29510), .ZN(n29511) );
  CLKNAND2HSV0 U33209 ( .A1(n56171), .A2(n56173), .ZN(n29512) );
  CLKNAND2HSV0 U33210 ( .A1(n29512), .A2(n29511), .ZN(n29513) );
  CLKNAND2HSV0 U33211 ( .A1(n48480), .A2(n42673), .ZN(n29516) );
  CLKNAND2HSV0 U33212 ( .A1(n53279), .A2(n59617), .ZN(n29519) );
  OAI21HSV0 U33213 ( .A1(n50752), .A2(n43457), .B(n29521), .ZN(n29522) );
  CLKNAND2HSV0 U33214 ( .A1(n56900), .A2(n59384), .ZN(n29524) );
  OAI21HSV0 U33215 ( .A1(n29524), .A2(n29523), .B(n29525), .ZN(\pe3/poht [6])
         );
  NOR2HSV0 U33216 ( .A1(n47905), .A2(n58013), .ZN(n29526) );
  CLKNAND2HSV0 U33217 ( .A1(n58219), .A2(n58254), .ZN(n29527) );
  CLKNAND2HSV0 U33218 ( .A1(n29527), .A2(n29526), .ZN(n29528) );
  OAI21HSV0 U33219 ( .A1(n29526), .A2(n29527), .B(n29528), .ZN(\pe4/poht [31])
         );
  XOR2HSV0 U33220 ( .A1(n49399), .A2(n49398), .Z(n29529) );
  CLKNAND2HSV0 U33221 ( .A1(n58480), .A2(n53101), .ZN(n29530) );
  CLKNAND2HSV0 U33222 ( .A1(n29530), .A2(n29529), .ZN(n29531) );
  OAI21HSV0 U33223 ( .A1(n29529), .A2(n29530), .B(n29531), .ZN(n29532) );
  CLKNAND2HSV0 U33224 ( .A1(n58934), .A2(n49096), .ZN(n29533) );
  CLKNAND2HSV0 U33225 ( .A1(n29533), .A2(n29532), .ZN(n29534) );
  OAI21HSV0 U33226 ( .A1(n29532), .A2(n29533), .B(n29534), .ZN(n29535) );
  CLKNAND2HSV0 U33227 ( .A1(n29753), .A2(n59029), .ZN(n29536) );
  CLKNAND2HSV0 U33228 ( .A1(n29536), .A2(n29535), .ZN(n29537) );
  OAI21HSV0 U33229 ( .A1(n29535), .A2(n29536), .B(n29537), .ZN(n29538) );
  CLKNAND2HSV0 U33230 ( .A1(n59172), .A2(\pe6/got [21]), .ZN(n29539) );
  CLKNAND2HSV0 U33231 ( .A1(n29539), .A2(n29538), .ZN(n29540) );
  OAI21HSV0 U33232 ( .A1(n29538), .A2(n29539), .B(n29540), .ZN(n29541) );
  CLKNAND2HSV0 U33233 ( .A1(n59170), .A2(n49825), .ZN(n29542) );
  CLKNAND2HSV0 U33234 ( .A1(n29542), .A2(n29541), .ZN(n29543) );
  OAI21HSV0 U33235 ( .A1(n29541), .A2(n29542), .B(n29543), .ZN(n29544) );
  CLKNAND2HSV0 U33236 ( .A1(n59027), .A2(n58575), .ZN(n29545) );
  CLKNAND2HSV0 U33237 ( .A1(n29545), .A2(n29544), .ZN(n29546) );
  OAI21HSV0 U33238 ( .A1(n29544), .A2(n29545), .B(n29546), .ZN(n29547) );
  CLKNAND2HSV0 U33239 ( .A1(n59021), .A2(n59165), .ZN(n29548) );
  CLKNAND2HSV0 U33240 ( .A1(n29548), .A2(n29547), .ZN(n29549) );
  OAI21HSV0 U33241 ( .A1(n29547), .A2(n29548), .B(n29549), .ZN(n29550) );
  CLKNAND2HSV0 U33242 ( .A1(n46283), .A2(n58476), .ZN(n29551) );
  CLKNAND2HSV0 U33243 ( .A1(n29551), .A2(n29550), .ZN(n29552) );
  OAI21HSV0 U33244 ( .A1(n29550), .A2(n29551), .B(n29552), .ZN(\pe6/poht [7])
         );
  XOR2HSV0 U33245 ( .A1(n52692), .A2(n52691), .Z(n29553) );
  CLKNAND2HSV0 U33246 ( .A1(n52693), .A2(n59355), .ZN(n29554) );
  CLKNAND2HSV0 U33247 ( .A1(n29554), .A2(n29553), .ZN(n29555) );
  OAI21HSV0 U33248 ( .A1(n29553), .A2(n29554), .B(n29555), .ZN(n29556) );
  CLKNAND2HSV0 U33249 ( .A1(n52835), .A2(n51418), .ZN(n29557) );
  CLKNAND2HSV0 U33250 ( .A1(n29557), .A2(n29556), .ZN(n29558) );
  OAI21HSV0 U33251 ( .A1(n29556), .A2(n29557), .B(n29558), .ZN(n29559) );
  CLKNAND2HSV0 U33252 ( .A1(n52669), .A2(n48841), .ZN(n29560) );
  CLKNAND2HSV0 U33253 ( .A1(n29560), .A2(n29559), .ZN(n29561) );
  OAI21HSV0 U33254 ( .A1(n29559), .A2(n29560), .B(n29561), .ZN(n29562) );
  CLKNAND2HSV0 U33255 ( .A1(n29778), .A2(n51200), .ZN(n29563) );
  CLKNAND2HSV0 U33256 ( .A1(n29563), .A2(n29562), .ZN(n29564) );
  OAI21HSV0 U33257 ( .A1(n29562), .A2(n29563), .B(n29564), .ZN(n29565) );
  CLKNAND2HSV0 U33258 ( .A1(n52668), .A2(n59905), .ZN(n29566) );
  CLKNAND2HSV0 U33259 ( .A1(n29566), .A2(n29565), .ZN(n29567) );
  OAI21HSV0 U33260 ( .A1(n29565), .A2(n29566), .B(n29567), .ZN(n29568) );
  NAND3HSV0 U33261 ( .A1(n50698), .A2(n53363), .A3(n53361), .ZN(n29569) );
  CLKNAND2HSV0 U33262 ( .A1(n29568), .A2(n29569), .ZN(n29570) );
  OAI21HSV0 U33263 ( .A1(n29568), .A2(n29569), .B(n29570), .ZN(\pe5/poht [24])
         );
  CLKNHSV0 U33264 ( .I(n51967), .ZN(n29571) );
  MUX2NHSV0 U33265 ( .I0(n29571), .I1(n51967), .S(n51813), .ZN(n29572) );
  XOR2HSV0 U33266 ( .A1(n48623), .A2(n29572), .Z(n29573) );
  CLKNAND2HSV0 U33267 ( .A1(n52901), .A2(n51797), .ZN(n29574) );
  CLKNAND2HSV0 U33268 ( .A1(n29574), .A2(n29573), .ZN(n29575) );
  OAI21HSV0 U33269 ( .A1(n29573), .A2(n29574), .B(n29575), .ZN(n29576) );
  CLKNAND2HSV0 U33270 ( .A1(n52895), .A2(n51120), .ZN(n29577) );
  CLKNAND2HSV0 U33271 ( .A1(n29577), .A2(n29576), .ZN(n29578) );
  OAI21HSV0 U33272 ( .A1(n29576), .A2(n29577), .B(n29578), .ZN(n29579) );
  CLKNAND2HSV0 U33273 ( .A1(n52902), .A2(n59351), .ZN(n29580) );
  CLKNAND2HSV0 U33274 ( .A1(n29580), .A2(n29579), .ZN(n29581) );
  OAI21HSV0 U33275 ( .A1(n29579), .A2(n29580), .B(n29581), .ZN(n29582) );
  CLKNAND2HSV0 U33276 ( .A1(n52840), .A2(n51896), .ZN(n29583) );
  CLKNAND2HSV0 U33277 ( .A1(n29583), .A2(n29582), .ZN(n29584) );
  CLKNAND2HSV0 U33278 ( .A1(n59778), .A2(n52558), .ZN(n29586) );
  CLKNAND2HSV0 U33279 ( .A1(n29586), .A2(n29585), .ZN(n29587) );
  OAI21HSV0 U33280 ( .A1(n29585), .A2(n29586), .B(n29587), .ZN(\pe2/poht [27])
         );
  CLKNAND2HSV0 U33281 ( .A1(n54541), .A2(n54728), .ZN(n29589) );
  OAI21HSV0 U33282 ( .A1(n29588), .A2(n29589), .B(n29590), .ZN(n29591) );
  CLKNAND2HSV0 U33283 ( .A1(n55228), .A2(n44530), .ZN(n29592) );
  CLKNAND2HSV0 U33284 ( .A1(n29592), .A2(n29591), .ZN(n29593) );
  OAI21HSV0 U33285 ( .A1(n29591), .A2(n29592), .B(n29593), .ZN(n29594) );
  CLKNHSV0 U33286 ( .I(n54724), .ZN(n29595) );
  OAI21HSV0 U33287 ( .A1(n55330), .A2(n29595), .B(n29594), .ZN(n29596) );
  OAI31HSV0 U33288 ( .A1(n55330), .A2(n29594), .A3(n29595), .B(n29596), .ZN(
        n29597) );
  CLKNAND2HSV0 U33289 ( .A1(n54452), .A2(n55332), .ZN(n29598) );
  CLKNAND2HSV0 U33290 ( .A1(n29598), .A2(n29597), .ZN(n29599) );
  OAI21HSV0 U33291 ( .A1(n29597), .A2(n29598), .B(n29599), .ZN(n29600) );
  CLKNAND2HSV0 U33292 ( .A1(\pe1/got [23]), .A2(n55226), .ZN(n29601) );
  CLKNAND2HSV0 U33293 ( .A1(n29601), .A2(n29600), .ZN(n29602) );
  OAI21HSV0 U33294 ( .A1(n29600), .A2(n29601), .B(n29602), .ZN(n29603) );
  CLKNAND2HSV0 U33295 ( .A1(n55593), .A2(n40913), .ZN(n29604) );
  CLKNAND2HSV0 U33296 ( .A1(n29604), .A2(n29603), .ZN(n29605) );
  OAI21HSV0 U33297 ( .A1(n29603), .A2(n29604), .B(n29605), .ZN(n29606) );
  CLKNAND2HSV0 U33298 ( .A1(n59428), .A2(\pe1/got [25]), .ZN(n29607) );
  CLKNAND2HSV0 U33299 ( .A1(n29607), .A2(n29606), .ZN(n29608) );
  OAI21HSV0 U33300 ( .A1(n29606), .A2(n29607), .B(n29608), .ZN(n29609) );
  CLKNAND2HSV0 U33301 ( .A1(n29610), .A2(n29609), .ZN(n29611) );
  OAI21HSV0 U33302 ( .A1(n29609), .A2(n29610), .B(n29611), .ZN(\pe1/poht [6])
         );
  CLKNHSV0 U33303 ( .I(\pe6/pq ), .ZN(n29612) );
  MUX2NHSV0 U33304 ( .I0(n29612), .I1(n31269), .S(n48025), .ZN(\pe6/ti_1t ) );
  CLKNAND2HSV0 U33305 ( .A1(n59393), .A2(n52694), .ZN(n29613) );
  CLKNAND2HSV0 U33306 ( .A1(n29613), .A2(n52695), .ZN(n29614) );
  OAI21HSV0 U33307 ( .A1(n52695), .A2(n29613), .B(n29614), .ZN(n60076) );
  NAND3HSV0 U33308 ( .A1(n52819), .A2(n52817), .A3(n52818), .ZN(n29615) );
  CLKNAND2HSV0 U33309 ( .A1(n29615), .A2(n52816), .ZN(n29616) );
  OAI21HSV0 U33310 ( .A1(n52816), .A2(n29615), .B(n29616), .ZN(n60032) );
  CLKNHSV0 U33311 ( .I(\pe5/pq ), .ZN(n29617) );
  MUX2NHSV0 U33312 ( .I0(n29617), .I1(n48040), .S(n53215), .ZN(\pe5/ti_1t ) );
  CLKNHSV0 U33313 ( .I(n46594), .ZN(n29618) );
  MUX2NHSV0 U33314 ( .I0(n29618), .I1(n46594), .S(n46593), .ZN(n60064) );
  CLKNHSV0 U33315 ( .I(\pe4/pq ), .ZN(n29619) );
  NAND3HSV0 U33316 ( .A1(n45798), .A2(n45796), .A3(n45797), .ZN(n29620) );
  CLKNAND2HSV0 U33317 ( .A1(n29620), .A2(n45799), .ZN(n29621) );
  OAI21HSV0 U33318 ( .A1(n45799), .A2(n29620), .B(n29621), .ZN(n60056) );
  CLKNHSV0 U33319 ( .I(n53375), .ZN(n29622) );
  CLKNHSV0 U33320 ( .I(n53373), .ZN(n29623) );
  MUX2NHSV0 U33321 ( .I0(n29623), .I1(n53373), .S(n53374), .ZN(n29624) );
  MUX2NHSV0 U33322 ( .I0(n53375), .I1(n29622), .S(n29624), .ZN(n60101) );
  AOI21HSV0 U33323 ( .A1(n52809), .A2(n52808), .B(n52810), .ZN(n29625) );
  AO31HSV0 U33324 ( .A1(n52809), .A2(n52808), .A3(n52810), .B(n29625), .Z(
        n60052) );
  INAND3HSV0 U33325 ( .A1(n25884), .B1(n52824), .B2(n52825), .ZN(n29626) );
  CLKNAND2HSV0 U33326 ( .A1(n29626), .A2(n52822), .ZN(n29627) );
  OAI21HSV0 U33327 ( .A1(n52822), .A2(n29626), .B(n29627), .ZN(n60062) );
  CLKNHSV0 U33328 ( .I(\pe2/pq ), .ZN(n29628) );
  MUX2NHSV0 U33329 ( .I0(n29628), .I1(n38126), .S(n38576), .ZN(\pe2/ti_1t ) );
  CLKNHSV0 U33330 ( .I(n48006), .ZN(n29629) );
  MUX2NHSV0 U33331 ( .I0(n29629), .I1(n48006), .S(n48005), .ZN(n29630) );
  XOR2HSV0 U33332 ( .A1(n29630), .A2(n48008), .Z(n60065) );
  OAI21HSV0 U33333 ( .A1(n52760), .A2(n52761), .B(n52762), .ZN(n29631) );
  OAI31HSV0 U33334 ( .A1(n52760), .A2(n52762), .A3(n52761), .B(n29631), .ZN(
        n60039) );
  INHSV8 U33335 ( .I(\pe4/aot [22]), .ZN(n50134) );
  INHSV8 U33336 ( .I(n50134), .ZN(n33965) );
  INHSV6 U33337 ( .I(\pe3/bq[28] ), .ZN(n45649) );
  INHSV2 U33338 ( .I(n45649), .ZN(n55867) );
  INHSV2 U33339 ( .I(n45649), .ZN(n43539) );
  INHSV4 U33340 ( .I(n45649), .ZN(n42634) );
  INHSV4 U33341 ( .I(n35058), .ZN(n47692) );
  INHSV4 U33342 ( .I(n34501), .ZN(n35201) );
  INHSV8 U33343 ( .I(\pe4/bq[24] ), .ZN(n34276) );
  INHSV4 U33344 ( .I(n34276), .ZN(n34120) );
  INHSV6 U33345 ( .I(n34276), .ZN(n50007) );
  INHSV4 U33346 ( .I(n34276), .ZN(n33712) );
  BUFHSV4 U33347 ( .I(\pe3/aot [24]), .Z(n43034) );
  BUFHSV4 U33348 ( .I(\pe3/aot [24]), .Z(n45695) );
  INHSV6 U33349 ( .I(\pe4/bq[22] ), .ZN(n50129) );
  INHSV4 U33350 ( .I(n50129), .ZN(n33711) );
  INHSV6 U33351 ( .I(n50129), .ZN(n34044) );
  INHSV8 U33352 ( .I(\pe6/bq[13] ), .ZN(n46853) );
  INHSV4 U33353 ( .I(n46853), .ZN(n59265) );
  INHSV2 U33354 ( .I(n46853), .ZN(n36143) );
  INHSV2 U33355 ( .I(n41870), .ZN(n41964) );
  INHSV4 U33356 ( .I(n41870), .ZN(n59985) );
  INHSV2 U33357 ( .I(n45461), .ZN(n39130) );
  INHSV4 U33358 ( .I(n45461), .ZN(n48755) );
  INHSV4 U33359 ( .I(n56295), .ZN(n56349) );
  CLKNHSV6 U33360 ( .I(n56295), .ZN(n42950) );
  CLKNHSV6 U33361 ( .I(\pe3/aot [18]), .ZN(n56295) );
  INHSV6 U33362 ( .I(\pe4/aot [4]), .ZN(n57011) );
  INHSV6 U33363 ( .I(\pe1/aot [9]), .ZN(n54472) );
  INHSV2 U33364 ( .I(n54472), .ZN(n54978) );
  BUFHSV4 U33365 ( .I(\pe3/bq[25] ), .Z(n42527) );
  INHSV8 U33366 ( .I(\pe4/aot [20]), .ZN(n49982) );
  INHSV6 U33367 ( .I(n49982), .ZN(n59839) );
  INHSV6 U33368 ( .I(n49982), .ZN(n34743) );
  INHSV8 U33369 ( .I(\pe5/bq[24] ), .ZN(n30452) );
  INHSV4 U33370 ( .I(n30452), .ZN(n30341) );
  INHSV6 U33371 ( .I(n30452), .ZN(n30891) );
  INHSV2 U33372 ( .I(n34249), .ZN(n47658) );
  INHSV6 U33373 ( .I(\pe2/bq[26] ), .ZN(n49518) );
  INHSV6 U33374 ( .I(n49518), .ZN(n38064) );
  INHSV8 U33375 ( .I(\pe1/bq[25] ), .ZN(n42264) );
  INHSV4 U33376 ( .I(n47661), .ZN(n35533) );
  CLKNHSV6 U33377 ( .I(\pe3/aot [20]), .ZN(n37357) );
  INHSV12 U33378 ( .I(n37357), .ZN(n56204) );
  INHSV4 U33379 ( .I(n38418), .ZN(n36590) );
  INHSV4 U33380 ( .I(n38418), .ZN(n53015) );
  INHSV2 U33381 ( .I(n38418), .ZN(n38303) );
  INHSV8 U33382 ( .I(\pe2/aot [29]), .ZN(n38787) );
  INHSV8 U33383 ( .I(\pe6/bq[25] ), .ZN(n36132) );
  INHSV4 U33384 ( .I(n36132), .ZN(n46624) );
  CLKNHSV6 U33385 ( .I(n36132), .ZN(n59206) );
  INHSV6 U33386 ( .I(n41442), .ZN(n40898) );
  INHSV8 U33387 ( .I(\pe2/aot [26]), .ZN(n44049) );
  INHSV6 U33388 ( .I(n44049), .ZN(n52974) );
  INHSV6 U33389 ( .I(\pe1/aot [21]), .ZN(n41944) );
  INHSV4 U33390 ( .I(n41944), .ZN(n59987) );
  INHSV4 U33391 ( .I(\pe4/aot [24]), .ZN(n57326) );
  INHSV4 U33392 ( .I(n57326), .ZN(n57727) );
  INHSV4 U33393 ( .I(n33467), .ZN(n33726) );
  INHSV6 U33394 ( .I(n59105), .ZN(n36150) );
  CLKNHSV6 U33395 ( .I(n59105), .ZN(n33023) );
  CLKNHSV6 U33396 ( .I(n50008), .ZN(n59951) );
  INHSV2 U33397 ( .I(n36123), .ZN(n59251) );
  INHSV2 U33398 ( .I(n36123), .ZN(n35760) );
  INHSV6 U33399 ( .I(n35175), .ZN(n57014) );
  INHSV4 U33400 ( .I(n40236), .ZN(n39629) );
  INHSV8 U33401 ( .I(\pe3/bq[21] ), .ZN(n43039) );
  INHSV2 U33402 ( .I(n43039), .ZN(n56218) );
  INHSV4 U33403 ( .I(n43039), .ZN(n56106) );
  INHSV4 U33404 ( .I(n43039), .ZN(n49439) );
  INHSV4 U33405 ( .I(n55714), .ZN(n48530) );
  INHSV8 U33406 ( .I(\pe5/bq[25] ), .ZN(n30287) );
  INHSV4 U33407 ( .I(n30287), .ZN(n30526) );
  INHSV4 U33408 ( .I(n30287), .ZN(n52585) );
  INHSV6 U33409 ( .I(\pe6/bq[16] ), .ZN(n58984) );
  INHSV4 U33410 ( .I(n58984), .ZN(n58833) );
  INHSV4 U33411 ( .I(n58984), .ZN(n49844) );
  CLKNHSV6 U33412 ( .I(n51736), .ZN(n53005) );
  INHSV4 U33413 ( .I(n35653), .ZN(n59247) );
  INHSV4 U33414 ( .I(n35647), .ZN(n59267) );
  CLKNHSV6 U33415 ( .I(n57030), .ZN(n57234) );
  CLKNHSV6 U33416 ( .I(n57030), .ZN(n59952) );
  INHSV6 U33417 ( .I(\pe6/aot [12]), .ZN(n49188) );
  INHSV2 U33418 ( .I(n49188), .ZN(n58631) );
  INHSV4 U33419 ( .I(n49188), .ZN(n53115) );
  INHSV4 U33420 ( .I(n49188), .ZN(n32972) );
  BUFHSV4 U33421 ( .I(\pe4/bq[21] ), .Z(n57505) );
  BUFHSV8 U33422 ( .I(n34254), .Z(n33969) );
  BUFHSV8 U33423 ( .I(\pe4/bq[21] ), .Z(n34254) );
  BUFHSV4 U33424 ( .I(n36574), .Z(n36560) );
  BUFHSV4 U33425 ( .I(n36560), .Z(n38454) );
  CLKNHSV0 U33426 ( .I(n48015), .ZN(n59490) );
  BUFHSV2 U33427 ( .I(n37017), .Z(n37177) );
  INHSV8 U33428 ( .I(\pe2/aot [21]), .ZN(n47575) );
  INHSV6 U33429 ( .I(n47575), .ZN(n59758) );
  INHSV4 U33430 ( .I(n47575), .ZN(n52104) );
  INHSV4 U33431 ( .I(n44889), .ZN(n36603) );
  INHSV6 U33432 ( .I(\pe5/ti_1 ), .ZN(n29826) );
  BUFHSV8 U33433 ( .I(n47499), .Z(n49606) );
  INHSV4 U33434 ( .I(n49606), .ZN(n51893) );
  INHSV4 U33435 ( .I(n49606), .ZN(n51798) );
  BUFHSV4 U33436 ( .I(n32193), .Z(n32714) );
  INHSV4 U33437 ( .I(n33113), .ZN(n33611) );
  INHSV4 U33438 ( .I(\pe3/aot [32]), .ZN(n42821) );
  INHSV6 U33439 ( .I(\pe5/bq[21] ), .ZN(n45460) );
  INHSV6 U33440 ( .I(\pe4/aot [19]), .ZN(n57605) );
  INHSV4 U33441 ( .I(n46126), .ZN(n37007) );
  INHSV4 U33442 ( .I(n46126), .ZN(n37051) );
  INHSV6 U33443 ( .I(ctro3), .ZN(n36682) );
  INHSV2 U33444 ( .I(\pe6/got [32]), .ZN(n31256) );
  INHSV6 U33445 ( .I(\pe2/bq[22] ), .ZN(n52430) );
  INHSV4 U33446 ( .I(n52430), .ZN(n38054) );
  CLKNHSV6 U33447 ( .I(ctro4), .ZN(n33097) );
  CLKNHSV6 U33448 ( .I(n33339), .ZN(n33848) );
  INHSV6 U33449 ( .I(\pe6/aot [28]), .ZN(n35816) );
  INHSV6 U33450 ( .I(n44053), .ZN(n39061) );
  INHSV4 U33451 ( .I(n44053), .ZN(n36409) );
  BUFHSV4 U33452 ( .I(n50400), .Z(n57819) );
  BUFHSV8 U33453 ( .I(n50400), .Z(n47841) );
  INHSV4 U33454 ( .I(n35092), .ZN(n35194) );
  INHSV6 U33455 ( .I(n35092), .ZN(n33966) );
  INHSV6 U33456 ( .I(n35092), .ZN(n48069) );
  INHSV6 U33457 ( .I(\pe4/bq[27] ), .ZN(n35084) );
  INHSV4 U33458 ( .I(n35084), .ZN(n33427) );
  INHSV8 U33459 ( .I(\pe4/bq[16] ), .ZN(n48024) );
  INHSV4 U33460 ( .I(n48024), .ZN(n49943) );
  INHSV4 U33461 ( .I(n34485), .ZN(n57134) );
  INHSV4 U33462 ( .I(n34485), .ZN(n34021) );
  INHSV4 U33463 ( .I(n34485), .ZN(n46617) );
  INHSV6 U33464 ( .I(n48934), .ZN(n52998) );
  BUFHSV8 U33465 ( .I(n41334), .Z(n41967) );
  INHSV6 U33466 ( .I(n41334), .ZN(n40890) );
  INHSV4 U33467 ( .I(n41967), .ZN(n40684) );
  INHSV2 U33468 ( .I(n42264), .ZN(n41173) );
  INHSV2 U33469 ( .I(n43623), .ZN(n37180) );
  INHSV4 U33470 ( .I(n43623), .ZN(n46614) );
  INHSV6 U33471 ( .I(\pe2/bq[24] ), .ZN(n38687) );
  INHSV4 U33472 ( .I(n38687), .ZN(n38053) );
  INHSV6 U33473 ( .I(n40501), .ZN(n41334) );
  INHSV4 U33474 ( .I(n41334), .ZN(n41083) );
  INHSV6 U33475 ( .I(\pe1/bq[22] ), .ZN(n41947) );
  INHSV4 U33476 ( .I(n48393), .ZN(n54465) );
  INHSV4 U33477 ( .I(n41947), .ZN(n54302) );
  INHSV4 U33478 ( .I(ctro4), .ZN(n33687) );
  INHSV4 U33479 ( .I(n33093), .ZN(n33094) );
  INHSV8 U33480 ( .I(n48450), .ZN(n40873) );
  INHSV8 U33481 ( .I(\pe1/aot [15]), .ZN(n42361) );
  INHSV4 U33482 ( .I(n42361), .ZN(n55186) );
  INHSV6 U33483 ( .I(n48056), .ZN(n57476) );
  INHSV8 U33484 ( .I(\pe1/got [29]), .ZN(n40719) );
  BUFHSV4 U33485 ( .I(\pe5/bq[11] ), .Z(n39592) );
  INHSV8 U33486 ( .I(\pe6/aot [22]), .ZN(n32373) );
  INHSV4 U33487 ( .I(n32373), .ZN(n49831) );
  INHSV4 U33488 ( .I(n39166), .ZN(n31192) );
  INHSV4 U33489 ( .I(n39166), .ZN(n30789) );
  INHSV4 U33490 ( .I(n39166), .ZN(n30616) );
  INHSV6 U33491 ( .I(\pe5/aot [19]), .ZN(n31029) );
  INHSV6 U33492 ( .I(n38946), .ZN(n51759) );
  INHSV2 U33493 ( .I(\pe3/aot [13]), .ZN(n56382) );
  INHSV4 U33494 ( .I(n43151), .ZN(n43280) );
  INHSV8 U33495 ( .I(\pe5/bq[20] ), .ZN(n45426) );
  INHSV4 U33496 ( .I(n45426), .ZN(n48237) );
  INHSV4 U33497 ( .I(n45426), .ZN(n39487) );
  INHSV6 U33498 ( .I(\pe4/bq[7] ), .ZN(n50114) );
  INHSV4 U33499 ( .I(n50114), .ZN(n58003) );
  INHSV4 U33500 ( .I(n50114), .ZN(n58197) );
  INHSV2 U33501 ( .I(n50837), .ZN(n33022) );
  INHSV2 U33502 ( .I(n50837), .ZN(n59239) );
  INHSV8 U33503 ( .I(\pe2/aot [18]), .ZN(n52103) );
  INHSV8 U33504 ( .I(\pe6/bq[15] ), .ZN(n48047) );
  INHSV4 U33505 ( .I(n48047), .ZN(n35751) );
  INHSV4 U33506 ( .I(n48047), .ZN(n58682) );
  INHSV4 U33507 ( .I(n48047), .ZN(n59045) );
  INHSV6 U33508 ( .I(\pe5/bq[22] ), .ZN(n45844) );
  INHSV2 U33509 ( .I(n45844), .ZN(n47059) );
  BUFHSV2 U33510 ( .I(n32053), .Z(n31624) );
  INHSV8 U33511 ( .I(\pe6/bq[12] ), .ZN(n59094) );
  INHSV6 U33512 ( .I(n59094), .ZN(n48051) );
  INHSV6 U33513 ( .I(n59094), .ZN(n58976) );
  INHSV8 U33514 ( .I(\pe5/bq[9] ), .ZN(n47162) );
  INHSV6 U33515 ( .I(n47162), .ZN(n48775) );
  INHSV4 U33516 ( .I(n47162), .ZN(n51307) );
  INHSV4 U33517 ( .I(n47162), .ZN(n50533) );
  INHSV4 U33518 ( .I(n43392), .ZN(n43265) );
  INHSV2 U33519 ( .I(n43392), .ZN(n43547) );
  INHSV2 U33520 ( .I(n37933), .ZN(n45149) );
  BUFHSV4 U33521 ( .I(n45149), .Z(n39011) );
  BUFHSV4 U33522 ( .I(n45149), .Z(n44185) );
  BUFHSV4 U33523 ( .I(n36575), .Z(n45267) );
  BUFHSV4 U33524 ( .I(n36575), .Z(n36319) );
  INHSV6 U33525 ( .I(\pe2/bq[25] ), .ZN(n44854) );
  INHSV6 U33526 ( .I(n44854), .ZN(n44987) );
  INHSV6 U33527 ( .I(n44854), .ZN(n52950) );
  INHSV8 U33528 ( .I(\pe1/bq[12] ), .ZN(n53691) );
  INHSV12 U33529 ( .I(n53691), .ZN(n42373) );
  INHSV6 U33530 ( .I(\pe1/aot [13]), .ZN(n53672) );
  INHSV2 U33531 ( .I(n53672), .ZN(n59990) );
  INHSV2 U33532 ( .I(n53672), .ZN(n44541) );
  BUFHSV8 U33533 ( .I(\pe6/bq[14] ), .Z(n58668) );
  INHSV6 U33534 ( .I(n59869), .ZN(n52600) );
  INHSV6 U33535 ( .I(\pe3/bq[9] ), .ZN(n56277) );
  INHSV4 U33536 ( .I(n56277), .ZN(n56785) );
  INHSV4 U33537 ( .I(n56277), .ZN(n53232) );
  INHSV6 U33538 ( .I(\pe5/aot [24]), .ZN(n44704) );
  INHSV2 U33539 ( .I(n44704), .ZN(n39499) );
  INHSV2 U33540 ( .I(n44704), .ZN(n37660) );
  INHSV6 U33541 ( .I(\pe1/bq[27] ), .ZN(n41425) );
  CLKNHSV6 U33542 ( .I(n41425), .ZN(n41771) );
  INHSV4 U33543 ( .I(n41425), .ZN(n40494) );
  INHSV8 U33544 ( .I(n42835), .ZN(n56464) );
  BUFHSV4 U33545 ( .I(n40547), .Z(n40952) );
  INHSV6 U33546 ( .I(\pe5/bq[13] ), .ZN(n48050) );
  INHSV4 U33547 ( .I(n48050), .ZN(n39471) );
  INHSV8 U33548 ( .I(n48050), .ZN(n50668) );
  BUFHSV4 U33549 ( .I(\pe4/bq[4] ), .Z(n57498) );
  BUFHSV8 U33550 ( .I(\pe4/bq[4] ), .Z(n57595) );
  INHSV4 U33551 ( .I(n39796), .ZN(n52610) );
  INHSV8 U33552 ( .I(\pe3/aot [21]), .ZN(n42539) );
  INHSV6 U33553 ( .I(n42539), .ZN(n42940) );
  INHSV4 U33554 ( .I(n42539), .ZN(n56182) );
  INHSV2 U33555 ( .I(n37265), .ZN(n36671) );
  INHSV4 U33556 ( .I(\pe2/bq[14] ), .ZN(n47580) );
  INHSV2 U33557 ( .I(\pe1/bq[9] ), .ZN(n55385) );
  BUFHSV8 U33558 ( .I(\pe1/bq[4] ), .Z(n55544) );
  BUFHSV4 U33559 ( .I(n38899), .Z(n38630) );
  BUFHSV4 U33560 ( .I(n38195), .Z(n45099) );
  INHSV6 U33561 ( .I(n38630), .ZN(n44309) );
  INHSV4 U33562 ( .I(n35487), .ZN(n34416) );
  INHSV4 U33563 ( .I(n40969), .ZN(n40466) );
  BUFHSV8 U33564 ( .I(ctro2), .Z(n38899) );
  INHSV6 U33565 ( .I(n36553), .ZN(n36377) );
  INHSV4 U33566 ( .I(n36397), .ZN(n36398) );
  INHSV4 U33567 ( .I(n54829), .ZN(n54900) );
  INHSV4 U33568 ( .I(n57918), .ZN(n57852) );
  INHSV4 U33569 ( .I(n57918), .ZN(n59953) );
  INHSV6 U33570 ( .I(\pe3/got [27]), .ZN(n42683) );
  INHSV2 U33571 ( .I(n37784), .ZN(n59963) );
  INHSV6 U33572 ( .I(\pe2/aot [15]), .ZN(n47503) );
  CLKNHSV6 U33573 ( .I(n47503), .ZN(n59974) );
  INHSV4 U33574 ( .I(n47503), .ZN(n52070) );
  INHSV4 U33575 ( .I(n44532), .ZN(n41802) );
  BUFHSV4 U33576 ( .I(\pe1/ctrq ), .Z(n48054) );
  BUFHSV4 U33577 ( .I(\pe1/ctrq ), .Z(n48080) );
  BUFHSV8 U33578 ( .I(\pe1/ctrq ), .Z(n48061) );
  CLKNHSV0 U33579 ( .I(n48015), .ZN(n59492) );
  BUFHSV2 U33580 ( .I(n59582), .Z(n44892) );
  BUFHSV4 U33581 ( .I(n44832), .Z(n52920) );
  INHSV4 U33582 ( .I(n51121), .ZN(n44968) );
  BUFHSV4 U33583 ( .I(n46825), .Z(n46769) );
  BUFHSV4 U33584 ( .I(n46825), .Z(n58718) );
  CLKNAND2HSV4 U33585 ( .A1(n35784), .A2(n35778), .ZN(n46825) );
  INHSV4 U33586 ( .I(n38119), .ZN(n45150) );
  INHSV2 U33587 ( .I(n38119), .ZN(n52288) );
  INHSV6 U33588 ( .I(\pe1/bq[24] ), .ZN(n54185) );
  INHSV4 U33589 ( .I(n44095), .ZN(n49530) );
  INHSV4 U33590 ( .I(n44095), .ZN(n52310) );
  BUFHSV8 U33591 ( .I(n32286), .Z(n59038) );
  BUFHSV4 U33592 ( .I(n49726), .Z(n58601) );
  INHSV2 U33593 ( .I(n47394), .ZN(n51273) );
  INHSV4 U33594 ( .I(n38213), .ZN(n38401) );
  BUFHSV4 U33595 ( .I(n57308), .Z(n58096) );
  BUFHSV4 U33596 ( .I(n57308), .Z(n58029) );
  BUFHSV4 U33597 ( .I(n59665), .Z(n35577) );
  BUFHSV4 U33598 ( .I(n59526), .Z(n57550) );
  INHSV2 U33599 ( .I(n43372), .ZN(n56562) );
  BUFHSV8 U33600 ( .I(n32167), .Z(n35813) );
  BUFHSV8 U33601 ( .I(n35813), .Z(n59183) );
  BUFHSV8 U33602 ( .I(n35813), .Z(n59597) );
  BUFHSV8 U33603 ( .I(n35917), .Z(n35796) );
  INHSV6 U33604 ( .I(\pe6/got [31]), .ZN(n35917) );
  INHSV4 U33605 ( .I(n59339), .ZN(n32530) );
  INHSV4 U33606 ( .I(n31269), .ZN(n59236) );
  INHSV4 U33607 ( .I(n31269), .ZN(n33016) );
  BUFHSV4 U33608 ( .I(n49667), .Z(n46632) );
  INHSV4 U33609 ( .I(n46145), .ZN(n49316) );
  INHSV4 U33610 ( .I(n49316), .ZN(n59024) );
  INHSV4 U33611 ( .I(n49316), .ZN(n58575) );
  INHSV2 U33612 ( .I(n45924), .ZN(n29778) );
  INHSV2 U33613 ( .I(n45924), .ZN(n29779) );
  BUFHSV4 U33614 ( .I(n53979), .Z(n41549) );
  BUFHSV4 U33615 ( .I(n41549), .Z(n42210) );
  INHSV4 U33616 ( .I(n56420), .ZN(n56340) );
  BUFHSV4 U33617 ( .I(n53228), .Z(n55947) );
  BUFHSV4 U33618 ( .I(n53228), .Z(n56624) );
  BUFHSV4 U33619 ( .I(n47770), .Z(n50298) );
  INHSV4 U33620 ( .I(n47770), .ZN(n59574) );
  INHSV4 U33621 ( .I(n46823), .ZN(n53109) );
  INHSV2 U33622 ( .I(n46532), .ZN(n43463) );
  INHSV6 U33623 ( .I(\pe2/bq[17] ), .ZN(n44844) );
  INHSV6 U33624 ( .I(n44844), .ZN(n44074) );
  INHSV4 U33625 ( .I(n37555), .ZN(n40172) );
  INHSV4 U33626 ( .I(n37555), .ZN(n48624) );
  INHSV4 U33627 ( .I(n44520), .ZN(n39230) );
  BUFHSV4 U33628 ( .I(n40567), .Z(n41333) );
  INHSV6 U33629 ( .I(n41333), .ZN(n41160) );
  INHSV6 U33630 ( .I(\pe5/got [29]), .ZN(n40130) );
  INHSV4 U33631 ( .I(n48023), .ZN(n57785) );
  BUFHSV4 U33632 ( .I(n45794), .Z(n43869) );
  INHSV2 U33633 ( .I(n30887), .ZN(n39466) );
  INHSV4 U33634 ( .I(n32723), .ZN(n44446) );
  INHSV6 U33635 ( .I(\pe6/bq[24] ), .ZN(n59194) );
  INHSV4 U33636 ( .I(n59194), .ZN(n59050) );
  BUFHSV2 U33637 ( .I(n53218), .Z(n48072) );
  BUFHSV4 U33638 ( .I(n45517), .Z(n43755) );
  BUFHSV8 U33639 ( .I(n46156), .Z(n49181) );
  NAND2HSV4 U33640 ( .A1(n45791), .A2(n45790), .ZN(n46156) );
  BUFHSV4 U33641 ( .I(n49181), .Z(n58576) );
  INHSV4 U33642 ( .I(n49401), .ZN(n59514) );
  INHSV4 U33643 ( .I(n47145), .ZN(n59903) );
  INHSV4 U33644 ( .I(n51217), .ZN(n48745) );
  INHSV8 U33645 ( .I(\pe6/aot [27]), .ZN(n32589) );
  INHSV4 U33646 ( .I(n53227), .ZN(n50757) );
  INHSV4 U33647 ( .I(n54631), .ZN(n54154) );
  INHSV2 U33648 ( .I(n54631), .ZN(n53513) );
  INHSV8 U33649 ( .I(\pe4/aot [23]), .ZN(n46143) );
  INHSV4 U33650 ( .I(n46143), .ZN(n33716) );
  INHSV4 U33651 ( .I(n39716), .ZN(n39992) );
  AND2HSV2 U33652 ( .A1(n45273), .A2(n47997), .Z(n29633) );
  INHSV6 U33653 ( .I(\pe4/aot [25]), .ZN(n57026) );
  BUFHSV4 U33654 ( .I(\pe2/ctrq ), .Z(n37952) );
  INHSV2 U33655 ( .I(n44884), .ZN(n36380) );
  BUFHSV4 U33656 ( .I(n39745), .Z(n40171) );
  BUFHSV4 U33657 ( .I(n25854), .Z(n39745) );
  INHSV4 U33658 ( .I(n47920), .ZN(n59348) );
  BUFHSV8 U33659 ( .I(\pe5/got [32]), .Z(n37544) );
  INHSV6 U33660 ( .I(n37544), .ZN(n39733) );
  INHSV6 U33661 ( .I(\pe2/aot [24]), .ZN(n38655) );
  INHSV4 U33662 ( .I(n38655), .ZN(n59972) );
  INHSV4 U33663 ( .I(\pe4/bq[18] ), .ZN(n48026) );
  INHSV4 U33664 ( .I(n39143), .ZN(n39278) );
  INHSV2 U33665 ( .I(n39143), .ZN(n30806) );
  INHSV6 U33666 ( .I(n30106), .ZN(n59393) );
  INHSV4 U33667 ( .I(n39143), .ZN(n30377) );
  INHSV8 U33668 ( .I(n50947), .ZN(n39052) );
  INHSV6 U33669 ( .I(\pe1/aot [28]), .ZN(n53447) );
  INHSV12 U33670 ( .I(n53447), .ZN(n40683) );
  INHSV6 U33671 ( .I(\pe6/bq[21] ), .ZN(n59205) );
  INHSV4 U33672 ( .I(n59205), .ZN(n32568) );
  INHSV4 U33673 ( .I(n59205), .ZN(n32172) );
  INHSV8 U33674 ( .I(\pe6/bq[1] ), .ZN(n48887) );
  INHSV2 U33675 ( .I(n48887), .ZN(n58990) );
  INHSV4 U33676 ( .I(n35817), .ZN(n31829) );
  BUFHSV6 U33677 ( .I(n30255), .Z(n39583) );
  BUFHSV8 U33678 ( .I(n39583), .Z(n31151) );
  INHSV2 U33679 ( .I(n50822), .ZN(n44435) );
  INHSV2 U33680 ( .I(n50822), .ZN(n59100) );
  INHSV6 U33681 ( .I(\pe2/bq[16] ), .ZN(n48063) );
  INHSV6 U33682 ( .I(n48063), .ZN(n38803) );
  BUFHSV8 U33683 ( .I(\pe3/aot [23]), .Z(n42818) );
  BUFHSV4 U33684 ( .I(\pe3/aot [23]), .Z(n59612) );
  INHSV6 U33685 ( .I(\pe1/aot [20]), .ZN(n41650) );
  INHSV6 U33686 ( .I(n41650), .ZN(n54669) );
  BUFHSV4 U33687 ( .I(n36574), .Z(n38629) );
  INHSV4 U33688 ( .I(n48331), .ZN(n40654) );
  INHSV2 U33689 ( .I(n57025), .ZN(n33867) );
  INHSV4 U33690 ( .I(n57025), .ZN(n59605) );
  INHSV6 U33691 ( .I(n57025), .ZN(n57218) );
  INHSV2 U33692 ( .I(n40785), .ZN(n41609) );
  INHSV4 U33693 ( .I(n40785), .ZN(n41144) );
  INHSV2 U33694 ( .I(n43757), .ZN(n37362) );
  INHSV2 U33695 ( .I(n43757), .ZN(n48496) );
  BUFHSV4 U33696 ( .I(n37659), .Z(n37558) );
  INHSV8 U33697 ( .I(\pe5/bq[28] ), .ZN(n30116) );
  INHSV2 U33698 ( .I(n30116), .ZN(n48802) );
  INHSV8 U33699 ( .I(\pe2/bq[29] ), .ZN(n36389) );
  INHSV8 U33700 ( .I(n36389), .ZN(n36608) );
  INHSV8 U33701 ( .I(\pe1/aot [31]), .ZN(n40445) );
  INHSV2 U33702 ( .I(n46192), .ZN(n59217) );
  INHSV4 U33703 ( .I(n46192), .ZN(n32252) );
  BUFHSV4 U33704 ( .I(n31791), .Z(n46192) );
  INHSV6 U33705 ( .I(\pe6/bq[26] ), .ZN(n31791) );
  INHSV4 U33706 ( .I(\pe2/aot [8]), .ZN(n47518) );
  INHSV4 U33707 ( .I(n47518), .ZN(n52951) );
  INHSV8 U33708 ( .I(\pe6/bq[20] ), .ZN(n35837) );
  INHSV4 U33709 ( .I(n35837), .ZN(n33005) );
  INHSV4 U33710 ( .I(n35837), .ZN(n59098) );
  INHSV4 U33711 ( .I(n35837), .ZN(n32606) );
  INHSV2 U33712 ( .I(n31560), .ZN(n32576) );
  INHSV6 U33713 ( .I(\pe3/aot [26]), .ZN(n45564) );
  INHSV4 U33714 ( .I(n45564), .ZN(n55988) );
  INHSV4 U33715 ( .I(n45564), .ZN(n42743) );
  INHSV6 U33716 ( .I(\pe1/aot [24]), .ZN(n41974) );
  INHSV8 U33717 ( .I(n41974), .ZN(n54307) );
  INHSV2 U33718 ( .I(n57605), .ZN(n57140) );
  INHSV4 U33719 ( .I(n57605), .ZN(n50215) );
  BUFHSV2 U33720 ( .I(n46123), .Z(n32218) );
  INHSV6 U33721 ( .I(\pe1/bq[26] ), .ZN(n53553) );
  INHSV6 U33722 ( .I(n53553), .ZN(n41644) );
  INHSV4 U33723 ( .I(n53553), .ZN(n40557) );
  INHSV8 U33724 ( .I(\pe1/aot [22]), .ZN(n41885) );
  INHSV6 U33725 ( .I(n41885), .ZN(n54078) );
  INHSV6 U33726 ( .I(n41885), .ZN(n41169) );
  INHSV6 U33727 ( .I(\pe2/aot [11]), .ZN(n47524) );
  INHSV6 U33728 ( .I(n47524), .ZN(n59976) );
  INHSV4 U33729 ( .I(n31667), .ZN(n31373) );
  INHSV6 U33730 ( .I(\pe2/aot [23]), .ZN(n47574) );
  INHSV4 U33731 ( .I(n47574), .ZN(n50930) );
  INHSV4 U33732 ( .I(n47574), .ZN(n59585) );
  INHSV8 U33733 ( .I(\pe5/bq[23] ), .ZN(n37564) );
  INHSV4 U33734 ( .I(n37564), .ZN(n31160) );
  INHSV4 U33735 ( .I(n30452), .ZN(n30692) );
  INHSV4 U33736 ( .I(n44332), .ZN(n39654) );
  INHSV2 U33737 ( .I(n38418), .ZN(n38549) );
  INHSV4 U33738 ( .I(n45460), .ZN(n46933) );
  INHSV2 U33739 ( .I(n45460), .ZN(n39445) );
  BUFHSV4 U33740 ( .I(n54814), .Z(n53392) );
  BUFHSV4 U33741 ( .I(n41847), .Z(n54814) );
  BUFHSV4 U33742 ( .I(n54814), .Z(n42358) );
  INHSV6 U33743 ( .I(\pe6/bq[18] ), .ZN(n59105) );
  BUFHSV2 U33744 ( .I(n33111), .Z(n35068) );
  INHSV4 U33745 ( .I(n33111), .ZN(n34738) );
  INHSV6 U33746 ( .I(n33111), .ZN(n33103) );
  BUFHSV4 U33747 ( .I(\pe5/bq[10] ), .Z(n48170) );
  INHSV6 U33748 ( .I(\pe6/bq[4] ), .ZN(n46642) );
  INHSV6 U33749 ( .I(n46642), .ZN(n59062) );
  INHSV4 U33750 ( .I(n46642), .ZN(n49106) );
  INHSV6 U33751 ( .I(\pe1/bq[15] ), .ZN(n54973) );
  INHSV4 U33752 ( .I(n29826), .ZN(n37584) );
  INHSV2 U33753 ( .I(n48040), .ZN(n30693) );
  INHSV6 U33754 ( .I(\pe2/aot [14]), .ZN(n45165) );
  INHSV4 U33755 ( .I(n45165), .ZN(n44745) );
  INHSV4 U33756 ( .I(n45165), .ZN(n59636) );
  INHSV4 U33757 ( .I(n45165), .ZN(n51920) );
  INHSV4 U33758 ( .I(n44403), .ZN(n59054) );
  INHSV4 U33759 ( .I(n43527), .ZN(n46363) );
  BUFHSV4 U33760 ( .I(n40411), .Z(n41622) );
  BUFHSV4 U33761 ( .I(n59379), .Z(n59033) );
  INHSV4 U33762 ( .I(\pe6/got [18]), .ZN(n46270) );
  INHSV4 U33763 ( .I(n48347), .ZN(n53805) );
  INHSV2 U33764 ( .I(n48347), .ZN(n41623) );
  INHSV2 U33765 ( .I(n34537), .ZN(n57183) );
  INHSV4 U33766 ( .I(n34537), .ZN(n34405) );
  BUFHSV4 U33767 ( .I(\pe3/bq[24] ), .Z(n42530) );
  INHSV6 U33768 ( .I(\pe6/bq[17] ), .ZN(n46688) );
  INHSV8 U33769 ( .I(n46688), .ZN(n32982) );
  BUFHSV4 U33770 ( .I(n44185), .Z(n52932) );
  CLKNHSV0 U33771 ( .I(n32970), .ZN(n32631) );
  BUFHSV4 U33772 ( .I(\pe6/got [24]), .Z(n31717) );
  BUFHSV6 U33773 ( .I(\pe6/got [24]), .Z(n32970) );
  BUFHSV4 U33774 ( .I(n49318), .Z(n53113) );
  BUFHSV4 U33775 ( .I(n49318), .Z(n58938) );
  BUFHSV4 U33776 ( .I(n49318), .Z(n58664) );
  INHSV6 U33777 ( .I(\pe3/aot [2]), .ZN(n56956) );
  INHSV2 U33778 ( .I(n36530), .ZN(n39032) );
  INHSV4 U33779 ( .I(n36530), .ZN(n38394) );
  INHSV4 U33780 ( .I(n36530), .ZN(n38047) );
  INHSV8 U33781 ( .I(\pe1/bq[11] ), .ZN(n48030) );
  INHSV4 U33782 ( .I(n48030), .ZN(n54311) );
  INHSV4 U33783 ( .I(n48030), .ZN(n55166) );
  INHSV4 U33784 ( .I(n49265), .ZN(n56508) );
  INHSV4 U33785 ( .I(n43178), .ZN(n45645) );
  INHSV4 U33786 ( .I(n45662), .ZN(n59816) );
  INHSV8 U33787 ( .I(\pe3/aot [5]), .ZN(n45662) );
  INHSV6 U33788 ( .I(\pe6/aot [23]), .ZN(n49699) );
  INHSV4 U33789 ( .I(n49699), .ZN(n36153) );
  INHSV4 U33790 ( .I(\pe3/got [32]), .ZN(n43467) );
  INHSV4 U33791 ( .I(n36704), .ZN(n59962) );
  INHSV8 U33792 ( .I(\pe3/aot [10]), .ZN(n47447) );
  INHSV4 U33793 ( .I(n47447), .ZN(n56740) );
  INHSV4 U33794 ( .I(n47447), .ZN(n59960) );
  BUFHSV8 U33795 ( .I(\pe3/aot [14]), .Z(n56188) );
  BUFHSV2 U33796 ( .I(n40525), .Z(n42067) );
  INHSV4 U33797 ( .I(n41701), .ZN(n40668) );
  INHSV8 U33798 ( .I(\pe2/bq[8] ), .ZN(n51567) );
  CLKNHSV6 U33799 ( .I(n51057), .ZN(n39914) );
  INHSV4 U33800 ( .I(n51057), .ZN(n53314) );
  INHSV4 U33801 ( .I(n44699), .ZN(n38393) );
  BUFHSV4 U33802 ( .I(n38823), .Z(n44699) );
  INHSV6 U33803 ( .I(n38823), .ZN(n39020) );
  INHSV4 U33804 ( .I(\pe3/bq[14] ), .ZN(n49281) );
  INHSV6 U33805 ( .I(n49281), .ZN(n48499) );
  INHSV4 U33806 ( .I(\pe1/bq[14] ), .ZN(n54281) );
  INHSV4 U33807 ( .I(n54281), .ZN(n41641) );
  INHSV6 U33808 ( .I(\pe5/aot [15]), .ZN(n48823) );
  INHSV6 U33809 ( .I(\pe5/got [22]), .ZN(n47140) );
  INHSV6 U33810 ( .I(n54879), .ZN(n55337) );
  INHSV4 U33811 ( .I(\pe2/bq[6] ), .ZN(n44718) );
  INHSV2 U33812 ( .I(\pe4/aot [14]), .ZN(n34470) );
  INHSV4 U33813 ( .I(n46609), .ZN(n42360) );
  INHSV4 U33814 ( .I(n40952), .ZN(n41712) );
  INHSV4 U33815 ( .I(n40437), .ZN(n48331) );
  INHSV6 U33816 ( .I(\pe2/aot [13]), .ZN(n38822) );
  INHSV4 U33817 ( .I(n48032), .ZN(n57837) );
  INHSV4 U33818 ( .I(n30223), .ZN(n39436) );
  INHSV4 U33819 ( .I(n30223), .ZN(n30698) );
  INHSV6 U33820 ( .I(\pe1/aot [2]), .ZN(n55504) );
  INHSV2 U33821 ( .I(n55504), .ZN(n55595) );
  BUFHSV8 U33822 ( .I(n33097), .Z(n33779) );
  BUFHSV4 U33823 ( .I(n41701), .Z(n48320) );
  INHSV6 U33824 ( .I(\pe1/got [31]), .ZN(n40335) );
  BUFHSV4 U33825 ( .I(n40525), .Z(n41701) );
  BUFHSV8 U33826 ( .I(\pe6/got [4]), .Z(n46173) );
  INHSV8 U33827 ( .I(\pe5/bq[17] ), .ZN(n45821) );
  INHSV6 U33828 ( .I(n45821), .ZN(n51176) );
  INHSV4 U33829 ( .I(n45821), .ZN(n48236) );
  INHSV6 U33830 ( .I(\pe2/bq[18] ), .ZN(n48064) );
  INHSV12 U33831 ( .I(n48064), .ZN(n52988) );
  INHSV6 U33832 ( .I(\pe2/got [31]), .ZN(n36575) );
  BUFHSV4 U33833 ( .I(n36575), .Z(n39105) );
  INHSV4 U33834 ( .I(n49929), .ZN(n58306) );
  INHSV4 U33835 ( .I(n45421), .ZN(n52581) );
  BUFHSV2 U33836 ( .I(n36665), .Z(n44030) );
  INHSV2 U33837 ( .I(n31900), .ZN(n32329) );
  INHSV4 U33838 ( .I(n57011), .ZN(n57230) );
  INHSV8 U33839 ( .I(\pe5/bq[19] ), .ZN(n46134) );
  INHSV4 U33840 ( .I(n46134), .ZN(n39454) );
  INHSV6 U33841 ( .I(\pe4/got [1]), .ZN(n49967) );
  INHSV6 U33842 ( .I(\pe6/got [25]), .ZN(n46750) );
  INHSV6 U33843 ( .I(\pe4/got [18]), .ZN(n33830) );
  INHSV8 U33844 ( .I(\pe1/bq[16] ), .ZN(n45814) );
  INHSV6 U33845 ( .I(n45814), .ZN(n54836) );
  INHSV4 U33846 ( .I(n45814), .ZN(n55100) );
  INHSV2 U33847 ( .I(n32466), .ZN(n31590) );
  INHSV6 U33848 ( .I(n35907), .ZN(n59022) );
  INHSV2 U33849 ( .I(n32239), .ZN(n32422) );
  INHSV2 U33850 ( .I(n35796), .ZN(n46567) );
  INHSV6 U33851 ( .I(\pe4/got [28]), .ZN(n33564) );
  INHSV4 U33852 ( .I(n48028), .ZN(n35184) );
  INHSV6 U33853 ( .I(n48028), .ZN(n58130) );
  BUFHSV4 U33854 ( .I(n36719), .Z(n43880) );
  INHSV4 U33855 ( .I(n43468), .ZN(n43469) );
  INHSV4 U33856 ( .I(n37348), .ZN(n37161) );
  INHSV8 U33857 ( .I(\pe3/bq[3] ), .ZN(n50722) );
  INHSV12 U33858 ( .I(n50722), .ZN(n56529) );
  INHSV4 U33859 ( .I(\pe2/got [17]), .ZN(n44002) );
  INHSV4 U33860 ( .I(n44002), .ZN(n59983) );
  INHSV4 U33861 ( .I(n44002), .ZN(n38782) );
  INHSV6 U33862 ( .I(n38163), .ZN(n38327) );
  INHSV8 U33863 ( .I(\pe2/aot [1]), .ZN(n52095) );
  INHSV2 U33864 ( .I(n52095), .ZN(n59783) );
  INHSV4 U33865 ( .I(n52095), .ZN(n51547) );
  INHSV6 U33866 ( .I(\pe2/bq[3] ), .ZN(n47893) );
  CLKNHSV6 U33867 ( .I(n47893), .ZN(n52484) );
  INHSV4 U33868 ( .I(\pe3/got [26]), .ZN(n42895) );
  INHSV4 U33869 ( .I(n43457), .ZN(n59616) );
  INHSV4 U33870 ( .I(n42895), .ZN(n36955) );
  INHSV6 U33871 ( .I(n42895), .ZN(n46311) );
  BUFHSV4 U33872 ( .I(n51336), .Z(n51370) );
  CLKNHSV6 U33873 ( .I(n55376), .ZN(n54455) );
  INHSV2 U33874 ( .I(n48545), .ZN(n56507) );
  INHSV2 U33875 ( .I(n48545), .ZN(n56688) );
  BUFHSV4 U33876 ( .I(n38099), .Z(n44821) );
  INHSV6 U33877 ( .I(\pe2/got [30]), .ZN(n38733) );
  INHSV8 U33878 ( .I(\pe2/got [25]), .ZN(n39088) );
  INHSV8 U33879 ( .I(n39088), .ZN(n44711) );
  INHSV6 U33880 ( .I(n39088), .ZN(n38324) );
  BUFHSV4 U33881 ( .I(n40719), .Z(n41228) );
  BUFHSV2 U33882 ( .I(n40719), .Z(n41507) );
  INHSV6 U33883 ( .I(\pe5/got [19]), .ZN(n30686) );
  INHSV6 U33884 ( .I(\pe3/got [20]), .ZN(n45635) );
  INHSV4 U33885 ( .I(n45635), .ZN(n42996) );
  INHSV2 U33886 ( .I(n43235), .ZN(n37516) );
  INHSV4 U33887 ( .I(n43235), .ZN(n37107) );
  INHSV4 U33888 ( .I(n43235), .ZN(n36958) );
  INHSV4 U33889 ( .I(n50910), .ZN(n59767) );
  INHSV4 U33890 ( .I(n50910), .ZN(n52896) );
  INHSV2 U33891 ( .I(n43866), .ZN(n43868) );
  INHSV6 U33892 ( .I(n52723), .ZN(n35007) );
  INHSV8 U33893 ( .I(n35007), .ZN(n47772) );
  INHSV8 U33894 ( .I(\pe1/got [17]), .ZN(n53911) );
  INHSV4 U33895 ( .I(n44337), .ZN(n40923) );
  INHSV6 U33896 ( .I(n44337), .ZN(n59374) );
  CLKNHSV0 U33897 ( .I(n48472), .ZN(n59496) );
  CLKNHSV0 U33898 ( .I(n48083), .ZN(n59494) );
  CLKNHSV0 U33899 ( .I(n48472), .ZN(n59424) );
  CLKNHSV0 U33900 ( .I(n48472), .ZN(n59425) );
  BUFHSV4 U33901 ( .I(n41557), .Z(n53602) );
  INHSV4 U33902 ( .I(n48060), .ZN(n41760) );
  INHSV6 U33903 ( .I(n48060), .ZN(n54565) );
  INHSV4 U33904 ( .I(n46960), .ZN(n52653) );
  INHSV2 U33905 ( .I(n46960), .ZN(n51211) );
  BUFHSV4 U33906 ( .I(n29907), .Z(n30864) );
  BUFHSV2 U33907 ( .I(n58717), .Z(n58611) );
  INHSV4 U33908 ( .I(n47199), .ZN(n52564) );
  BUFHSV4 U33909 ( .I(n58718), .Z(n58936) );
  INHSV4 U33910 ( .I(n46977), .ZN(n53293) );
  INHSV4 U33911 ( .I(n45416), .ZN(n48166) );
  INHSV6 U33912 ( .I(\pe1/aot [29]), .ZN(n40787) );
  BUFHSV4 U33913 ( .I(n40787), .Z(n53957) );
  BUFHSV4 U33914 ( .I(n40787), .Z(n40412) );
  INHSV4 U33915 ( .I(n49099), .ZN(n53114) );
  BUFHSV4 U33916 ( .I(n44833), .Z(n47500) );
  BUFHSV4 U33917 ( .I(n59525), .Z(n51018) );
  BUFHSV4 U33918 ( .I(n31147), .Z(n52574) );
  BUFHSV4 U33919 ( .I(n59916), .Z(n53112) );
  INHSV4 U33920 ( .I(n50094), .ZN(n57755) );
  INHSV4 U33921 ( .I(n50094), .ZN(n58185) );
  NAND2HSV4 U33922 ( .A1(n36371), .A2(n36370), .ZN(n36614) );
  BUFHSV4 U33923 ( .I(n36614), .Z(n59349) );
  INHSV4 U33924 ( .I(n36434), .ZN(n36588) );
  INHSV4 U33925 ( .I(n36434), .ZN(n52987) );
  INHSV6 U33926 ( .I(\pe3/aot [27]), .ZN(n42843) );
  BUFHSV8 U33927 ( .I(n43222), .Z(n59380) );
  INHSV4 U33928 ( .I(n59380), .ZN(n45728) );
  INHSV2 U33929 ( .I(n59380), .ZN(n56391) );
  INHSV4 U33930 ( .I(n59380), .ZN(n43840) );
  BUFHSV4 U33931 ( .I(n35668), .Z(n36183) );
  BUFHSV4 U33932 ( .I(n35668), .Z(n32293) );
  INHSV2 U33933 ( .I(n54146), .ZN(n55529) );
  AND3HSV2 U33934 ( .A1(n30780), .A2(n52834), .A3(n39871), .Z(n29634) );
  BUFHSV8 U33935 ( .I(n37274), .Z(n37017) );
  OA21HSV2 U33936 ( .A1(n35447), .A2(n35448), .B(n35449), .Z(n29635) );
  INHSV4 U33937 ( .I(n29915), .ZN(n40293) );
  CLKAND2HSV2 U33938 ( .A1(n34711), .A2(n34419), .Z(n29636) );
  INHSV6 U33939 ( .I(\pe5/aot [29]), .ZN(n30163) );
  INHSV4 U33940 ( .I(n39431), .ZN(n51158) );
  BUFHSV4 U33941 ( .I(n51158), .Z(n52570) );
  INHSV2 U33942 ( .I(n34814), .ZN(n29758) );
  INHSV2 U33943 ( .I(n34814), .ZN(n29759) );
  BUFHSV4 U33944 ( .I(n45801), .Z(n34459) );
  NAND2HSV4 U33945 ( .A1(n33524), .A2(n33523), .ZN(n45801) );
  INHSV8 U33946 ( .I(\pe4/bq[17] ), .ZN(n47809) );
  CLKAND2HSV2 U33947 ( .A1(n32198), .A2(\pe6/pvq [7]), .Z(n29638) );
  INHSV6 U33948 ( .I(\pe4/bq[30] ), .ZN(n34485) );
  INHSV6 U33949 ( .I(\pe4/aot [28]), .ZN(n47661) );
  CLKAND2HSV2 U33950 ( .A1(n53524), .A2(n53786), .Z(n29639) );
  CLKNHSV0 U33951 ( .I(n32436), .ZN(n32340) );
  INHSV6 U33952 ( .I(\pe4/bq[31] ), .ZN(n33111) );
  INHSV2 U33953 ( .I(n33687), .ZN(n33156) );
  NAND2HSV4 U33954 ( .A1(n31284), .A2(n31283), .ZN(n31303) );
  INHSV8 U33955 ( .I(\pe6/aot [32]), .ZN(n31253) );
  BUFHSV2 U33956 ( .I(n41243), .Z(n41734) );
  BUFHSV4 U33957 ( .I(n42088), .Z(n53913) );
  INHSV4 U33958 ( .I(n37953), .ZN(n36480) );
  INHSV2 U33959 ( .I(n37953), .ZN(n38046) );
  CLKNHSV0 U33960 ( .I(n33240), .ZN(n29738) );
  BUFHSV2 U33961 ( .I(n59662), .Z(n34396) );
  BUFHSV2 U33962 ( .I(n33224), .Z(n59662) );
  AO21HSV1 U33963 ( .A1(n39871), .A2(n29842), .B(n29855), .Z(n29642) );
  INHSV2 U33964 ( .I(n40491), .ZN(n41256) );
  INHSV4 U33965 ( .I(n33218), .ZN(n57166) );
  AND2HSV2 U33966 ( .A1(n43133), .A2(n43234), .Z(n29643) );
  INHSV6 U33967 ( .I(\pe6/aot [31]), .ZN(n31487) );
  BUFHSV4 U33968 ( .I(n31487), .Z(n32723) );
  BUFHSV4 U33969 ( .I(n30458), .Z(n39143) );
  CLKAND2HSV2 U33970 ( .A1(n25911), .A2(n32133), .Z(n29644) );
  INHSV4 U33971 ( .I(n33750), .ZN(n47742) );
  INHSV6 U33972 ( .I(\pe5/aot [26]), .ZN(n48219) );
  INHSV4 U33973 ( .I(n48219), .ZN(n39473) );
  INHSV8 U33974 ( .I(n41963), .ZN(n42092) );
  INHSV4 U33975 ( .I(n50847), .ZN(n59084) );
  BUFHSV4 U33976 ( .I(n46123), .Z(n59678) );
  BUFHSV4 U33977 ( .I(n46123), .Z(n32841) );
  INHSV2 U33978 ( .I(n52251), .ZN(n53065) );
  INHSV2 U33979 ( .I(n38368), .ZN(n45071) );
  INHSV6 U33980 ( .I(\pe6/got [30]), .ZN(n32443) );
  BUFHSV4 U33981 ( .I(n32443), .Z(n32651) );
  INHSV4 U33982 ( .I(\pe6/got [30]), .ZN(n35710) );
  INHSV6 U33983 ( .I(ctro6), .ZN(n31298) );
  BUFHSV4 U33984 ( .I(n31461), .Z(n32961) );
  BUFHSV4 U33985 ( .I(\pe1/aot [25]), .Z(n59589) );
  INHSV4 U33986 ( .I(n51567), .ZN(n51825) );
  INHSV6 U33987 ( .I(\pe5/bq[27] ), .ZN(n30113) );
  BUFHSV4 U33988 ( .I(n31461), .Z(n32822) );
  INHSV4 U33989 ( .I(n31873), .ZN(n31261) );
  INHSV6 U33990 ( .I(\pe6/got [23]), .ZN(n49315) );
  INHSV8 U33991 ( .I(\pe6/bq[8] ), .ZN(n48042) );
  INHSV4 U33992 ( .I(n48042), .ZN(n59246) );
  INHSV6 U33993 ( .I(n48042), .ZN(n58619) );
  INHSV2 U33994 ( .I(n35740), .ZN(n32484) );
  INHSV2 U33995 ( .I(n40365), .ZN(n40366) );
  BUFHSV8 U33996 ( .I(n59646), .Z(n56788) );
  BUFHSV4 U33997 ( .I(n39398), .Z(n30667) );
  INHSV4 U33998 ( .I(n38711), .ZN(n52922) );
  INHSV4 U33999 ( .I(n38711), .ZN(n52167) );
  INHSV6 U34000 ( .I(\pe3/aot [22]), .ZN(n45567) );
  INHSV6 U34001 ( .I(n45567), .ZN(n59618) );
  INHSV6 U34002 ( .I(\pe3/aot [17]), .ZN(n43527) );
  INHSV2 U34003 ( .I(n43527), .ZN(n56113) );
  INHSV4 U34004 ( .I(n38823), .ZN(n38043) );
  BUFHSV4 U34005 ( .I(n43870), .Z(n36979) );
  INHSV4 U34006 ( .I(n36979), .ZN(n47428) );
  INHSV4 U34007 ( .I(n57260), .ZN(n34598) );
  INHSV6 U34008 ( .I(\pe2/aot [3]), .ZN(n51538) );
  INHSV4 U34009 ( .I(n51538), .ZN(n52344) );
  INHSV4 U34010 ( .I(n51538), .ZN(n59792) );
  INHSV6 U34011 ( .I(\pe1/aot [18]), .ZN(n41931) );
  INHSV6 U34012 ( .I(\pe1/got [30]), .ZN(n40649) );
  INHSV4 U34013 ( .I(n53518), .ZN(n42196) );
  INHSV2 U34014 ( .I(n40933), .ZN(n40936) );
  INHSV6 U34015 ( .I(\pe3/aot [9]), .ZN(n56567) );
  INHSV4 U34016 ( .I(n56567), .ZN(n59808) );
  BUFHSV4 U34017 ( .I(\pe5/aot [21]), .Z(n51187) );
  INHSV4 U34018 ( .I(n36434), .ZN(n38565) );
  BUFHSV4 U34019 ( .I(n30206), .Z(n37645) );
  INHSV8 U34020 ( .I(\pe3/aot [29]), .ZN(n36989) );
  INHSV2 U34021 ( .I(n36989), .ZN(n48500) );
  INHSV4 U34022 ( .I(n52430), .ZN(n45033) );
  INHSV4 U34023 ( .I(n52430), .ZN(n52299) );
  BUFHSV2 U34024 ( .I(n42067), .Z(n42070) );
  BUFHSV8 U34025 ( .I(n54263), .Z(n54039) );
  INHSV6 U34026 ( .I(n54039), .ZN(n41550) );
  INHSV6 U34027 ( .I(\pe5/aot [12]), .ZN(n50507) );
  INHSV6 U34028 ( .I(\pe2/aot [12]), .ZN(n51736) );
  INHSV2 U34029 ( .I(n42899), .ZN(n42689) );
  BUFHSV8 U34030 ( .I(n48036), .Z(n48025) );
  INHSV2 U34031 ( .I(n59094), .ZN(n59240) );
  INHSV6 U34032 ( .I(\pe2/got [26]), .ZN(n38042) );
  BUFHSV4 U34033 ( .I(n38042), .Z(n52285) );
  INHSV6 U34034 ( .I(\pe6/bq[5] ), .ZN(n46146) );
  INHSV2 U34035 ( .I(n35710), .ZN(n35808) );
  BUFHSV8 U34036 ( .I(\pe5/aot [10]), .Z(n51313) );
  BUFHSV4 U34037 ( .I(\pe5/aot [10]), .Z(n59642) );
  BUFHSV8 U34038 ( .I(\pe5/aot [16]), .Z(n59640) );
  INHSV6 U34039 ( .I(\pe6/bq[6] ), .ZN(n46147) );
  CLKNHSV6 U34040 ( .I(n42230), .ZN(n54578) );
  BUFHSV8 U34041 ( .I(\pe3/bq[7] ), .Z(n45639) );
  INHSV6 U34042 ( .I(\pe6/aot [3]), .ZN(n49681) );
  INHSV2 U34043 ( .I(n49681), .ZN(n58353) );
  INHSV4 U34044 ( .I(n49681), .ZN(n59252) );
  INHSV6 U34045 ( .I(\pe2/bq[19] ), .ZN(n45199) );
  INHSV4 U34046 ( .I(n45199), .ZN(n43961) );
  INHSV4 U34047 ( .I(n45199), .ZN(n38792) );
  BUFHSV4 U34048 ( .I(n33897), .Z(n47679) );
  INHSV4 U34049 ( .I(n46618), .ZN(n35370) );
  INHSV6 U34050 ( .I(\pe1/bq[19] ), .ZN(n41963) );
  INHSV2 U34051 ( .I(\pe5/aot [18]), .ZN(n45858) );
  INHSV6 U34052 ( .I(\pe5/aot [30]), .ZN(n30212) );
  BUFHSV4 U34053 ( .I(n40236), .Z(n39123) );
  INHSV4 U34054 ( .I(n49423), .ZN(n55975) );
  INHSV4 U34055 ( .I(n49423), .ZN(n45534) );
  INHSV4 U34056 ( .I(n32373), .ZN(n33004) );
  INHSV2 U34057 ( .I(n33588), .ZN(n47788) );
  INHSV4 U34058 ( .I(n32858), .ZN(n58943) );
  INHSV4 U34059 ( .I(n32858), .ZN(n49208) );
  INHSV8 U34060 ( .I(\pe5/aot [14]), .ZN(n59641) );
  INHSV6 U34061 ( .I(n59641), .ZN(n39490) );
  INHSV8 U34062 ( .I(\pe6/bq[10] ), .ZN(n49680) );
  INHSV4 U34063 ( .I(n49680), .ZN(n44336) );
  INHSV6 U34064 ( .I(n49680), .ZN(n58962) );
  BUFHSV8 U34065 ( .I(\pe1/bq[5] ), .Z(n54289) );
  INHSV4 U34066 ( .I(n46916), .ZN(n48760) );
  INHSV8 U34067 ( .I(\pe5/bq[16] ), .ZN(n39796) );
  INHSV4 U34068 ( .I(n39796), .ZN(n48181) );
  INHSV4 U34069 ( .I(n43059), .ZN(n46613) );
  BUFHSV4 U34070 ( .I(\pe3/aot [11]), .Z(n56354) );
  INHSV6 U34071 ( .I(\pe5/bq[6] ), .ZN(n46136) );
  CLKNHSV6 U34072 ( .I(n46136), .ZN(n50526) );
  INHSV6 U34073 ( .I(n46136), .ZN(n51191) );
  INHSV6 U34074 ( .I(\pe5/bq[12] ), .ZN(n50428) );
  INHSV4 U34075 ( .I(n50428), .ZN(n52619) );
  INHSV2 U34076 ( .I(n50428), .ZN(n31045) );
  INHSV4 U34077 ( .I(n47230), .ZN(n59944) );
  INHSV6 U34078 ( .I(n47230), .ZN(n51247) );
  INHSV6 U34079 ( .I(\pe6/bq[3] ), .ZN(n49327) );
  BUFHSV12 U34080 ( .I(\pe2/aot [7]), .Z(n59633) );
  INHSV6 U34081 ( .I(\pe4/bq[12] ), .ZN(n57841) );
  INHSV6 U34082 ( .I(\pe4/aot [16]), .ZN(n57030) );
  INHSV8 U34083 ( .I(\pe1/bq[13] ), .ZN(n48059) );
  INHSV4 U34084 ( .I(n48059), .ZN(n41645) );
  INHSV6 U34085 ( .I(n48059), .ZN(n54179) );
  INHSV6 U34086 ( .I(\pe1/aot [5]), .ZN(n55430) );
  INHSV4 U34087 ( .I(n55430), .ZN(n54303) );
  INHSV6 U34088 ( .I(n55430), .ZN(n59993) );
  INHSV4 U34089 ( .I(n55430), .ZN(n55553) );
  INHSV4 U34090 ( .I(n52431), .ZN(n51460) );
  INHSV6 U34091 ( .I(\pe4/aot [12]), .ZN(n34498) );
  CLKNHSV6 U34092 ( .I(n34498), .ZN(n34873) );
  INHSV6 U34093 ( .I(n34498), .ZN(n59343) );
  INHSV2 U34094 ( .I(n40973), .ZN(n40438) );
  INHSV4 U34095 ( .I(n44521), .ZN(n48468) );
  INHSV8 U34096 ( .I(\pe5/bq[18] ), .ZN(n48822) );
  OR2HSV2 U34097 ( .A1(n37871), .A2(n38195), .Z(n38335) );
  BUFHSV4 U34098 ( .I(n45409), .Z(n44312) );
  INHSV4 U34099 ( .I(n38335), .ZN(n36562) );
  INHSV4 U34100 ( .I(n56904), .ZN(n56781) );
  INHSV4 U34101 ( .I(n56904), .ZN(n56684) );
  INHSV8 U34102 ( .I(\pe2/bq[20] ), .ZN(n47599) );
  INHSV4 U34103 ( .I(n47599), .ZN(n52965) );
  INHSV2 U34104 ( .I(n47599), .ZN(n44197) );
  INHSV4 U34105 ( .I(n53292), .ZN(n48841) );
  INHSV6 U34106 ( .I(n53292), .ZN(n52576) );
  CLKNHSV6 U34107 ( .I(n50926), .ZN(n51932) );
  INHSV6 U34108 ( .I(n50926), .ZN(n52895) );
  INHSV6 U34109 ( .I(\pe4/got [25]), .ZN(n33859) );
  INHSV4 U34110 ( .I(n33859), .ZN(n57190) );
  INHSV4 U34111 ( .I(n33859), .ZN(n35318) );
  BUFHSV4 U34112 ( .I(\pe2/aot [6]), .Z(n51636) );
  BUFHSV6 U34113 ( .I(\pe2/aot [6]), .Z(n52456) );
  INHSV6 U34114 ( .I(\pe2/got [24]), .ZN(n38205) );
  INHSV4 U34115 ( .I(n38205), .ZN(n59584) );
  INHSV8 U34116 ( .I(n38205), .ZN(n52416) );
  BUFHSV8 U34117 ( .I(\pe4/aot [10]), .Z(n47718) );
  INHSV12 U34118 ( .I(n54884), .ZN(n54969) );
  INHSV8 U34119 ( .I(\pe1/got [18]), .ZN(n54248) );
  INHSV6 U34120 ( .I(n54248), .ZN(n42359) );
  INHSV8 U34121 ( .I(n54248), .ZN(n54716) );
  INHSV8 U34122 ( .I(\pe4/bq[15] ), .ZN(n47818) );
  INHSV4 U34123 ( .I(n47818), .ZN(n34879) );
  INHSV8 U34124 ( .I(\pe1/bq[20] ), .ZN(n48060) );
  INHSV4 U34125 ( .I(n48060), .ZN(n42238) );
  INHSV4 U34126 ( .I(\pe2/got [23]), .ZN(n38275) );
  INHSV4 U34127 ( .I(n38275), .ZN(n45249) );
  INHSV6 U34128 ( .I(\pe5/bq[15] ), .ZN(n51057) );
  INHSV8 U34129 ( .I(\pe1/got [13]), .ZN(n54957) );
  INHSV6 U34130 ( .I(n54957), .ZN(n42155) );
  INHSV4 U34131 ( .I(n54957), .ZN(n55086) );
  INHSV6 U34132 ( .I(\pe1/aot [16]), .ZN(n54673) );
  INHSV6 U34133 ( .I(n54673), .ZN(n59989) );
  INHSV2 U34134 ( .I(n52226), .ZN(n59973) );
  INHSV4 U34135 ( .I(n52226), .ZN(n51743) );
  BUFHSV4 U34136 ( .I(n40439), .Z(n41418) );
  INHSV4 U34137 ( .I(n46143), .ZN(n57384) );
  CLKNHSV0 U34138 ( .I(\pe6/got [20]), .ZN(n32125) );
  INHSV6 U34139 ( .I(n49739), .ZN(n46818) );
  BUFHSV4 U34140 ( .I(n45091), .Z(n45276) );
  INHSV6 U34141 ( .I(\pe2/bq[15] ), .ZN(n48066) );
  INHSV4 U34142 ( .I(n48066), .ZN(n49619) );
  OR2HSV1 U34143 ( .A1(n30874), .A2(n39733), .Z(n29645) );
  INHSV6 U34144 ( .I(n30202), .ZN(n30046) );
  INHSV6 U34145 ( .I(n47555), .ZN(n52172) );
  BUFHSV4 U34146 ( .I(n53936), .Z(n54913) );
  BUFHSV2 U34147 ( .I(\pe2/aot [5]), .Z(n59499) );
  INHSV6 U34148 ( .I(n48622), .ZN(n52056) );
  INHSV4 U34149 ( .I(n48622), .ZN(n29736) );
  INHSV4 U34150 ( .I(n45662), .ZN(n55873) );
  INHSV4 U34151 ( .I(n45662), .ZN(n56439) );
  INHSV4 U34152 ( .I(n54672), .ZN(n55113) );
  INHSV4 U34153 ( .I(n41653), .ZN(n44533) );
  BUFHSV4 U34154 ( .I(\pe5/aot [8]), .Z(n59880) );
  BUFHSV4 U34155 ( .I(\pe5/aot [8]), .Z(n50511) );
  INHSV4 U34156 ( .I(n49529), .ZN(n51457) );
  INHSV6 U34157 ( .I(n54879), .ZN(n55087) );
  INHSV2 U34158 ( .I(n49967), .ZN(n58219) );
  BUFHSV4 U34159 ( .I(n33184), .Z(n52696) );
  BUFHSV4 U34160 ( .I(n33184), .Z(n47777) );
  INHSV8 U34161 ( .I(n49826), .ZN(n59328) );
  INHSV8 U34162 ( .I(\pe1/bq[10] ), .ZN(n53723) );
  INHSV2 U34163 ( .I(n53723), .ZN(n55352) );
  INHSV8 U34164 ( .I(\pe6/aot [5]), .ZN(n58359) );
  INHSV4 U34165 ( .I(n58359), .ZN(n58378) );
  INHSV4 U34166 ( .I(n58359), .ZN(n59250) );
  INHSV8 U34167 ( .I(\pe1/bq[3] ), .ZN(n54399) );
  INHSV2 U34168 ( .I(n54399), .ZN(n55518) );
  INHSV6 U34169 ( .I(\pe5/got [1]), .ZN(n48625) );
  INHSV12 U34170 ( .I(n48625), .ZN(n51362) );
  BUFHSV2 U34171 ( .I(n55523), .Z(n54735) );
  INHSV4 U34172 ( .I(n55523), .ZN(n54911) );
  INHSV8 U34173 ( .I(n55523), .ZN(n55231) );
  BUFHSV8 U34174 ( .I(\pe6/got [12]), .Z(n33039) );
  BUFHSV4 U34175 ( .I(\pe6/got [14]), .Z(n58713) );
  BUFHSV6 U34176 ( .I(\pe6/got [14]), .Z(n58810) );
  INHSV2 U34177 ( .I(n48740), .ZN(n31122) );
  INHSV4 U34178 ( .I(n50550), .ZN(n51302) );
  INHSV2 U34179 ( .I(n32422), .ZN(n32457) );
  INHSV2 U34180 ( .I(n41228), .ZN(n42084) );
  INHSV6 U34181 ( .I(\pe3/bq[15] ), .ZN(n46615) );
  INHSV4 U34182 ( .I(n46615), .ZN(n56641) );
  CLKNHSV6 U34183 ( .I(n55364), .ZN(n55319) );
  INHSV6 U34184 ( .I(\pe5/aot [9]), .ZN(n48246) );
  CLKNHSV6 U34185 ( .I(n48246), .ZN(n39887) );
  INHSV6 U34186 ( .I(\pe1/got [5]), .ZN(n55542) );
  INHSV8 U34187 ( .I(n55542), .ZN(n55475) );
  INHSV8 U34188 ( .I(\pe3/got [19]), .ZN(n49250) );
  INHSV4 U34189 ( .I(n49250), .ZN(n42937) );
  INHSV4 U34190 ( .I(n49250), .ZN(n56489) );
  INHSV6 U34191 ( .I(n49250), .ZN(n59965) );
  INHSV4 U34192 ( .I(n56956), .ZN(n56972) );
  INHSV8 U34193 ( .I(n56956), .ZN(n59961) );
  INHSV4 U34194 ( .I(n35796), .ZN(n59339) );
  BUFHSV4 U34195 ( .I(n25344), .Z(n30048) );
  BUFHSV4 U34196 ( .I(n30089), .Z(n29950) );
  INHSV4 U34197 ( .I(n29825), .ZN(n30075) );
  INHSV6 U34198 ( .I(\pe4/aot [5]), .ZN(n49929) );
  INHSV4 U34199 ( .I(n49929), .ZN(n59831) );
  INHSV4 U34200 ( .I(n47570), .ZN(n59982) );
  INHSV4 U34201 ( .I(n47570), .ZN(n39075) );
  INHSV4 U34202 ( .I(n39250), .ZN(n30976) );
  INHSV4 U34203 ( .I(n29907), .ZN(n39702) );
  INHSV4 U34204 ( .I(n57453), .ZN(n59956) );
  INHSV6 U34205 ( .I(\pe5/got [16]), .ZN(n30888) );
  INHSV4 U34206 ( .I(n33997), .ZN(n33696) );
  INHSV6 U34207 ( .I(\pe4/aot [13]), .ZN(n44338) );
  INHSV2 U34208 ( .I(n44378), .ZN(n36050) );
  INHSV4 U34209 ( .I(n39403), .ZN(n39241) );
  INHSV8 U34210 ( .I(\pe3/got [5]), .ZN(n56859) );
  INHSV6 U34211 ( .I(\pe5/aot [1]), .ZN(n45904) );
  INHSV6 U34212 ( .I(\pe3/got [21]), .ZN(n37275) );
  INHSV4 U34213 ( .I(n48186), .ZN(n52632) );
  INHSV12 U34214 ( .I(n34460), .ZN(n58153) );
  INHSV6 U34215 ( .I(\pe5/got [14]), .ZN(n31199) );
  INHSV4 U34216 ( .I(n48026), .ZN(n57906) );
  INHSV4 U34217 ( .I(\pe3/got [18]), .ZN(n49251) );
  INHSV6 U34218 ( .I(n49251), .ZN(n43374) );
  INHSV4 U34219 ( .I(\pe4/aot [1]), .ZN(n47905) );
  INHSV8 U34220 ( .I(\pe3/got [24]), .ZN(n42817) );
  INHSV4 U34221 ( .I(n42817), .ZN(n43452) );
  INHSV6 U34222 ( .I(n42817), .ZN(n59617) );
  INHSV2 U34223 ( .I(n32815), .ZN(n31971) );
  INHSV6 U34224 ( .I(\pe3/got [23]), .ZN(n42827) );
  INHSV6 U34225 ( .I(n42827), .ZN(n42673) );
  BUFHSV4 U34226 ( .I(\pe6/got [26]), .Z(n32242) );
  INHSV6 U34227 ( .I(\pe1/aot [3]), .ZN(n55515) );
  INHSV6 U34228 ( .I(n55515), .ZN(n55496) );
  INHSV4 U34229 ( .I(n32439), .ZN(n32783) );
  INHSV8 U34230 ( .I(\pe2/got [15]), .ZN(n47573) );
  INHSV8 U34231 ( .I(\pe2/got [20]), .ZN(n44327) );
  INHSV4 U34232 ( .I(n34566), .ZN(n34571) );
  INHSV6 U34233 ( .I(\pe3/bq[10] ), .ZN(n56269) );
  INHSV8 U34234 ( .I(n56269), .ZN(n56627) );
  BUFHSV4 U34235 ( .I(n34328), .Z(n34727) );
  INHSV8 U34236 ( .I(\pe4/bq[13] ), .ZN(n53219) );
  INHSV6 U34237 ( .I(n53219), .ZN(n34480) );
  INHSV6 U34238 ( .I(n53219), .ZN(n58127) );
  INHSV8 U34239 ( .I(\pe5/got [3]), .ZN(n51231) );
  INHSV6 U34240 ( .I(\pe5/got [21]), .ZN(n30516) );
  INHSV4 U34241 ( .I(n59615), .ZN(n46107) );
  INHSV8 U34242 ( .I(\pe4/bq[1] ), .ZN(n58013) );
  INHSV8 U34243 ( .I(\pe3/bq[2] ), .ZN(n48495) );
  INHSV2 U34244 ( .I(n48495), .ZN(n56348) );
  INHSV6 U34245 ( .I(\pe3/got [15]), .ZN(n45727) );
  INHSV6 U34246 ( .I(\pe2/got [28]), .ZN(n45411) );
  INHSV4 U34247 ( .I(n31003), .ZN(n40008) );
  INHSV12 U34248 ( .I(n46042), .ZN(n56493) );
  INHSV2 U34249 ( .I(n49003), .ZN(n49825) );
  INHSV2 U34250 ( .I(n54691), .ZN(n54521) );
  INHSV2 U34251 ( .I(n54691), .ZN(n54600) );
  INHSV4 U34252 ( .I(n54691), .ZN(n41850) );
  INHSV2 U34253 ( .I(n30320), .ZN(n40007) );
  INHSV6 U34254 ( .I(\pe1/got [20]), .ZN(n48338) );
  INHSV6 U34255 ( .I(n48338), .ZN(n44530) );
  INHSV4 U34256 ( .I(n58253), .ZN(n58111) );
  INHSV6 U34257 ( .I(\pe3/got [17]), .ZN(n44693) );
  INHSV4 U34258 ( .I(n44693), .ZN(n56064) );
  INHSV8 U34259 ( .I(n44693), .ZN(n56335) );
  BUFHSV4 U34260 ( .I(\pe6/got [1]), .Z(n58403) );
  BUFHSV4 U34261 ( .I(\pe6/got [1]), .Z(n58817) );
  BUFHSV4 U34262 ( .I(\pe6/got [1]), .Z(n59235) );
  BUFHSV8 U34263 ( .I(n34452), .Z(n34591) );
  INHSV4 U34264 ( .I(n34452), .ZN(n33748) );
  INHSV12 U34265 ( .I(n34591), .ZN(n59350) );
  INHSV4 U34266 ( .I(n42344), .ZN(n40541) );
  INHSV2 U34267 ( .I(n38523), .ZN(n38890) );
  INHSV4 U34268 ( .I(n39105), .ZN(n44827) );
  INHSV2 U34269 ( .I(n36319), .ZN(n59979) );
  INHSV2 U34270 ( .I(n46438), .ZN(n29750) );
  INHSV4 U34271 ( .I(n43744), .ZN(n43898) );
  INHSV4 U34272 ( .I(n53834), .ZN(n55110) );
  INHSV6 U34273 ( .I(n53834), .ZN(n55605) );
  BUFHSV4 U34274 ( .I(\pe6/got [7]), .Z(n58562) );
  BUFHSV4 U34275 ( .I(\pe6/got [7]), .Z(n36109) );
  BUFHSV4 U34276 ( .I(n34328), .Z(n57204) );
  INHSV4 U34277 ( .I(n33694), .ZN(n34718) );
  INHSV6 U34278 ( .I(\pe2/aot [4]), .ZN(n51537) );
  INHSV2 U34279 ( .I(n51537), .ZN(n51824) );
  INHSV4 U34280 ( .I(n47143), .ZN(n59643) );
  INHSV4 U34281 ( .I(n47143), .ZN(n51305) );
  INHSV8 U34282 ( .I(\pe3/got [12]), .ZN(n50802) );
  INHSV4 U34283 ( .I(n35488), .ZN(n34239) );
  INHSV4 U34284 ( .I(n35488), .ZN(n59369) );
  INHSV2 U34285 ( .I(n46270), .ZN(n58715) );
  INHSV4 U34286 ( .I(n46270), .ZN(n36104) );
  INHSV4 U34287 ( .I(n46270), .ZN(n53101) );
  INHSV8 U34288 ( .I(\pe5/got [10]), .ZN(n46961) );
  INHSV2 U34289 ( .I(n46961), .ZN(n51210) );
  INHSV6 U34290 ( .I(\pe6/aot [8]), .ZN(n58483) );
  CLKNHSV6 U34291 ( .I(n58483), .ZN(n58857) );
  INHSV4 U34292 ( .I(n58483), .ZN(n35632) );
  INHSV6 U34293 ( .I(\pe3/aot [3]), .ZN(n56704) );
  INHSV6 U34294 ( .I(n56704), .ZN(n56434) );
  INHSV6 U34295 ( .I(n56704), .ZN(n53250) );
  BUFHSV4 U34296 ( .I(n35311), .Z(n35011) );
  INHSV4 U34297 ( .I(n40394), .ZN(n42471) );
  INHSV2 U34298 ( .I(n41701), .ZN(n40407) );
  INHSV4 U34299 ( .I(n40525), .ZN(n53787) );
  INHSV4 U34300 ( .I(n40393), .ZN(n40957) );
  CLKNHSV6 U34301 ( .I(\pe3/got [9]), .ZN(n56680) );
  INHSV2 U34302 ( .I(n56680), .ZN(n59645) );
  INHSV6 U34303 ( .I(\pe5/got [8]), .ZN(n45901) );
  INHSV12 U34304 ( .I(n45901), .ZN(n50698) );
  INHSV6 U34305 ( .I(\pe2/bq[4] ), .ZN(n48621) );
  INHSV4 U34306 ( .I(n48621), .ZN(n51803) );
  NAND2HSV2 U34307 ( .A1(n42689), .A2(\pe3/ti_7t [23]), .ZN(n43871) );
  INHSV4 U34308 ( .I(n43604), .ZN(n36967) );
  INHSV4 U34309 ( .I(n36979), .ZN(n36980) );
  BUFHSV2 U34310 ( .I(n36682), .Z(n43021) );
  BUFHSV4 U34311 ( .I(n37168), .Z(n45625) );
  BUFHSV4 U34312 ( .I(n43870), .Z(n36873) );
  INHSV2 U34313 ( .I(ctro2), .ZN(n45399) );
  INHSV4 U34314 ( .I(n35035), .ZN(n34864) );
  INHSV2 U34315 ( .I(n35035), .ZN(n33708) );
  INHSV4 U34316 ( .I(n31590), .ZN(n32241) );
  INHSV8 U34317 ( .I(\pe4/bq[5] ), .ZN(n48032) );
  INHSV4 U34318 ( .I(n48032), .ZN(n58155) );
  INHSV4 U34319 ( .I(n48032), .ZN(n58010) );
  INHSV4 U34320 ( .I(n53098), .ZN(n38264) );
  INHSV4 U34321 ( .I(n44030), .ZN(n44322) );
  INHSV4 U34322 ( .I(n50756), .ZN(n56558) );
  INHSV4 U34323 ( .I(n50756), .ZN(n59644) );
  INHSV4 U34324 ( .I(n46119), .ZN(n40257) );
  INHSV4 U34325 ( .I(n46119), .ZN(n52641) );
  INHSV4 U34326 ( .I(n30210), .ZN(n37630) );
  INHSV8 U34327 ( .I(\pe1/got [22]), .ZN(n42209) );
  INHSV4 U34328 ( .I(n55575), .ZN(n54104) );
  CLKNHSV6 U34329 ( .I(n49494), .ZN(n52052) );
  INHSV8 U34330 ( .I(\pe2/got [4]), .ZN(n50909) );
  INHSV4 U34331 ( .I(n50909), .ZN(n59984) );
  INHSV6 U34332 ( .I(\pe1/got [19]), .ZN(n41928) );
  INHSV4 U34333 ( .I(n56906), .ZN(n56823) );
  INHSV4 U34334 ( .I(n47140), .ZN(n48744) );
  INHSV4 U34335 ( .I(n47140), .ZN(n47267) );
  INHSV8 U34336 ( .I(\pe4/got [2]), .ZN(n58325) );
  INHSV6 U34337 ( .I(n58325), .ZN(n58314) );
  INHSV6 U34338 ( .I(n58325), .ZN(n59346) );
  INHSV2 U34339 ( .I(n43484), .ZN(n45607) );
  INHSV4 U34340 ( .I(\pe5/got [23]), .ZN(n39743) );
  INHSV4 U34341 ( .I(n39743), .ZN(n47200) );
  INHSV4 U34342 ( .I(n40520), .ZN(n53650) );
  INHSV4 U34343 ( .I(n39366), .ZN(n39730) );
  INHSV4 U34344 ( .I(n44188), .ZN(n59371) );
  BUFHSV2 U34345 ( .I(n47793), .Z(n50294) );
  INHSV4 U34346 ( .I(n47793), .ZN(n57189) );
  INHSV4 U34347 ( .I(n47793), .ZN(n47656) );
  INHSV6 U34348 ( .I(n52696), .ZN(n52723) );
  INHSV8 U34349 ( .I(\pe4/got [17]), .ZN(n47861) );
  BUFHSV4 U34350 ( .I(n38013), .Z(n38375) );
  INHSV2 U34351 ( .I(n52745), .ZN(n36519) );
  INHSV2 U34352 ( .I(n44494), .ZN(n58807) );
  INHSV4 U34353 ( .I(n32696), .ZN(n35922) );
  INHSV2 U34354 ( .I(n43868), .ZN(n43371) );
  INHSV6 U34355 ( .I(\pe5/got [27]), .ZN(n30431) );
  BUFHSV4 U34356 ( .I(n32961), .Z(n52710) );
  INHSV8 U34357 ( .I(\pe2/got [11]), .ZN(n49656) );
  INHSV4 U34358 ( .I(n43483), .ZN(n43484) );
  INHSV4 U34359 ( .I(n30686), .ZN(n47056) );
  INHSV4 U34360 ( .I(n30686), .ZN(n51103) );
  INHSV8 U34361 ( .I(\pe3/got [11]), .ZN(n50799) );
  INHSV4 U34362 ( .I(n40169), .ZN(n59946) );
  INHSV6 U34363 ( .I(\pe5/got [6]), .ZN(n45903) );
  INHSV12 U34364 ( .I(n45903), .ZN(n51200) );
  INHSV8 U34365 ( .I(n39119), .ZN(n45816) );
  INHSV6 U34366 ( .I(\pe1/got [7]), .ZN(n55019) );
  INHSV6 U34367 ( .I(\pe2/got [18]), .ZN(n47648) );
  INHSV4 U34368 ( .I(n47648), .ZN(n52050) );
  INHSV4 U34369 ( .I(n47648), .ZN(n44712) );
  BUFHSV2 U34370 ( .I(\pe1/ctrq ), .Z(n48053) );
  BUFHSV6 U34371 ( .I(n59486), .Z(n48073) );
  BUFHSV8 U34372 ( .I(n48049), .Z(n48077) );
  BUFHSV4 U34373 ( .I(n48049), .Z(n48034) );
  BUFHSV4 U34374 ( .I(n46623), .Z(n38576) );
  INHSV6 U34375 ( .I(\pe1/aot [26]), .ZN(n46629) );
  INHSV2 U34376 ( .I(n46629), .ZN(n41153) );
  CLKNHSV0 U34377 ( .I(n59660), .ZN(n59493) );
  CLKNHSV0 U34378 ( .I(n48479), .ZN(n59488) );
  BUFHSV2 U34379 ( .I(n59412), .Z(n59925) );
  CLKNHSV0 U34380 ( .I(n48472), .ZN(n59512) );
  CLKNHSV0 U34381 ( .I(n48015), .ZN(n59491) );
  INHSV4 U34382 ( .I(n36719), .ZN(n45755) );
  BUFHSV8 U34383 ( .I(n59615), .Z(n36719) );
  BUFHSV4 U34384 ( .I(n36719), .Z(n37268) );
  BUFHSV8 U34385 ( .I(\pe2/bq[23] ), .Z(n52179) );
  BUFHSV4 U34386 ( .I(n52179), .Z(n52300) );
  INHSV2 U34387 ( .I(n35798), .ZN(n46549) );
  INHSV6 U34388 ( .I(\pe3/bq[22] ), .ZN(n37196) );
  BUFHSV4 U34389 ( .I(n59317), .Z(n58901) );
  BUFHSV4 U34390 ( .I(n29741), .Z(n55230) );
  BUFHSV4 U34391 ( .I(n59811), .Z(n55912) );
  INHSV4 U34392 ( .I(n32723), .ZN(n32973) );
  INHSV4 U34393 ( .I(n32086), .ZN(n36114) );
  INHSV4 U34394 ( .I(n54431), .ZN(n54872) );
  INHSV4 U34395 ( .I(n54431), .ZN(n54946) );
  INHSV4 U34396 ( .I(n55018), .ZN(n53768) );
  INHSV6 U34397 ( .I(\pe4/aot [29]), .ZN(n34479) );
  BUFHSV4 U34398 ( .I(n43467), .Z(n45931) );
  INHSV6 U34399 ( .I(\pe4/aot [15]), .ZN(n57918) );
  BUFHSV4 U34400 ( .I(n35712), .Z(n58480) );
  INHSV6 U34401 ( .I(\pe6/aot [19]), .ZN(n46637) );
  BUFHSV4 U34402 ( .I(n35036), .Z(n57404) );
  BUFHSV4 U34403 ( .I(n35036), .Z(n57530) );
  BUFHSV4 U34404 ( .I(n34888), .Z(n33934) );
  OAI21HSV2 U34405 ( .A1(n33196), .A2(n33195), .B(n25876), .ZN(n29781) );
  BUFHSV4 U34406 ( .I(n54362), .Z(n54041) );
  BUFHSV4 U34407 ( .I(n31527), .Z(n35797) );
  INHSV6 U34408 ( .I(\pe5/bq[30] ), .ZN(n29892) );
  BUFHSV4 U34409 ( .I(n34967), .Z(n50213) );
  INHSV4 U34410 ( .I(n35317), .ZN(n50065) );
  BUFHSV4 U34411 ( .I(n34285), .Z(n59382) );
  INHSV2 U34412 ( .I(n33463), .ZN(n34285) );
  BUFHSV4 U34413 ( .I(n25218), .Z(n59295) );
  INHSV4 U34414 ( .I(n45416), .ZN(n51361) );
  INHSV4 U34415 ( .I(n54635), .ZN(n55489) );
  INHSV4 U34416 ( .I(n47926), .ZN(n59933) );
  INHSV4 U34417 ( .I(n47926), .ZN(n51155) );
  INHSV6 U34418 ( .I(\pe3/aot [28]), .ZN(n45555) );
  BUFHSV4 U34419 ( .I(n34459), .Z(n57209) );
  CLKNHSV0 U34420 ( .I(n33277), .ZN(n35010) );
  NOR2HSV4 U34421 ( .A1(n47777), .A2(n33156), .ZN(n33277) );
  INHSV6 U34422 ( .I(\pe2/bq[27] ), .ZN(n36530) );
  INHSV4 U34423 ( .I(n55162), .ZN(n55449) );
  AND2HSV2 U34424 ( .A1(n41061), .A2(n42484), .Z(n29648) );
  INHSV2 U34425 ( .I(n42512), .ZN(n37528) );
  BUFHSV4 U34426 ( .I(n59775), .Z(n52923) );
  AND3HSV4 U34427 ( .A1(n33161), .A2(n33160), .A3(n33277), .Z(n29650) );
  BUFHSV2 U34428 ( .I(n45800), .Z(n48748) );
  INHSV2 U34429 ( .I(n35816), .ZN(n59065) );
  INHSV6 U34430 ( .I(\pe3/bq[29] ), .ZN(n36694) );
  INHSV6 U34431 ( .I(\pe6/bq[30] ), .ZN(n31425) );
  BUFHSV2 U34432 ( .I(n44212), .Z(n37940) );
  INHSV2 U34433 ( .I(n44212), .ZN(n52995) );
  AND2HSV4 U34434 ( .A1(n47983), .A2(n41410), .Z(n29653) );
  INHSV4 U34435 ( .I(n43029), .ZN(n42810) );
  INHSV4 U34436 ( .I(n43029), .ZN(n42918) );
  INHSV4 U34437 ( .I(n43919), .ZN(n36320) );
  BUFHSV8 U34438 ( .I(n30075), .Z(n30421) );
  NAND2HSV4 U34439 ( .A1(n33094), .A2(n34203), .ZN(n33095) );
  INHSV2 U34440 ( .I(\pe5/ti_1 ), .ZN(n29900) );
  INHSV2 U34441 ( .I(n29826), .ZN(n29827) );
  BUFHSV4 U34442 ( .I(n38195), .Z(n38886) );
  XOR3HSV2 U34443 ( .A1(n44517), .A2(n44516), .A3(n44515), .Z(n29655) );
  BUFHSV4 U34444 ( .I(n45517), .Z(n55948) );
  CLKNAND2HSV2 U34445 ( .A1(n35294), .A2(\pe4/ti_7t [5]), .ZN(n33170) );
  AND2HSV2 U34446 ( .A1(n52754), .A2(n30322), .Z(n29656) );
  INHSV2 U34447 ( .I(n34819), .ZN(n35317) );
  INHSV4 U34448 ( .I(\pe2/pvq [1]), .ZN(n36252) );
  OR2HSV1 U34449 ( .A1(n33655), .A2(n34452), .Z(n29658) );
  INHSV2 U34450 ( .I(n37020), .ZN(n37312) );
  XNOR3HSV2 U34451 ( .A1(n43229), .A2(n43228), .A3(n43227), .ZN(n29659) );
  AND2HSV2 U34452 ( .A1(n30505), .A2(n30504), .Z(n29660) );
  AO21HSV1 U34453 ( .A1(n30303), .A2(n52732), .B(n30302), .Z(n29662) );
  INHSV6 U34454 ( .I(\pe4/aot [27]), .ZN(n33250) );
  AND2HSV2 U34455 ( .A1(n37774), .A2(n37773), .Z(n29664) );
  AND2HSV2 U34456 ( .A1(n59596), .A2(n59166), .Z(n29665) );
  INHSV4 U34457 ( .I(n37335), .ZN(n47992) );
  NAND2HSV2 U34458 ( .A1(n52717), .A2(n29841), .ZN(n29666) );
  INHSV6 U34459 ( .I(\pe4/aot [30]), .ZN(n34631) );
  BUFHSV4 U34460 ( .I(n32976), .Z(n32877) );
  INHSV2 U34461 ( .I(n33224), .ZN(n33240) );
  CLKAND2HSV2 U34462 ( .A1(n31364), .A2(n32783), .Z(n29670) );
  XNOR2HSV4 U34463 ( .A1(n30494), .A2(n30493), .ZN(n29672) );
  CLKAND2HSV2 U34464 ( .A1(n52288), .A2(n36377), .Z(n29673) );
  XOR2HSV0 U34465 ( .A1(n29877), .A2(n29876), .Z(n29675) );
  AND2HSV2 U34466 ( .A1(n33388), .A2(n33389), .Z(n29676) );
  INHSV2 U34467 ( .I(n39824), .ZN(n44332) );
  CLKAND2HSV2 U34468 ( .A1(n36570), .A2(n36565), .Z(n29678) );
  INHSV6 U34469 ( .I(\pe4/bq[26] ), .ZN(n33350) );
  CLKXOR2HSV2 U34470 ( .A1(n40574), .A2(n40573), .Z(n29679) );
  INHSV6 U34471 ( .I(\pe6/aot [24]), .ZN(n50837) );
  INHSV6 U34472 ( .I(\pe6/aot [25]), .ZN(n46663) );
  INHSV6 U34473 ( .I(\pe5/aot [25]), .ZN(n30150) );
  INHSV6 U34474 ( .I(\pe4/aot [21]), .ZN(n50008) );
  INHSV6 U34475 ( .I(\pe3/aot [25]), .ZN(n55714) );
  INHSV6 U34476 ( .I(\pe2/aot [20]), .ZN(n50947) );
  NAND2HSV4 U34477 ( .A1(n36843), .A2(n36846), .ZN(n36847) );
  INHSV6 U34478 ( .I(n36385), .ZN(n37953) );
  INHSV4 U34479 ( .I(n36237), .ZN(n52444) );
  INHSV4 U34480 ( .I(n37953), .ZN(n36607) );
  BUFHSV4 U34481 ( .I(n31140), .Z(n31141) );
  CLKAND2HSV2 U34482 ( .A1(n44323), .A2(n36250), .Z(n29681) );
  CLKAND2HSV2 U34483 ( .A1(n36880), .A2(n36879), .Z(n29682) );
  CLKXOR2HSV2 U34484 ( .A1(n42577), .A2(n42576), .Z(n29683) );
  INHSV2 U34485 ( .I(n41706), .ZN(n42031) );
  INHSV6 U34486 ( .I(\pe3/aot [30]), .ZN(n42643) );
  INHSV8 U34487 ( .I(\pe1/bq[29] ), .ZN(n40455) );
  NOR2HSV2 U34488 ( .A1(n44180), .A2(n44170), .ZN(n45113) );
  AND2HSV2 U34489 ( .A1(n35462), .A2(n35472), .Z(n29685) );
  AND3HSV2 U34490 ( .A1(n44301), .A2(n44300), .A3(n45409), .Z(n29686) );
  INHSV2 U34491 ( .I(n34712), .ZN(n33450) );
  BUFHSV4 U34492 ( .I(n33282), .Z(n34226) );
  CLKXOR2HSV4 U34493 ( .A1(n36247), .A2(n36246), .Z(n29687) );
  BUFHSV4 U34494 ( .I(n52738), .Z(n55825) );
  INHSV6 U34495 ( .I(\pe6/bq[32] ), .ZN(n31844) );
  INHSV4 U34496 ( .I(n31418), .ZN(n31560) );
  INHSV4 U34497 ( .I(n31844), .ZN(n31418) );
  INHSV4 U34498 ( .I(n31560), .ZN(n46627) );
  INHSV2 U34499 ( .I(n45418), .ZN(n30781) );
  INHSV4 U34500 ( .I(\pe4/bq[28] ), .ZN(n33538) );
  BUFHSV8 U34501 ( .I(n33538), .Z(n35092) );
  NAND2HSV0 U34502 ( .A1(n44508), .A2(n46760), .ZN(n29690) );
  XOR2HSV4 U34503 ( .A1(n40855), .A2(n40854), .Z(n29692) );
  INHSV4 U34504 ( .I(\pe4/bq[29] ), .ZN(n33112) );
  CLKAND2HSV2 U34505 ( .A1(n37649), .A2(n37648), .Z(n29693) );
  CLKAND2HSV2 U34506 ( .A1(n36655), .A2(n36654), .Z(n29694) );
  CLKAND2HSV2 U34507 ( .A1(n36887), .A2(n36886), .Z(n29695) );
  CLKNHSV0 U34508 ( .I(n43896), .ZN(n44666) );
  INHSV6 U34509 ( .I(\pe2/bq[28] ), .ZN(n36434) );
  INHSV2 U34510 ( .I(n39992), .ZN(n39860) );
  INHSV4 U34511 ( .I(n39992), .ZN(n53344) );
  INHSV4 U34512 ( .I(n35454), .ZN(n35465) );
  INHSV4 U34513 ( .I(n44531), .ZN(n41849) );
  CLKAND2HSV2 U34514 ( .A1(n30507), .A2(n59946), .Z(n29699) );
  INHSV6 U34515 ( .I(\pe5/bq[31] ), .ZN(n39163) );
  OR2HSV1 U34516 ( .A1(n34580), .A2(n33095), .Z(n29700) );
  BUFHSV4 U34517 ( .I(n36299), .Z(n36587) );
  CLKAND2HSV2 U34518 ( .A1(n36899), .A2(n43905), .Z(n29701) );
  CLKNHSV0 U34519 ( .I(n35479), .ZN(n46565) );
  INHSV6 U34520 ( .I(\pe6/ti_1 ), .ZN(n31424) );
  AND2HSV2 U34521 ( .A1(n52803), .A2(n30872), .Z(n29702) );
  CLKAND2HSV2 U34522 ( .A1(n36408), .A2(n36562), .Z(n29703) );
  CLKXOR2HSV4 U34523 ( .A1(n37166), .A2(n37165), .Z(n29704) );
  CLKNAND2HSV4 U34524 ( .A1(n31271), .A2(n31270), .ZN(n31288) );
  XNOR2HSV1 U34525 ( .A1(n34192), .A2(n34191), .ZN(n34235) );
  BUFHSV4 U34526 ( .I(n40437), .Z(n41134) );
  BUFHSV2 U34527 ( .I(n42212), .Z(n41076) );
  INHSV4 U34528 ( .I(n36898), .ZN(n36844) );
  OR2HSV1 U34529 ( .A1(n42791), .A2(n42790), .Z(n29705) );
  NAND2HSV4 U34530 ( .A1(n38016), .A2(n38098), .ZN(n38206) );
  INHSV2 U34531 ( .I(n39734), .ZN(n39713) );
  INHSV2 U34532 ( .I(n38787), .ZN(n59588) );
  OR2HSV1 U34533 ( .A1(n39676), .A2(n39675), .Z(n29706) );
  CLKAND2HSV2 U34534 ( .A1(n31502), .A2(n31501), .Z(n29708) );
  CLKAND2HSV2 U34535 ( .A1(n36090), .A2(n36089), .Z(n29710) );
  INHSV4 U34536 ( .I(n51121), .ZN(n59522) );
  CLKAND2HSV4 U34537 ( .A1(n37762), .A2(n31241), .Z(n29711) );
  INHSV4 U34538 ( .I(\pe5/got [32]), .ZN(n30051) );
  CLKNHSV0 U34539 ( .I(n37223), .ZN(n37229) );
  XNOR2HSV4 U34540 ( .A1(n37172), .A2(n37171), .ZN(n37223) );
  CLKAND2HSV2 U34541 ( .A1(n30137), .A2(n39558), .Z(n29714) );
  INHSV2 U34542 ( .I(n40556), .ZN(n40491) );
  BUFHSV4 U34543 ( .I(n40556), .Z(n41870) );
  INHSV6 U34544 ( .I(\pe1/aot [30]), .ZN(n40556) );
  CLKNHSV0 U34545 ( .I(n39365), .ZN(n39360) );
  BUFHSV4 U34546 ( .I(n33498), .Z(n57526) );
  INHSV2 U34547 ( .I(n38655), .ZN(n38479) );
  INHSV12 U34548 ( .I(n55227), .ZN(n55339) );
  INHSV6 U34549 ( .I(\pe6/aot [18]), .ZN(n32245) );
  INHSV2 U34550 ( .I(n32245), .ZN(n59088) );
  INHSV2 U34551 ( .I(n32245), .ZN(n58760) );
  INHSV8 U34552 ( .I(\pe5/aot [28]), .ZN(n40235) );
  INHSV4 U34553 ( .I(n40235), .ZN(n40234) );
  INHSV4 U34554 ( .I(n40235), .ZN(n39266) );
  INHSV4 U34555 ( .I(n44411), .ZN(n46658) );
  INHSV2 U34556 ( .I(n35631), .ZN(n31990) );
  INHSV2 U34557 ( .I(n32269), .ZN(n32992) );
  BUFHSV8 U34558 ( .I(\pe3/bq[23] ), .Z(n56213) );
  INHSV2 U34559 ( .I(n48063), .ZN(n51732) );
  INHSV4 U34560 ( .I(n48063), .ZN(n52984) );
  INHSV6 U34561 ( .I(\pe5/got [28]), .ZN(n30297) );
  INHSV8 U34562 ( .I(\pe2/aot [27]), .ZN(n44095) );
  INHSV4 U34563 ( .I(n44095), .ZN(n45295) );
  BUFHSV8 U34564 ( .I(n59519), .Z(n56180) );
  INHSV6 U34565 ( .I(\pe3/bq[27] ), .ZN(n45525) );
  INHSV4 U34566 ( .I(n45525), .ZN(n55960) );
  INHSV4 U34567 ( .I(n38664), .ZN(n59971) );
  INHSV4 U34568 ( .I(n38664), .ZN(n38048) );
  BUFHSV4 U34569 ( .I(n29742), .Z(n46587) );
  INHSV6 U34570 ( .I(\pe6/aot [20]), .ZN(n35607) );
  BUFHSV8 U34571 ( .I(n31958), .Z(n44476) );
  BUFHSV4 U34572 ( .I(n59917), .Z(n58886) );
  INHSV4 U34573 ( .I(n52080), .ZN(n52294) );
  INHSV4 U34574 ( .I(n42361), .ZN(n42132) );
  BUFHSV8 U34575 ( .I(\pe4/bq[4] ), .Z(n58156) );
  INHSV6 U34576 ( .I(n55082), .ZN(n55214) );
  INHSV6 U34577 ( .I(\pe2/aot [22]), .ZN(n44871) );
  INHSV6 U34578 ( .I(n44871), .ZN(n37801) );
  OR2HSV4 U34579 ( .A1(n44322), .A2(n45099), .Z(n36277) );
  INHSV4 U34580 ( .I(\pe4/bq[14] ), .ZN(n53217) );
  INHSV4 U34581 ( .I(n53217), .ZN(n58069) );
  INHSV4 U34582 ( .I(n40412), .ZN(n44569) );
  INHSV2 U34583 ( .I(n53957), .ZN(n59385) );
  INHSV2 U34584 ( .I(n40787), .ZN(n41145) );
  BUFHSV8 U34585 ( .I(\pe3/aot [4]), .Z(n59646) );
  INHSV4 U34586 ( .I(n39405), .ZN(n39245) );
  INHSV2 U34587 ( .I(n39741), .ZN(n39239) );
  INHSV4 U34588 ( .I(n41453), .ZN(n42231) );
  INHSV8 U34589 ( .I(n58530), .ZN(n58459) );
  CLKNHSV0 U34590 ( .I(n36512), .ZN(n36514) );
  INHSV4 U34591 ( .I(n41418), .ZN(n41230) );
  BUFHSV4 U34592 ( .I(n32198), .Z(n36161) );
  BUFHSV4 U34593 ( .I(n53214), .Z(n48046) );
  BUFHSV4 U34594 ( .I(n52727), .Z(n55826) );
  INHSV4 U34595 ( .I(n54973), .ZN(n48380) );
  BUFHSV4 U34596 ( .I(n37659), .Z(n48168) );
  INHSV4 U34597 ( .I(n36901), .ZN(n45622) );
  INHSV8 U34598 ( .I(\pe6/bq[19] ), .ZN(n44397) );
  INHSV4 U34599 ( .I(n44397), .ZN(n59224) );
  INHSV4 U34600 ( .I(n44397), .ZN(n59051) );
  INHSV4 U34601 ( .I(n33522), .ZN(n35295) );
  BUFHSV4 U34602 ( .I(\pe1/aot [25]), .Z(n53848) );
  BUFHSV4 U34603 ( .I(\pe1/aot [25]), .Z(n41743) );
  BUFHSV4 U34604 ( .I(n42938), .Z(n48488) );
  BUFHSV8 U34605 ( .I(n37176), .Z(n42938) );
  INHSV4 U34606 ( .I(n40012), .ZN(n37551) );
  BUFHSV4 U34607 ( .I(n48043), .Z(n59902) );
  BUFHSV4 U34608 ( .I(\pe3/bq[24] ), .Z(n55872) );
  BUFHSV4 U34609 ( .I(\pe3/bq[24] ), .Z(n43052) );
  INHSV2 U34610 ( .I(n41931), .ZN(n54500) );
  INHSV2 U34611 ( .I(n33282), .ZN(n33694) );
  INHSV4 U34612 ( .I(n35303), .ZN(n34843) );
  INHSV6 U34613 ( .I(\pe6/aot [15]), .ZN(n44396) );
  INHSV8 U34614 ( .I(n44396), .ZN(n58842) );
  INHSV2 U34615 ( .I(n53672), .ZN(n55103) );
  INHSV6 U34616 ( .I(\pe1/got [27]), .ZN(n44337) );
  INHSV6 U34617 ( .I(\pe5/aot [7]), .ZN(n47230) );
  INHSV4 U34618 ( .I(n39772), .ZN(n30222) );
  INHSV4 U34619 ( .I(n39772), .ZN(n30542) );
  BUFHSV8 U34620 ( .I(n56071), .Z(n55976) );
  BUFHSV4 U34621 ( .I(n56071), .Z(n48520) );
  BUFHSV8 U34622 ( .I(\pe3/bq[25] ), .Z(n56071) );
  BUFHSV4 U34623 ( .I(\pe6/aot [6]), .Z(n53134) );
  INHSV6 U34624 ( .I(\pe4/bq[8] ), .ZN(n48028) );
  INHSV12 U34625 ( .I(n45810), .ZN(n42971) );
  BUFHSV8 U34626 ( .I(\pe3/aot [6]), .Z(n45973) );
  INHSV4 U34627 ( .I(n47575), .ZN(n39029) );
  BUFHSV2 U34628 ( .I(\pe3/bq[7] ), .Z(n56832) );
  BUFHSV4 U34629 ( .I(n43211), .Z(n46313) );
  INHSV6 U34630 ( .I(\pe6/bq[11] ), .ZN(n46850) );
  INHSV4 U34631 ( .I(n46850), .ZN(n35750) );
  INHSV4 U34632 ( .I(n46850), .ZN(n46210) );
  BUFHSV4 U34633 ( .I(n59725), .Z(n54557) );
  INHSV4 U34634 ( .I(n34571), .ZN(n34565) );
  INHSV4 U34635 ( .I(n49003), .ZN(n32009) );
  INHSV4 U34636 ( .I(n58463), .ZN(n58488) );
  BUFHSV8 U34637 ( .I(n49966), .Z(n57675) );
  BUFHSV4 U34638 ( .I(\pe3/aot [15]), .Z(n55864) );
  BUFHSV4 U34639 ( .I(\pe3/aot [15]), .Z(n56651) );
  BUFHSV4 U34640 ( .I(\pe3/aot [15]), .Z(n56378) );
  INHSV4 U34641 ( .I(n50428), .ZN(n39615) );
  INHSV6 U34642 ( .I(\pe3/bq[20] ), .ZN(n45810) );
  INHSV6 U34643 ( .I(\pe1/aot [1]), .ZN(n55524) );
  BUFHSV4 U34644 ( .I(n47058), .Z(n47338) );
  INHSV6 U34645 ( .I(\pe5/aot [17]), .ZN(n50518) );
  INHSV4 U34646 ( .I(\pe4/got [20]), .ZN(n33860) );
  INHSV6 U34647 ( .I(n33860), .ZN(n59386) );
  INHSV6 U34648 ( .I(\pe6/aot [14]), .ZN(n32858) );
  BUFHSV4 U34649 ( .I(n32466), .Z(n35907) );
  INHSV6 U34650 ( .I(\pe1/aot [19]), .ZN(n44705) );
  NOR2HSV0 U34651 ( .A1(n40542), .A2(n40541), .ZN(n29715) );
  INHSV6 U34652 ( .I(\pe5/aot [11]), .ZN(n48204) );
  INHSV6 U34653 ( .I(\pe1/aot [17]), .ZN(n54829) );
  INHSV6 U34654 ( .I(\pe1/aot [10]), .ZN(n54846) );
  INHSV6 U34655 ( .I(\pe3/aot [12]), .ZN(n53229) );
  XNOR3HSV2 U34656 ( .A1(n30295), .A2(n30294), .A3(n30293), .ZN(n29716) );
  INHSV4 U34657 ( .I(n54281), .ZN(n53571) );
  INHSV4 U34658 ( .I(n47524), .ZN(n39019) );
  CLKNHSV0 U34659 ( .I(n30207), .ZN(n30203) );
  BUFHSV4 U34660 ( .I(n30297), .Z(n30595) );
  INHSV4 U34661 ( .I(n39163), .ZN(n30029) );
  INHSV4 U34662 ( .I(n40169), .ZN(n52799) );
  INHSV8 U34663 ( .I(\pe4/bq[19] ), .ZN(n48022) );
  INHSV4 U34664 ( .I(n48022), .ZN(n50250) );
  INHSV6 U34665 ( .I(n48022), .ZN(n57929) );
  INHSV4 U34666 ( .I(n48022), .ZN(n57368) );
  BUFHSV4 U34667 ( .I(\pe6/aot [2]), .Z(n58464) );
  INHSV4 U34668 ( .I(n42196), .ZN(n40781) );
  BUFHSV4 U34669 ( .I(\pe1/bq[8] ), .Z(n53708) );
  INHSV2 U34670 ( .I(n30320), .ZN(n30874) );
  INHSV4 U34671 ( .I(\pe2/got [16]), .ZN(n43999) );
  INHSV8 U34672 ( .I(n52526), .ZN(n51796) );
  INHSV2 U34673 ( .I(\pe4/aot [6]), .ZN(n47802) );
  INHSV4 U34674 ( .I(n47802), .ZN(n57338) );
  INHSV4 U34675 ( .I(n47809), .ZN(n57926) );
  INHSV6 U34676 ( .I(n47809), .ZN(n57850) );
  INHSV8 U34677 ( .I(\pe3/bq[16] ), .ZN(n46138) );
  INHSV4 U34678 ( .I(n46138), .ZN(n43544) );
  INHSV8 U34679 ( .I(\pe3/bq[17] ), .ZN(n55755) );
  INHSV6 U34680 ( .I(n55755), .ZN(n56433) );
  INHSV2 U34681 ( .I(n55755), .ZN(n56519) );
  INHSV4 U34682 ( .I(n49315), .ZN(n59174) );
  INHSV4 U34683 ( .I(n49315), .ZN(n35812) );
  INHSV4 U34684 ( .I(n31029), .ZN(n40190) );
  INHSV4 U34685 ( .I(n39733), .ZN(n30322) );
  INHSV6 U34686 ( .I(\pe6/aot [16]), .ZN(n46789) );
  INHSV4 U34687 ( .I(n46789), .ZN(n35732) );
  CLKNHSV6 U34688 ( .I(n58433), .ZN(n59182) );
  INHSV6 U34689 ( .I(\pe5/aot [20]), .ZN(n45815) );
  INHSV6 U34690 ( .I(n45815), .ZN(n52591) );
  INHSV6 U34691 ( .I(n45815), .ZN(n30788) );
  CLKAND2HSV2 U34692 ( .A1(n42507), .A2(n59964), .Z(n29717) );
  BUFHSV4 U34693 ( .I(\pe1/bq[17] ), .Z(n54995) );
  BUFHSV4 U34694 ( .I(n54995), .Z(n42098) );
  INHSV4 U34695 ( .I(n57841), .ZN(n58077) );
  INHSV4 U34696 ( .I(n57841), .ZN(n57986) );
  BUFHSV4 U34697 ( .I(\pe6/got [14]), .Z(n35991) );
  OA21HSV4 U34698 ( .A1(n33779), .A2(\pe4/ti_7t [12]), .B(n33676), .Z(n29718)
         );
  INHSV6 U34699 ( .I(\pe1/aot [23]), .ZN(n46142) );
  INHSV4 U34700 ( .I(n46142), .ZN(n53954) );
  INHSV2 U34701 ( .I(n46142), .ZN(n42255) );
  BUFHSV4 U34702 ( .I(n58661), .Z(n58478) );
  BUFHSV8 U34703 ( .I(\pe4/aot [11]), .Z(n59683) );
  BUFHSV4 U34704 ( .I(\pe6/bq[2] ), .Z(n58360) );
  BUFHSV4 U34705 ( .I(\pe6/bq[2] ), .Z(n59041) );
  INHSV2 U34706 ( .I(n52200), .ZN(n53019) );
  INHSV6 U34707 ( .I(n52200), .ZN(n59768) );
  INHSV6 U34708 ( .I(\pe3/got [28]), .ZN(n37273) );
  INHSV4 U34709 ( .I(n37041), .ZN(n45941) );
  BUFHSV4 U34710 ( .I(n37273), .Z(n36799) );
  INHSV4 U34711 ( .I(n49327), .ZN(n49205) );
  INHSV4 U34712 ( .I(n46750), .ZN(n46283) );
  INHSV4 U34713 ( .I(n46750), .ZN(n31710) );
  INHSV6 U34714 ( .I(\pe5/aot [22]), .ZN(n45451) );
  INHSV2 U34715 ( .I(n46283), .ZN(n44507) );
  CLKNHSV0 U34716 ( .I(n30590), .ZN(n30589) );
  CLKNHSV0 U34717 ( .I(n39669), .ZN(n47946) );
  CLKAND2HSV2 U34718 ( .A1(n32025), .A2(n49736), .Z(n29719) );
  INHSV4 U34719 ( .I(n51306), .ZN(n51161) );
  INHSV4 U34720 ( .I(n36574), .ZN(n38108) );
  INHSV4 U34721 ( .I(n35777), .ZN(n35705) );
  CLKNHSV6 U34722 ( .I(n58194), .ZN(n58283) );
  INHSV6 U34723 ( .I(\pe2/bq[11] ), .ZN(n47508) );
  INHSV6 U34724 ( .I(n47508), .ZN(n51900) );
  INHSV6 U34725 ( .I(n47508), .ZN(n52073) );
  INHSV2 U34726 ( .I(n38195), .ZN(n36654) );
  INHSV6 U34727 ( .I(\pe6/got [8]), .ZN(n58433) );
  INHSV4 U34728 ( .I(n58433), .ZN(n58526) );
  INHSV6 U34729 ( .I(\pe1/aot [6]), .ZN(n54901) );
  INHSV2 U34730 ( .I(n54901), .ZN(n55234) );
  INHSV6 U34731 ( .I(\pe2/bq[13] ), .ZN(n49628) );
  INHSV2 U34732 ( .I(n43469), .ZN(n42815) );
  INHSV8 U34733 ( .I(\pe5/got [26]), .ZN(n31081) );
  INHSV4 U34734 ( .I(n31081), .ZN(n30685) );
  INHSV12 U34735 ( .I(n31081), .ZN(n48742) );
  BUFHSV8 U34736 ( .I(\pe4/bq[10] ), .Z(n58116) );
  INHSV4 U34737 ( .I(n39743), .ZN(n59948) );
  INHSV4 U34738 ( .I(n59641), .ZN(n48681) );
  BUFHSV4 U34739 ( .I(n35991), .Z(n49741) );
  INHSV4 U34740 ( .I(n30583), .ZN(n39382) );
  AND2HSV2 U34741 ( .A1(n37645), .A2(n59507), .Z(n30063) );
  INHSV4 U34742 ( .I(n57776), .ZN(n59954) );
  BUFHSV8 U34743 ( .I(\pe6/got [12]), .Z(n59180) );
  BUFHSV4 U34744 ( .I(n52694), .Z(n52767) );
  BUFHSV8 U34745 ( .I(n59507), .Z(n52694) );
  INHSV6 U34746 ( .I(\pe2/bq[10] ), .ZN(n49515) );
  INHSV4 U34747 ( .I(n49515), .ZN(n52063) );
  INHSV4 U34748 ( .I(n49515), .ZN(n51997) );
  BUFHSV4 U34749 ( .I(\pe3/aot [7]), .Z(n56864) );
  BUFHSV4 U34750 ( .I(\pe3/aot [7]), .Z(n56221) );
  BUFHSV4 U34751 ( .I(\pe3/aot [7]), .Z(n59627) );
  INHSV2 U34752 ( .I(n34019), .ZN(n33928) );
  INHSV4 U34753 ( .I(n32640), .ZN(n33061) );
  CLKNHSV0 U34754 ( .I(n41218), .ZN(n41135) );
  BUFHSV4 U34755 ( .I(\pe5/aot [8]), .Z(n52675) );
  BUFHSV4 U34756 ( .I(n59880), .Z(n53296) );
  BUFHSV4 U34757 ( .I(\pe1/aot [4]), .Z(n55433) );
  BUFHSV4 U34758 ( .I(\pe1/aot [4]), .Z(n59619) );
  INHSV2 U34759 ( .I(n33848), .ZN(n33993) );
  INHSV4 U34760 ( .I(n34220), .ZN(n34221) );
  INHSV4 U34761 ( .I(n33522), .ZN(n35483) );
  INHSV4 U34762 ( .I(n41712), .ZN(n42488) );
  BUFHSV4 U34763 ( .I(\pe4/aot [7]), .Z(n59632) );
  INHSV6 U34764 ( .I(n35042), .ZN(n58198) );
  BUFHSV4 U34765 ( .I(n42362), .Z(n55307) );
  INHSV6 U34766 ( .I(\pe2/bq[9] ), .ZN(n47511) );
  INHSV4 U34767 ( .I(n47511), .ZN(n51623) );
  INHSV8 U34768 ( .I(\pe3/bq[6] ), .ZN(n49258) );
  INHSV6 U34769 ( .I(n49258), .ZN(n56915) );
  INHSV2 U34770 ( .I(n49258), .ZN(n56272) );
  INHSV6 U34771 ( .I(\pe4/bq[6] ), .ZN(n50351) );
  INHSV4 U34772 ( .I(n50351), .ZN(n58265) );
  BUFHSV4 U34773 ( .I(\pe1/aot [8]), .Z(n55452) );
  BUFHSV4 U34774 ( .I(\pe1/aot [8]), .Z(n54904) );
  INHSV4 U34775 ( .I(n53723), .ZN(n54847) );
  INHSV2 U34776 ( .I(n53723), .ZN(n55379) );
  INHSV4 U34777 ( .I(n34423), .ZN(n34419) );
  INHSV2 U34778 ( .I(n36671), .ZN(n43483) );
  OR2HSV1 U34779 ( .A1(n42798), .A2(n43880), .Z(n29720) );
  INHSV4 U34780 ( .I(\pe6/aot [4]), .ZN(n58530) );
  INHSV2 U34781 ( .I(n30864), .ZN(n37638) );
  INHSV4 U34782 ( .I(n49272), .ZN(n56827) );
  INHSV4 U34783 ( .I(n49272), .ZN(n56454) );
  INHSV4 U34784 ( .I(n52285), .ZN(n38778) );
  INHSV4 U34785 ( .I(n30966), .ZN(n39692) );
  INHSV4 U34786 ( .I(n41650), .ZN(n42093) );
  INHSV4 U34787 ( .I(n41650), .ZN(n41768) );
  INHSV2 U34788 ( .I(n39693), .ZN(n40009) );
  INHSV6 U34789 ( .I(\pe4/bq[3] ), .ZN(n57010) );
  INHSV6 U34790 ( .I(n57010), .ZN(n58196) );
  INHSV8 U34791 ( .I(n57010), .ZN(n58301) );
  INHSV4 U34792 ( .I(n40719), .ZN(n59994) );
  INHSV6 U34793 ( .I(\pe3/got [13]), .ZN(n46406) );
  INHSV4 U34794 ( .I(n46406), .ZN(n43829) );
  INHSV4 U34795 ( .I(n46406), .ZN(n56421) );
  INHSV2 U34796 ( .I(n45755), .ZN(n43361) );
  INHSV2 U34797 ( .I(n47963), .ZN(n34233) );
  INHSV2 U34798 ( .I(n32344), .ZN(n47970) );
  INHSV4 U34799 ( .I(n39222), .ZN(n40006) );
  BUFHSV4 U34800 ( .I(n33097), .Z(n33785) );
  INHSV4 U34801 ( .I(n33403), .ZN(n33588) );
  INHSV4 U34802 ( .I(n32053), .ZN(n51438) );
  INHSV2 U34803 ( .I(n29742), .ZN(n36066) );
  BUFHSV6 U34804 ( .I(\pe5/aot [4]), .Z(n50501) );
  INHSV4 U34805 ( .I(n30431), .ZN(n31225) );
  INHSV4 U34806 ( .I(n32044), .ZN(n33079) );
  INHSV4 U34807 ( .I(n31298), .ZN(n32941) );
  INHSV8 U34808 ( .I(n42086), .ZN(n41689) );
  INHSV4 U34809 ( .I(n42086), .ZN(n40605) );
  INHSV6 U34810 ( .I(\pe6/aot [9]), .ZN(n58537) );
  INHSV2 U34811 ( .I(n58537), .ZN(n58999) );
  INHSV6 U34812 ( .I(\pe6/got [17]), .ZN(n53103) );
  INHSV4 U34813 ( .I(n53103), .ZN(n49098) );
  INHSV4 U34814 ( .I(\pe2/aot [9]), .ZN(n52200) );
  INHSV6 U34815 ( .I(n49922), .ZN(n59663) );
  INHSV4 U34816 ( .I(n38902), .ZN(n38723) );
  INHSV6 U34817 ( .I(n49603), .ZN(n44944) );
  INHSV6 U34818 ( .I(n57830), .ZN(n57564) );
  INHSV4 U34819 ( .I(n31101), .ZN(n31102) );
  INHSV6 U34820 ( .I(\pe3/got [16]), .ZN(n45576) );
  INHSV4 U34821 ( .I(n45576), .ZN(n49252) );
  INHSV4 U34822 ( .I(n41928), .ZN(n59995) );
  INHSV4 U34823 ( .I(\pe5/aot [3]), .ZN(n59869) );
  INHSV4 U34824 ( .I(\pe2/aot [2]), .ZN(n49618) );
  INHSV4 U34825 ( .I(n43021), .ZN(n43132) );
  BUFHSV4 U34826 ( .I(n32242), .Z(n59025) );
  INHSV8 U34827 ( .I(\pe4/got [23]), .ZN(n35488) );
  INHSV6 U34828 ( .I(\pe4/got [27]), .ZN(n34452) );
  INHSV2 U34829 ( .I(n33748), .ZN(n33749) );
  INHSV4 U34830 ( .I(n46146), .ZN(n58731) );
  BUFHSV4 U34831 ( .I(n32970), .Z(n59165) );
  INHSV6 U34832 ( .I(\pe4/aot [8]), .ZN(n57775) );
  INHSV2 U34833 ( .I(n57775), .ZN(n57993) );
  BUFHSV2 U34834 ( .I(\pe6/got [9]), .Z(n58658) );
  INHSV6 U34835 ( .I(\pe5/got [13]), .ZN(n45817) );
  BUFHSV4 U34836 ( .I(n58562), .Z(n58709) );
  INHSV2 U34837 ( .I(n29825), .ZN(n39246) );
  BUFHSV8 U34838 ( .I(n40437), .Z(n42335) );
  BUFHSV4 U34839 ( .I(\pe6/got [15]), .Z(n32596) );
  INHSV6 U34840 ( .I(\pe5/aot [2]), .ZN(n51232) );
  INHSV4 U34841 ( .I(n51232), .ZN(n53203) );
  INHSV4 U34842 ( .I(n51235), .ZN(n51276) );
  INHSV4 U34843 ( .I(n51235), .ZN(n53199) );
  INHSV2 U34844 ( .I(n38603), .ZN(n44156) );
  BUFHSV4 U34845 ( .I(\pe6/got [3]), .Z(n58527) );
  BUFHSV4 U34846 ( .I(\pe6/got [3]), .Z(n48891) );
  INHSV4 U34847 ( .I(n54399), .ZN(n55577) );
  INHSV8 U34848 ( .I(\pe3/bq[8] ), .ZN(n49272) );
  INHSV2 U34849 ( .I(n49272), .ZN(n55970) );
  INHSV4 U34850 ( .I(n47905), .ZN(n58230) );
  INHSV6 U34851 ( .I(\pe2/bq[5] ), .ZN(n51131) );
  INHSV6 U34852 ( .I(n51131), .ZN(n51897) );
  INHSV2 U34853 ( .I(n51131), .ZN(n52857) );
  OR2HSV1 U34854 ( .A1(n43477), .A2(n42806), .Z(n29721) );
  INHSV4 U34855 ( .I(n48495), .ZN(n56892) );
  INHSV6 U34856 ( .I(\pe5/aot [5]), .ZN(n47409) );
  INHSV4 U34857 ( .I(n47409), .ZN(n59945) );
  INHSV8 U34858 ( .I(\pe3/bq[5] ), .ZN(n56914) );
  INHSV4 U34859 ( .I(n56914), .ZN(n56937) );
  INHSV2 U34860 ( .I(n42683), .ZN(n43234) );
  INHSV6 U34861 ( .I(\pe1/bq[7] ), .ZN(n54093) );
  INHSV6 U34862 ( .I(\pe1/bq[6] ), .ZN(n55523) );
  INHSV8 U34863 ( .I(\pe5/bq[5] ), .ZN(n51021) );
  INHSV4 U34864 ( .I(n51021), .ZN(n52671) );
  INHSV2 U34865 ( .I(n51021), .ZN(n51373) );
  INHSV4 U34866 ( .I(\pe6/got [21]), .ZN(n49826) );
  INHSV6 U34867 ( .I(\pe2/bq[7] ), .ZN(n49529) );
  INHSV4 U34868 ( .I(n49529), .ZN(n51832) );
  INHSV2 U34869 ( .I(n49529), .ZN(n52859) );
  INHSV2 U34870 ( .I(n58174), .ZN(n58070) );
  INHSV4 U34871 ( .I(n58174), .ZN(n59352) );
  AND2HSV2 U34872 ( .A1(\pe5/ti_7t [21]), .A2(n39730), .Z(n29722) );
  INHSV6 U34873 ( .I(\pe5/bq[8] ), .ZN(n46916) );
  INHSV4 U34874 ( .I(n46916), .ZN(n50675) );
  INHSV2 U34875 ( .I(n46916), .ZN(n52672) );
  OA21HSV2 U34876 ( .A1(n39007), .A2(n39102), .B(n59980), .Z(n29723) );
  INHSV4 U34877 ( .I(n44184), .ZN(n44145) );
  INHSV2 U34878 ( .I(n49000), .ZN(n45388) );
  CLKNHSV0 U34879 ( .I(n43139), .ZN(n43466) );
  NAND2HSV2 U34880 ( .A1(\pe3/ti_7t [22]), .A2(n43743), .ZN(n43139) );
  NAND2HSV2 U34881 ( .A1(n37771), .A2(n52799), .ZN(n29724) );
  INHSV4 U34882 ( .I(n52916), .ZN(n49000) );
  INHSV2 U34883 ( .I(n31381), .ZN(n35908) );
  INHSV4 U34884 ( .I(n35303), .ZN(n52755) );
  INHSV4 U34885 ( .I(n41835), .ZN(n41831) );
  CLKNHSV0 U34886 ( .I(n34837), .ZN(n34705) );
  CLKNAND2HSV2 U34887 ( .A1(n35806), .A2(\pe6/ti_7t [20]), .ZN(n29725) );
  INHSV2 U34888 ( .I(n47977), .ZN(n32156) );
  OR2HSV1 U34889 ( .A1(n41835), .A2(n41217), .Z(n29726) );
  INHSV4 U34890 ( .I(n37275), .ZN(n55945) );
  BUFHSV4 U34891 ( .I(n30992), .Z(n39741) );
  INHSV4 U34892 ( .I(n40130), .ZN(n30142) );
  INHSV8 U34893 ( .I(\pe1/bq[1] ), .ZN(n55185) );
  INHSV6 U34894 ( .I(n55185), .ZN(n55495) );
  INHSV8 U34895 ( .I(\pe3/bq[1] ), .ZN(n49275) );
  INHSV4 U34896 ( .I(n49275), .ZN(n56971) );
  INHSV4 U34897 ( .I(n49275), .ZN(n55857) );
  INHSV4 U34898 ( .I(n49275), .ZN(n56824) );
  INHSV4 U34899 ( .I(\pe3/aot [1]), .ZN(n56784) );
  BUFHSV8 U34900 ( .I(\pe3/aot [1]), .Z(n59511) );
  INHSV6 U34901 ( .I(n56784), .ZN(n56970) );
  BUFHSV4 U34902 ( .I(\pe6/got [4]), .Z(n58479) );
  INHSV4 U34903 ( .I(n45904), .ZN(n51339) );
  INHSV2 U34904 ( .I(n45904), .ZN(n51182) );
  INHSV6 U34905 ( .I(\pe6/got [22]), .ZN(n49003) );
  INHSV2 U34906 ( .I(n49003), .ZN(n59175) );
  INHSV6 U34907 ( .I(\pe5/got [24]), .ZN(n45900) );
  INHSV4 U34908 ( .I(n45900), .ZN(n59637) );
  INHSV4 U34909 ( .I(n45900), .ZN(n37631) );
  INHSV4 U34910 ( .I(n30888), .ZN(n52658) );
  INHSV8 U34911 ( .I(\pe3/got [22]), .ZN(n49314) );
  INHSV4 U34912 ( .I(n49314), .ZN(n48485) );
  INHSV4 U34913 ( .I(n49314), .ZN(n42770) );
  INHSV4 U34914 ( .I(n49314), .ZN(n55821) );
  INHSV4 U34915 ( .I(n49965), .ZN(n59601) );
  BUFHSV4 U34916 ( .I(n45091), .Z(n38514) );
  BUFHSV4 U34917 ( .I(n58527), .Z(n58423) );
  INHSV4 U34918 ( .I(n30516), .ZN(n40170) );
  INHSV6 U34919 ( .I(\pe4/got [13]), .ZN(n58189) );
  INHSV4 U34920 ( .I(n58189), .ZN(n35400) );
  INHSV2 U34921 ( .I(n58189), .ZN(n59629) );
  INHSV8 U34922 ( .I(\pe1/got [2]), .ZN(n55575) );
  INHSV4 U34923 ( .I(n55575), .ZN(n55340) );
  INHSV4 U34924 ( .I(n55575), .ZN(n59756) );
  INHSV6 U34925 ( .I(\pe3/got [25]), .ZN(n45948) );
  INHSV4 U34926 ( .I(n45948), .ZN(n46441) );
  INHSV4 U34927 ( .I(n42209), .ZN(n53390) );
  INHSV4 U34928 ( .I(n42209), .ZN(n54160) );
  INHSV8 U34929 ( .I(\pe2/got [22]), .ZN(n45248) );
  INHSV6 U34930 ( .I(\pe2/got [3]), .ZN(n53032) );
  INHSV2 U34931 ( .I(n57836), .ZN(n58041) );
  INHSV2 U34932 ( .I(n57836), .ZN(n57818) );
  INHSV2 U34933 ( .I(n57836), .ZN(n58140) );
  INHSV8 U34934 ( .I(\pe2/got [19]), .ZN(n47570) );
  INHSV6 U34935 ( .I(\pe4/got [10]), .ZN(n49922) );
  INHSV4 U34936 ( .I(n49922), .ZN(n57646) );
  BUFHSV4 U34937 ( .I(n44969), .Z(n49603) );
  INHSV8 U34938 ( .I(\pe4/got [12]), .ZN(n49954) );
  INHSV8 U34939 ( .I(\pe4/got [7]), .ZN(n50064) );
  INHSV8 U34940 ( .I(\pe2/bq[1] ), .ZN(n50920) );
  INHSV4 U34941 ( .I(n50920), .ZN(n51532) );
  INHSV4 U34942 ( .I(n50920), .ZN(n52851) );
  INHSV4 U34943 ( .I(n50920), .ZN(n51614) );
  INHSV6 U34944 ( .I(\pe4/got [16]), .ZN(n47793) );
  INHSV8 U34945 ( .I(\pe4/got [21]), .ZN(n50207) );
  BUFHSV8 U34946 ( .I(\pe6/got [10]), .Z(n44393) );
  BUFHSV4 U34947 ( .I(\pe6/got [10]), .Z(n58812) );
  INHSV6 U34948 ( .I(\pe6/got [11]), .ZN(n53110) );
  INHSV4 U34949 ( .I(n53110), .ZN(n49742) );
  INHSV2 U34950 ( .I(n36562), .ZN(n36563) );
  INHSV6 U34951 ( .I(\pe4/got [4]), .ZN(n50091) );
  INHSV4 U34952 ( .I(n49967), .ZN(n58300) );
  INHSV8 U34953 ( .I(\pe2/got [14]), .ZN(n47498) );
  INHSV6 U34954 ( .I(\pe4/got [22]), .ZN(n49965) );
  INHSV6 U34955 ( .I(\pe4/got [24]), .ZN(n50060) );
  INHSV2 U34956 ( .I(n59603), .ZN(n35319) );
  INHSV4 U34957 ( .I(n50060), .ZN(n33556) );
  INHSV8 U34958 ( .I(n50060), .ZN(n59603) );
  INHSV4 U34959 ( .I(n35319), .ZN(n57574) );
  INHSV6 U34960 ( .I(\pe4/got [15]), .ZN(n50212) );
  INHSV4 U34961 ( .I(n50212), .ZN(n57752) );
  INHSV4 U34962 ( .I(n50212), .ZN(n59664) );
  INHSV6 U34963 ( .I(\pe4/got [14]), .ZN(n50042) );
  BUFHSV4 U34964 ( .I(\pe6/got [13]), .Z(n58654) );
  BUFHSV4 U34965 ( .I(\pe6/got [13]), .Z(n58811) );
  BUFHSV8 U34966 ( .I(n58654), .Z(n58711) );
  INHSV4 U34967 ( .I(n48338), .ZN(n41676) );
  INHSV6 U34968 ( .I(\pe3/got [8]), .ZN(n56496) );
  INHSV12 U34969 ( .I(n56496), .ZN(n56855) );
  INHSV6 U34970 ( .I(\pe1/bq[2] ), .ZN(n53834) );
  INHSV4 U34971 ( .I(n47431), .ZN(n56975) );
  INHSV2 U34972 ( .I(n37766), .ZN(n37767) );
  INHSV8 U34973 ( .I(\pe4/got [19]), .ZN(n50052) );
  INHSV4 U34974 ( .I(n50052), .ZN(n50404) );
  INHSV4 U34975 ( .I(n50052), .ZN(n59602) );
  INHSV6 U34976 ( .I(\pe4/got [5]), .ZN(n50095) );
  INHSV4 U34977 ( .I(n50095), .ZN(n57677) );
  INHSV6 U34978 ( .I(n50095), .ZN(n58246) );
  INHSV4 U34979 ( .I(n58013), .ZN(n58322) );
  INHSV4 U34980 ( .I(n58013), .ZN(n57241) );
  INHSV6 U34981 ( .I(n48337), .ZN(n54724) );
  INHSV4 U34982 ( .I(n46583), .ZN(n52566) );
  INHSV4 U34983 ( .I(n46583), .ZN(n50495) );
  INHSV6 U34984 ( .I(\pe5/got [4]), .ZN(n50550) );
  INHSV4 U34985 ( .I(n50550), .ZN(n52577) );
  INHSV4 U34986 ( .I(n50550), .ZN(n51418) );
  INHSV4 U34987 ( .I(n52559), .ZN(n44709) );
  INHSV6 U34988 ( .I(\pe5/bq[3] ), .ZN(n48031) );
  INHSV2 U34989 ( .I(n48031), .ZN(n51281) );
  INHSV6 U34990 ( .I(\pe2/got [6]), .ZN(n52018) );
  INHSV4 U34991 ( .I(n52018), .ZN(n51939) );
  INHSV4 U34992 ( .I(n52018), .ZN(n59777) );
  INHSV4 U34993 ( .I(n58359), .ZN(n49847) );
  INHSV6 U34994 ( .I(\pe5/got [12]), .ZN(n46966) );
  INHSV12 U34995 ( .I(n46966), .ZN(n48167) );
  BUFHSV8 U34996 ( .I(\pe2/bq[2] ), .Z(n51805) );
  BUFHSV4 U34997 ( .I(n51805), .Z(n53226) );
  BUFHSV4 U34998 ( .I(n51493), .Z(n51919) );
  INHSV4 U34999 ( .I(n31199), .ZN(n53285) );
  INHSV8 U35000 ( .I(\pe1/got [10]), .ZN(n54636) );
  INHSV4 U35001 ( .I(n54636), .ZN(n55088) );
  INHSV4 U35002 ( .I(n54636), .ZN(n53473) );
  INHSV4 U35003 ( .I(n41392), .ZN(n53520) );
  INHSV4 U35004 ( .I(n33830), .ZN(n57754) );
  INHSV4 U35005 ( .I(n33830), .ZN(n57834) );
  INHSV4 U35006 ( .I(n46311), .ZN(n43457) );
  INHSV4 U35007 ( .I(\pe2/got [12]), .ZN(n47555) );
  INHSV6 U35008 ( .I(\pe5/got [20]), .ZN(n39119) );
  INHSV4 U35009 ( .I(n39119), .ZN(n40185) );
  INHSV4 U35010 ( .I(n32241), .ZN(n46289) );
  INHSV4 U35011 ( .I(n32949), .ZN(n46591) );
  INHSV2 U35012 ( .I(n35806), .ZN(n33089) );
  NAND2HSV0 U35013 ( .A1(n32949), .A2(\pe6/ti_7t [29]), .ZN(n29727) );
  INHSV4 U35014 ( .I(n36873), .ZN(n43743) );
  AND2HSV2 U35015 ( .A1(n33093), .A2(\pe4/ti_7t [30]), .Z(n29728) );
  CLKNHSV0 U35016 ( .I(n45760), .ZN(n46091) );
  BUFHSV4 U35017 ( .I(\pe4/ctrq ), .Z(n48082) );
  INHSV4 U35018 ( .I(n32047), .ZN(n46546) );
  INHSV4 U35019 ( .I(n47934), .ZN(n48013) );
  INHSV6 U35020 ( .I(\pe5/got [15]), .ZN(n48722) );
  INHSV4 U35021 ( .I(n48722), .ZN(n50643) );
  INHSV4 U35022 ( .I(n47935), .ZN(n52831) );
  INHSV6 U35023 ( .I(\pe1/got [15]), .ZN(n54263) );
  INHSV4 U35024 ( .I(n54263), .ZN(n54241) );
  INHSV4 U35025 ( .I(n54263), .ZN(n48339) );
  INHSV2 U35026 ( .I(n46613), .ZN(n48020) );
  BUFHSV4 U35027 ( .I(n46628), .Z(n30925) );
  INHSV4 U35028 ( .I(n47573), .ZN(n45289) );
  BUFHSV4 U35029 ( .I(n48029), .Z(n48039) );
  BUFHSV4 U35030 ( .I(n34496), .Z(n34054) );
  INHSV2 U35031 ( .I(n35493), .ZN(n47659) );
  BUFHSV4 U35032 ( .I(n48065), .Z(n53224) );
  BUFHSV4 U35033 ( .I(n48065), .Z(n48067) );
  BUFHSV4 U35034 ( .I(n48065), .Z(n53225) );
  INHSV6 U35035 ( .I(\pe1/got [9]), .ZN(n55163) );
  INHSV4 U35036 ( .I(n55163), .ZN(n55145) );
  INHSV4 U35037 ( .I(n55163), .ZN(n44605) );
  INHSV4 U35038 ( .I(n55163), .ZN(n55331) );
  BUFHSV4 U35039 ( .I(n48061), .Z(n48076) );
  BUFHSV4 U35040 ( .I(n46623), .Z(n48062) );
  BUFHSV4 U35041 ( .I(n48062), .Z(n53222) );
  BUFHSV4 U35042 ( .I(n48029), .Z(n53215) );
  INHSV6 U35043 ( .I(\pe1/got [8]), .ZN(n55227) );
  BUFHSV4 U35044 ( .I(n48078), .Z(n48079) );
  BUFHSV2 U35045 ( .I(n48043), .Z(n46621) );
  BUFHSV4 U35046 ( .I(n53218), .Z(n48068) );
  BUFHSV4 U35047 ( .I(n33808), .Z(n48058) );
  BUFHSV4 U35048 ( .I(n48036), .Z(n44701) );
  BUFHSV4 U35049 ( .I(n48036), .Z(n48043) );
  INHSV6 U35050 ( .I(\pe1/got [4]), .ZN(n55444) );
  INHSV4 U35051 ( .I(n55444), .ZN(n55410) );
  INHSV4 U35052 ( .I(n55444), .ZN(n53863) );
  INHSV4 U35053 ( .I(n55444), .ZN(n55267) );
  INHSV4 U35054 ( .I(n46750), .ZN(n59173) );
  INHSV6 U35055 ( .I(\pe1/got [11]), .ZN(n55082) );
  INHSV4 U35056 ( .I(n55082), .ZN(n54970) );
  INHSV2 U35057 ( .I(n51438), .ZN(n36029) );
  INHSV6 U35058 ( .I(\pe3/got [6]), .ZN(n56821) );
  INHSV4 U35059 ( .I(n56821), .ZN(n56779) );
  INHSV4 U35060 ( .I(n56821), .ZN(n56560) );
  INHSV4 U35061 ( .I(n50802), .ZN(n56618) );
  INHSV6 U35062 ( .I(\pe1/got [6]), .ZN(n55369) );
  INHSV6 U35063 ( .I(n55369), .ZN(n55448) );
  INHSV4 U35064 ( .I(n55369), .ZN(n53523) );
  INHSV6 U35065 ( .I(\pe3/got [4]), .ZN(n56904) );
  INHSV4 U35066 ( .I(n56904), .ZN(n56861) );
  INHSV6 U35067 ( .I(\pe1/got [3]), .ZN(n55364) );
  INHSV4 U35068 ( .I(n55364), .ZN(n55514) );
  INHSV4 U35069 ( .I(n30595), .ZN(n30779) );
  INHSV6 U35070 ( .I(\pe5/got [9]), .ZN(n46119) );
  INHSV4 U35071 ( .I(n46119), .ZN(n51358) );
  INHSV4 U35072 ( .I(n46119), .ZN(n59891) );
  INHSV6 U35073 ( .I(\pe3/got [3]), .ZN(n56906) );
  INHSV4 U35074 ( .I(n56906), .ZN(n56735) );
  INHSV6 U35075 ( .I(\pe5/got [7]), .ZN(n46978) );
  INHSV4 U35076 ( .I(n46978), .ZN(n59905) );
  INHSV4 U35077 ( .I(n56859), .ZN(n56822) );
  INHSV6 U35078 ( .I(\pe2/got [1]), .ZN(n50910) );
  INHSV4 U35079 ( .I(n50910), .ZN(n51688) );
  INHSV4 U35080 ( .I(\pe1/got [14]), .ZN(n54884) );
  INHSV6 U35081 ( .I(\pe3/got [2]), .ZN(n56936) );
  INHSV4 U35082 ( .I(n56936), .ZN(n56908) );
  INHSV6 U35083 ( .I(\pe2/got [13]), .ZN(n51607) );
  INHSV4 U35084 ( .I(n51607), .ZN(n52418) );
  INHSV6 U35085 ( .I(\pe3/got [7]), .ZN(n56778) );
  INHSV4 U35086 ( .I(n45727), .ZN(n56419) );
  INHSV8 U35087 ( .I(\pe4/got [6]), .ZN(n50214) );
  INHSV8 U35088 ( .I(n50214), .ZN(n58184) );
  INHSV6 U35089 ( .I(n50214), .ZN(n58137) );
  INHSV4 U35090 ( .I(n58253), .ZN(n57177) );
  INHSV6 U35091 ( .I(\pe3/got [10]), .ZN(n50756) );
  INHSV4 U35092 ( .I(n50756), .ZN(n56495) );
  INHSV6 U35093 ( .I(\pe2/got [2]), .ZN(n50926) );
  INHSV4 U35094 ( .I(n50799), .ZN(n56342) );
  INHSV6 U35095 ( .I(\pe5/got [17]), .ZN(n50422) );
  INHSV4 U35096 ( .I(n50422), .ZN(n59949) );
  INHSV6 U35097 ( .I(\pe2/got [7]), .ZN(n50928) );
  INHSV4 U35098 ( .I(n50928), .ZN(n52890) );
  INHSV6 U35099 ( .I(\pe6/got [20]), .ZN(n49739) );
  INHSV2 U35100 ( .I(n49739), .ZN(n59176) );
  INHSV6 U35101 ( .I(\pe5/got [5]), .ZN(n53292) );
  INHSV4 U35102 ( .I(n53292), .ZN(n51334) );
  INHSV6 U35103 ( .I(\pe2/got [5]), .ZN(n50908) );
  INHSV4 U35104 ( .I(n50908), .ZN(n59778) );
  INHSV4 U35105 ( .I(n54957), .ZN(n54812) );
  INHSV4 U35106 ( .I(n50909), .ZN(n52855) );
  INHSV4 U35107 ( .I(n50909), .ZN(n51896) );
  INHSV4 U35108 ( .I(n45281), .ZN(n59980) );
  INHSV4 U35109 ( .I(n45281), .ZN(n38873) );
  INHSV2 U35110 ( .I(n38873), .ZN(n38874) );
  INHSV6 U35111 ( .I(\pe5/got [11]), .ZN(n47143) );
  INHSV4 U35112 ( .I(n31883), .ZN(n36023) );
  INHSV2 U35113 ( .I(n31883), .ZN(n32148) );
  BUFHSV2 U35114 ( .I(n35797), .Z(n44519) );
  BUFHSV4 U35115 ( .I(n31461), .Z(n32463) );
  INHSV4 U35116 ( .I(n46961), .ZN(n53289) );
  INHSV4 U35117 ( .I(n48887), .ZN(n58336) );
  INHSV6 U35118 ( .I(\pe6/bq[29] ), .ZN(n46620) );
  INHSV2 U35119 ( .I(n35653), .ZN(n35768) );
  INHSV6 U35120 ( .I(\pe6/bq[7] ), .ZN(n48041) );
  CLKNHSV0 U35121 ( .I(n42603), .ZN(n52790) );
  CLKNHSV0 U35122 ( .I(n29734), .ZN(n48015) );
  CLKNHSV0 U35123 ( .I(n59400), .ZN(n48083) );
  CLKNHSV0 U35124 ( .I(n59397), .ZN(n59660) );
  CLKNHSV0 U35125 ( .I(n59660), .ZN(n29729) );
  CLKNHSV0 U35126 ( .I(n59660), .ZN(n29730) );
  OAI21HSV2 U35127 ( .A1(n57131), .A2(n33946), .B(n33945), .ZN(n33952) );
  INHSV4 U35128 ( .I(n35153), .ZN(n46581) );
  INHSV2 U35129 ( .I(n34463), .ZN(n35377) );
  NOR2HSV4 U35130 ( .A1(n34485), .A2(n34463), .ZN(n33115) );
  CLKNHSV0 U35131 ( .I(n59660), .ZN(n29731) );
  CLKNHSV0 U35132 ( .I(n48478), .ZN(n29732) );
  CLKNHSV0 U35133 ( .I(n48015), .ZN(n29733) );
  CLKNHSV0 U35134 ( .I(n48477), .ZN(n29734) );
  AOI21HSV0 U35135 ( .A1(n35316), .A2(n34327), .B(n33457), .ZN(n47963) );
  NOR2HSV0 U35136 ( .A1(n34970), .A2(n47777), .ZN(n34333) );
  INHSV4 U35137 ( .I(n42706), .ZN(n46519) );
  INHSV4 U35138 ( .I(n31440), .ZN(n52706) );
  NAND2HSV4 U35139 ( .A1(n41845), .A2(n41844), .ZN(n42317) );
  INHSV4 U35140 ( .I(\pe2/aot [5]), .ZN(n48622) );
  CLKNHSV0 U35141 ( .I(n31705), .ZN(n29737) );
  NAND2HSV4 U35142 ( .A1(n30994), .A2(n31126), .ZN(n31005) );
  NAND2HSV0 U35143 ( .A1(\pe4/bq[31] ), .A2(n34110), .ZN(n33253) );
  NAND2HSV2 U35144 ( .A1(n34110), .A2(n57476), .ZN(n33812) );
  INHSV4 U35145 ( .I(n33250), .ZN(n34110) );
  CLKNAND2HSV2 U35146 ( .A1(n37430), .A2(n37349), .ZN(n42584) );
  NAND2HSV2 U35147 ( .A1(n36579), .A2(n37918), .ZN(n36580) );
  NAND2HSV2 U35148 ( .A1(n56172), .A2(n56171), .ZN(n56259) );
  CLKNHSV0 U35149 ( .I(n37275), .ZN(n56171) );
  NOR2HSV0 U35150 ( .A1(n30106), .A2(n37635), .ZN(n30014) );
  NAND2HSV0 U35151 ( .A1(n29649), .A2(n44359), .ZN(n36097) );
  NAND2HSV2 U35152 ( .A1(n60028), .A2(n29681), .ZN(n44962) );
  CLKNHSV0 U35153 ( .I(n35462), .ZN(n29739) );
  INHSV2 U35154 ( .I(n47928), .ZN(n35462) );
  XNOR2HSV4 U35155 ( .A1(n33179), .A2(n33178), .ZN(n29740) );
  CLKNHSV0 U35156 ( .I(n44529), .ZN(n29741) );
  BUFHSV2 U35157 ( .I(n25463), .Z(n29742) );
  NAND2HSV4 U35158 ( .A1(n36415), .A2(n36414), .ZN(n29743) );
  NAND2HSV2 U35159 ( .A1(n38872), .A2(n38871), .ZN(n47539) );
  CLKNHSV0 U35160 ( .I(n42924), .ZN(n42919) );
  BUFHSV2 U35161 ( .I(n43344), .Z(n55917) );
  BUFHSV4 U35162 ( .I(n38163), .Z(n44143) );
  NOR2HSV2 U35163 ( .A1(n38164), .A2(n38163), .ZN(n38162) );
  BUFHSV4 U35164 ( .I(n45411), .Z(n38163) );
  NOR2HSV2 U35165 ( .A1(n45264), .A2(n45263), .ZN(n45272) );
  NOR2HSV2 U35166 ( .A1(n45401), .A2(n52411), .ZN(n45403) );
  NAND2HSV2 U35167 ( .A1(n45401), .A2(n38874), .ZN(n45405) );
  INHSV4 U35168 ( .I(n43598), .ZN(n29747) );
  INHSV4 U35169 ( .I(n43609), .ZN(n43598) );
  NAND2HSV2 U35170 ( .A1(n37528), .A2(n42509), .ZN(n59620) );
  CLKNAND2HSV2 U35171 ( .A1(n42510), .A2(n42509), .ZN(n42511) );
  CLKNHSV0 U35172 ( .I(n31894), .ZN(n29748) );
  NOR2HSV2 U35173 ( .A1(n37241), .A2(n37454), .ZN(n36840) );
  MUX2NHSV2 U35174 ( .I0(n33850), .I1(n33854), .S(n33851), .ZN(n60042) );
  CLKNHSV0 U35175 ( .I(n59347), .ZN(n46438) );
  INHSV2 U35176 ( .I(n45615), .ZN(n45618) );
  OAI21HSV2 U35177 ( .A1(n37162), .A2(n37161), .B(n45615), .ZN(n37248) );
  NAND2HSV0 U35178 ( .A1(n45615), .A2(n36892), .ZN(n36893) );
  BUFHSV6 U35179 ( .I(n37168), .Z(n45615) );
  AND2HSV2 U35180 ( .A1(n38629), .A2(\pe2/ti_7t [6]), .Z(n36520) );
  NAND2HSV0 U35181 ( .A1(n43453), .A2(n42936), .ZN(n43012) );
  NAND2HSV0 U35182 ( .A1(n37520), .A2(n42936), .ZN(n37521) );
  CLKNAND2HSV2 U35183 ( .A1(n44183), .A2(n44300), .ZN(n44155) );
  XNOR2HSV4 U35184 ( .A1(n32227), .A2(n32226), .ZN(n29751) );
  CLKNHSV2 U35185 ( .I(n49400), .ZN(n29753) );
  AOI21HSV2 U35186 ( .A1(n44029), .A2(n44034), .B(n44028), .ZN(n44036) );
  NAND2HSV2 U35187 ( .A1(n42052), .A2(n42041), .ZN(n29754) );
  NAND2HSV2 U35188 ( .A1(n42052), .A2(n42041), .ZN(n42049) );
  INHSV4 U35189 ( .I(n32960), .ZN(n29755) );
  INHSV2 U35190 ( .I(n32960), .ZN(n35921) );
  INHSV4 U35191 ( .I(n52831), .ZN(n41414) );
  CLKAND2HSV2 U35192 ( .A1(n48313), .A2(n48312), .Z(n48315) );
  CLKNAND2HSV4 U35193 ( .A1(n48313), .A2(n42341), .ZN(n42476) );
  CLKNHSV0 U35194 ( .I(n36631), .ZN(n29756) );
  CLKNAND2HSV8 U35195 ( .A1(n36469), .A2(n36468), .ZN(n36630) );
  OAI21HSV0 U35196 ( .A1(n43240), .A2(n45755), .B(n45615), .ZN(n43130) );
  NAND2HSV0 U35197 ( .A1(n39122), .A2(n30037), .ZN(n29961) );
  NAND2HSV0 U35198 ( .A1(n39122), .A2(n30547), .ZN(n30036) );
  NAND2HSV2 U35199 ( .A1(n39122), .A2(n30164), .ZN(n39889) );
  NAND2HSV0 U35200 ( .A1(n39122), .A2(n30222), .ZN(n30168) );
  OAI21HSV0 U35201 ( .A1(n29722), .A2(n39548), .B(n30142), .ZN(n39549) );
  CLKNHSV0 U35202 ( .I(n39548), .ZN(n39379) );
  INHSV2 U35203 ( .I(n39548), .ZN(n30755) );
  NAND2HSV2 U35204 ( .A1(n29995), .A2(n39548), .ZN(n29996) );
  BUFHSV8 U35205 ( .I(n30992), .Z(n39548) );
  CLKNHSV0 U35206 ( .I(n38444), .ZN(n38446) );
  INHSV2 U35207 ( .I(n34447), .ZN(n34814) );
  XNOR2HSV4 U35208 ( .A1(n41918), .A2(n29754), .ZN(n29760) );
  XNOR2HSV4 U35209 ( .A1(n40322), .A2(n40321), .ZN(n29761) );
  INHSV4 U35210 ( .I(n38972), .ZN(n38024) );
  INHSV2 U35211 ( .I(n41484), .ZN(n29762) );
  INHSV2 U35212 ( .I(n41484), .ZN(n29763) );
  CLKNHSV0 U35213 ( .I(n41484), .ZN(n41677) );
  CLKNHSV0 U35214 ( .I(n44311), .ZN(n29764) );
  NAND2HSV0 U35215 ( .A1(n39415), .A2(n39365), .ZN(n39361) );
  INHSV2 U35216 ( .I(n39415), .ZN(n39364) );
  NOR2HSV2 U35217 ( .A1(n37649), .A2(n39415), .ZN(n39234) );
  INHSV6 U35218 ( .I(n37547), .ZN(n39415) );
  INHSV2 U35219 ( .I(\pe4/aot [31]), .ZN(n34463) );
  CLKNHSV0 U35220 ( .I(n35004), .ZN(n29768) );
  CLKNHSV0 U35221 ( .I(n48892), .ZN(n33918) );
  CLKNHSV0 U35222 ( .I(n48892), .ZN(n34949) );
  XNOR2HSV1 U35223 ( .A1(n37527), .A2(n42617), .ZN(pov3[16]) );
  NAND2HSV0 U35224 ( .A1(n42502), .A2(n42690), .ZN(n42503) );
  XNOR2HSV4 U35225 ( .A1(n37345), .A2(n42690), .ZN(n60088) );
  NAND2HSV2 U35226 ( .A1(n42690), .A2(n37447), .ZN(n37449) );
  CLKNAND2HSV4 U35227 ( .A1(n39005), .A2(n39004), .ZN(n29769) );
  DELHS4 U35228 ( .I(n59513), .Z(n29770) );
  NAND2HSV2 U35229 ( .A1(n47427), .A2(n47426), .ZN(n29771) );
  NAND2HSV2 U35230 ( .A1(n47427), .A2(n47426), .ZN(n53210) );
  NAND2HSV4 U35231 ( .A1(n29765), .A2(n58383), .ZN(n59023) );
  CLKNHSV0 U35232 ( .I(n25326), .ZN(n59845) );
  CLKNHSV0 U35233 ( .I(n47972), .ZN(n59932) );
  BUFHSV2 U35234 ( .I(n47972), .Z(n57816) );
  INHSV4 U35235 ( .I(n49400), .ZN(n59528) );
  INHSV2 U35236 ( .I(n41484), .ZN(n29773) );
  CLKNHSV0 U35237 ( .I(n40874), .ZN(n41484) );
  INHSV4 U35238 ( .I(n44377), .ZN(n44387) );
  CLKNAND2HSV2 U35239 ( .A1(n40786), .A2(n40427), .ZN(n40431) );
  CLKNAND2HSV4 U35240 ( .A1(n43480), .A2(n43481), .ZN(n43609) );
  CLKNAND2HSV2 U35241 ( .A1(n31689), .A2(n31688), .ZN(n31693) );
  INHSV4 U35242 ( .I(n31402), .ZN(n48012) );
  NOR2HSV4 U35243 ( .A1(n42052), .A2(n42051), .ZN(n42062) );
  XNOR2HSV2 U35244 ( .A1(n43910), .A2(n43913), .ZN(n46089) );
  IOA21HSV2 U35245 ( .A1(n35434), .A2(n35437), .B(n35002), .ZN(n35003) );
  AOI21HSV4 U35246 ( .A1(n48335), .A2(n48334), .B(n48333), .ZN(n48459) );
  NAND2HSV2 U35247 ( .A1(n38323), .A2(n38389), .ZN(n38156) );
  INHSV2 U35248 ( .I(n31383), .ZN(n31325) );
  INHSV6 U35249 ( .I(n31383), .ZN(n31440) );
  CLKNAND2HSV4 U35250 ( .A1(n36412), .A2(n36413), .ZN(n36619) );
  CLKNAND2HSV8 U35251 ( .A1(n36335), .A2(n36334), .ZN(n36412) );
  INHSV4 U35252 ( .I(n39415), .ZN(n39671) );
  MUX2NHSV2 U35253 ( .I0(n36631), .I1(n29756), .S(n36629), .ZN(n60004) );
  NAND3HSV4 U35254 ( .A1(n42316), .A2(n42317), .A3(n48468), .ZN(n42186) );
  AND2HSV4 U35255 ( .A1(n32816), .A2(n59171), .Z(n32819) );
  AOI21HSV0 U35256 ( .A1(n30651), .A2(n30649), .B(n30653), .ZN(n30429) );
  CLKNHSV2 U35257 ( .I(n45924), .ZN(n29775) );
  CLKNHSV2 U35258 ( .I(n45924), .ZN(n29776) );
  CLKNHSV2 U35259 ( .I(n45924), .ZN(n29777) );
  CLKNHSV0 U35260 ( .I(n34207), .ZN(n34211) );
  INHSV2 U35261 ( .I(n34207), .ZN(n34013) );
  CLKNHSV0 U35262 ( .I(n35570), .ZN(n34955) );
  INHSV2 U35263 ( .I(n35570), .ZN(n57547) );
  INHSV4 U35264 ( .I(n57816), .ZN(n57985) );
  NOR2HSV8 U35265 ( .A1(n29755), .A2(n32962), .ZN(n33068) );
  NOR2HSV4 U35266 ( .A1(n42342), .A2(n42343), .ZN(n42477) );
  CLKNAND2HSV2 U35267 ( .A1(n34696), .A2(n34697), .ZN(n34723) );
  CLKNAND2HSV4 U35268 ( .A1(n34696), .A2(n34968), .ZN(n34435) );
  NAND2HSV4 U35269 ( .A1(n34335), .A2(n34334), .ZN(n34696) );
  INHSV4 U35270 ( .I(n29937), .ZN(n30106) );
  NOR2HSV4 U35271 ( .A1(n38907), .A2(n49603), .ZN(n36494) );
  OAI22HSV4 U35272 ( .A1(n39423), .A2(n39422), .B1(n39421), .B2(n47948), .ZN(
        n39425) );
  NAND2HSV4 U35273 ( .A1(n33693), .A2(n33692), .ZN(n33802) );
  OAI21HSV2 U35274 ( .A1(n33196), .A2(n33195), .B(n25876), .ZN(n29780) );
  NAND2HSV2 U35275 ( .A1(n44355), .A2(n36092), .ZN(n36094) );
  NAND2HSV2 U35276 ( .A1(n36203), .A2(n46289), .ZN(n36205) );
  OAI22HSV2 U35277 ( .A1(n34680), .A2(n34685), .B1(n35598), .B2(n34679), .ZN(
        n34681) );
  OAI21HSV2 U35278 ( .A1(n32438), .A2(n32437), .B(n32340), .ZN(n32440) );
  BUFHSV4 U35279 ( .I(n35721), .Z(n49318) );
  NAND2HSV4 U35280 ( .A1(n45945), .A2(n45944), .ZN(n46071) );
  NAND2HSV2 U35281 ( .A1(n40003), .A2(n40002), .ZN(n40005) );
  NOR2HSV4 U35282 ( .A1(n46298), .A2(n46297), .ZN(n58438) );
  AOI21HSV4 U35283 ( .A1(n36905), .A2(n42924), .B(n36904), .ZN(n36906) );
  NAND2HSV4 U35284 ( .A1(n29882), .A2(n29881), .ZN(n29888) );
  NOR2HSV0 U35285 ( .A1(n42512), .A2(n42511), .ZN(n42517) );
  CLKNAND2HSV8 U35286 ( .A1(n60067), .A2(n45414), .ZN(n51230) );
  XNOR2HSV4 U35287 ( .A1(n36428), .A2(n36427), .ZN(n36513) );
  INHSV2 U35288 ( .I(go2[32]), .ZN(n59341) );
  INHSV6 U35290 ( .I(\pe5/aot [32]), .ZN(n29959) );
  INHSV4 U35291 ( .I(n29959), .ZN(n30155) );
  NAND2HSV2 U35292 ( .A1(n30155), .A2(n30526), .ZN(n29783) );
  INHSV2 U35293 ( .I(n37584), .ZN(n48040) );
  INHSV2 U35294 ( .I(n48040), .ZN(n48752) );
  INHSV2 U35295 ( .I(\pe5/got [25]), .ZN(n30210) );
  NAND2HSV2 U35296 ( .A1(n48752), .A2(\pe5/got [25]), .ZN(n29782) );
  XOR2HSV0 U35297 ( .A1(n29783), .A2(n29782), .Z(n29787) );
  INHSV2 U35298 ( .I(n30163), .ZN(n59938) );
  INHSV2 U35299 ( .I(n30116), .ZN(n30164) );
  CLKNAND2HSV1 U35300 ( .A1(n59938), .A2(n30164), .ZN(n29785) );
  INHSV2 U35301 ( .I(n40235), .ZN(n30165) );
  INHSV2 U35302 ( .I(\pe5/bq[29] ), .ZN(n30032) );
  INHSV2 U35303 ( .I(n30032), .ZN(n29965) );
  CLKNAND2HSV0 U35304 ( .A1(n30165), .A2(n29965), .ZN(n29784) );
  XOR2HSV0 U35305 ( .A1(n29785), .A2(n29784), .Z(n29786) );
  XOR2HSV0 U35306 ( .A1(n29787), .A2(n29786), .Z(n29793) );
  INHSV4 U35307 ( .I(\pe5/aot [31]), .ZN(n39779) );
  INHSV2 U35308 ( .I(n39779), .ZN(n59937) );
  INHSV2 U35309 ( .I(\pe5/bq[26] ), .ZN(n39772) );
  INHSV2 U35310 ( .I(n39772), .ZN(n52594) );
  NAND2HSV2 U35311 ( .A1(n59937), .A2(n52594), .ZN(n29789) );
  INHSV2 U35312 ( .I(n48219), .ZN(n30147) );
  BUFHSV8 U35313 ( .I(n39163), .Z(n30223) );
  INHSV2 U35314 ( .I(n30223), .ZN(n48785) );
  NAND2HSV2 U35315 ( .A1(n30147), .A2(n48785), .ZN(n29788) );
  XOR2HSV0 U35316 ( .A1(n29789), .A2(n29788), .Z(n29791) );
  INHSV2 U35317 ( .I(n30113), .ZN(n47234) );
  NAND2HSV2 U35318 ( .A1(n59427), .A2(n47234), .ZN(n29790) );
  XNOR2HSV1 U35319 ( .A1(n29791), .A2(n29790), .ZN(n29792) );
  XOR2HSV0 U35320 ( .A1(n29793), .A2(n29792), .Z(n29934) );
  INHSV6 U35321 ( .I(\pe5/bq[32] ), .ZN(n29890) );
  NAND2HSV2 U35322 ( .A1(n29815), .A2(\pe5/aot [32]), .ZN(n29796) );
  NOR2HSV2 U35323 ( .A1(n30051), .A2(n29826), .ZN(n29794) );
  OAI21HSV2 U35324 ( .A1(n29826), .A2(n30051), .B(n29796), .ZN(n29797) );
  CLKNAND2HSV2 U35325 ( .A1(n29798), .A2(n29797), .ZN(n29805) );
  CLKNAND2HSV1 U35326 ( .A1(\pe5/pvq [1]), .A2(\pe5/phq [1]), .ZN(n29799) );
  NAND2HSV4 U35327 ( .A1(n29804), .A2(n29803), .ZN(n29812) );
  INHSV4 U35328 ( .I(ctro5), .ZN(n29851) );
  CLKBUFHSV4 U35329 ( .I(n29851), .Z(n30199) );
  CLKBUFHSV4 U35330 ( .I(n30199), .Z(n44520) );
  BUFHSV3 U35331 ( .I(n29851), .Z(n29907) );
  NAND2HSV2 U35332 ( .A1(n39702), .A2(\pe5/ti_7t [1]), .ZN(n29806) );
  NAND2HSV4 U35333 ( .A1(n29849), .A2(n29806), .ZN(n29937) );
  CLKNAND2HSV1 U35334 ( .A1(n59393), .A2(n30685), .ZN(n29810) );
  INHSV2 U35335 ( .I(n30150), .ZN(n52590) );
  NAND2HSV2 U35336 ( .A1(n52590), .A2(n30146), .ZN(n29808) );
  INHSV2 U35337 ( .I(\pe5/aot [27]), .ZN(n30358) );
  INHSV2 U35338 ( .I(n30358), .ZN(n59939) );
  INHSV2 U35339 ( .I(n29892), .ZN(n30367) );
  NAND2HSV2 U35340 ( .A1(n59939), .A2(n30367), .ZN(n29807) );
  XOR2HSV0 U35341 ( .A1(n29808), .A2(n29807), .Z(n29809) );
  CLKNHSV0 U35342 ( .I(\pe5/ctrq ), .ZN(n30100) );
  CLKBUFHSV4 U35343 ( .I(n48029), .Z(n46628) );
  NAND2HSV4 U35344 ( .A1(n29812), .A2(n29811), .ZN(n59398) );
  CLKBUFHSV4 U35345 ( .I(n29851), .Z(n30992) );
  CLKAND2HSV2 U35346 ( .A1(n30992), .A2(n37544), .Z(n30196) );
  CLKNAND2HSV3 U35347 ( .A1(n59398), .A2(n30196), .ZN(n29916) );
  BUFHSV8 U35348 ( .I(n29848), .Z(n29914) );
  NOR2HSV4 U35349 ( .A1(n29900), .A2(n29914), .ZN(n29813) );
  INHSV2 U35350 ( .I(n29813), .ZN(n29814) );
  INHSV4 U35351 ( .I(n29815), .ZN(n39797) );
  NOR2HSV4 U35352 ( .A1(n39797), .A2(n39779), .ZN(n29816) );
  XNOR2HSV4 U35353 ( .A1(n29818), .A2(n29817), .ZN(n29946) );
  NOR2HSV2 U35354 ( .A1(n29916), .A2(n29946), .ZN(n29820) );
  BUFHSV2 U35355 ( .I(n30992), .Z(n30318) );
  INHSV2 U35356 ( .I(\pe5/ti_7t [2]), .ZN(n29843) );
  OR2HSV1 U35357 ( .A1(n30318), .A2(n29843), .Z(n29917) );
  INHSV2 U35358 ( .I(n29917), .ZN(n29819) );
  INHSV2 U35359 ( .I(ctro5), .ZN(n30206) );
  BUFHSV2 U35360 ( .I(n30206), .Z(n39558) );
  NAND2HSV2 U35361 ( .A1(n59398), .A2(n37544), .ZN(n29913) );
  INHSV2 U35362 ( .I(n30431), .ZN(n30254) );
  CLKNAND2HSV1 U35363 ( .A1(n29889), .A2(n30254), .ZN(n29823) );
  XNOR2HSV1 U35364 ( .A1(n29824), .A2(n29823), .ZN(n29865) );
  INHSV2 U35365 ( .I(n30297), .ZN(n59947) );
  CLKBUFHSV4 U35366 ( .I(n29849), .Z(n29856) );
  INHSV4 U35367 ( .I(n29856), .ZN(n29842) );
  INHSV2 U35368 ( .I(n29946), .ZN(n29944) );
  BUFHSV2 U35369 ( .I(n29851), .Z(n39250) );
  INAND2HSV2 U35370 ( .A1(n29842), .B1(n29940), .ZN(n52717) );
  INHSV4 U35371 ( .I(n29937), .ZN(n30458) );
  BUFHSV2 U35372 ( .I(\pe5/got [31]), .Z(n29825) );
  NOR2HSV2 U35373 ( .A1(n30458), .A2(n30089), .ZN(n52713) );
  INHSV4 U35374 ( .I(\pe5/got [30]), .ZN(n30682) );
  INHSV4 U35375 ( .I(n30682), .ZN(n30098) );
  CLKNAND2HSV4 U35376 ( .A1(n29827), .A2(n30098), .ZN(n29876) );
  CLKNAND2HSV2 U35377 ( .A1(\pe5/ctrq ), .A2(\pe5/pvq [3]), .ZN(n29871) );
  XNOR2HSV4 U35378 ( .A1(n29876), .A2(n29871), .ZN(n29829) );
  INHSV2 U35379 ( .I(n29890), .ZN(n30033) );
  INHSV2 U35380 ( .I(n30212), .ZN(n29828) );
  NAND2HSV4 U35381 ( .A1(n30033), .A2(n29828), .ZN(n29872) );
  INHSV2 U35382 ( .I(n29872), .ZN(n29891) );
  XNOR2HSV4 U35383 ( .A1(n29829), .A2(n29891), .ZN(n29840) );
  INHSV6 U35384 ( .I(\pe5/aot [31]), .ZN(n30365) );
  INHSV6 U35385 ( .I(n30365), .ZN(n29999) );
  CLKNAND2HSV2 U35386 ( .A1(n29830), .A2(\pe5/phq [3]), .ZN(n29834) );
  INHSV2 U35387 ( .I(\pe5/phq [3]), .ZN(n29831) );
  CLKNAND2HSV3 U35388 ( .A1(n29832), .A2(n29831), .ZN(n29833) );
  CLKNAND2HSV3 U35389 ( .A1(n29833), .A2(n29834), .ZN(n29835) );
  NAND2HSV2 U35390 ( .A1(n30155), .A2(n30367), .ZN(n29877) );
  INHSV3 U35391 ( .I(n29835), .ZN(n29837) );
  INHSV2 U35392 ( .I(n29877), .ZN(n29836) );
  CLKNAND2HSV3 U35393 ( .A1(n29837), .A2(n29836), .ZN(n29838) );
  CLKNAND2HSV4 U35394 ( .A1(n29838), .A2(n29839), .ZN(n29847) );
  XNOR2HSV4 U35395 ( .A1(n29840), .A2(n29847), .ZN(n29948) );
  BUFHSV8 U35396 ( .I(n29948), .Z(n29855) );
  NAND2HSV2 U35397 ( .A1(n52713), .A2(n29855), .ZN(n29841) );
  INHSV2 U35398 ( .I(n30421), .ZN(n39871) );
  INHSV1 U35399 ( .I(n29944), .ZN(n52695) );
  INHSV2 U35400 ( .I(n30199), .ZN(n40310) );
  AOI21HSV4 U35401 ( .A1(n29843), .A2(n40310), .B(n39733), .ZN(n52716) );
  INHSV2 U35402 ( .I(n52716), .ZN(n29947) );
  NOR2HSV2 U35403 ( .A1(n29947), .A2(n39383), .ZN(n29844) );
  CLKNAND2HSV2 U35404 ( .A1(n52715), .A2(n29844), .ZN(n29845) );
  INHSV2 U35405 ( .I(n29845), .ZN(n29846) );
  BUFHSV2 U35406 ( .I(n25344), .Z(n40169) );
  BUFHSV4 U35407 ( .I(n25344), .Z(n30089) );
  NOR2HSV2 U35408 ( .A1(n29849), .A2(n29950), .ZN(n29850) );
  NAND2HSV2 U35409 ( .A1(n29945), .A2(n29850), .ZN(n29853) );
  BUFHSV2 U35410 ( .I(n29851), .Z(n30320) );
  BUFHSV2 U35411 ( .I(n30320), .Z(n39366) );
  CLKNHSV1 U35412 ( .I(n37766), .ZN(n29852) );
  CLKNAND2HSV2 U35413 ( .A1(n29853), .A2(n29852), .ZN(n29854) );
  CLKNAND2HSV1 U35414 ( .A1(n29858), .A2(n29859), .ZN(n29864) );
  CLKAND2HSV1 U35415 ( .A1(n52716), .A2(n29859), .Z(n29860) );
  INHSV2 U35416 ( .I(n29861), .ZN(n29862) );
  BUFHSV2 U35417 ( .I(n45477), .Z(n29866) );
  NAND3HSV2 U35418 ( .A1(n29865), .A2(n59947), .A3(n29866), .ZN(n29870) );
  INHSV1 U35419 ( .I(n29865), .ZN(n29868) );
  INHSV2 U35420 ( .I(n30297), .ZN(n39430) );
  NAND2HSV2 U35421 ( .A1(n29868), .A2(n29867), .ZN(n29869) );
  INHSV2 U35422 ( .I(n59398), .ZN(n29886) );
  NOR2HSV2 U35423 ( .A1(n29886), .A2(n30089), .ZN(n29887) );
  XNOR2HSV4 U35424 ( .A1(n29872), .A2(n29871), .ZN(n29875) );
  NOR2HSV2 U35425 ( .A1(n39779), .A2(n39163), .ZN(n29874) );
  CLKNAND2HSV1 U35426 ( .A1(n29999), .A2(\pe5/phq [3]), .ZN(n29873) );
  NAND2HSV2 U35427 ( .A1(n29878), .A2(n29675), .ZN(n29882) );
  INHSV4 U35428 ( .I(n29878), .ZN(n29880) );
  INHSV2 U35429 ( .I(n29675), .ZN(n29879) );
  MUX2NHSV1 U35430 ( .I0(n29886), .I1(n29887), .S(n29888), .ZN(n29885) );
  CLKNHSV0 U35431 ( .I(n29888), .ZN(n29883) );
  CLKNAND2HSV1 U35432 ( .A1(n29883), .A2(n30048), .ZN(n29884) );
  INHSV2 U35433 ( .I(n39548), .ZN(n39383) );
  INHSV2 U35434 ( .I(n39383), .ZN(n30139) );
  NOR2HSV2 U35435 ( .A1(n30864), .A2(\pe5/ti_7t [3]), .ZN(n29951) );
  NOR2HSV2 U35436 ( .A1(n29951), .A2(n39733), .ZN(n29988) );
  NAND3HSV4 U35437 ( .A1(n29989), .A2(n29990), .A3(n29988), .ZN(n29929) );
  BUFHSV3 U35438 ( .I(n29890), .Z(n39166) );
  INHSV4 U35439 ( .I(n30212), .ZN(n39122) );
  CLKNAND2HSV2 U35440 ( .A1(n30029), .A2(n39122), .ZN(n37664) );
  NOR2HSV4 U35441 ( .A1(n30223), .A2(n30163), .ZN(n29960) );
  CLKNAND2HSV1 U35442 ( .A1(n29960), .A2(n29891), .ZN(n29895) );
  NAND2HSV2 U35443 ( .A1(n30155), .A2(n29965), .ZN(n29894) );
  INHSV3 U35444 ( .I(n29892), .ZN(n30037) );
  XNOR2HSV4 U35445 ( .A1(n29894), .A2(n29893), .ZN(n29897) );
  NAND3HSV2 U35446 ( .A1(n29897), .A2(n29896), .A3(n29895), .ZN(n29898) );
  NAND2HSV2 U35447 ( .A1(n29899), .A2(n29898), .ZN(n29906) );
  NOR2HSV4 U35448 ( .A1(n40130), .A2(n29900), .ZN(n29902) );
  INHSV2 U35449 ( .I(\pe5/phq [4]), .ZN(n29901) );
  XNOR2HSV4 U35450 ( .A1(n29902), .A2(n29901), .ZN(n29904) );
  XNOR2HSV4 U35451 ( .A1(n29904), .A2(n29903), .ZN(n29905) );
  XNOR2HSV4 U35452 ( .A1(n29906), .A2(n29905), .ZN(n29912) );
  INHSV2 U35453 ( .I(n29907), .ZN(n31101) );
  CLKNHSV0 U35454 ( .I(\pe5/ti_7t [1]), .ZN(n29908) );
  INHSV2 U35455 ( .I(\pe5/got [30]), .ZN(n31116) );
  AOI21HSV2 U35456 ( .A1(n31101), .A2(n29908), .B(n31116), .ZN(n29909) );
  OAI21HSV2 U35457 ( .A1(n29910), .A2(n39702), .B(n29909), .ZN(n29911) );
  XNOR2HSV4 U35458 ( .A1(n29912), .A2(n29911), .ZN(n29923) );
  NOR2HSV4 U35459 ( .A1(n30976), .A2(n29914), .ZN(n39718) );
  NAND2HSV0 U35460 ( .A1(n29946), .A2(n39718), .ZN(n29922) );
  CLKNHSV0 U35461 ( .I(n29913), .ZN(n29921) );
  CLKNHSV0 U35462 ( .I(n29914), .ZN(n29915) );
  NOR2HSV2 U35463 ( .A1(n29916), .A2(n40293), .ZN(n29919) );
  NOR2HSV2 U35464 ( .A1(n29917), .A2(n40293), .ZN(n29918) );
  AOI21HSV4 U35465 ( .A1(n29944), .A2(n29919), .B(n29918), .ZN(n29920) );
  CLKNAND2HSV1 U35466 ( .A1(n29923), .A2(n29924), .ZN(n29928) );
  INHSV4 U35467 ( .I(n29923), .ZN(n29926) );
  INHSV2 U35468 ( .I(n29924), .ZN(n29925) );
  CLKNAND2HSV3 U35469 ( .A1(n29926), .A2(n29925), .ZN(n29927) );
  NAND2HSV4 U35470 ( .A1(n29927), .A2(n29928), .ZN(n29995) );
  NAND2HSV2 U35471 ( .A1(n29995), .A2(n25861), .ZN(n29931) );
  INHSV4 U35472 ( .I(n29929), .ZN(n29994) );
  INHSV4 U35473 ( .I(n29995), .ZN(n29992) );
  CLKNAND2HSV3 U35474 ( .A1(n29994), .A2(n29992), .ZN(n29930) );
  INHSV2 U35475 ( .I(n31101), .ZN(n39417) );
  INHSV2 U35476 ( .I(\pe5/ti_7t [4]), .ZN(n29978) );
  NOR2HSV2 U35477 ( .A1(n39403), .A2(n29978), .ZN(n29991) );
  BUFHSV2 U35478 ( .I(n40130), .Z(n30202) );
  NAND2HSV2 U35479 ( .A1(n30255), .A2(n30142), .ZN(n29932) );
  XOR3HSV2 U35480 ( .A1(n29934), .A2(n29933), .A3(n29932), .Z(n29987) );
  NAND2HSV2 U35481 ( .A1(n59393), .A2(n30142), .ZN(n29936) );
  INHSV2 U35482 ( .I(n29936), .ZN(n29935) );
  CLKNHSV2 U35483 ( .I(n29948), .ZN(n52714) );
  INHSV2 U35484 ( .I(n30320), .ZN(n30204) );
  NOR2HSV2 U35485 ( .A1(n29937), .A2(n30204), .ZN(n29938) );
  OAI21HSV2 U35486 ( .A1(n29948), .A2(n52716), .B(n29938), .ZN(n29939) );
  INHSV2 U35487 ( .I(n29940), .ZN(n29942) );
  NOR2HSV2 U35488 ( .A1(n29945), .A2(n29947), .ZN(n29941) );
  CLKNAND2HSV2 U35489 ( .A1(n29942), .A2(n29941), .ZN(n29956) );
  INHSV2 U35490 ( .I(n39718), .ZN(n39704) );
  NOR2HSV3 U35491 ( .A1(n30458), .A2(n39704), .ZN(n29943) );
  OAI21HSV2 U35492 ( .A1(n29945), .A2(n29944), .B(n29943), .ZN(n29954) );
  NOR2HSV2 U35493 ( .A1(n29951), .A2(n29950), .ZN(n29952) );
  AOI21HSV4 U35494 ( .A1(n29957), .A2(n29956), .B(n29955), .ZN(n29958) );
  CLKBUFHSV2 U35495 ( .I(n29959), .Z(n31044) );
  NAND2HSV2 U35496 ( .A1(n30165), .A2(n30146), .ZN(n29962) );
  XOR2HSV0 U35497 ( .A1(n29962), .A2(n29961), .Z(n29963) );
  XOR2HSV0 U35498 ( .A1(n29964), .A2(n29963), .Z(n29972) );
  NOR2HSV2 U35499 ( .A1(n30297), .A2(n48040), .ZN(n29967) );
  CLKNAND2HSV1 U35500 ( .A1(n29999), .A2(n29965), .ZN(n29966) );
  XOR2HSV0 U35501 ( .A1(n29967), .A2(n29966), .Z(n29970) );
  NAND2HSV2 U35502 ( .A1(n48049), .A2(\pe5/pvq [5]), .ZN(n29968) );
  XOR2HSV0 U35503 ( .A1(n29968), .A2(\pe5/phq [5]), .Z(n29969) );
  XOR2HSV0 U35504 ( .A1(n29970), .A2(n29969), .Z(n29971) );
  XOR2HSV0 U35505 ( .A1(n29972), .A2(n29971), .Z(n29973) );
  BUFHSV2 U35506 ( .I(n31116), .Z(n39240) );
  XNOR2HSV4 U35507 ( .A1(n29973), .A2(n29651), .ZN(n29975) );
  INHSV2 U35508 ( .I(n29975), .ZN(n29976) );
  INHSV2 U35509 ( .I(n39250), .ZN(n37766) );
  INHSV2 U35510 ( .I(n39702), .ZN(n39403) );
  INHSV2 U35511 ( .I(n39733), .ZN(n47927) );
  INHSV2 U35512 ( .I(n47927), .ZN(n40309) );
  AOI21HSV2 U35513 ( .A1(n29978), .A2(n39241), .B(n40309), .ZN(n29979) );
  NAND2HSV2 U35514 ( .A1(n29980), .A2(n29981), .ZN(n29983) );
  CLKAND2HSV2 U35515 ( .A1(n39230), .A2(\pe5/ti_7t [5]), .Z(n30064) );
  INHSV2 U35516 ( .I(n30064), .ZN(n29984) );
  BUFHSV2 U35517 ( .I(n31116), .Z(n39995) );
  NOR2HSV4 U35518 ( .A1(n29985), .A2(n39995), .ZN(n29986) );
  BUFHSV2 U35519 ( .I(n30206), .Z(n39398) );
  CLKNHSV2 U35520 ( .I(n29994), .ZN(n29998) );
  INHSV2 U35521 ( .I(n29996), .ZN(n29997) );
  INHSV2 U35522 ( .I(n30682), .ZN(n30028) );
  INHSV2 U35523 ( .I(n30113), .ZN(n48787) );
  CLKNAND2HSV1 U35524 ( .A1(n29999), .A2(n48787), .ZN(n30001) );
  CLKNAND2HSV0 U35525 ( .A1(\pe5/got [26]), .A2(n30918), .ZN(n30000) );
  XOR2HSV0 U35526 ( .A1(n30001), .A2(n30000), .Z(n30004) );
  NAND2HSV2 U35527 ( .A1(n48029), .A2(\pe5/pvq [7]), .ZN(n30002) );
  NAND2HSV2 U35528 ( .A1(n30147), .A2(n30146), .ZN(n30006) );
  INHSV2 U35529 ( .I(n30358), .ZN(n30288) );
  XOR2HSV0 U35530 ( .A1(n30006), .A2(n30005), .Z(n30010) );
  CLKNAND2HSV1 U35531 ( .A1(n30165), .A2(n30037), .ZN(n30008) );
  CLKNAND2HSV0 U35532 ( .A1(n30155), .A2(\pe5/bq[26] ), .ZN(n30007) );
  XOR2HSV0 U35533 ( .A1(n30008), .A2(n30007), .Z(n30009) );
  XOR2HSV0 U35534 ( .A1(n30010), .A2(n30009), .Z(n30013) );
  INHSV1 U35535 ( .I(n30032), .ZN(n30230) );
  CLKNAND2HSV1 U35536 ( .A1(n59938), .A2(n30230), .ZN(n30011) );
  XOR2HSV0 U35537 ( .A1(n39889), .A2(n30011), .Z(n30012) );
  XNOR2HSV4 U35538 ( .A1(n30013), .A2(n30012), .ZN(n30015) );
  NAND2HSV2 U35539 ( .A1(n30017), .A2(n30016), .ZN(n30340) );
  INHSV2 U35540 ( .I(n30297), .ZN(n30513) );
  CLKNAND2HSV0 U35541 ( .A1(n30340), .A2(n30513), .ZN(n30018) );
  CLKXOR2HSV2 U35542 ( .A1(n30019), .A2(n30018), .Z(n30021) );
  CLKNAND2HSV1 U35543 ( .A1(n30020), .A2(n30021), .ZN(n30024) );
  INHSV2 U35544 ( .I(n30021), .ZN(n30022) );
  CLKNHSV2 U35545 ( .I(n45477), .ZN(n30887) );
  NAND2HSV2 U35546 ( .A1(n30783), .A2(n30046), .ZN(n30025) );
  XNOR2HSV4 U35547 ( .A1(n30026), .A2(n30025), .ZN(n30194) );
  OA21HSV1 U35548 ( .A1(n30064), .A2(n37645), .B(n52799), .Z(n30027) );
  XNOR2HSV4 U35549 ( .A1(n30194), .A2(n30181), .ZN(n30192) );
  INHSV2 U35550 ( .I(n30113), .ZN(n39449) );
  CLKNAND2HSV1 U35551 ( .A1(n39449), .A2(n30155), .ZN(n30031) );
  XOR2HSV0 U35552 ( .A1(n30031), .A2(n30030), .Z(n30045) );
  INHSV1 U35553 ( .I(n30032), .ZN(n30547) );
  INHSV4 U35554 ( .I(\pe5/aot [27]), .ZN(n48175) );
  INHSV2 U35555 ( .I(n48175), .ZN(n39801) );
  NAND2HSV2 U35556 ( .A1(n39801), .A2(n30033), .ZN(n30034) );
  CLKXOR2HSV2 U35557 ( .A1(n30034), .A2(\pe5/phq [6]), .Z(n30035) );
  XNOR2HSV4 U35558 ( .A1(n30036), .A2(n30035), .ZN(n30044) );
  INHSV2 U35559 ( .I(n30163), .ZN(n48816) );
  CLKNAND2HSV1 U35560 ( .A1(n48816), .A2(n30037), .ZN(n30038) );
  NOR2HSV2 U35561 ( .A1(n30431), .A2(n48040), .ZN(n30041) );
  INHSV2 U35562 ( .I(n30365), .ZN(n48817) );
  INHSV2 U35563 ( .I(n30116), .ZN(n45470) );
  NAND2HSV2 U35564 ( .A1(n48817), .A2(n45470), .ZN(n30040) );
  XOR2HSV0 U35565 ( .A1(n30041), .A2(n30040), .Z(n30042) );
  INHSV2 U35566 ( .I(n30048), .ZN(n39578) );
  CLKNAND2HSV1 U35567 ( .A1(n30130), .A2(n39578), .ZN(n30049) );
  XNOR2HSV4 U35568 ( .A1(n30050), .A2(n30049), .ZN(n30067) );
  CLKNHSV2 U35569 ( .I(n30067), .ZN(n30052) );
  BUFHSV2 U35570 ( .I(n30206), .Z(n39405) );
  INHSV2 U35571 ( .I(n30051), .ZN(n59507) );
  OAI21HSV2 U35572 ( .A1(n39405), .A2(\pe5/ti_7t [6]), .B(n59507), .ZN(n30188)
         );
  OR2HSV1 U35573 ( .A1(n30188), .A2(n30204), .Z(n30090) );
  NAND3HSV3 U35574 ( .A1(n30060), .A2(n30067), .A3(n39705), .ZN(n30193) );
  NAND2HSV2 U35575 ( .A1(n30053), .A2(n30193), .ZN(n30054) );
  NOR2HSV4 U35576 ( .A1(n30192), .A2(n30054), .ZN(n30059) );
  NOR2HSV4 U35577 ( .A1(n30184), .A2(n37638), .ZN(n30182) );
  NOR2HSV2 U35578 ( .A1(n37645), .A2(\pe5/ti_7t [7]), .ZN(n30183) );
  INHSV2 U35579 ( .I(n30183), .ZN(n30055) );
  NAND2HSV2 U35580 ( .A1(n30055), .A2(n30322), .ZN(n30056) );
  CLKNHSV1 U35581 ( .I(n30196), .ZN(n30583) );
  MOAI22HSV4 U35582 ( .A1(n30182), .A2(n30056), .B1(n30193), .B2(n39382), .ZN(
        n30057) );
  INHSV4 U35583 ( .I(n30057), .ZN(n30058) );
  NOR2HSV4 U35584 ( .A1(n30059), .A2(n30058), .ZN(n30077) );
  BUFHSV2 U35585 ( .I(n30667), .Z(n31086) );
  BUFHSV8 U35586 ( .I(n39121), .Z(n47269) );
  NOR2HSV2 U35587 ( .A1(n30067), .A2(n30204), .ZN(n30061) );
  CLKNAND2HSV4 U35588 ( .A1(n47269), .A2(n30061), .ZN(n30190) );
  BUFHSV2 U35589 ( .I(n47927), .Z(n31240) );
  CLKNAND2HSV1 U35590 ( .A1(n30064), .A2(n31240), .ZN(n30065) );
  INHSV2 U35591 ( .I(\pe5/ti_7t [6]), .ZN(n30069) );
  NOR2HSV2 U35592 ( .A1(n30318), .A2(n30069), .ZN(n30207) );
  CLKAND2HSV4 U35593 ( .A1(n30071), .A2(n39366), .Z(n30072) );
  BUFHSV2 U35594 ( .I(n30667), .Z(n40012) );
  CLKAND2HSV2 U35595 ( .A1(n30253), .A2(n40012), .Z(n30073) );
  NOR2HSV2 U35596 ( .A1(n39578), .A2(n30874), .ZN(n30083) );
  INHSV2 U35597 ( .I(n30076), .ZN(n30082) );
  INHSV2 U35598 ( .I(n30078), .ZN(n30079) );
  NOR2HSV4 U35599 ( .A1(n30080), .A2(n30079), .ZN(n30087) );
  INHSV2 U35600 ( .I(n30087), .ZN(n30081) );
  INHSV2 U35601 ( .I(n30083), .ZN(n30084) );
  NOR2HSV4 U35602 ( .A1(n30085), .A2(n30084), .ZN(n30086) );
  CLKNAND2HSV3 U35603 ( .A1(n30087), .A2(n30086), .ZN(n30137) );
  NAND2HSV2 U35604 ( .A1(n39245), .A2(\pe5/ti_7t [8]), .ZN(n30088) );
  BUFHSV2 U35605 ( .I(n30192), .Z(n52732) );
  INHSV2 U35606 ( .I(n52732), .ZN(n30097) );
  CLKNHSV0 U35607 ( .I(n30193), .ZN(n30091) );
  NOR2HSV2 U35608 ( .A1(n30091), .A2(n30090), .ZN(n30191) );
  NAND2HSV2 U35609 ( .A1(n30191), .A2(n30190), .ZN(n30298) );
  CLKNHSV0 U35610 ( .I(n30188), .ZN(n30092) );
  NAND2HSV0 U35611 ( .A1(n30193), .A2(n30092), .ZN(n30093) );
  NOR2HSV2 U35612 ( .A1(n30192), .A2(n39245), .ZN(n30095) );
  NAND2HSV2 U35613 ( .A1(\pe5/ti_7t [7]), .A2(n39230), .ZN(n30300) );
  INHSV2 U35614 ( .I(n30300), .ZN(n30094) );
  OAI21HSV4 U35615 ( .A1(n30097), .A2(n30298), .B(n30096), .ZN(n30485) );
  BUFHSV2 U35616 ( .I(n30098), .Z(n39249) );
  INHSV2 U35617 ( .I(n39121), .ZN(n30441) );
  NAND2HSV2 U35618 ( .A1(n30515), .A2(n59947), .ZN(n30134) );
  CLKNAND2HSV0 U35619 ( .A1(n59937), .A2(n30341), .ZN(n30214) );
  CLKNHSV2 U35620 ( .I(n30100), .ZN(n44335) );
  NAND2HSV2 U35621 ( .A1(n44335), .A2(\pe5/pvq [10]), .ZN(n30101) );
  XNOR2HSV1 U35622 ( .A1(n30101), .A2(\pe5/phq [10]), .ZN(n30105) );
  INHSV2 U35623 ( .I(\pe5/aot [23]), .ZN(n40043) );
  CLKNAND2HSV1 U35624 ( .A1(\pe5/aot [23]), .A2(n30616), .ZN(n30103) );
  INHSV2 U35625 ( .I(n30150), .ZN(n59387) );
  NAND2HSV0 U35626 ( .A1(n59387), .A2(n30367), .ZN(n30102) );
  XOR2HSV0 U35627 ( .A1(n30103), .A2(n30102), .Z(n30104) );
  XOR3HSV2 U35628 ( .A1(n30214), .A2(n30105), .A3(n30104), .Z(n30125) );
  NAND2HSV2 U35629 ( .A1(n30377), .A2(n59637), .ZN(n30124) );
  CLKNAND2HSV0 U35630 ( .A1(n47200), .A2(n48752), .ZN(n30108) );
  INHSV2 U35631 ( .I(n44704), .ZN(n30799) );
  NAND2HSV0 U35632 ( .A1(n30799), .A2(n48785), .ZN(n30107) );
  XOR2HSV0 U35633 ( .A1(n30108), .A2(n30107), .Z(n30112) );
  INHSV2 U35634 ( .I(n31044), .ZN(n30538) );
  INHSV2 U35635 ( .I(n37564), .ZN(n30825) );
  NAND2HSV2 U35636 ( .A1(n30538), .A2(n30825), .ZN(n30110) );
  INHSV1 U35637 ( .I(n30163), .ZN(n30529) );
  NAND2HSV0 U35638 ( .A1(n30529), .A2(n30222), .ZN(n30109) );
  XOR2HSV0 U35639 ( .A1(n30110), .A2(n30109), .Z(n30111) );
  XOR2HSV0 U35640 ( .A1(n30112), .A2(n30111), .Z(n30122) );
  INHSV2 U35641 ( .I(n48219), .ZN(n30257) );
  CLKNAND2HSV0 U35642 ( .A1(n30257), .A2(n30230), .ZN(n30115) );
  INHSV2 U35643 ( .I(n30113), .ZN(n30256) );
  NAND2HSV0 U35644 ( .A1(n30165), .A2(n30256), .ZN(n30114) );
  XOR2HSV0 U35645 ( .A1(n30115), .A2(n30114), .Z(n30120) );
  INHSV2 U35646 ( .I(n30116), .ZN(n30357) );
  CLKNAND2HSV0 U35647 ( .A1(n30288), .A2(n30357), .ZN(n30118) );
  NAND2HSV0 U35648 ( .A1(n39122), .A2(n52585), .ZN(n30117) );
  XOR2HSV0 U35649 ( .A1(n30118), .A2(n30117), .Z(n30119) );
  XOR2HSV0 U35650 ( .A1(n30120), .A2(n30119), .Z(n30121) );
  XOR2HSV0 U35651 ( .A1(n30122), .A2(n30121), .Z(n30123) );
  XOR3HSV2 U35652 ( .A1(n30125), .A2(n30124), .A3(n30123), .Z(n30127) );
  BUFHSV2 U35653 ( .I(n30340), .Z(n30270) );
  CLKNAND2HSV1 U35654 ( .A1(n30270), .A2(n37630), .ZN(n30126) );
  XNOR2HSV1 U35655 ( .A1(n30127), .A2(n30126), .ZN(n30129) );
  CLKNAND2HSV1 U35656 ( .A1(n40187), .A2(n30685), .ZN(n30128) );
  XNOR2HSV1 U35657 ( .A1(n30129), .A2(n30128), .ZN(n30132) );
  NAND2HSV0 U35658 ( .A1(n30130), .A2(n30254), .ZN(n30131) );
  XNOR2HSV1 U35659 ( .A1(n30132), .A2(n30131), .ZN(n30133) );
  XNOR2HSV1 U35660 ( .A1(n30134), .A2(n30133), .ZN(n30135) );
  NOR2HSV2 U35661 ( .A1(n59507), .A2(n30874), .ZN(n31133) );
  INHSV2 U35662 ( .I(n31133), .ZN(n39222) );
  CLKAND2HSV2 U35663 ( .A1(n30143), .A2(n30142), .Z(n30180) );
  CLKNAND2HSV1 U35664 ( .A1(n30255), .A2(n59947), .ZN(n30178) );
  AND2HSV1 U35665 ( .A1(n37608), .A2(n30685), .Z(n30144) );
  XNOR2HSV4 U35666 ( .A1(n30145), .A2(n30144), .ZN(n30176) );
  CLKNAND2HSV1 U35667 ( .A1(n30799), .A2(n30146), .ZN(n30149) );
  CLKNAND2HSV0 U35668 ( .A1(n30147), .A2(n30367), .ZN(n30148) );
  XOR2HSV0 U35669 ( .A1(n30149), .A2(n30148), .Z(n30154) );
  INHSV2 U35670 ( .I(n45900), .ZN(n45500) );
  CLKNAND2HSV1 U35671 ( .A1(n45500), .A2(n48752), .ZN(n30152) );
  INHSV2 U35672 ( .I(n30150), .ZN(n30543) );
  CLKNAND2HSV0 U35673 ( .A1(n30543), .A2(n48785), .ZN(n30151) );
  XOR2HSV0 U35674 ( .A1(n30152), .A2(n30151), .Z(n30153) );
  XOR2HSV0 U35675 ( .A1(n30154), .A2(n30153), .Z(n30162) );
  CLKNAND2HSV0 U35676 ( .A1(n30155), .A2(\pe5/bq[24] ), .ZN(n30157) );
  INHSV2 U35677 ( .I(n30287), .ZN(n46622) );
  CLKNAND2HSV0 U35678 ( .A1(n59937), .A2(n46622), .ZN(n30156) );
  XOR2HSV0 U35679 ( .A1(n30157), .A2(n30156), .Z(n30160) );
  NAND2HSV2 U35680 ( .A1(n48034), .A2(\pe5/pvq [9]), .ZN(n30158) );
  XOR2HSV0 U35681 ( .A1(n30158), .A2(\pe5/phq [9]), .Z(n30159) );
  XOR2HSV0 U35682 ( .A1(n30160), .A2(n30159), .Z(n30161) );
  XOR2HSV0 U35683 ( .A1(n30162), .A2(n30161), .Z(n30172) );
  NOR2HSV1 U35684 ( .A1(n30163), .A2(n30113), .ZN(n30167) );
  NAND2HSV0 U35685 ( .A1(n30165), .A2(n30164), .ZN(n30166) );
  XOR2HSV0 U35686 ( .A1(n30167), .A2(n30166), .Z(n30170) );
  NAND2HSV2 U35687 ( .A1(n59939), .A2(n30230), .ZN(n37665) );
  XOR2HSV0 U35688 ( .A1(n37665), .A2(n30168), .Z(n30169) );
  XNOR2HSV1 U35689 ( .A1(n30170), .A2(n30169), .ZN(n30171) );
  XNOR2HSV1 U35690 ( .A1(n30172), .A2(n30171), .ZN(n30174) );
  INHSV2 U35691 ( .I(n30210), .ZN(n48739) );
  CLKNAND2HSV0 U35692 ( .A1(n59393), .A2(n48739), .ZN(n30173) );
  XNOR2HSV1 U35693 ( .A1(n30174), .A2(n30173), .ZN(n30175) );
  XNOR2HSV4 U35694 ( .A1(n30176), .A2(n30175), .ZN(n30177) );
  XNOR2HSV4 U35695 ( .A1(n30178), .A2(n30177), .ZN(n30179) );
  INHSV2 U35696 ( .I(n39249), .ZN(n40142) );
  CLKNHSV0 U35697 ( .I(n30181), .ZN(n30187) );
  NOR2HSV1 U35698 ( .A1(n30183), .A2(n25344), .ZN(n30186) );
  NAND3HSV1 U35699 ( .A1(n30187), .A2(n30184), .A3(n39398), .ZN(n30185) );
  NOR2HSV1 U35700 ( .A1(n39704), .A2(n30188), .ZN(n30189) );
  NAND2HSV2 U35701 ( .A1(n30190), .A2(n30189), .ZN(n30195) );
  NAND2HSV2 U35702 ( .A1(n30874), .A2(\pe5/ti_7t [9]), .ZN(n30327) );
  INHSV2 U35703 ( .I(n30327), .ZN(n30198) );
  CLKNHSV0 U35704 ( .I(\pe5/ti_7t [10]), .ZN(n30201) );
  AOI21HSV2 U35705 ( .A1(n30201), .A2(n31101), .B(n40309), .ZN(n30396) );
  INHSV2 U35706 ( .I(n30075), .ZN(n37554) );
  NOR2HSV2 U35707 ( .A1(n25852), .A2(n39995), .ZN(n30250) );
  CLKBUFHSV4 U35708 ( .I(n30485), .Z(n37724) );
  CLKNAND2HSV3 U35709 ( .A1(n37724), .A2(n30046), .ZN(n30248) );
  NOR2HSV0 U35710 ( .A1(n60074), .A2(n30207), .ZN(n30205) );
  NOR2HSV0 U35711 ( .A1(n30297), .A2(n30204), .ZN(n30299) );
  BUFHSV2 U35712 ( .I(n30206), .Z(n39705) );
  OAI21HSV0 U35713 ( .A1(n30207), .A2(n39705), .B(n59947), .ZN(n30209) );
  AND2HSV2 U35714 ( .A1(n30207), .A2(n59947), .Z(n30208) );
  NAND2HSV0 U35715 ( .A1(n30255), .A2(\pe5/got [26]), .ZN(n30244) );
  CLKNAND2HSV1 U35716 ( .A1(n30270), .A2(n37631), .ZN(n30242) );
  NAND2HSV2 U35717 ( .A1(n39466), .A2(n37630), .ZN(n30241) );
  BUFHSV2 U35718 ( .I(n48049), .Z(n37707) );
  NAND2HSV2 U35719 ( .A1(n37707), .A2(\pe5/pvq [11]), .ZN(n30211) );
  XOR2HSV0 U35720 ( .A1(n30211), .A2(\pe5/phq [11]), .Z(n30216) );
  BUFHSV2 U35721 ( .I(n30212), .Z(n40236) );
  INHSV2 U35722 ( .I(n40236), .ZN(n30519) );
  INHSV2 U35723 ( .I(n37564), .ZN(n30607) );
  NAND2HSV2 U35724 ( .A1(n30519), .A2(n30607), .ZN(n30265) );
  INHSV2 U35725 ( .I(n37564), .ZN(n47305) );
  IOA22HSV1 U35726 ( .B1(n40236), .B2(n30452), .A1(n59937), .A2(n47305), .ZN(
        n30213) );
  OAI21HSV1 U35727 ( .A1(n30214), .A2(n30265), .B(n30213), .ZN(n30215) );
  XNOR2HSV1 U35728 ( .A1(n30216), .A2(n30215), .ZN(n30219) );
  CLKNAND2HSV1 U35729 ( .A1(n30288), .A2(n30256), .ZN(n48177) );
  CLKNAND2HSV1 U35730 ( .A1(n30257), .A2(n30357), .ZN(n30217) );
  XOR2HSV0 U35731 ( .A1(n48177), .A2(n30217), .Z(n30218) );
  XNOR2HSV1 U35732 ( .A1(n30219), .A2(n30218), .ZN(n30239) );
  NAND2HSV2 U35733 ( .A1(n30377), .A2(n47200), .ZN(n30238) );
  INHSV2 U35734 ( .I(n45451), .ZN(n30701) );
  CLKNAND2HSV0 U35735 ( .A1(n30701), .A2(n30616), .ZN(n30221) );
  NAND2HSV0 U35736 ( .A1(n30799), .A2(n30367), .ZN(n30220) );
  XOR2HSV0 U35737 ( .A1(n30221), .A2(n30220), .Z(n30227) );
  CLKNAND2HSV0 U35738 ( .A1(n31048), .A2(n30222), .ZN(n30225) );
  INHSV2 U35739 ( .I(n30223), .ZN(n30344) );
  CLKNAND2HSV0 U35740 ( .A1(\pe5/aot [23]), .A2(n30344), .ZN(n30224) );
  XOR2HSV0 U35741 ( .A1(n30225), .A2(n30224), .Z(n30226) );
  XOR2HSV0 U35742 ( .A1(n30227), .A2(n30226), .Z(n30236) );
  BUFHSV2 U35743 ( .I(n30163), .Z(n37595) );
  NOR2HSV2 U35744 ( .A1(n37595), .A2(n30287), .ZN(n30229) );
  CLKNAND2HSV1 U35745 ( .A1(n48744), .A2(n30693), .ZN(n30228) );
  XOR2HSV0 U35746 ( .A1(n30229), .A2(n30228), .Z(n30234) );
  NAND2HSV0 U35747 ( .A1(n59387), .A2(n30230), .ZN(n30232) );
  INHSV2 U35748 ( .I(n45844), .ZN(n30798) );
  CLKNAND2HSV1 U35749 ( .A1(n30538), .A2(n30798), .ZN(n30231) );
  XOR2HSV0 U35750 ( .A1(n30232), .A2(n30231), .Z(n30233) );
  XOR2HSV0 U35751 ( .A1(n30234), .A2(n30233), .Z(n30235) );
  XOR2HSV0 U35752 ( .A1(n30236), .A2(n30235), .Z(n30237) );
  XOR3HSV2 U35753 ( .A1(n30239), .A2(n30238), .A3(n30237), .Z(n30240) );
  XOR3HSV2 U35754 ( .A1(n30242), .A2(n30241), .A3(n30240), .Z(n30243) );
  XNOR2HSV1 U35755 ( .A1(n30244), .A2(n30243), .ZN(n30245) );
  XNOR2HSV1 U35756 ( .A1(n30246), .A2(n30245), .ZN(n30247) );
  XNOR2HSV4 U35757 ( .A1(n30248), .A2(n30247), .ZN(n30249) );
  NAND2HSV4 U35758 ( .A1(n30568), .A2(n30251), .ZN(n30422) );
  CLKNAND2HSV4 U35759 ( .A1(n30423), .A2(n30422), .ZN(n30428) );
  INHSV2 U35760 ( .I(n30428), .ZN(n30316) );
  CLKNHSV0 U35761 ( .I(n25862), .ZN(n30684) );
  BUFHSV4 U35762 ( .I(n30253), .Z(n31065) );
  INHSV4 U35763 ( .I(n31065), .ZN(n39824) );
  NAND2HSV2 U35764 ( .A1(n39583), .A2(n48739), .ZN(n30276) );
  INHSV2 U35765 ( .I(n47140), .ZN(n39532) );
  CLKNAND2HSV1 U35766 ( .A1(n30377), .A2(n39532), .ZN(n30269) );
  CLKNAND2HSV1 U35767 ( .A1(n30257), .A2(n30256), .ZN(n30259) );
  INHSV2 U35768 ( .I(n30516), .ZN(n30782) );
  CLKNAND2HSV1 U35769 ( .A1(n30782), .A2(n30693), .ZN(n30258) );
  XOR2HSV0 U35770 ( .A1(n30259), .A2(n30258), .Z(n30263) );
  INHSV2 U35771 ( .I(n45460), .ZN(n30366) );
  CLKNAND2HSV0 U35772 ( .A1(n30543), .A2(n30366), .ZN(n30931) );
  OAI22HSV0 U35773 ( .A1(n31044), .A2(n45460), .B1(n30150), .B2(n30116), .ZN(
        n30260) );
  OAI21HSV0 U35774 ( .A1(n30931), .A2(n30261), .B(n30260), .ZN(n30262) );
  XNOR2HSV1 U35775 ( .A1(n30263), .A2(n30262), .ZN(n30267) );
  NAND2HSV0 U35776 ( .A1(n48243), .A2(n30547), .ZN(n30264) );
  XOR2HSV0 U35777 ( .A1(n30265), .A2(n30264), .Z(n30266) );
  XNOR2HSV1 U35778 ( .A1(n30267), .A2(n30266), .ZN(n30268) );
  XNOR2HSV1 U35779 ( .A1(n30269), .A2(n30268), .ZN(n30272) );
  CLKNAND2HSV0 U35780 ( .A1(n30270), .A2(n47200), .ZN(n30271) );
  XNOR2HSV1 U35781 ( .A1(n30272), .A2(n30271), .ZN(n30274) );
  CLKNAND2HSV1 U35782 ( .A1(n30783), .A2(n59637), .ZN(n30273) );
  XNOR2HSV1 U35783 ( .A1(n30274), .A2(n30273), .ZN(n30275) );
  XNOR2HSV4 U35784 ( .A1(n30276), .A2(n30275), .ZN(n30278) );
  INHSV2 U35785 ( .I(n30278), .ZN(n30277) );
  NOR2HSV2 U35786 ( .A1(n30277), .A2(n31081), .ZN(n30280) );
  CLKBUFHSV4 U35787 ( .I(n47269), .Z(n59936) );
  AOI21HSV2 U35788 ( .A1(n59936), .A2(n30685), .B(n30278), .ZN(n30279) );
  CLKNAND2HSV1 U35789 ( .A1(\pe5/aot [23]), .A2(n30367), .ZN(n30282) );
  NAND2HSV2 U35790 ( .A1(n30701), .A2(n30344), .ZN(n30281) );
  XOR2HSV0 U35791 ( .A1(n30282), .A2(n30281), .Z(n30295) );
  NAND2HSV2 U35792 ( .A1(n48034), .A2(\pe5/pvq [12]), .ZN(n30283) );
  XNOR2HSV1 U35793 ( .A1(n30283), .A2(\pe5/phq [12]), .ZN(n30284) );
  NAND2HSV2 U35794 ( .A1(n30529), .A2(n30341), .ZN(n48665) );
  XNOR2HSV1 U35795 ( .A1(n30284), .A2(n48665), .ZN(n30294) );
  CLKNAND2HSV0 U35796 ( .A1(n59937), .A2(n30798), .ZN(n30286) );
  CLKNAND2HSV1 U35797 ( .A1(\pe5/aot [21]), .A2(n30616), .ZN(n30285) );
  XOR2HSV0 U35798 ( .A1(n30286), .A2(n30285), .Z(n30292) );
  NAND2HSV2 U35799 ( .A1(n31048), .A2(n30526), .ZN(n30290) );
  CLKNAND2HSV1 U35800 ( .A1(n30288), .A2(n30542), .ZN(n30289) );
  XOR2HSV0 U35801 ( .A1(n30290), .A2(n30289), .Z(n30291) );
  XOR2HSV0 U35802 ( .A1(n30292), .A2(n30291), .Z(n30293) );
  NOR2HSV1 U35803 ( .A1(n30298), .A2(n30297), .ZN(n30303) );
  NAND2HSV0 U35804 ( .A1(n52733), .A2(n30299), .ZN(n30301) );
  OAI22HSV0 U35805 ( .A1(n52732), .A2(n30301), .B1(n30297), .B2(n30300), .ZN(
        n30302) );
  OAI21HSV2 U35806 ( .A1(n30684), .A2(n31003), .B(n30311), .ZN(n30307) );
  INHSV4 U35807 ( .I(n25862), .ZN(n30440) );
  CLKNAND2HSV2 U35808 ( .A1(n30306), .A2(n30305), .ZN(n30313) );
  INHSV4 U35809 ( .I(n30308), .ZN(n30309) );
  NOR2HSV4 U35810 ( .A1(n30309), .A2(n40007), .ZN(n30310) );
  INHSV4 U35811 ( .I(n30310), .ZN(n30426) );
  INHSV4 U35812 ( .I(n30440), .ZN(n30514) );
  NAND2HSV2 U35813 ( .A1(n30514), .A2(n59395), .ZN(n30312) );
  CLKNAND2HSV4 U35814 ( .A1(n30314), .A2(n30313), .ZN(n30334) );
  CLKNAND2HSV3 U35815 ( .A1(n30334), .A2(n52834), .ZN(n30319) );
  CLKNAND2HSV1 U35816 ( .A1(n30316), .A2(n30315), .ZN(n30324) );
  INHSV2 U35817 ( .I(\pe5/ti_7t [12]), .ZN(n30317) );
  NOR2HSV1 U35818 ( .A1(n30318), .A2(n30317), .ZN(n30653) );
  INHSV4 U35819 ( .I(n30319), .ZN(n30427) );
  BUFHSV2 U35820 ( .I(n47927), .Z(n52834) );
  NOR2HSV4 U35821 ( .A1(n30427), .A2(n29645), .ZN(n30321) );
  CLKNAND2HSV1 U35822 ( .A1(n30324), .A2(n30323), .ZN(n30333) );
  CLKNHSV0 U35823 ( .I(n30325), .ZN(n30326) );
  INHSV2 U35824 ( .I(n30326), .ZN(n30329) );
  INHSV2 U35825 ( .I(n40162), .ZN(n30330) );
  CLKAND2HSV2 U35826 ( .A1(n40162), .A2(\pe5/ti_7t [10]), .Z(n30331) );
  INHSV1 U35827 ( .I(n30653), .ZN(n30509) );
  NAND3HSV2 U35828 ( .A1(n25854), .A2(n59946), .A3(n30509), .ZN(n30332) );
  CLKNAND2HSV2 U35829 ( .A1(n30333), .A2(n30332), .ZN(n30338) );
  NAND2HSV4 U35830 ( .A1(n30423), .A2(n30422), .ZN(n59426) );
  NOR2HSV4 U35831 ( .A1(n59426), .A2(n52754), .ZN(n30506) );
  INHSV2 U35832 ( .I(n30506), .ZN(n30336) );
  CLKNAND2HSV4 U35833 ( .A1(n59426), .A2(n29656), .ZN(n30505) );
  AOI21HSV2 U35834 ( .A1(n30334), .A2(n39733), .B(n30755), .ZN(n30504) );
  CLKAND2HSV4 U35835 ( .A1(n29634), .A2(n30504), .Z(n30335) );
  NAND3HSV4 U35836 ( .A1(n30336), .A2(n30505), .A3(n30335), .ZN(n30337) );
  NAND2HSV2 U35837 ( .A1(n30514), .A2(n30142), .ZN(n30393) );
  INAND2HSV4 U35838 ( .A1(n30339), .B1(n29663), .ZN(n30885) );
  NAND2HSV2 U35839 ( .A1(n30885), .A2(n30513), .ZN(n30391) );
  CLKNAND2HSV0 U35840 ( .A1(n30515), .A2(n37630), .ZN(n30386) );
  NAND2HSV2 U35841 ( .A1(n31151), .A2(n59637), .ZN(n30384) );
  BUFHSV2 U35842 ( .I(n30340), .Z(n37608) );
  BUFHSV2 U35843 ( .I(n37608), .Z(n30785) );
  CLKNAND2HSV1 U35844 ( .A1(n30785), .A2(n47267), .ZN(n30382) );
  CLKNAND2HSV1 U35845 ( .A1(n30783), .A2(n59948), .ZN(n30381) );
  NAND2HSV0 U35846 ( .A1(n39266), .A2(n30341), .ZN(n30343) );
  NAND2HSV0 U35847 ( .A1(\pe5/aot [23]), .A2(n30547), .ZN(n30342) );
  XOR2HSV0 U35848 ( .A1(n30343), .A2(n30342), .Z(n30348) );
  NAND2HSV0 U35849 ( .A1(n30529), .A2(n30607), .ZN(n30346) );
  NAND2HSV0 U35850 ( .A1(\pe5/aot [21]), .A2(n30344), .ZN(n30345) );
  XOR2HSV0 U35851 ( .A1(n30346), .A2(n30345), .Z(n30347) );
  XOR2HSV0 U35852 ( .A1(n30348), .A2(n30347), .Z(n30356) );
  CLKNAND2HSV0 U35853 ( .A1(n30543), .A2(n47234), .ZN(n30350) );
  NAND2HSV0 U35854 ( .A1(\pe5/got [20]), .A2(n30693), .ZN(n30349) );
  XOR2HSV0 U35855 ( .A1(n30350), .A2(n30349), .Z(n30354) );
  NAND2HSV0 U35856 ( .A1(\pe5/aot [20]), .A2(n30616), .ZN(n30352) );
  NAND2HSV0 U35857 ( .A1(n48796), .A2(n30542), .ZN(n30351) );
  XOR2HSV0 U35858 ( .A1(n30352), .A2(n30351), .Z(n30353) );
  XOR2HSV0 U35859 ( .A1(n30354), .A2(n30353), .Z(n30355) );
  XOR2HSV0 U35860 ( .A1(n30356), .A2(n30355), .Z(n30376) );
  NAND2HSV0 U35861 ( .A1(n59940), .A2(n30357), .ZN(n30360) );
  CLKNHSV0 U35862 ( .I(n30358), .ZN(n30702) );
  NAND2HSV0 U35863 ( .A1(n30702), .A2(n30526), .ZN(n30359) );
  XOR2HSV0 U35864 ( .A1(n30360), .A2(n30359), .Z(n30364) );
  NAND2HSV0 U35865 ( .A1(n30519), .A2(n30798), .ZN(n30362) );
  INHSV2 U35866 ( .I(n45426), .ZN(n51048) );
  CLKNAND2HSV0 U35867 ( .A1(n30538), .A2(n51048), .ZN(n30361) );
  XOR2HSV0 U35868 ( .A1(n30362), .A2(n30361), .Z(n30363) );
  XOR2HSV0 U35869 ( .A1(n30364), .A2(n30363), .Z(n30374) );
  INHSV2 U35870 ( .I(n39779), .ZN(n39601) );
  NAND2HSV2 U35871 ( .A1(n39601), .A2(n30366), .ZN(n30369) );
  NAND2HSV0 U35872 ( .A1(n30701), .A2(n30367), .ZN(n30368) );
  XOR2HSV0 U35873 ( .A1(n30369), .A2(n30368), .Z(n30372) );
  NAND2HSV0 U35874 ( .A1(n46628), .A2(\pe5/pvq [13]), .ZN(n30370) );
  XOR2HSV0 U35875 ( .A1(n30370), .A2(\pe5/phq [13]), .Z(n30371) );
  XOR2HSV0 U35876 ( .A1(n30372), .A2(n30371), .Z(n30373) );
  XOR2HSV0 U35877 ( .A1(n30374), .A2(n30373), .Z(n30375) );
  XOR2HSV0 U35878 ( .A1(n30376), .A2(n30375), .Z(n30379) );
  INHSV2 U35879 ( .I(n30516), .ZN(n31149) );
  CLKNAND2HSV0 U35880 ( .A1(n30377), .A2(n31149), .ZN(n30378) );
  XNOR2HSV1 U35881 ( .A1(n30379), .A2(n30378), .ZN(n30380) );
  XOR3HSV2 U35882 ( .A1(n30382), .A2(n30381), .A3(n30380), .Z(n30383) );
  XNOR2HSV1 U35883 ( .A1(n30384), .A2(n30383), .ZN(n30385) );
  XNOR2HSV1 U35884 ( .A1(n30386), .A2(n30385), .ZN(n30389) );
  NAND2HSV2 U35885 ( .A1(n39824), .A2(n48742), .ZN(n30388) );
  INHSV1 U35886 ( .I(n30431), .ZN(n30596) );
  NAND2HSV2 U35887 ( .A1(n37724), .A2(n30596), .ZN(n30387) );
  XOR3HSV2 U35888 ( .A1(n30389), .A2(n30388), .A3(n30387), .Z(n30390) );
  XNOR2HSV1 U35889 ( .A1(n30391), .A2(n30390), .ZN(n30392) );
  XNOR2HSV4 U35890 ( .A1(n30395), .A2(n30394), .ZN(n30411) );
  CLKNAND2HSV2 U35891 ( .A1(n30397), .A2(n30396), .ZN(n30432) );
  NOR2HSV0 U35892 ( .A1(n30404), .A2(n39246), .ZN(n30400) );
  NAND2HSV0 U35893 ( .A1(n30405), .A2(n30404), .ZN(n30398) );
  CLKNHSV2 U35894 ( .I(n30398), .ZN(n30399) );
  CLKNHSV0 U35895 ( .I(n30404), .ZN(n30401) );
  BUFHSV2 U35896 ( .I(n44520), .Z(n40305) );
  CLKNAND2HSV3 U35897 ( .A1(n30402), .A2(n40305), .ZN(n30435) );
  NAND2HSV0 U35898 ( .A1(n30440), .A2(n30404), .ZN(n30403) );
  MUX2NHSV1 U35899 ( .I0(n30405), .I1(n39578), .S(n30404), .ZN(n30406) );
  INHSV2 U35900 ( .I(n30406), .ZN(n30436) );
  NAND2HSV2 U35901 ( .A1(n39245), .A2(\pe5/ti_7t [11]), .ZN(n30572) );
  OR2HSV1 U35902 ( .A1(n30572), .A2(n30075), .Z(n30407) );
  OAI21HSV2 U35903 ( .A1(n30408), .A2(n30432), .B(n30407), .ZN(n30409) );
  AOI21HSV2 U35904 ( .A1(n30432), .A2(n30410), .B(n30409), .ZN(n30412) );
  NAND2HSV2 U35905 ( .A1(n30411), .A2(n30412), .ZN(n30416) );
  INHSV2 U35906 ( .I(n30411), .ZN(n30414) );
  INHSV2 U35907 ( .I(n30412), .ZN(n30413) );
  NAND2HSV2 U35908 ( .A1(n30414), .A2(n30413), .ZN(n30415) );
  NAND2HSV4 U35909 ( .A1(n30416), .A2(n30415), .ZN(n30662) );
  XNOR2HSV4 U35910 ( .A1(n30661), .A2(n30662), .ZN(n60041) );
  CLKNAND2HSV2 U35911 ( .A1(n60041), .A2(n30864), .ZN(n30418) );
  NAND2HSV2 U35912 ( .A1(\pe5/ti_7t [13]), .A2(n39730), .ZN(n30417) );
  NAND2HSV4 U35913 ( .A1(n30418), .A2(n30417), .ZN(n30884) );
  INHSV2 U35914 ( .I(n30504), .ZN(n30419) );
  CLKNAND2HSV2 U35915 ( .A1(n30420), .A2(n30505), .ZN(n30657) );
  INHSV2 U35916 ( .I(n30423), .ZN(n30424) );
  INHSV4 U35917 ( .I(n30507), .ZN(n52753) );
  NOR2HSV2 U35918 ( .A1(n30508), .A2(n52753), .ZN(n30651) );
  AOI21HSV4 U35919 ( .A1(n30428), .A2(n30427), .B(n30426), .ZN(n30649) );
  OAI21HSV2 U35920 ( .A1(n30657), .A2(n30507), .B(n30429), .ZN(n30430) );
  INHSV3 U35921 ( .I(n30430), .ZN(n30496) );
  INHSV2 U35922 ( .I(n30432), .ZN(n30574) );
  INHSV4 U35923 ( .I(n30433), .ZN(n30434) );
  INAND2HSV4 U35924 ( .A1(n30435), .B1(n30434), .ZN(n30570) );
  NAND2HSV2 U35925 ( .A1(n29671), .A2(n30436), .ZN(n30573) );
  INHSV2 U35926 ( .I(n30573), .ZN(n30438) );
  INHSV2 U35927 ( .I(n30572), .ZN(n30437) );
  AOI21HSV4 U35928 ( .A1(n30574), .A2(n30438), .B(n30437), .ZN(n30439) );
  OAI21HSV4 U35929 ( .A1(n30574), .A2(n30570), .B(n30439), .ZN(n45800) );
  BUFHSV4 U35930 ( .I(n45800), .Z(n37657) );
  NAND2HSV2 U35931 ( .A1(n37657), .A2(n48742), .ZN(n30495) );
  NAND2HSV2 U35932 ( .A1(n39745), .A2(n37630), .ZN(n30494) );
  BUFHSV2 U35933 ( .I(n30440), .Z(n37555) );
  NAND2HSV2 U35934 ( .A1(n52578), .A2(n37631), .ZN(n30492) );
  BUFHSV2 U35935 ( .I(n30885), .Z(n59381) );
  CLKBUFHSV4 U35936 ( .I(n59381), .Z(n39882) );
  INHSV2 U35937 ( .I(n39743), .ZN(n30840) );
  CLKNAND2HSV1 U35938 ( .A1(n39882), .A2(n30840), .ZN(n30490) );
  NAND2HSV0 U35939 ( .A1(n37659), .A2(\pe5/got [20]), .ZN(n30484) );
  INHSV2 U35940 ( .I(n30686), .ZN(n30886) );
  NAND2HSV0 U35941 ( .A1(n31151), .A2(n30886), .ZN(n30482) );
  INHSV2 U35942 ( .I(\pe5/got [18]), .ZN(n30784) );
  INHSV2 U35943 ( .I(n30784), .ZN(n31150) );
  CLKNAND2HSV0 U35944 ( .A1(n30783), .A2(n31150), .ZN(n30443) );
  INHSV2 U35945 ( .I(n50422), .ZN(n37725) );
  NAND2HSV0 U35946 ( .A1(n30785), .A2(n37725), .ZN(n30442) );
  XNOR2HSV1 U35947 ( .A1(n30443), .A2(n30442), .ZN(n30480) );
  BUFHSV2 U35948 ( .I(\pe5/aot [21]), .Z(n59638) );
  CLKNHSV0 U35949 ( .I(n39772), .ZN(n40207) );
  NAND2HSV0 U35950 ( .A1(n59638), .A2(n40207), .ZN(n30445) );
  CLKNHSV0 U35951 ( .I(\pe5/bq[29] ), .ZN(n45461) );
  CLKNAND2HSV0 U35952 ( .A1(\pe5/aot [18]), .A2(n39130), .ZN(n30444) );
  XOR2HSV0 U35953 ( .A1(n30445), .A2(n30444), .Z(n30449) );
  INHSV2 U35954 ( .I(n31029), .ZN(n39446) );
  CLKNAND2HSV0 U35955 ( .A1(n39446), .A2(n48802), .ZN(n30447) );
  NAND2HSV0 U35956 ( .A1(n30788), .A2(n47234), .ZN(n30446) );
  XOR2HSV0 U35957 ( .A1(n30447), .A2(n30446), .Z(n30448) );
  XOR2HSV0 U35958 ( .A1(n30449), .A2(n30448), .Z(n30457) );
  INHSV2 U35959 ( .I(n48822), .ZN(n30900) );
  CLKNAND2HSV0 U35960 ( .A1(n30529), .A2(n30900), .ZN(n30451) );
  INHSV2 U35961 ( .I(n45460), .ZN(n31190) );
  NAND2HSV0 U35962 ( .A1(n59879), .A2(n31190), .ZN(n30450) );
  XOR2HSV0 U35963 ( .A1(n30451), .A2(n30450), .Z(n30455) );
  INHSV1 U35964 ( .I(n30365), .ZN(n31039) );
  CLKNAND2HSV1 U35965 ( .A1(n31039), .A2(n48181), .ZN(n30816) );
  CLKNAND2HSV0 U35966 ( .A1(\pe5/aot [23]), .A2(n30891), .ZN(n30453) );
  XOR2HSV0 U35967 ( .A1(n30816), .A2(n30453), .Z(n30454) );
  XOR2HSV0 U35968 ( .A1(n30455), .A2(n30454), .Z(n30456) );
  XOR2HSV0 U35969 ( .A1(n30457), .A2(n30456), .Z(n30460) );
  INHSV2 U35970 ( .I(n30888), .ZN(n39434) );
  NAND2HSV2 U35971 ( .A1(n30806), .A2(n39434), .ZN(n30459) );
  XNOR2HSV1 U35972 ( .A1(n30460), .A2(n30459), .ZN(n30478) );
  CLKNHSV0 U35973 ( .I(n40235), .ZN(n31048) );
  NAND2HSV2 U35974 ( .A1(n31048), .A2(n39454), .ZN(n31177) );
  CLKNHSV0 U35975 ( .I(n31044), .ZN(n39496) );
  CLKNAND2HSV0 U35976 ( .A1(n39496), .A2(n53314), .ZN(n39586) );
  XOR2HSV0 U35977 ( .A1(n31177), .A2(n39586), .Z(n30476) );
  NAND2HSV0 U35978 ( .A1(n30925), .A2(\pe5/pvq [18]), .ZN(n30461) );
  XOR2HSV0 U35979 ( .A1(n30461), .A2(\pe5/phq [18]), .Z(n30464) );
  CLKNHSV0 U35980 ( .I(n29892), .ZN(n48198) );
  CLKNAND2HSV1 U35981 ( .A1(n59640), .A2(n48198), .ZN(n30930) );
  INHSV2 U35982 ( .I(n50518), .ZN(n39616) );
  NAND2HSV2 U35983 ( .A1(n39616), .A2(n30698), .ZN(n30824) );
  NAND2HSV0 U35984 ( .A1(n59640), .A2(n30698), .ZN(n48182) );
  OAI21HSV0 U35985 ( .A1(n50518), .A2(n29892), .B(n48182), .ZN(n30462) );
  OAI21HSV1 U35986 ( .A1(n30930), .A2(n30824), .B(n30462), .ZN(n30463) );
  XOR2HSV0 U35987 ( .A1(n30464), .A2(n30463), .Z(n30475) );
  CLKNHSV0 U35988 ( .I(n48175), .ZN(n31161) );
  INHSV1 U35989 ( .I(n45821), .ZN(n51041) );
  CLKNAND2HSV1 U35990 ( .A1(n31161), .A2(n51041), .ZN(n31040) );
  INHSV2 U35991 ( .I(n45426), .ZN(n30911) );
  NAND2HSV0 U35992 ( .A1(n30519), .A2(n30911), .ZN(n30622) );
  OAI22HSV0 U35993 ( .A1(n39123), .A2(n45821), .B1(n48175), .B2(n45426), .ZN(
        n30465) );
  OAI21HSV0 U35994 ( .A1(n31040), .A2(n30622), .B(n30465), .ZN(n30466) );
  CLKNHSV0 U35995 ( .I(n45844), .ZN(n31178) );
  NAND2HSV0 U35996 ( .A1(n59387), .A2(n31178), .ZN(n31032) );
  XNOR2HSV1 U35997 ( .A1(n30466), .A2(n31032), .ZN(n30474) );
  NOR2HSV0 U35998 ( .A1(n45451), .A2(n30287), .ZN(n30468) );
  NAND2HSV0 U35999 ( .A1(\pe5/aot [15]), .A2(n30789), .ZN(n30467) );
  XOR2HSV0 U36000 ( .A1(n30468), .A2(n30467), .Z(n30472) );
  NAND2HSV0 U36001 ( .A1(n30799), .A2(n30825), .ZN(n30470) );
  INHSV1 U36002 ( .I(n48722), .ZN(n31007) );
  CLKNAND2HSV0 U36003 ( .A1(n31007), .A2(n30918), .ZN(n30469) );
  XOR2HSV0 U36004 ( .A1(n30470), .A2(n30469), .Z(n30471) );
  XOR2HSV0 U36005 ( .A1(n30472), .A2(n30471), .Z(n30473) );
  XOR4HSV1 U36006 ( .A1(n30476), .A2(n30475), .A3(n30474), .A4(n30473), .Z(
        n30477) );
  XNOR2HSV1 U36007 ( .A1(n30478), .A2(n30477), .ZN(n30479) );
  XNOR2HSV1 U36008 ( .A1(n30480), .A2(n30479), .ZN(n30481) );
  XNOR2HSV1 U36009 ( .A1(n30482), .A2(n30481), .ZN(n30483) );
  XNOR2HSV1 U36010 ( .A1(n30484), .A2(n30483), .ZN(n30488) );
  CLKNHSV1 U36011 ( .I(n31065), .ZN(n30944) );
  CLKNAND2HSV1 U36012 ( .A1(n30944), .A2(n31149), .ZN(n30487) );
  CLKNAND2HSV1 U36013 ( .A1(n47058), .A2(n47267), .ZN(n30486) );
  XOR3HSV2 U36014 ( .A1(n30488), .A2(n30487), .A3(n30486), .Z(n30489) );
  XNOR2HSV1 U36015 ( .A1(n30490), .A2(n30489), .ZN(n30491) );
  XNOR2HSV1 U36016 ( .A1(n30492), .A2(n30491), .ZN(n30493) );
  XNOR2HSV4 U36017 ( .A1(n30495), .A2(n29672), .ZN(n30497) );
  AO21HSV0 U36018 ( .A1(n39744), .A2(n31225), .B(n30497), .Z(n30501) );
  INHSV4 U36019 ( .I(n30496), .ZN(n39120) );
  INAND2HSV2 U36020 ( .A1(n37635), .B1(n30497), .ZN(n30498) );
  INHSV2 U36021 ( .I(n30498), .ZN(n30499) );
  NAND2HSV2 U36022 ( .A1(n39744), .A2(n30499), .ZN(n30500) );
  NAND2HSV2 U36023 ( .A1(n30501), .A2(n30500), .ZN(n30502) );
  NOR2HSV4 U36024 ( .A1(n60041), .A2(n30976), .ZN(n30764) );
  INHSV2 U36025 ( .I(\pe5/ti_7t [14]), .ZN(n30503) );
  NOR2HSV2 U36026 ( .A1(n37645), .A2(n30503), .ZN(n30590) );
  INAND2HSV0 U36027 ( .A1(n30590), .B1(n39222), .ZN(n30582) );
  NOR2HSV0 U36028 ( .A1(n30507), .A2(n30506), .ZN(n30512) );
  OR2HSV1 U36029 ( .A1(n30509), .A2(n30075), .Z(n30510) );
  AOI21HSV4 U36030 ( .A1(n29660), .A2(n30512), .B(n30511), .ZN(n30581) );
  NAND2HSV2 U36031 ( .A1(n30780), .A2(n30142), .ZN(n30567) );
  NAND2HSV2 U36032 ( .A1(n30514), .A2(n30513), .ZN(n30565) );
  CLKNAND2HSV1 U36033 ( .A1(n30885), .A2(n30596), .ZN(n30564) );
  NAND2HSV0 U36034 ( .A1(n30515), .A2(n59637), .ZN(n30562) );
  CLKNAND2HSV1 U36035 ( .A1(n31151), .A2(n59948), .ZN(n30560) );
  NAND2HSV0 U36036 ( .A1(n39466), .A2(n47267), .ZN(n30518) );
  INHSV2 U36037 ( .I(n30516), .ZN(n37656) );
  CLKNAND2HSV1 U36038 ( .A1(n30785), .A2(n37656), .ZN(n30517) );
  XNOR2HSV1 U36039 ( .A1(n30518), .A2(n30517), .ZN(n30558) );
  INHSV2 U36040 ( .I(n45460), .ZN(n48206) );
  CLKNAND2HSV0 U36041 ( .A1(n30519), .A2(n48206), .ZN(n30521) );
  CLKNAND2HSV1 U36042 ( .A1(n39601), .A2(n30911), .ZN(n30520) );
  XOR2HSV0 U36043 ( .A1(n30521), .A2(n30520), .Z(n30525) );
  CLKNAND2HSV1 U36044 ( .A1(\pe5/aot [23]), .A2(n30357), .ZN(n30523) );
  INHSV2 U36045 ( .I(n40235), .ZN(n30689) );
  NAND2HSV0 U36046 ( .A1(n30689), .A2(n30607), .ZN(n30522) );
  XOR2HSV0 U36047 ( .A1(n30523), .A2(n30522), .Z(n30524) );
  XOR2HSV0 U36048 ( .A1(n30525), .A2(n30524), .Z(n30535) );
  NAND2HSV0 U36049 ( .A1(n39473), .A2(n30526), .ZN(n30528) );
  NAND2HSV0 U36050 ( .A1(n37660), .A2(n30256), .ZN(n30527) );
  XOR2HSV0 U36051 ( .A1(n30528), .A2(n30527), .Z(n30533) );
  CLKNAND2HSV1 U36052 ( .A1(n30702), .A2(n30692), .ZN(n30531) );
  NAND2HSV0 U36053 ( .A1(n30529), .A2(n30798), .ZN(n30530) );
  XOR2HSV0 U36054 ( .A1(n30531), .A2(n30530), .Z(n30532) );
  XOR2HSV0 U36055 ( .A1(n30533), .A2(n30532), .Z(n30534) );
  XOR2HSV0 U36056 ( .A1(n30535), .A2(n30534), .Z(n30537) );
  CLKNAND2HSV1 U36057 ( .A1(n30806), .A2(n40185), .ZN(n30536) );
  XNOR2HSV1 U36058 ( .A1(n30537), .A2(n30536), .ZN(n30556) );
  CLKNAND2HSV0 U36059 ( .A1(n30538), .A2(\pe5/bq[19] ), .ZN(n30540) );
  NAND2HSV0 U36060 ( .A1(n30788), .A2(n48785), .ZN(n30539) );
  XOR2HSV0 U36061 ( .A1(n30540), .A2(n30539), .Z(n30554) );
  NAND2HSV0 U36062 ( .A1(n30925), .A2(\pe5/pvq [14]), .ZN(n30541) );
  XNOR2HSV1 U36063 ( .A1(n30541), .A2(\pe5/phq [14]), .ZN(n30544) );
  CLKNAND2HSV0 U36064 ( .A1(n30543), .A2(n30542), .ZN(n30619) );
  XNOR2HSV1 U36065 ( .A1(n30544), .A2(n30619), .ZN(n30553) );
  INHSV2 U36066 ( .I(n31029), .ZN(n48199) );
  NAND2HSV0 U36067 ( .A1(n48199), .A2(n30616), .ZN(n30546) );
  NAND2HSV0 U36068 ( .A1(n30886), .A2(n30693), .ZN(n30545) );
  XOR2HSV0 U36069 ( .A1(n30546), .A2(n30545), .Z(n30551) );
  NAND2HSV0 U36070 ( .A1(n30701), .A2(n30547), .ZN(n30549) );
  INHSV2 U36071 ( .I(n29892), .ZN(n39495) );
  NAND2HSV2 U36072 ( .A1(n59638), .A2(n39495), .ZN(n30548) );
  XOR2HSV0 U36073 ( .A1(n30549), .A2(n30548), .Z(n30550) );
  XOR2HSV0 U36074 ( .A1(n30551), .A2(n30550), .Z(n30552) );
  XOR3HSV2 U36075 ( .A1(n30554), .A2(n30553), .A3(n30552), .Z(n30555) );
  XNOR2HSV1 U36076 ( .A1(n30556), .A2(n30555), .ZN(n30557) );
  XNOR2HSV1 U36077 ( .A1(n30558), .A2(n30557), .ZN(n30559) );
  XNOR2HSV1 U36078 ( .A1(n30560), .A2(n30559), .ZN(n30561) );
  NAND2HSV2 U36079 ( .A1(n39824), .A2(n37630), .ZN(n30563) );
  BUFHSV2 U36080 ( .I(n37724), .Z(n30734) );
  CLKXOR2HSV4 U36081 ( .A1(n30567), .A2(n30566), .Z(n30579) );
  NAND2HSV0 U36082 ( .A1(n30572), .A2(n30568), .ZN(n30569) );
  INHSV2 U36083 ( .I(n30569), .ZN(n30571) );
  AOI21HSV4 U36084 ( .A1(n30571), .A2(n30570), .B(n39240), .ZN(n30577) );
  CLKAND2HSV1 U36085 ( .A1(n30573), .A2(n30572), .Z(n30575) );
  CLKNAND2HSV1 U36086 ( .A1(n30575), .A2(n30574), .ZN(n30576) );
  CLKNAND2HSV2 U36087 ( .A1(n30577), .A2(n30576), .ZN(n30578) );
  XNOR2HSV4 U36088 ( .A1(n30579), .A2(n30578), .ZN(n30580) );
  XNOR2HSV4 U36089 ( .A1(n30581), .A2(n30580), .ZN(n30591) );
  OAI22HSV2 U36090 ( .A1(n30764), .A2(n30582), .B1(n30591), .B2(n30590), .ZN(
        n30586) );
  CLKNAND2HSV3 U36091 ( .A1(n60041), .A2(n39382), .ZN(n30765) );
  INHSV2 U36092 ( .I(n30765), .ZN(n30584) );
  INHSV4 U36093 ( .I(n30591), .ZN(n52768) );
  CLKNAND2HSV2 U36094 ( .A1(n30584), .A2(n52768), .ZN(n30585) );
  INHSV2 U36095 ( .I(n30753), .ZN(n37653) );
  INHSV4 U36096 ( .I(n37653), .ZN(n30752) );
  NAND2HSV2 U36097 ( .A1(n30752), .A2(\pe5/got [29]), .ZN(n30587) );
  NAND2HSV2 U36098 ( .A1(n30591), .A2(n30589), .ZN(n30594) );
  NOR2HSV2 U36099 ( .A1(n30591), .A2(n30590), .ZN(n30592) );
  AOI21HSV2 U36100 ( .A1(n30592), .A2(n30765), .B(n40309), .ZN(n30593) );
  OAI21HSV2 U36101 ( .A1(n30764), .A2(n30594), .B(n30593), .ZN(n30670) );
  NAND2HSV2 U36102 ( .A1(n45800), .A2(n30142), .ZN(n30648) );
  NAND2HSV2 U36103 ( .A1(n25854), .A2(n30779), .ZN(n30646) );
  INHSV2 U36104 ( .I(n30684), .ZN(n51162) );
  CLKNAND2HSV2 U36105 ( .A1(n51162), .A2(n30596), .ZN(n30644) );
  CLKNAND2HSV1 U36106 ( .A1(n30885), .A2(n30685), .ZN(n30642) );
  CLKNAND2HSV1 U36107 ( .A1(n37659), .A2(n30840), .ZN(n30637) );
  BUFHSV2 U36108 ( .I(n31151), .Z(n59639) );
  CLKNAND2HSV1 U36109 ( .A1(n30783), .A2(n30782), .ZN(n30598) );
  CLKNAND2HSV0 U36110 ( .A1(n30785), .A2(n40185), .ZN(n30597) );
  XNOR2HSV1 U36111 ( .A1(n30598), .A2(n30597), .ZN(n30633) );
  CLKNAND2HSV1 U36112 ( .A1(n39496), .A2(n30900), .ZN(n30600) );
  CLKNAND2HSV0 U36113 ( .A1(n39601), .A2(\pe5/bq[19] ), .ZN(n30599) );
  XOR2HSV0 U36114 ( .A1(n30600), .A2(n30599), .Z(n30604) );
  CLKNAND2HSV0 U36115 ( .A1(n52591), .A2(n39495), .ZN(n30602) );
  NAND2HSV0 U36116 ( .A1(n39446), .A2(n48785), .ZN(n30601) );
  XOR2HSV0 U36117 ( .A1(n30602), .A2(n30601), .Z(n30603) );
  XOR2HSV0 U36118 ( .A1(n30604), .A2(n30603), .Z(n30613) );
  CLKNAND2HSV0 U36119 ( .A1(\pe5/aot [23]), .A2(n30256), .ZN(n30606) );
  NAND2HSV0 U36120 ( .A1(n30689), .A2(n30798), .ZN(n30605) );
  XOR2HSV0 U36121 ( .A1(n30606), .A2(n30605), .Z(n30611) );
  NAND2HSV0 U36122 ( .A1(n30702), .A2(n30607), .ZN(n30609) );
  CLKNAND2HSV0 U36123 ( .A1(n31175), .A2(n30692), .ZN(n30608) );
  XOR2HSV0 U36124 ( .A1(n30609), .A2(n30608), .Z(n30610) );
  XOR2HSV0 U36125 ( .A1(n30611), .A2(n30610), .Z(n30612) );
  XOR2HSV0 U36126 ( .A1(n30613), .A2(n30612), .Z(n30615) );
  INHSV2 U36127 ( .I(n30686), .ZN(n37556) );
  CLKNAND2HSV0 U36128 ( .A1(n30806), .A2(n37556), .ZN(n30614) );
  XNOR2HSV1 U36129 ( .A1(n30615), .A2(n30614), .ZN(n30631) );
  NOR2HSV1 U36130 ( .A1(n37595), .A2(n45460), .ZN(n48208) );
  NAND2HSV0 U36131 ( .A1(\pe5/aot [18]), .A2(n30616), .ZN(n39799) );
  XOR2HSV0 U36132 ( .A1(n48208), .A2(n39799), .Z(n30629) );
  NAND2HSV0 U36133 ( .A1(n48029), .A2(\pe5/pvq [15]), .ZN(n30617) );
  XOR2HSV0 U36134 ( .A1(n30617), .A2(\pe5/phq [15]), .Z(n30621) );
  NAND2HSV0 U36135 ( .A1(n30799), .A2(n52585), .ZN(n30721) );
  NAND2HSV0 U36136 ( .A1(n59387), .A2(n52585), .ZN(n48193) );
  OAI21HSV0 U36137 ( .A1(n44704), .A2(n39772), .B(n48193), .ZN(n30618) );
  OAI21HSV1 U36138 ( .A1(n30619), .A2(n30721), .B(n30618), .ZN(n30620) );
  XNOR2HSV1 U36139 ( .A1(n30621), .A2(n30620), .ZN(n30628) );
  NAND2HSV2 U36140 ( .A1(n59638), .A2(n48755), .ZN(n48666) );
  XOR2HSV0 U36141 ( .A1(n30622), .A2(n48666), .Z(n30626) );
  NAND2HSV0 U36142 ( .A1(n31150), .A2(n30693), .ZN(n30624) );
  NAND2HSV0 U36143 ( .A1(n30701), .A2(n30357), .ZN(n30623) );
  XOR2HSV0 U36144 ( .A1(n30624), .A2(n30623), .Z(n30625) );
  XOR2HSV0 U36145 ( .A1(n30626), .A2(n30625), .Z(n30627) );
  XOR3HSV2 U36146 ( .A1(n30629), .A2(n30628), .A3(n30627), .Z(n30630) );
  XNOR2HSV1 U36147 ( .A1(n30631), .A2(n30630), .ZN(n30632) );
  XNOR2HSV1 U36148 ( .A1(n30633), .A2(n30632), .ZN(n30634) );
  XNOR2HSV1 U36149 ( .A1(n30635), .A2(n30634), .ZN(n30636) );
  XNOR2HSV1 U36150 ( .A1(n30637), .A2(n30636), .ZN(n30640) );
  CLKNHSV1 U36151 ( .I(n45900), .ZN(n37654) );
  CLKNAND2HSV1 U36152 ( .A1(n39824), .A2(n37654), .ZN(n30639) );
  NAND2HSV2 U36153 ( .A1(n30734), .A2(n37630), .ZN(n30638) );
  XOR3HSV2 U36154 ( .A1(n30640), .A2(n30639), .A3(n30638), .Z(n30641) );
  XNOR2HSV1 U36155 ( .A1(n30642), .A2(n30641), .ZN(n30643) );
  XNOR2HSV1 U36156 ( .A1(n30644), .A2(n30643), .ZN(n30645) );
  XOR2HSV0 U36157 ( .A1(n30646), .A2(n30645), .Z(n30647) );
  XNOR2HSV4 U36158 ( .A1(n30648), .A2(n30647), .ZN(n30659) );
  INHSV3 U36159 ( .I(n30682), .ZN(n48885) );
  NAND2HSV2 U36160 ( .A1(n52753), .A2(n48885), .ZN(n30656) );
  CLKNHSV0 U36161 ( .I(n31116), .ZN(n59395) );
  CLKNAND2HSV2 U36162 ( .A1(n30649), .A2(n59395), .ZN(n30650) );
  INHSV2 U36163 ( .I(n30650), .ZN(n30652) );
  NAND2HSV2 U36164 ( .A1(n30652), .A2(n30651), .ZN(n30655) );
  CLKNAND2HSV0 U36165 ( .A1(n30653), .A2(n48885), .ZN(n30654) );
  OAI211HSV2 U36166 ( .A1(n30657), .A2(n30656), .B(n30655), .C(n30654), .ZN(
        n30658) );
  XNOR2HSV4 U36167 ( .A1(n30659), .A2(n30658), .ZN(n30669) );
  INHSV1 U36168 ( .I(n30662), .ZN(n30660) );
  NAND2HSV2 U36169 ( .A1(n30661), .A2(n30660), .ZN(n30665) );
  INHSV2 U36170 ( .I(n30661), .ZN(n30663) );
  OAI21HSV2 U36171 ( .A1(n39405), .A2(\pe5/ti_7t [13]), .B(n39871), .ZN(n30666) );
  XNOR2HSV4 U36172 ( .A1(n30669), .A2(n30668), .ZN(n30678) );
  XNOR2HSV4 U36173 ( .A1(n30670), .A2(n30678), .ZN(n60035) );
  NOR2HSV4 U36174 ( .A1(n60035), .A2(n30204), .ZN(n30673) );
  CLKNHSV0 U36175 ( .I(\pe5/ti_7t [15]), .ZN(n30671) );
  CLKNAND2HSV1 U36176 ( .A1(n30671), .A2(n30755), .ZN(n30675) );
  CLKNHSV2 U36177 ( .I(n48885), .ZN(n31003) );
  NAND2HSV2 U36178 ( .A1(n30675), .A2(n40008), .ZN(n30672) );
  NOR2HSV8 U36179 ( .A1(n30673), .A2(n30672), .ZN(n30995) );
  NAND2HSV0 U36180 ( .A1(n30675), .A2(n30322), .ZN(n30756) );
  CLKNHSV0 U36181 ( .I(n30756), .ZN(n52786) );
  NAND2HSV0 U36182 ( .A1(n52786), .A2(n30753), .ZN(n30676) );
  NOR2HSV2 U36183 ( .A1(n30751), .A2(n30676), .ZN(n30677) );
  INHSV3 U36184 ( .I(n30677), .ZN(n31085) );
  NOR2HSV0 U36185 ( .A1(n30753), .A2(n30756), .ZN(n30680) );
  NOR2HSV4 U36186 ( .A1(n30678), .A2(n30755), .ZN(n30754) );
  INHSV2 U36187 ( .I(n30754), .ZN(n30679) );
  CLKNAND2HSV2 U36188 ( .A1(n30680), .A2(n30679), .ZN(n31087) );
  CLKNHSV0 U36189 ( .I(n39704), .ZN(n30681) );
  INHSV4 U36190 ( .I(n30753), .ZN(n30856) );
  NOR2HSV4 U36191 ( .A1(n30856), .A2(n30089), .ZN(n30750) );
  BUFHSV2 U36192 ( .I(n30682), .Z(n30966) );
  CLKNAND2HSV2 U36193 ( .A1(n30884), .A2(n39692), .ZN(n30771) );
  NAND2HSV2 U36194 ( .A1(n30884), .A2(n40008), .ZN(n30683) );
  INHSV2 U36195 ( .I(n30683), .ZN(n30748) );
  CLKNAND2HSV3 U36196 ( .A1(n39120), .A2(\pe5/got [29]), .ZN(n30747) );
  CLKNAND2HSV1 U36197 ( .A1(n45800), .A2(n30779), .ZN(n30745) );
  NAND2HSV2 U36198 ( .A1(n30781), .A2(n31225), .ZN(n30743) );
  INHSV2 U36199 ( .I(n30684), .ZN(n52578) );
  NAND2HSV2 U36200 ( .A1(n52578), .A2(n30685), .ZN(n30741) );
  NAND2HSV2 U36201 ( .A1(n39882), .A2(n37630), .ZN(n30739) );
  CLKNAND2HSV0 U36202 ( .A1(n37659), .A2(n47267), .ZN(n30733) );
  CLKNAND2HSV1 U36203 ( .A1(n59639), .A2(n30782), .ZN(n30731) );
  CLKNAND2HSV0 U36204 ( .A1(n30783), .A2(n40185), .ZN(n30688) );
  INHSV2 U36205 ( .I(n30686), .ZN(n39432) );
  NAND2HSV0 U36206 ( .A1(n30785), .A2(n39432), .ZN(n30687) );
  XNOR2HSV1 U36207 ( .A1(n30688), .A2(n30687), .ZN(n30729) );
  CLKNAND2HSV0 U36208 ( .A1(n30689), .A2(n48206), .ZN(n30691) );
  CLKNAND2HSV1 U36209 ( .A1(n30788), .A2(n39130), .ZN(n30690) );
  XOR2HSV0 U36210 ( .A1(n30691), .A2(n30690), .Z(n30697) );
  NAND2HSV0 U36211 ( .A1(n59387), .A2(n30692), .ZN(n30695) );
  NAND2HSV0 U36212 ( .A1(n37725), .A2(n30693), .ZN(n30694) );
  XOR2HSV0 U36213 ( .A1(n30695), .A2(n30694), .Z(n30696) );
  XOR2HSV0 U36214 ( .A1(n30697), .A2(n30696), .Z(n30708) );
  NAND2HSV0 U36215 ( .A1(n59879), .A2(n30825), .ZN(n30700) );
  CLKNAND2HSV1 U36216 ( .A1(\pe5/aot [18]), .A2(n30698), .ZN(n30699) );
  XOR2HSV0 U36217 ( .A1(n30700), .A2(n30699), .Z(n30706) );
  NAND2HSV0 U36218 ( .A1(n30701), .A2(n47234), .ZN(n30704) );
  NAND2HSV0 U36219 ( .A1(n30702), .A2(n30798), .ZN(n30703) );
  XOR2HSV0 U36220 ( .A1(n30704), .A2(n30703), .Z(n30705) );
  XOR2HSV0 U36221 ( .A1(n30706), .A2(n30705), .Z(n30707) );
  XOR2HSV0 U36222 ( .A1(n30708), .A2(n30707), .Z(n30710) );
  INHSV2 U36223 ( .I(n30784), .ZN(n37658) );
  NAND2HSV0 U36224 ( .A1(n30806), .A2(n37658), .ZN(n30709) );
  XNOR2HSV1 U36225 ( .A1(n30710), .A2(n30709), .ZN(n30727) );
  INHSV2 U36226 ( .I(n50518), .ZN(n51022) );
  NAND2HSV2 U36227 ( .A1(n51022), .A2(n30789), .ZN(n30712) );
  CLKNAND2HSV1 U36228 ( .A1(n31039), .A2(n30900), .ZN(n30711) );
  XOR2HSV0 U36229 ( .A1(n30712), .A2(n30711), .Z(n30716) );
  NAND2HSV2 U36230 ( .A1(\pe5/aot [23]), .A2(n40207), .ZN(n30714) );
  CLKNAND2HSV1 U36231 ( .A1(n39629), .A2(\pe5/bq[19] ), .ZN(n30713) );
  XOR2HSV0 U36232 ( .A1(n30714), .A2(n30713), .Z(n30715) );
  XOR2HSV0 U36233 ( .A1(n30716), .A2(n30715), .Z(n30720) );
  NAND2HSV0 U36234 ( .A1(n30925), .A2(\pe5/pvq [16]), .ZN(n30717) );
  XNOR2HSV1 U36235 ( .A1(n30717), .A2(\pe5/phq [16]), .ZN(n30718) );
  NOR2HSV0 U36236 ( .A1(n37595), .A2(n45426), .ZN(n30817) );
  XNOR2HSV1 U36237 ( .A1(n30718), .A2(n30817), .ZN(n30719) );
  XNOR2HSV1 U36238 ( .A1(n30720), .A2(n30719), .ZN(n30725) );
  INHSV2 U36239 ( .I(n45821), .ZN(n52595) );
  CLKNAND2HSV1 U36240 ( .A1(n39496), .A2(n52595), .ZN(n30815) );
  XOR2HSV0 U36241 ( .A1(n30721), .A2(n30815), .Z(n30723) );
  INHSV1 U36242 ( .I(n31029), .ZN(n59942) );
  CLKNHSV0 U36243 ( .I(n29892), .ZN(n40074) );
  NAND2HSV2 U36244 ( .A1(n59942), .A2(n40074), .ZN(n48197) );
  CLKNAND2HSV0 U36245 ( .A1(n59638), .A2(n30357), .ZN(n48801) );
  XOR2HSV0 U36246 ( .A1(n48197), .A2(n48801), .Z(n30722) );
  XOR2HSV0 U36247 ( .A1(n30723), .A2(n30722), .Z(n30724) );
  XNOR2HSV1 U36248 ( .A1(n30725), .A2(n30724), .ZN(n30726) );
  XNOR2HSV1 U36249 ( .A1(n30727), .A2(n30726), .ZN(n30728) );
  XNOR2HSV1 U36250 ( .A1(n30729), .A2(n30728), .ZN(n30730) );
  XNOR2HSV1 U36251 ( .A1(n30731), .A2(n30730), .ZN(n30732) );
  XNOR2HSV1 U36252 ( .A1(n30733), .A2(n30732), .ZN(n30737) );
  NAND2HSV2 U36253 ( .A1(n30944), .A2(n30840), .ZN(n30736) );
  NAND2HSV2 U36254 ( .A1(n30734), .A2(n37654), .ZN(n30735) );
  XOR3HSV2 U36255 ( .A1(n30737), .A2(n30736), .A3(n30735), .Z(n30738) );
  XNOR2HSV1 U36256 ( .A1(n30739), .A2(n30738), .ZN(n30740) );
  XNOR2HSV1 U36257 ( .A1(n30741), .A2(n30740), .ZN(n30742) );
  XOR2HSV0 U36258 ( .A1(n30743), .A2(n30742), .Z(n30744) );
  XOR2HSV0 U36259 ( .A1(n30745), .A2(n30744), .Z(n30746) );
  XNOR2HSV4 U36260 ( .A1(n30747), .A2(n30746), .ZN(n30772) );
  MUX2NHSV2 U36261 ( .I0(n30771), .I1(n30748), .S(n30772), .ZN(n30749) );
  INHSV2 U36262 ( .I(n30753), .ZN(n30960) );
  NOR2HSV2 U36263 ( .A1(n30756), .A2(n30755), .ZN(n30757) );
  INHSV2 U36264 ( .I(\pe5/ti_7t [16]), .ZN(n30758) );
  NOR2HSV2 U36265 ( .A1(n37645), .A2(n30758), .ZN(n31089) );
  CLKNAND2HSV0 U36266 ( .A1(n31089), .A2(n39578), .ZN(n30759) );
  NAND2HSV2 U36267 ( .A1(n30975), .A2(n30997), .ZN(n30762) );
  CLKNHSV2 U36268 ( .I(n30997), .ZN(n30760) );
  CLKNHSV4 U36269 ( .I(n30965), .ZN(n31091) );
  CLKNHSV2 U36270 ( .I(n30763), .ZN(n30770) );
  OAI21HSV2 U36271 ( .A1(n52768), .A2(n30764), .B(n59946), .ZN(n30768) );
  NAND2HSV2 U36272 ( .A1(n30765), .A2(n52768), .ZN(n30766) );
  INHSV2 U36273 ( .I(n30766), .ZN(n30767) );
  NOR2HSV4 U36274 ( .A1(n30768), .A2(n30767), .ZN(n30769) );
  MUX2NHSV4 U36275 ( .I0(n30771), .I1(n30770), .S(n30769), .ZN(n30774) );
  INHSV2 U36276 ( .I(n30772), .ZN(n30773) );
  XNOR2HSV4 U36277 ( .A1(n30774), .A2(n30773), .ZN(n30860) );
  CLKNAND2HSV2 U36278 ( .A1(n31091), .A2(n30860), .ZN(n52804) );
  INHSV2 U36279 ( .I(n30860), .ZN(n30776) );
  CLKNAND2HSV3 U36280 ( .A1(n30776), .A2(n30775), .ZN(n52803) );
  OAI21HSV0 U36281 ( .A1(n39405), .A2(\pe5/ti_7t [16]), .B(n52694), .ZN(n30777) );
  INHSV2 U36282 ( .I(n30777), .ZN(n52802) );
  NOR2HSV2 U36283 ( .A1(n30777), .A2(n39379), .ZN(n30872) );
  NAND3HSV4 U36284 ( .A1(n52804), .A2(n52803), .A3(n30872), .ZN(n30778) );
  INHSV4 U36285 ( .I(n30778), .ZN(n31117) );
  NAND2HSV2 U36286 ( .A1(n30884), .A2(n30046), .ZN(n30855) );
  CLKNAND2HSV1 U36287 ( .A1(n45800), .A2(n31225), .ZN(n30851) );
  CLKNHSV0 U36288 ( .I(n30780), .ZN(n45418) );
  NAND2HSV2 U36289 ( .A1(n59513), .A2(n48742), .ZN(n30849) );
  NAND2HSV2 U36290 ( .A1(n48624), .A2(n37630), .ZN(n30847) );
  CLKNAND2HSV1 U36291 ( .A1(n39882), .A2(n37654), .ZN(n30845) );
  NAND2HSV0 U36292 ( .A1(n37659), .A2(n30782), .ZN(n30839) );
  CLKNAND2HSV0 U36293 ( .A1(n59639), .A2(n40185), .ZN(n30837) );
  CLKNAND2HSV0 U36294 ( .A1(n30783), .A2(n30886), .ZN(n30787) );
  INHSV2 U36295 ( .I(n30784), .ZN(n39433) );
  NAND2HSV0 U36296 ( .A1(n30785), .A2(n39433), .ZN(n30786) );
  XNOR2HSV1 U36297 ( .A1(n30787), .A2(n30786), .ZN(n30835) );
  CLKNAND2HSV0 U36298 ( .A1(n30788), .A2(n48802), .ZN(n30791) );
  CLKNAND2HSV0 U36299 ( .A1(\pe5/aot [16]), .A2(n30789), .ZN(n30790) );
  XOR2HSV0 U36300 ( .A1(n30791), .A2(n30790), .Z(n30795) );
  INHSV2 U36301 ( .I(n30888), .ZN(n37557) );
  CLKNAND2HSV1 U36302 ( .A1(n37557), .A2(n30918), .ZN(n30793) );
  CLKNAND2HSV0 U36303 ( .A1(n59942), .A2(n48755), .ZN(n30792) );
  XOR2HSV0 U36304 ( .A1(n30793), .A2(n30792), .Z(n30794) );
  XOR2HSV0 U36305 ( .A1(n30795), .A2(n30794), .Z(n30805) );
  INHSV2 U36306 ( .I(n45451), .ZN(n39444) );
  CLKNAND2HSV0 U36307 ( .A1(n39444), .A2(n40207), .ZN(n30797) );
  NAND2HSV0 U36308 ( .A1(\pe5/aot [23]), .A2(n52585), .ZN(n30796) );
  XOR2HSV0 U36309 ( .A1(n30797), .A2(n30796), .Z(n30803) );
  NAND2HSV0 U36310 ( .A1(n59879), .A2(n30798), .ZN(n30801) );
  NAND2HSV0 U36311 ( .A1(n30799), .A2(n30891), .ZN(n30800) );
  XOR2HSV0 U36312 ( .A1(n30801), .A2(n30800), .Z(n30802) );
  XOR2HSV0 U36313 ( .A1(n30803), .A2(n30802), .Z(n30804) );
  XOR2HSV0 U36314 ( .A1(n30805), .A2(n30804), .Z(n30808) );
  NAND2HSV0 U36315 ( .A1(n30806), .A2(n37725), .ZN(n30807) );
  XNOR2HSV1 U36316 ( .A1(n30808), .A2(n30807), .ZN(n30833) );
  NOR2HSV2 U36317 ( .A1(n39123), .A2(n48822), .ZN(n30810) );
  NAND2HSV0 U36318 ( .A1(n59638), .A2(n47234), .ZN(n30809) );
  XOR2HSV0 U36319 ( .A1(n30810), .A2(n30809), .Z(n30813) );
  NAND2HSV0 U36320 ( .A1(n48049), .A2(\pe5/pvq [17]), .ZN(n30811) );
  XOR2HSV0 U36321 ( .A1(n30811), .A2(\pe5/phq [17]), .Z(n30812) );
  XOR2HSV0 U36322 ( .A1(n30813), .A2(n30812), .Z(n30823) );
  OAI22HSV0 U36323 ( .A1(n30365), .A2(n45821), .B1(n31044), .B2(n39796), .ZN(
        n30814) );
  OAI21HSV1 U36324 ( .A1(n30816), .A2(n30815), .B(n30814), .ZN(n30821) );
  CLKNHSV0 U36325 ( .I(n30817), .ZN(n30819) );
  OAI22HSV0 U36326 ( .A1(n30163), .A2(n46134), .B1(n40235), .B2(n45426), .ZN(
        n30818) );
  OAI21HSV2 U36327 ( .A1(n30819), .A2(n31177), .B(n30818), .ZN(n30820) );
  XOR2HSV0 U36328 ( .A1(n30821), .A2(n30820), .Z(n30822) );
  XOR2HSV0 U36329 ( .A1(n30823), .A2(n30822), .Z(n30831) );
  NAND2HSV2 U36330 ( .A1(\pe5/aot [18]), .A2(n48198), .ZN(n48803) );
  XOR2HSV0 U36331 ( .A1(n30824), .A2(n48803), .Z(n30829) );
  NAND2HSV0 U36332 ( .A1(n59387), .A2(n30825), .ZN(n30827) );
  CLKNAND2HSV0 U36333 ( .A1(n31161), .A2(n48206), .ZN(n30826) );
  XOR2HSV0 U36334 ( .A1(n30827), .A2(n30826), .Z(n30828) );
  XOR2HSV0 U36335 ( .A1(n30829), .A2(n30828), .Z(n30830) );
  XNOR2HSV1 U36336 ( .A1(n30831), .A2(n30830), .ZN(n30832) );
  XNOR2HSV1 U36337 ( .A1(n30833), .A2(n30832), .ZN(n30834) );
  XNOR2HSV1 U36338 ( .A1(n30835), .A2(n30834), .ZN(n30836) );
  XNOR2HSV1 U36339 ( .A1(n30837), .A2(n30836), .ZN(n30838) );
  XNOR2HSV1 U36340 ( .A1(n30839), .A2(n30838), .ZN(n30843) );
  CLKNAND2HSV1 U36341 ( .A1(n30944), .A2(n47267), .ZN(n30842) );
  NAND2HSV2 U36342 ( .A1(n47058), .A2(n30840), .ZN(n30841) );
  XOR3HSV2 U36343 ( .A1(n30843), .A2(n30842), .A3(n30841), .Z(n30844) );
  XNOR2HSV1 U36344 ( .A1(n30845), .A2(n30844), .ZN(n30846) );
  XNOR2HSV1 U36345 ( .A1(n30847), .A2(n30846), .ZN(n30848) );
  XOR2HSV0 U36346 ( .A1(n30849), .A2(n30848), .Z(n30850) );
  XOR2HSV0 U36347 ( .A1(n30851), .A2(n30850), .Z(n30852) );
  XNOR2HSV4 U36348 ( .A1(n30853), .A2(n30852), .ZN(n30854) );
  XNOR2HSV4 U36349 ( .A1(n30855), .A2(n30854), .ZN(n30858) );
  NOR2HSV4 U36350 ( .A1(n30856), .A2(n30966), .ZN(n30857) );
  XNOR2HSV4 U36351 ( .A1(n30858), .A2(n30857), .ZN(n52800) );
  NAND2HSV4 U36352 ( .A1(n60035), .A2(n37554), .ZN(n30862) );
  INHSV4 U36353 ( .I(n30870), .ZN(n30863) );
  NAND2HSV4 U36354 ( .A1(n31117), .A2(n30863), .ZN(n31006) );
  NAND3HSV2 U36355 ( .A1(n52785), .A2(n52787), .A3(n52802), .ZN(n30859) );
  NAND2HSV2 U36356 ( .A1(n30860), .A2(n52802), .ZN(n30861) );
  XOR2HSV4 U36357 ( .A1(n52800), .A2(n30862), .Z(n31126) );
  NAND2HSV4 U36358 ( .A1(n31006), .A2(n31005), .ZN(n31107) );
  INHSV2 U36359 ( .I(n52819), .ZN(n30869) );
  INHSV4 U36360 ( .I(n31135), .ZN(n31106) );
  INHSV2 U36361 ( .I(n30978), .ZN(n30865) );
  CLKNAND2HSV3 U36362 ( .A1(n31106), .A2(n30865), .ZN(n52818) );
  NOR2HSV0 U36363 ( .A1(n31102), .A2(\pe5/ti_7t [18]), .ZN(n31130) );
  NOR2HSV0 U36364 ( .A1(n31130), .A2(n39733), .ZN(n52817) );
  CLKNHSV0 U36365 ( .I(n52817), .ZN(n30866) );
  NOR2HSV2 U36366 ( .A1(n30866), .A2(n39379), .ZN(n30867) );
  CLKNHSV0 U36367 ( .I(n52804), .ZN(n30871) );
  INHSV2 U36368 ( .I(n40169), .ZN(n48741) );
  NOR2HSV2 U36369 ( .A1(n30871), .A2(n29950), .ZN(n30873) );
  NAND3HSV2 U36370 ( .A1(n30993), .A2(n30873), .A3(n29702), .ZN(n30876) );
  CLKNAND2HSV1 U36371 ( .A1(n30874), .A2(\pe5/ti_7t [17]), .ZN(n30990) );
  OR2HSV1 U36372 ( .A1(n30990), .A2(n40169), .Z(n30875) );
  CLKNAND2HSV3 U36373 ( .A1(n30876), .A2(n30875), .ZN(n30880) );
  NOR2HSV4 U36374 ( .A1(n30993), .A2(n30048), .ZN(n30877) );
  INHSV4 U36375 ( .I(n30878), .ZN(n30879) );
  NOR2HSV8 U36376 ( .A1(n30880), .A2(n30879), .ZN(n30982) );
  INHSV4 U36377 ( .I(n30982), .ZN(n30985) );
  CLKNHSV0 U36378 ( .I(n39379), .ZN(n30881) );
  NAND2HSV2 U36379 ( .A1(n60035), .A2(n30881), .ZN(n30883) );
  NAND2HSV2 U36380 ( .A1(n37638), .A2(\pe5/ti_7t [15]), .ZN(n30882) );
  NAND2HSV4 U36381 ( .A1(n30883), .A2(n30882), .ZN(n31146) );
  CLKNAND2HSV2 U36382 ( .A1(n31146), .A2(n30046), .ZN(n30964) );
  BUFHSV4 U36383 ( .I(n30884), .Z(n45819) );
  NAND2HSV2 U36384 ( .A1(n45819), .A2(n31225), .ZN(n30959) );
  CLKBUFHSV4 U36385 ( .I(n39120), .Z(n31147) );
  NAND2HSV2 U36386 ( .A1(n31147), .A2(n48742), .ZN(n30957) );
  CLKNAND2HSV1 U36387 ( .A1(n37657), .A2(n37630), .ZN(n30955) );
  NAND2HSV2 U36388 ( .A1(n40171), .A2(n37631), .ZN(n30953) );
  CLKNHSV0 U36389 ( .I(n39743), .ZN(n31148) );
  CLKNAND2HSV1 U36390 ( .A1(n40172), .A2(n31148), .ZN(n30951) );
  BUFHSV2 U36391 ( .I(n30885), .Z(n39258) );
  NAND2HSV2 U36392 ( .A1(n39258), .A2(n47267), .ZN(n30949) );
  CLKNAND2HSV1 U36393 ( .A1(n37558), .A2(n30886), .ZN(n30943) );
  NAND2HSV0 U36394 ( .A1(n31151), .A2(n31150), .ZN(n30941) );
  INHSV2 U36395 ( .I(n30887), .ZN(n40187) );
  CLKNAND2HSV1 U36396 ( .A1(n40187), .A2(n37725), .ZN(n30890) );
  INHSV2 U36397 ( .I(n30888), .ZN(n39881) );
  NAND2HSV0 U36398 ( .A1(n37608), .A2(n39881), .ZN(n30889) );
  XOR2HSV0 U36399 ( .A1(n30890), .A2(n30889), .Z(n30939) );
  NAND2HSV0 U36400 ( .A1(n39446), .A2(n47234), .ZN(n30893) );
  NAND2HSV0 U36401 ( .A1(n39444), .A2(n30891), .ZN(n30892) );
  XOR2HSV0 U36402 ( .A1(n30893), .A2(n30892), .Z(n30897) );
  CLKNAND2HSV0 U36403 ( .A1(n30529), .A2(n51041), .ZN(n30895) );
  NAND2HSV0 U36404 ( .A1(\pe5/aot [18]), .A2(n48802), .ZN(n30894) );
  XOR2HSV0 U36405 ( .A1(n30895), .A2(n30894), .Z(n30896) );
  XOR2HSV0 U36406 ( .A1(n30897), .A2(n30896), .Z(n30906) );
  BUFHSV2 U36407 ( .I(n59638), .Z(n37700) );
  NAND2HSV0 U36408 ( .A1(n37700), .A2(n30526), .ZN(n30899) );
  NAND2HSV0 U36409 ( .A1(n37660), .A2(n31178), .ZN(n30898) );
  XOR2HSV0 U36410 ( .A1(n30899), .A2(n30898), .Z(n30904) );
  NAND2HSV0 U36411 ( .A1(n31048), .A2(n30900), .ZN(n30902) );
  CLKNHSV1 U36412 ( .I(n50518), .ZN(n40210) );
  NAND2HSV0 U36413 ( .A1(n40210), .A2(n39130), .ZN(n30901) );
  XOR2HSV0 U36414 ( .A1(n30902), .A2(n30901), .Z(n30903) );
  XOR2HSV0 U36415 ( .A1(n30904), .A2(n30903), .Z(n30905) );
  XOR2HSV0 U36416 ( .A1(n30906), .A2(n30905), .Z(n30908) );
  CLKNAND2HSV0 U36417 ( .A1(n30806), .A2(n31007), .ZN(n30907) );
  XNOR2HSV1 U36418 ( .A1(n30908), .A2(n30907), .ZN(n30937) );
  NAND2HSV0 U36419 ( .A1(\pe5/aot [23]), .A2(n31160), .ZN(n30910) );
  NAND2HSV0 U36420 ( .A1(n30788), .A2(n40207), .ZN(n30909) );
  XOR2HSV0 U36421 ( .A1(n30910), .A2(n30909), .Z(n30915) );
  NAND2HSV0 U36422 ( .A1(n31161), .A2(\pe5/bq[19] ), .ZN(n30913) );
  CLKNHSV0 U36423 ( .I(n48219), .ZN(n31175) );
  NAND2HSV0 U36424 ( .A1(n31175), .A2(n30911), .ZN(n30912) );
  XOR2HSV0 U36425 ( .A1(n30913), .A2(n30912), .Z(n30914) );
  XOR2HSV0 U36426 ( .A1(n30915), .A2(n30914), .Z(n30924) );
  CLKNAND2HSV1 U36427 ( .A1(n48681), .A2(n31192), .ZN(n30917) );
  INHSV2 U36428 ( .I(n48823), .ZN(n50653) );
  CLKNAND2HSV0 U36429 ( .A1(n50653), .A2(n39436), .ZN(n30916) );
  XOR2HSV0 U36430 ( .A1(n30917), .A2(n30916), .Z(n30922) );
  NAND2HSV0 U36431 ( .A1(n39629), .A2(n52610), .ZN(n30920) );
  INHSV2 U36432 ( .I(n31199), .ZN(n39259) );
  CLKNAND2HSV0 U36433 ( .A1(n39259), .A2(n30918), .ZN(n30919) );
  XOR2HSV0 U36434 ( .A1(n30920), .A2(n30919), .Z(n30921) );
  XOR2HSV0 U36435 ( .A1(n30922), .A2(n30921), .Z(n30923) );
  XOR2HSV0 U36436 ( .A1(n30924), .A2(n30923), .Z(n30935) );
  NAND2HSV0 U36437 ( .A1(n30925), .A2(\pe5/pvq [19]), .ZN(n30926) );
  XOR2HSV0 U36438 ( .A1(n30926), .A2(\pe5/phq [19]), .Z(n30929) );
  INHSV2 U36439 ( .I(\pe5/bq[14] ), .ZN(n31041) );
  INHSV2 U36440 ( .I(n31041), .ZN(n39472) );
  CLKNAND2HSV0 U36441 ( .A1(n31039), .A2(n39472), .ZN(n31194) );
  INHSV2 U36442 ( .I(\pe5/bq[14] ), .ZN(n48186) );
  OAI22HSV0 U36443 ( .A1(n39779), .A2(n51057), .B1(n31044), .B2(n48186), .ZN(
        n30927) );
  OAI21HSV1 U36444 ( .A1(n31194), .A2(n39586), .B(n30927), .ZN(n30928) );
  XNOR2HSV1 U36445 ( .A1(n30929), .A2(n30928), .ZN(n30933) );
  XOR2HSV0 U36446 ( .A1(n30931), .A2(n30930), .Z(n30932) );
  XNOR2HSV1 U36447 ( .A1(n30933), .A2(n30932), .ZN(n30934) );
  XNOR2HSV1 U36448 ( .A1(n30935), .A2(n30934), .ZN(n30936) );
  XOR2HSV0 U36449 ( .A1(n30937), .A2(n30936), .Z(n30938) );
  XOR2HSV0 U36450 ( .A1(n30939), .A2(n30938), .Z(n30940) );
  XOR2HSV0 U36451 ( .A1(n30941), .A2(n30940), .Z(n30942) );
  XOR2HSV0 U36452 ( .A1(n30943), .A2(n30942), .Z(n30947) );
  CLKNAND2HSV0 U36453 ( .A1(n30944), .A2(\pe5/got [20]), .ZN(n30946) );
  CLKNAND2HSV0 U36454 ( .A1(n47338), .A2(n31149), .ZN(n30945) );
  XOR3HSV2 U36455 ( .A1(n30947), .A2(n30946), .A3(n30945), .Z(n30948) );
  XNOR2HSV1 U36456 ( .A1(n30949), .A2(n30948), .ZN(n30950) );
  XOR2HSV0 U36457 ( .A1(n30951), .A2(n30950), .Z(n30952) );
  XOR2HSV0 U36458 ( .A1(n30953), .A2(n30952), .Z(n30954) );
  XOR2HSV0 U36459 ( .A1(n30955), .A2(n30954), .Z(n30956) );
  XOR2HSV0 U36460 ( .A1(n30957), .A2(n30956), .Z(n30958) );
  CLKXOR2HSV4 U36461 ( .A1(n30959), .A2(n30958), .Z(n30962) );
  XNOR2HSV4 U36462 ( .A1(n30962), .A2(n30961), .ZN(n30963) );
  INAND2HSV2 U36463 ( .A1(n30965), .B1(n59395), .ZN(n30971) );
  INHSV4 U36464 ( .I(n31140), .ZN(n52788) );
  NAND2HSV2 U36465 ( .A1(n31087), .A2(n31085), .ZN(n30967) );
  INHSV2 U36466 ( .I(n30966), .ZN(n48740) );
  NAND2HSV2 U36467 ( .A1(n39741), .A2(n48740), .ZN(n39247) );
  NOR2HSV2 U36468 ( .A1(n30967), .A2(n39247), .ZN(n30968) );
  NAND2HSV0 U36469 ( .A1(n30968), .A2(n52788), .ZN(n30970) );
  CLKNAND2HSV1 U36470 ( .A1(n31089), .A2(n48740), .ZN(n30969) );
  OAI211HSV2 U36471 ( .A1(n30971), .A2(n52788), .B(n30970), .C(n30969), .ZN(
        n30972) );
  INHSV4 U36472 ( .I(n30984), .ZN(n30983) );
  NAND2HSV2 U36473 ( .A1(n30985), .A2(n30983), .ZN(n30974) );
  NAND2HSV2 U36474 ( .A1(n30982), .A2(n30984), .ZN(n30973) );
  INHSV2 U36475 ( .I(n31107), .ZN(n30977) );
  XNOR2HSV4 U36476 ( .A1(n30975), .A2(n30997), .ZN(n31111) );
  AOI31HSV2 U36477 ( .A1(n30977), .A2(n31111), .A3(n52817), .B(n30976), .ZN(
        n30980) );
  NAND2HSV2 U36478 ( .A1(n30980), .A2(n30979), .ZN(n30981) );
  INHSV4 U36479 ( .I(n30981), .ZN(n31242) );
  CLKNAND2HSV2 U36480 ( .A1(n30983), .A2(n30982), .ZN(n30987) );
  CLKNAND2HSV4 U36481 ( .A1(n30986), .A2(n30987), .ZN(n52816) );
  INHSV2 U36482 ( .I(\pe5/ti_7t [19]), .ZN(n30988) );
  NOR2HSV2 U36483 ( .A1(n39705), .A2(n30988), .ZN(n37753) );
  INHSV2 U36484 ( .I(n37753), .ZN(n37540) );
  NAND3HSV2 U36485 ( .A1(n37550), .A2(n37549), .A3(n37540), .ZN(n30989) );
  NAND2HSV2 U36486 ( .A1(n30989), .A2(n29825), .ZN(n31098) );
  INHSV2 U36487 ( .I(n30990), .ZN(n31119) );
  BUFHSV2 U36488 ( .I(n30992), .Z(n39693) );
  NOR2HSV2 U36489 ( .A1(n37534), .A2(n40009), .ZN(n30999) );
  CLKNHSV2 U36490 ( .I(n30995), .ZN(n30996) );
  AND2HSV2 U36491 ( .A1(\pe5/ti_7t [18]), .A2(n39245), .Z(n37639) );
  INHSV2 U36492 ( .I(n37639), .ZN(n31001) );
  CLKNAND2HSV1 U36493 ( .A1(n31000), .A2(n31001), .ZN(n31002) );
  INHSV0 U36494 ( .I(n31119), .ZN(n31004) );
  NAND3HSV3 U36495 ( .A1(n31006), .A2(n31005), .A3(n31004), .ZN(n37652) );
  CLKNAND2HSV1 U36496 ( .A1(n31146), .A2(n31225), .ZN(n31084) );
  NAND2HSV2 U36497 ( .A1(n45819), .A2(n37630), .ZN(n31080) );
  CLKNAND2HSV1 U36498 ( .A1(n31147), .A2(n45500), .ZN(n31078) );
  CLKNAND2HSV0 U36499 ( .A1(n37657), .A2(n31148), .ZN(n31076) );
  NAND2HSV2 U36500 ( .A1(n30781), .A2(n48744), .ZN(n31074) );
  CLKNAND2HSV0 U36501 ( .A1(n40172), .A2(n37656), .ZN(n31072) );
  CLKNAND2HSV0 U36502 ( .A1(n39258), .A2(n45816), .ZN(n31070) );
  CLKNAND2HSV0 U36503 ( .A1(n37558), .A2(n37725), .ZN(n31064) );
  NAND2HSV0 U36504 ( .A1(n39583), .A2(n37557), .ZN(n31062) );
  CLKNAND2HSV0 U36505 ( .A1(n40187), .A2(n31007), .ZN(n31009) );
  INHSV2 U36506 ( .I(n31199), .ZN(n40186) );
  NAND2HSV0 U36507 ( .A1(n37608), .A2(n40186), .ZN(n31008) );
  XOR2HSV0 U36508 ( .A1(n31009), .A2(n31008), .Z(n31060) );
  NAND2HSV0 U36509 ( .A1(n39490), .A2(n39495), .ZN(n31011) );
  NAND2HSV0 U36510 ( .A1(\pe5/got [12]), .A2(n37584), .ZN(n31010) );
  XOR2HSV0 U36511 ( .A1(n31011), .A2(n31010), .Z(n31015) );
  NAND2HSV0 U36512 ( .A1(n51022), .A2(n48787), .ZN(n31013) );
  NAND2HSV0 U36513 ( .A1(n59640), .A2(n45470), .ZN(n31012) );
  XOR2HSV0 U36514 ( .A1(n31013), .A2(n31012), .Z(n31014) );
  XOR2HSV0 U36515 ( .A1(n31015), .A2(n31014), .Z(n31023) );
  NOR2HSV0 U36516 ( .A1(n44704), .A2(n45426), .ZN(n31017) );
  NAND2HSV0 U36517 ( .A1(n30529), .A2(n53314), .ZN(n31016) );
  XOR2HSV0 U36518 ( .A1(n31017), .A2(n31016), .Z(n31021) );
  INHSV2 U36519 ( .I(n50507), .ZN(n48658) );
  CLKNAND2HSV0 U36520 ( .A1(n48658), .A2(n31192), .ZN(n31019) );
  NAND2HSV0 U36521 ( .A1(\pe5/aot [13]), .A2(n39436), .ZN(n31018) );
  XOR2HSV0 U36522 ( .A1(n31019), .A2(n31018), .Z(n31020) );
  XOR2HSV0 U36523 ( .A1(n31021), .A2(n31020), .Z(n31022) );
  XOR2HSV0 U36524 ( .A1(n31023), .A2(n31022), .Z(n31038) );
  NOR2HSV0 U36525 ( .A1(n45815), .A2(n30452), .ZN(n31025) );
  NAND2HSV0 U36526 ( .A1(\pe5/aot [23]), .A2(n31190), .ZN(n31024) );
  XOR2HSV0 U36527 ( .A1(n31025), .A2(n31024), .Z(n31028) );
  NAND2HSV0 U36528 ( .A1(n37707), .A2(\pe5/pvq [21]), .ZN(n31026) );
  XOR2HSV0 U36529 ( .A1(n31026), .A2(\pe5/phq [21]), .Z(n31027) );
  XOR2HSV0 U36530 ( .A1(n31028), .A2(n31027), .Z(n31036) );
  NAND2HSV0 U36531 ( .A1(n39446), .A2(n40207), .ZN(n31191) );
  NAND2HSV0 U36532 ( .A1(\pe5/aot [18]), .A2(n30526), .ZN(n37559) );
  OAI22HSV0 U36533 ( .A1(n39772), .A2(n45858), .B1(n31029), .B2(n30287), .ZN(
        n31030) );
  OAI21HSV1 U36534 ( .A1(n31191), .A2(n37559), .B(n31030), .ZN(n31034) );
  CLKNAND2HSV0 U36535 ( .A1(n39444), .A2(n39454), .ZN(n39263) );
  OAI22HSV0 U36536 ( .A1(n30150), .A2(n46134), .B1(n45451), .B2(n45844), .ZN(
        n31031) );
  OAI21HSV0 U36537 ( .A1(n39263), .A2(n31032), .B(n31031), .ZN(n31033) );
  XOR2HSV0 U36538 ( .A1(n31034), .A2(n31033), .Z(n31035) );
  XOR2HSV0 U36539 ( .A1(n31036), .A2(n31035), .Z(n31037) );
  XNOR2HSV1 U36540 ( .A1(n31038), .A2(n31037), .ZN(n31058) );
  NAND2HSV0 U36541 ( .A1(n31039), .A2(\pe5/bq[13] ), .ZN(n40045) );
  XOR2HSV0 U36542 ( .A1(n31040), .A2(n40045), .Z(n31043) );
  CLKNAND2HSV0 U36543 ( .A1(n37700), .A2(n31160), .ZN(n47304) );
  INHSV2 U36544 ( .I(n31041), .ZN(n40221) );
  CLKNAND2HSV1 U36545 ( .A1(n39629), .A2(n40221), .ZN(n48185) );
  XOR2HSV0 U36546 ( .A1(n47304), .A2(n48185), .Z(n31042) );
  XOR2HSV0 U36547 ( .A1(n31043), .A2(n31042), .Z(n31054) );
  CLKNAND2HSV0 U36548 ( .A1(n31175), .A2(n50444), .ZN(n31047) );
  CLKNHSV0 U36549 ( .I(n31044), .ZN(n59366) );
  CLKNAND2HSV0 U36550 ( .A1(n59366), .A2(n31045), .ZN(n31046) );
  XOR2HSV0 U36551 ( .A1(n31047), .A2(n31046), .Z(n31052) );
  INHSV2 U36552 ( .I(n48823), .ZN(n59943) );
  CLKNAND2HSV0 U36553 ( .A1(n59943), .A2(n48755), .ZN(n31050) );
  NAND2HSV0 U36554 ( .A1(n31048), .A2(n48181), .ZN(n31049) );
  XOR2HSV0 U36555 ( .A1(n31050), .A2(n31049), .Z(n31051) );
  XOR2HSV0 U36556 ( .A1(n31052), .A2(n31051), .Z(n31053) );
  XOR2HSV0 U36557 ( .A1(n31054), .A2(n31053), .Z(n31056) );
  INHSV2 U36558 ( .I(n45817), .ZN(n59367) );
  NAND2HSV0 U36559 ( .A1(n39278), .A2(n59367), .ZN(n31055) );
  XNOR2HSV1 U36560 ( .A1(n31056), .A2(n31055), .ZN(n31057) );
  XOR2HSV0 U36561 ( .A1(n31058), .A2(n31057), .Z(n31059) );
  XNOR2HSV1 U36562 ( .A1(n31060), .A2(n31059), .ZN(n31061) );
  XNOR2HSV1 U36563 ( .A1(n31062), .A2(n31061), .ZN(n31063) );
  XNOR2HSV1 U36564 ( .A1(n31064), .A2(n31063), .ZN(n31068) );
  INHSV2 U36565 ( .I(n44332), .ZN(n37723) );
  CLKNAND2HSV1 U36566 ( .A1(n37723), .A2(n37658), .ZN(n31067) );
  CLKNAND2HSV0 U36567 ( .A1(n47058), .A2(n37556), .ZN(n31066) );
  XOR3HSV2 U36568 ( .A1(n31068), .A2(n31067), .A3(n31066), .Z(n31069) );
  XNOR2HSV1 U36569 ( .A1(n31070), .A2(n31069), .ZN(n31071) );
  XNOR2HSV1 U36570 ( .A1(n31072), .A2(n31071), .ZN(n31073) );
  XOR2HSV0 U36571 ( .A1(n31074), .A2(n31073), .Z(n31075) );
  XOR2HSV0 U36572 ( .A1(n31076), .A2(n31075), .Z(n31077) );
  XOR2HSV0 U36573 ( .A1(n31078), .A2(n31077), .Z(n31079) );
  XNOR2HSV1 U36574 ( .A1(n31080), .A2(n31079), .ZN(n31083) );
  NAND2HSV0 U36575 ( .A1(n44694), .A2(n48742), .ZN(n31082) );
  INHSV2 U36576 ( .I(n31089), .ZN(n31142) );
  CLKNHSV1 U36577 ( .I(n31142), .ZN(n31090) );
  NAND2HSV2 U36578 ( .A1(n31092), .A2(n31143), .ZN(n39341) );
  NAND2HSV2 U36579 ( .A1(n39341), .A2(n39430), .ZN(n31093) );
  XOR2HSV2 U36580 ( .A1(n31094), .A2(n31093), .Z(n31095) );
  XNOR2HSV4 U36581 ( .A1(n31097), .A2(n37531), .ZN(n37760) );
  XNOR2HSV4 U36582 ( .A1(n31098), .A2(n37760), .ZN(n31252) );
  NAND2HSV4 U36583 ( .A1(n31100), .A2(n31099), .ZN(n31243) );
  CLKNHSV1 U36584 ( .I(n31243), .ZN(n31104) );
  NAND2HSV0 U36585 ( .A1(n39718), .A2(n39995), .ZN(n31105) );
  CLKNAND2HSV2 U36586 ( .A1(n31106), .A2(n31105), .ZN(n31110) );
  INHSV2 U36587 ( .I(n31113), .ZN(n31109) );
  CLKNAND2HSV1 U36588 ( .A1(n31111), .A2(n39247), .ZN(n31108) );
  NAND3HSV3 U36589 ( .A1(n31109), .A2(n31110), .A3(n31108), .ZN(n31236) );
  NAND2HSV2 U36590 ( .A1(n37652), .A2(n39692), .ZN(n31114) );
  NAND3HSV4 U36591 ( .A1(n31115), .A2(n31114), .A3(n31113), .ZN(n39216) );
  NOR2HSV4 U36592 ( .A1(n31126), .A2(n31116), .ZN(n31118) );
  CLKNAND2HSV2 U36593 ( .A1(n31118), .A2(n31117), .ZN(n31129) );
  NAND2HSV0 U36594 ( .A1(n31119), .A2(n48740), .ZN(n31128) );
  NAND2HSV0 U36595 ( .A1(n37639), .A2(n48741), .ZN(n31120) );
  AND2HSV2 U36596 ( .A1(n31128), .A2(n31120), .Z(n31127) );
  CLKNHSV0 U36597 ( .I(n31121), .ZN(n31125) );
  NAND3HSV3 U36598 ( .A1(n31126), .A2(n31125), .A3(n31124), .ZN(n31134) );
  NAND3HSV2 U36599 ( .A1(n31129), .A2(n31127), .A3(n31134), .ZN(n31138) );
  NOR2HSV0 U36600 ( .A1(n31130), .A2(n40169), .ZN(n31131) );
  CLKNAND2HSV3 U36601 ( .A1(n31132), .A2(n31131), .ZN(n31137) );
  NOR2HSV2 U36602 ( .A1(n31136), .A2(n31135), .ZN(n39215) );
  AOI21HSV4 U36603 ( .A1(n31137), .A2(n31138), .B(n39215), .ZN(n31139) );
  INHSV2 U36604 ( .I(n31141), .ZN(n31144) );
  INHSV2 U36605 ( .I(n31146), .ZN(n39118) );
  CLKNAND2HSV1 U36606 ( .A1(n31146), .A2(n30513), .ZN(n31229) );
  NAND2HSV2 U36607 ( .A1(n45819), .A2(n48742), .ZN(n31224) );
  NAND2HSV2 U36608 ( .A1(n31147), .A2(n48739), .ZN(n31222) );
  NAND2HSV2 U36609 ( .A1(n37657), .A2(n37631), .ZN(n31220) );
  NAND2HSV2 U36610 ( .A1(n25854), .A2(n31148), .ZN(n31218) );
  NAND2HSV2 U36611 ( .A1(n40172), .A2(\pe5/got [22]), .ZN(n31216) );
  NAND2HSV2 U36612 ( .A1(n39258), .A2(n31149), .ZN(n31214) );
  NAND2HSV2 U36613 ( .A1(n37558), .A2(n31150), .ZN(n31209) );
  NAND2HSV0 U36614 ( .A1(n31151), .A2(n37725), .ZN(n31207) );
  NAND2HSV2 U36615 ( .A1(n40187), .A2(n37557), .ZN(n31153) );
  INHSV2 U36616 ( .I(n48722), .ZN(n39516) );
  NAND2HSV0 U36617 ( .A1(n37608), .A2(n39516), .ZN(n31152) );
  XOR2HSV0 U36618 ( .A1(n31153), .A2(n31152), .Z(n31205) );
  CLKNAND2HSV0 U36619 ( .A1(n59938), .A2(n48181), .ZN(n31155) );
  CLKNAND2HSV0 U36620 ( .A1(n39490), .A2(n39436), .ZN(n31154) );
  XOR2HSV0 U36621 ( .A1(n31155), .A2(n31154), .Z(n31159) );
  CLKNAND2HSV1 U36622 ( .A1(n59366), .A2(\pe5/bq[13] ), .ZN(n31157) );
  NAND2HSV0 U36623 ( .A1(n59367), .A2(n37584), .ZN(n31156) );
  XOR2HSV0 U36624 ( .A1(n31157), .A2(n31156), .Z(n31158) );
  XOR2HSV0 U36625 ( .A1(n31159), .A2(n31158), .Z(n31169) );
  CLKNAND2HSV1 U36626 ( .A1(n39444), .A2(n31160), .ZN(n31163) );
  NAND2HSV0 U36627 ( .A1(n31161), .A2(n39443), .ZN(n31162) );
  XOR2HSV0 U36628 ( .A1(n31163), .A2(n31162), .Z(n31167) );
  NAND2HSV0 U36629 ( .A1(n30788), .A2(n30526), .ZN(n31165) );
  CLKNHSV0 U36630 ( .I(n30150), .ZN(n39269) );
  CLKNHSV0 U36631 ( .I(n45426), .ZN(n37685) );
  CLKNAND2HSV1 U36632 ( .A1(n39269), .A2(n37685), .ZN(n31164) );
  XOR2HSV0 U36633 ( .A1(n31165), .A2(n31164), .Z(n31166) );
  XOR2HSV0 U36634 ( .A1(n31167), .A2(n31166), .Z(n31168) );
  XOR2HSV0 U36635 ( .A1(n31169), .A2(n31168), .Z(n31183) );
  CLKNAND2HSV1 U36636 ( .A1(n59640), .A2(n39130), .ZN(n31171) );
  NAND2HSV0 U36637 ( .A1(n59943), .A2(n48198), .ZN(n31170) );
  XOR2HSV0 U36638 ( .A1(n31171), .A2(n31170), .Z(n31174) );
  NAND2HSV0 U36639 ( .A1(n44335), .A2(\pe5/pvq [20]), .ZN(n31172) );
  XNOR2HSV1 U36640 ( .A1(n31172), .A2(\pe5/phq [20]), .ZN(n31173) );
  XNOR2HSV1 U36641 ( .A1(n31174), .A2(n31173), .ZN(n31181) );
  CLKNAND2HSV1 U36642 ( .A1(n31175), .A2(n51041), .ZN(n37560) );
  OAI22HSV0 U36643 ( .A1(n40235), .A2(n45821), .B1(n48219), .B2(n46134), .ZN(
        n31176) );
  OAI21HSV2 U36644 ( .A1(n37560), .A2(n31177), .B(n31176), .ZN(n31179) );
  CLKNAND2HSV0 U36645 ( .A1(\pe5/aot [23]), .A2(n31178), .ZN(n52624) );
  XNOR2HSV1 U36646 ( .A1(n31179), .A2(n52624), .ZN(n31180) );
  XNOR2HSV1 U36647 ( .A1(n31181), .A2(n31180), .ZN(n31182) );
  XNOR2HSV1 U36648 ( .A1(n31183), .A2(n31182), .ZN(n31203) );
  NAND2HSV0 U36649 ( .A1(n39629), .A2(n53314), .ZN(n31185) );
  NAND2HSV0 U36650 ( .A1(\pe5/aot [18]), .A2(n47234), .ZN(n31184) );
  XOR2HSV0 U36651 ( .A1(n31185), .A2(n31184), .Z(n31189) );
  NAND2HSV2 U36652 ( .A1(n37700), .A2(n30891), .ZN(n31187) );
  NAND2HSV0 U36653 ( .A1(n51022), .A2(n45470), .ZN(n31186) );
  XOR2HSV0 U36654 ( .A1(n31187), .A2(n31186), .Z(n31188) );
  XOR2HSV0 U36655 ( .A1(n31189), .A2(n31188), .Z(n31198) );
  NAND2HSV2 U36656 ( .A1(n37660), .A2(n31190), .ZN(n37562) );
  XOR2HSV0 U36657 ( .A1(n37562), .A2(n31191), .Z(n31196) );
  CLKNAND2HSV1 U36658 ( .A1(\pe5/aot [13]), .A2(n31192), .ZN(n31193) );
  XOR2HSV0 U36659 ( .A1(n31194), .A2(n31193), .Z(n31195) );
  XOR2HSV0 U36660 ( .A1(n31196), .A2(n31195), .Z(n31197) );
  XOR2HSV0 U36661 ( .A1(n31198), .A2(n31197), .Z(n31201) );
  INHSV2 U36662 ( .I(n31199), .ZN(n39582) );
  CLKNAND2HSV1 U36663 ( .A1(n59393), .A2(n39582), .ZN(n31200) );
  XNOR2HSV1 U36664 ( .A1(n31201), .A2(n31200), .ZN(n31202) );
  XOR2HSV0 U36665 ( .A1(n31203), .A2(n31202), .Z(n31204) );
  XNOR2HSV1 U36666 ( .A1(n31205), .A2(n31204), .ZN(n31206) );
  XNOR2HSV1 U36667 ( .A1(n31207), .A2(n31206), .ZN(n31208) );
  XNOR2HSV1 U36668 ( .A1(n31209), .A2(n31208), .ZN(n31212) );
  NAND2HSV2 U36669 ( .A1(n37723), .A2(n37556), .ZN(n31211) );
  CLKNAND2HSV0 U36670 ( .A1(n48848), .A2(\pe5/got [20]), .ZN(n31210) );
  XOR3HSV2 U36671 ( .A1(n31212), .A2(n31211), .A3(n31210), .Z(n31213) );
  XNOR2HSV1 U36672 ( .A1(n31214), .A2(n31213), .ZN(n31215) );
  XNOR2HSV1 U36673 ( .A1(n31216), .A2(n31215), .ZN(n31217) );
  XOR2HSV0 U36674 ( .A1(n31218), .A2(n31217), .Z(n31219) );
  XNOR2HSV1 U36675 ( .A1(n31220), .A2(n31219), .ZN(n31221) );
  XOR2HSV0 U36676 ( .A1(n31222), .A2(n31221), .Z(n31223) );
  XNOR2HSV1 U36677 ( .A1(n31224), .A2(n31223), .ZN(n31227) );
  NAND2HSV2 U36678 ( .A1(n44694), .A2(n31225), .ZN(n31226) );
  XOR2HSV0 U36679 ( .A1(n31227), .A2(n31226), .Z(n31228) );
  XNOR2HSV1 U36680 ( .A1(n31229), .A2(n31228), .ZN(n31230) );
  CLKXOR2HSV4 U36681 ( .A1(n31231), .A2(n31230), .Z(n31233) );
  INHSV2 U36682 ( .I(n31233), .ZN(n39223) );
  OAI21HSV4 U36683 ( .A1(n31232), .A2(n31235), .B(n39223), .ZN(n31247) );
  INHSV2 U36684 ( .I(n31233), .ZN(n31234) );
  NOR2HSV4 U36685 ( .A1(n31235), .A2(n31234), .ZN(n31237) );
  NAND2HSV4 U36686 ( .A1(n31237), .A2(n31236), .ZN(n31246) );
  CLKNAND2HSV4 U36687 ( .A1(n31247), .A2(n31246), .ZN(n37756) );
  INHSV2 U36688 ( .I(\pe5/ti_7t [20]), .ZN(n31239) );
  NAND2HSV2 U36689 ( .A1(n31239), .A2(n39239), .ZN(n39251) );
  NAND2HSV0 U36690 ( .A1(n39251), .A2(n31240), .ZN(n37529) );
  INHSV2 U36691 ( .I(n37529), .ZN(n31241) );
  NAND2HSV2 U36692 ( .A1(n31242), .A2(n52816), .ZN(n31244) );
  CLKNHSV0 U36693 ( .I(n37642), .ZN(n31245) );
  INHSV2 U36694 ( .I(n31245), .ZN(n31249) );
  CLKNAND2HSV4 U36695 ( .A1(n31247), .A2(n31246), .ZN(n39117) );
  NOR2HSV4 U36696 ( .A1(n39117), .A2(n37551), .ZN(n31248) );
  CLKNAND2HSV4 U36697 ( .A1(n31248), .A2(n31249), .ZN(n37765) );
  CLKNAND2HSV2 U36698 ( .A1(n29711), .A2(n37765), .ZN(n31251) );
  CLKNAND2HSV3 U36699 ( .A1(n31252), .A2(n31251), .ZN(n31250) );
  OAI21HSV4 U36700 ( .A1(n31252), .A2(n31251), .B(n31250), .ZN(n60025) );
  INHSV2 U36701 ( .I(\pe6/pvq [1]), .ZN(n31254) );
  CLKBUFHSV4 U36702 ( .I(n31298), .Z(n31893) );
  INHSV2 U36703 ( .I(n31893), .ZN(n31873) );
  INHSV2 U36704 ( .I(ctro6), .ZN(n31461) );
  INHSV2 U36705 ( .I(n31461), .ZN(n47950) );
  NAND2HSV2 U36706 ( .A1(\pe6/ti_7t [1]), .A2(n47950), .ZN(n31258) );
  CLKBUFHSV4 U36707 ( .I(n31260), .Z(n31302) );
  NAND2HSV2 U36708 ( .A1(n31283), .A2(n31284), .ZN(n31262) );
  NOR2HSV4 U36709 ( .A1(n31263), .A2(n31262), .ZN(n31264) );
  NOR2HSV4 U36710 ( .A1(n31265), .A2(n31264), .ZN(n31383) );
  INHSV2 U36711 ( .I(n31440), .ZN(n31366) );
  INHSV4 U36712 ( .I(n31366), .ZN(n35725) );
  NOR2HSV1 U36713 ( .A1(n31424), .A2(n35917), .ZN(n31267) );
  BUFHSV8 U36714 ( .I(n31844), .Z(n31312) );
  NOR2HSV4 U36715 ( .A1(n31312), .A2(n31487), .ZN(n31268) );
  INHSV2 U36716 ( .I(n31268), .ZN(n31266) );
  OAI21HSV2 U36717 ( .A1(n31424), .A2(n35917), .B(n31268), .ZN(n31270) );
  NAND2HSV2 U36718 ( .A1(\pe6/phq [2]), .A2(\pe6/pvq [2]), .ZN(n31272) );
  NOR2HSV4 U36719 ( .A1(n31255), .A2(n31272), .ZN(n31278) );
  INHSV2 U36720 ( .I(n31278), .ZN(n31274) );
  AOI21HSV4 U36721 ( .A1(n32881), .A2(\pe6/pvq [2]), .B(\pe6/phq [2]), .ZN(
        n31277) );
  INHSV2 U36722 ( .I(\pe6/bq[31] ), .ZN(n35631) );
  INHSV2 U36723 ( .I(n35631), .ZN(n46625) );
  NAND3HSV4 U36724 ( .A1(n31275), .A2(n31273), .A3(n31274), .ZN(n31290) );
  OAI21HSV4 U36725 ( .A1(n31278), .A2(n31277), .B(n31276), .ZN(n31292) );
  CLKNAND2HSV1 U36726 ( .A1(n31290), .A2(n31292), .ZN(n31279) );
  INHSV4 U36727 ( .I(n31324), .ZN(n31326) );
  INHSV4 U36728 ( .I(n31326), .ZN(n31441) );
  BUFHSV2 U36729 ( .I(n25463), .Z(n33063) );
  NAND2HSV2 U36730 ( .A1(n32822), .A2(n29742), .ZN(n31381) );
  NOR2HSV4 U36731 ( .A1(n31441), .A2(n31381), .ZN(n31282) );
  CLKNAND2HSV3 U36732 ( .A1(n31282), .A2(n35725), .ZN(n31476) );
  NOR2HSV0 U36733 ( .A1(n31303), .A2(n31302), .ZN(n31285) );
  INHSV2 U36734 ( .I(n31285), .ZN(n31287) );
  NAND2HSV2 U36735 ( .A1(n31302), .A2(n31303), .ZN(n31286) );
  CLKNAND2HSV1 U36736 ( .A1(n31353), .A2(n44378), .ZN(n31296) );
  CLKNAND2HSV1 U36737 ( .A1(n31292), .A2(n31290), .ZN(n31289) );
  INHSV2 U36738 ( .I(n31382), .ZN(n31295) );
  NOR2HSV4 U36739 ( .A1(n31296), .A2(n31295), .ZN(n31474) );
  BUFHSV2 U36740 ( .I(n25463), .Z(n32348) );
  CLKBUFHSV4 U36741 ( .I(n31298), .Z(n31900) );
  INHSV2 U36742 ( .I(n31900), .ZN(n36055) );
  OR2HSV1 U36743 ( .A1(n32053), .A2(n36055), .Z(n31377) );
  CLKNHSV0 U36744 ( .I(n31377), .ZN(n31297) );
  NAND2HSV2 U36745 ( .A1(n31324), .A2(n31297), .ZN(n31300) );
  INHSV2 U36746 ( .I(\pe6/ti_7t [2]), .ZN(n31575) );
  CLKBUFHSV4 U36747 ( .I(n31298), .Z(n31883) );
  NAND2HSV2 U36748 ( .A1(n31575), .A2(n36023), .ZN(n31500) );
  INHSV2 U36749 ( .I(n35796), .ZN(n36089) );
  CLKAND2HSV2 U36750 ( .A1(n31500), .A2(n36089), .Z(n31299) );
  CLKNAND2HSV3 U36751 ( .A1(n31300), .A2(n31299), .ZN(n31473) );
  NOR2HSV2 U36752 ( .A1(n26485), .A2(n31303), .ZN(n31304) );
  AOI21HSV4 U36753 ( .A1(n31303), .A2(n26485), .B(n31304), .ZN(n48017) );
  CLKNAND2HSV3 U36754 ( .A1(n48017), .A2(n32961), .ZN(n31307) );
  CLKNHSV0 U36755 ( .I(\pe6/ti_7t [1]), .ZN(n31305) );
  AOI21HSV2 U36756 ( .A1(n31305), .A2(n32329), .B(n44376), .ZN(n31306) );
  CLKNAND2HSV3 U36757 ( .A1(n31307), .A2(n31306), .ZN(n31318) );
  CLKNAND2HSV1 U36758 ( .A1(\pe6/bq[31] ), .A2(\pe6/aot [30]), .ZN(n31308) );
  XNOR2HSV1 U36759 ( .A1(n31308), .A2(\pe6/phq [4]), .ZN(n31316) );
  INHSV2 U36760 ( .I(n31487), .ZN(n59278) );
  CLKNAND2HSV0 U36761 ( .A1(\pe6/pvq [4]), .A2(\pe6/ctrq ), .ZN(n31309) );
  CLKXOR2HSV4 U36762 ( .A1(n31310), .A2(n31309), .Z(n31315) );
  INHSV4 U36763 ( .I(\pe6/aot [29]), .ZN(n31924) );
  INHSV4 U36764 ( .I(n31924), .ZN(n31491) );
  INHSV4 U36765 ( .I(n31491), .ZN(n31311) );
  NOR2HSV8 U36766 ( .A1(n31312), .A2(n31311), .ZN(n32101) );
  CLKAND2HSV2 U36767 ( .A1(\pe6/ti_1 ), .A2(\pe6/got [29]), .Z(n31313) );
  XNOR2HSV4 U36768 ( .A1(n32101), .A2(n31313), .ZN(n31314) );
  CLKNAND2HSV1 U36769 ( .A1(n31319), .A2(n31477), .ZN(n31323) );
  INHSV2 U36770 ( .I(n31319), .ZN(n31321) );
  INHSV2 U36771 ( .I(n31477), .ZN(n31320) );
  CLKNAND2HSV2 U36772 ( .A1(n31321), .A2(n31320), .ZN(n31322) );
  INHSV4 U36773 ( .I(n31326), .ZN(n31389) );
  NAND2HSV2 U36774 ( .A1(n31328), .A2(n31388), .ZN(n31348) );
  CLKBUFHSV4 U36775 ( .I(n31900), .Z(n31527) );
  INHSV2 U36776 ( .I(\pe6/ti_7t [3]), .ZN(n31329) );
  NOR2HSV2 U36777 ( .A1(n31527), .A2(n31329), .ZN(n31443) );
  INHSV2 U36778 ( .I(n31443), .ZN(n31358) );
  INHSV2 U36779 ( .I(n36089), .ZN(n31442) );
  NOR2HSV1 U36780 ( .A1(n31353), .A2(n31442), .ZN(n31342) );
  NAND3HSV2 U36781 ( .A1(n31369), .A2(n31368), .A3(n31330), .ZN(n31333) );
  INHSV2 U36782 ( .I(n31330), .ZN(n31331) );
  OAI21HSV2 U36783 ( .A1(n31253), .A2(n31425), .B(n31331), .ZN(n31332) );
  NAND2HSV2 U36784 ( .A1(n31333), .A2(n31332), .ZN(n31338) );
  INHSV3 U36785 ( .I(\pe6/aot [30]), .ZN(n31334) );
  INHSV2 U36786 ( .I(n31334), .ZN(n31367) );
  CLKNAND2HSV1 U36787 ( .A1(n26514), .A2(\pe6/phq [3]), .ZN(n31336) );
  XNOR2HSV4 U36788 ( .A1(n31338), .A2(n31337), .ZN(n31344) );
  CLKBUFHSV4 U36789 ( .I(\pe6/ctrq ), .Z(n31593) );
  NAND2HSV2 U36790 ( .A1(n31593), .A2(\pe6/pvq [3]), .ZN(n31341) );
  INHSV4 U36791 ( .I(n32443), .ZN(n59168) );
  CLKNAND2HSV1 U36792 ( .A1(n59168), .A2(n31339), .ZN(n31340) );
  XOR2HSV2 U36793 ( .A1(n31341), .A2(n31340), .Z(n31343) );
  XNOR2HSV4 U36794 ( .A1(n31344), .A2(n31343), .ZN(n31445) );
  INHSV4 U36795 ( .I(n31445), .ZN(n31352) );
  XNOR2HSV4 U36796 ( .A1(n31344), .A2(n31343), .ZN(n52704) );
  BUFHSV2 U36797 ( .I(n35796), .Z(n44372) );
  INHSV2 U36798 ( .I(n44372), .ZN(n31345) );
  INHSV2 U36799 ( .I(n31893), .ZN(n44380) );
  CLKNAND2HSV2 U36800 ( .A1(n31347), .A2(n31346), .ZN(n31392) );
  CLKNHSV0 U36801 ( .I(n36089), .ZN(n31349) );
  NOR2HSV2 U36802 ( .A1(n48017), .A2(n31349), .ZN(n31351) );
  INHSV2 U36803 ( .I(n32463), .ZN(n31350) );
  AOI21HSV4 U36804 ( .A1(n31352), .A2(n31351), .B(n31350), .ZN(n31357) );
  BUFHSV2 U36805 ( .I(n35796), .Z(n36229) );
  INHSV4 U36806 ( .I(n36229), .ZN(n46765) );
  CLKNAND2HSV1 U36807 ( .A1(n31354), .A2(n46765), .ZN(n31355) );
  NAND2HSV2 U36808 ( .A1(n31355), .A2(n52704), .ZN(n31356) );
  NOR2HSV2 U36809 ( .A1(n31497), .A2(n31441), .ZN(n31360) );
  CLKNAND2HSV1 U36810 ( .A1(n31388), .A2(n31358), .ZN(n31359) );
  NOR2HSV2 U36811 ( .A1(n31360), .A2(n31359), .ZN(n31361) );
  CLKNAND2HSV3 U36812 ( .A1(n31456), .A2(n31361), .ZN(n31364) );
  BUFHSV2 U36813 ( .I(n25463), .Z(n32053) );
  NAND2HSV4 U36814 ( .A1(n31363), .A2(n31362), .ZN(n31578) );
  NAND3HSV2 U36815 ( .A1(n31578), .A2(n31579), .A3(n35908), .ZN(n31521) );
  CLKNHSV0 U36816 ( .I(n31521), .ZN(n31398) );
  INHSV2 U36817 ( .I(\pe6/got [29]), .ZN(n31903) );
  INHSV2 U36818 ( .I(n31903), .ZN(n31667) );
  NOR2HSV2 U36819 ( .A1(n31366), .A2(n31373), .ZN(n31371) );
  CLKNAND2HSV1 U36820 ( .A1(\pe6/aot [28]), .A2(\pe6/bq[32] ), .ZN(n31370) );
  INHSV2 U36821 ( .I(n31372), .ZN(n31374) );
  CLKNAND2HSV2 U36822 ( .A1(n31376), .A2(n31375), .ZN(n31387) );
  INHSV2 U36823 ( .I(n31377), .ZN(n35914) );
  CLKNAND2HSV4 U36824 ( .A1(n31572), .A2(n35914), .ZN(n31502) );
  CLKNHSV0 U36825 ( .I(n31500), .ZN(n31378) );
  BUFHSV2 U36826 ( .I(n35710), .Z(n44376) );
  NOR2HSV2 U36827 ( .A1(n31378), .A2(n44376), .ZN(n31379) );
  CLKNAND2HSV3 U36828 ( .A1(n31502), .A2(n31379), .ZN(n31380) );
  INHSV2 U36829 ( .I(n31380), .ZN(n31385) );
  INHSV2 U36830 ( .I(n31893), .ZN(n44369) );
  INHSV2 U36831 ( .I(n44369), .ZN(n32044) );
  CLKNAND2HSV2 U36832 ( .A1(n31382), .A2(n32044), .ZN(n31451) );
  INHSV3 U36833 ( .I(n31451), .ZN(n31410) );
  NOR2HSV2 U36834 ( .A1(n31382), .A2(n31381), .ZN(n31384) );
  INHSV6 U36835 ( .I(n52706), .ZN(n31592) );
  MUX2NHSV4 U36836 ( .I0(n31410), .I1(n31384), .S(n31592), .ZN(n31503) );
  CLKNAND2HSV3 U36837 ( .A1(n31385), .A2(n31503), .ZN(n31386) );
  XNOR2HSV4 U36838 ( .A1(n31387), .A2(n31386), .ZN(n31397) );
  AND2HSV2 U36839 ( .A1(n31500), .A2(n32348), .Z(n52709) );
  CLKNAND2HSV3 U36840 ( .A1(n31388), .A2(n52709), .ZN(n31391) );
  NOR2HSV4 U36841 ( .A1(n31389), .A2(n31497), .ZN(n31390) );
  NOR2HSV8 U36842 ( .A1(n31391), .A2(n31390), .ZN(n31457) );
  INHSV2 U36843 ( .I(n31443), .ZN(n31449) );
  BUFHSV2 U36844 ( .I(n35917), .Z(n32239) );
  AOI31HSV2 U36845 ( .A1(n31457), .A2(n31456), .A3(n31449), .B(n32239), .ZN(
        n31395) );
  INHSV2 U36846 ( .I(n31449), .ZN(n31453) );
  NOR2HSV4 U36847 ( .A1(n31457), .A2(n31453), .ZN(n31393) );
  CLKNAND2HSV1 U36848 ( .A1(n31393), .A2(n31392), .ZN(n31394) );
  NAND3HSV2 U36849 ( .A1(n31398), .A2(n31402), .A3(n46765), .ZN(n31407) );
  INHSV2 U36850 ( .I(n31578), .ZN(n31400) );
  CLKNAND2HSV2 U36851 ( .A1(n31579), .A2(n32348), .ZN(n31399) );
  NOR2HSV2 U36852 ( .A1(n31400), .A2(n31399), .ZN(n31401) );
  INHSV2 U36853 ( .I(n31401), .ZN(n31524) );
  NOR2HSV2 U36854 ( .A1(n32239), .A2(n36023), .ZN(n31816) );
  INHSV2 U36855 ( .I(n31816), .ZN(n36081) );
  INHSV2 U36856 ( .I(n36081), .ZN(n36065) );
  INHSV2 U36857 ( .I(\pe6/ti_7t [5]), .ZN(n31403) );
  NOR2HSV2 U36858 ( .A1(n31527), .A2(n31403), .ZN(n31534) );
  CLKNHSV0 U36859 ( .I(n31534), .ZN(n31404) );
  BUFHSV2 U36860 ( .I(n35917), .Z(n52705) );
  NOR2HSV2 U36861 ( .A1(n31404), .A2(n52705), .ZN(n31405) );
  INHSV2 U36862 ( .I(n33063), .ZN(n46159) );
  NOR2HSV4 U36863 ( .A1(n31434), .A2(n46159), .ZN(n31573) );
  INHSV2 U36864 ( .I(n31573), .ZN(n31411) );
  INHSV2 U36865 ( .I(n47950), .ZN(n32047) );
  NOR2HSV2 U36866 ( .A1(n31572), .A2(n44380), .ZN(n31408) );
  NAND2HSV2 U36867 ( .A1(n31573), .A2(n31408), .ZN(n31413) );
  INHSV2 U36868 ( .I(\pe6/got [28]), .ZN(n32466) );
  NAND2HSV0 U36869 ( .A1(n31500), .A2(n31590), .ZN(n31409) );
  AOI21HSV2 U36870 ( .A1(n31411), .A2(n31410), .B(n31409), .ZN(n31412) );
  CLKNAND2HSV1 U36871 ( .A1(n31413), .A2(n31412), .ZN(n31439) );
  NAND2HSV2 U36872 ( .A1(n31413), .A2(n31412), .ZN(n31414) );
  INHSV2 U36873 ( .I(n31414), .ZN(n31438) );
  BUFHSV2 U36874 ( .I(n46620), .Z(n31928) );
  INHSV2 U36875 ( .I(n31928), .ZN(n31718) );
  CLKNHSV1 U36876 ( .I(n31924), .ZN(n46677) );
  NAND2HSV2 U36877 ( .A1(n31718), .A2(n46677), .ZN(n31416) );
  INHSV2 U36878 ( .I(\pe6/bq[27] ), .ZN(n31908) );
  INHSV2 U36879 ( .I(n31908), .ZN(n31644) );
  CLKNAND2HSV3 U36880 ( .A1(n44446), .A2(n31644), .ZN(n31415) );
  INHSV4 U36881 ( .I(\pe6/aot [26]), .ZN(n32079) );
  CLKNHSV1 U36882 ( .I(n32079), .ZN(n31417) );
  NAND2HSV2 U36883 ( .A1(n31418), .A2(n31417), .ZN(n31420) );
  INHSV2 U36884 ( .I(n31791), .ZN(n31831) );
  CLKNAND2HSV1 U36885 ( .A1(n32740), .A2(n31831), .ZN(n31419) );
  BUFHSV2 U36886 ( .I(\pe6/ctrq ), .Z(n32198) );
  XNOR2HSV4 U36887 ( .A1(n31421), .A2(n29638), .ZN(n31422) );
  XNOR2HSV4 U36888 ( .A1(n31423), .A2(n31422), .ZN(n31433) );
  INHSV2 U36889 ( .I(n32166), .ZN(n36101) );
  CLKNHSV2 U36890 ( .I(n31269), .ZN(n46176) );
  CLKNAND2HSV1 U36891 ( .A1(n36101), .A2(n46176), .ZN(n31427) );
  INHSV4 U36892 ( .I(n31425), .ZN(n31776) );
  INHSV2 U36893 ( .I(n35816), .ZN(n46643) );
  CLKNAND2HSV1 U36894 ( .A1(n31776), .A2(n46643), .ZN(n31426) );
  XNOR2HSV1 U36895 ( .A1(n31427), .A2(n31426), .ZN(n31431) );
  INHSV2 U36896 ( .I(\pe6/bq[28] ), .ZN(n31561) );
  INHSV2 U36897 ( .I(n31561), .ZN(n31595) );
  INHSV2 U36898 ( .I(\pe6/aot [30]), .ZN(n32193) );
  CLKNAND2HSV1 U36899 ( .A1(n31595), .A2(n31910), .ZN(n31429) );
  INHSV2 U36900 ( .I(n32589), .ZN(n59061) );
  CLKNAND2HSV1 U36901 ( .A1(n31990), .A2(n59061), .ZN(n31428) );
  XOR2HSV0 U36902 ( .A1(n31429), .A2(n31428), .Z(n31430) );
  XNOR2HSV1 U36903 ( .A1(n31431), .A2(n31430), .ZN(n31432) );
  XNOR2HSV4 U36904 ( .A1(n31433), .A2(n31432), .ZN(n31436) );
  CLKNAND2HSV0 U36905 ( .A1(n44426), .A2(\pe6/got [27]), .ZN(n31435) );
  XNOR2HSV4 U36906 ( .A1(n31436), .A2(n31435), .ZN(n31437) );
  MUX2NHSV4 U36907 ( .I0(n31439), .I1(n31438), .S(n31437), .ZN(n31460) );
  INHSV2 U36908 ( .I(n31903), .ZN(n49736) );
  INHSV2 U36909 ( .I(n52706), .ZN(n31454) );
  NOR2HSV0 U36910 ( .A1(n31443), .A2(n48010), .ZN(n31450) );
  NOR2HSV0 U36911 ( .A1(n31443), .A2(n31442), .ZN(n31444) );
  NAND2HSV2 U36912 ( .A1(n31445), .A2(n31444), .ZN(n31446) );
  CLKNAND2HSV2 U36913 ( .A1(n31447), .A2(n31446), .ZN(n31448) );
  CLKNAND2HSV1 U36914 ( .A1(n31451), .A2(n31450), .ZN(n31452) );
  OAI21HSV2 U36915 ( .A1(n31453), .A2(n52704), .B(n31452), .ZN(n31455) );
  NAND2HSV2 U36916 ( .A1(n31455), .A2(n31366), .ZN(n31506) );
  NAND2HSV2 U36917 ( .A1(n31472), .A2(n31510), .ZN(n31591) );
  NAND2HSV2 U36918 ( .A1(n49736), .A2(n31591), .ZN(n31459) );
  NAND2HSV2 U36919 ( .A1(n31578), .A2(n31579), .ZN(n48009) );
  INHSV2 U36920 ( .I(n36055), .ZN(n31817) );
  CLKNAND2HSV1 U36921 ( .A1(n48009), .A2(n31817), .ZN(n31465) );
  INHSV2 U36922 ( .I(\pe6/ti_7t [4]), .ZN(n31462) );
  INHSV2 U36923 ( .I(n32463), .ZN(n46584) );
  NAND2HSV2 U36924 ( .A1(n31462), .A2(n46584), .ZN(n31479) );
  CLKNHSV1 U36925 ( .I(n31479), .ZN(n31463) );
  NOR2HSV2 U36926 ( .A1(n31463), .A2(n32651), .ZN(n31464) );
  NAND2HSV2 U36927 ( .A1(n31465), .A2(n31464), .ZN(n31467) );
  NAND2HSV2 U36928 ( .A1(n31466), .A2(n31467), .ZN(n31471) );
  INHSV2 U36929 ( .I(n31466), .ZN(n31469) );
  INHSV2 U36930 ( .I(n31467), .ZN(n31468) );
  CLKNAND2HSV1 U36931 ( .A1(n31469), .A2(n31468), .ZN(n31470) );
  NOR2HSV2 U36932 ( .A1(n32697), .A2(n32148), .ZN(n31517) );
  NOR2HSV2 U36933 ( .A1(n31474), .A2(n31473), .ZN(n31475) );
  CLKBUFHSV4 U36934 ( .I(n31478), .Z(n31516) );
  CLKAND2HSV2 U36935 ( .A1(n31479), .A2(n46154), .Z(n31480) );
  NAND2HSV0 U36936 ( .A1(n35908), .A2(n32697), .ZN(n31481) );
  INHSV2 U36937 ( .I(n31481), .ZN(n31483) );
  INHSV2 U36938 ( .I(n31516), .ZN(n31482) );
  NAND2HSV4 U36939 ( .A1(n31483), .A2(n31482), .ZN(n31518) );
  CLKNAND2HSV2 U36940 ( .A1(n31484), .A2(n31518), .ZN(n31514) );
  NOR2HSV2 U36941 ( .A1(n32193), .A2(n31928), .ZN(n31486) );
  CLKNHSV2 U36942 ( .I(\pe6/bq[31] ), .ZN(n44411) );
  NOR2HSV2 U36943 ( .A1(n35816), .A2(n44411), .ZN(n31489) );
  NAND2HSV2 U36944 ( .A1(n31595), .A2(\pe6/aot [31]), .ZN(n31488) );
  XOR2HSV2 U36945 ( .A1(n31489), .A2(n31488), .Z(n31490) );
  NOR2HSV2 U36946 ( .A1(n31425), .A2(n32589), .ZN(n31609) );
  CLKNHSV0 U36947 ( .I(n31609), .ZN(n31494) );
  CLKNHSV0 U36948 ( .I(n32101), .ZN(n31493) );
  INHSV2 U36949 ( .I(n32589), .ZN(n46662) );
  OAI21HSV2 U36950 ( .A1(n31494), .A2(n31493), .B(n31492), .ZN(n31496) );
  CLKNAND2HSV1 U36951 ( .A1(n31644), .A2(n59276), .ZN(n31495) );
  NOR2HSV4 U36952 ( .A1(n31497), .A2(n35907), .ZN(n31498) );
  XNOR2HSV4 U36953 ( .A1(n31499), .A2(n31498), .ZN(n31505) );
  AND2HSV2 U36954 ( .A1(n31500), .A2(n31667), .Z(n31501) );
  NAND2HSV2 U36955 ( .A1(n31503), .A2(n29708), .ZN(n31504) );
  XNOR2HSV4 U36956 ( .A1(n31505), .A2(n31504), .ZN(n31512) );
  INHSV2 U36957 ( .I(n35710), .ZN(n32647) );
  CLKNAND2HSV1 U36958 ( .A1(n31506), .A2(n32647), .ZN(n31509) );
  INHSV2 U36959 ( .I(n31507), .ZN(n31508) );
  OAI22HSV4 U36960 ( .A1(n32651), .A2(n31510), .B1(n31509), .B2(n31508), .ZN(
        n31511) );
  XNOR2HSV4 U36961 ( .A1(n31512), .A2(n31511), .ZN(n31519) );
  CLKNAND2HSV3 U36962 ( .A1(n31514), .A2(n31513), .ZN(n31627) );
  AOI21HSV2 U36963 ( .A1(n31517), .A2(n31516), .B(n31515), .ZN(n31520) );
  NAND3HSV4 U36964 ( .A1(n31520), .A2(n31519), .A3(n31518), .ZN(n31628) );
  NOR2HSV2 U36965 ( .A1(n31521), .A2(n31522), .ZN(n31535) );
  BUFHSV2 U36966 ( .I(n31900), .Z(n31690) );
  INHSV2 U36967 ( .I(n31690), .ZN(n32057) );
  NAND2HSV2 U36968 ( .A1(n31522), .A2(n31690), .ZN(n31523) );
  INHSV2 U36969 ( .I(n31523), .ZN(n31525) );
  BUFHSV2 U36970 ( .I(n31527), .Z(n52701) );
  NAND3HSV2 U36971 ( .A1(n31627), .A2(n36083), .A3(n31628), .ZN(n31537) );
  INHSV2 U36972 ( .I(\pe6/ti_7t [6]), .ZN(n31528) );
  CLKBUFHSV4 U36973 ( .I(n31883), .Z(n44378) );
  INHSV2 U36974 ( .I(n44378), .ZN(n48001) );
  NAND2HSV2 U36975 ( .A1(n31528), .A2(n48001), .ZN(n31673) );
  INHSV1 U36976 ( .I(n31673), .ZN(n31529) );
  NOR2HSV2 U36977 ( .A1(n31529), .A2(n32439), .ZN(n31532) );
  CLKNAND2HSV0 U36978 ( .A1(n31537), .A2(n31532), .ZN(n31530) );
  INHSV1 U36979 ( .I(n31530), .ZN(n31531) );
  INHSV2 U36980 ( .I(n31532), .ZN(n31685) );
  INHSV2 U36981 ( .I(n31685), .ZN(n31533) );
  NOR2HSV4 U36982 ( .A1(n31535), .A2(n31534), .ZN(n31541) );
  CLKNAND2HSV3 U36983 ( .A1(n31540), .A2(n31541), .ZN(n31621) );
  CLKBUFHSV4 U36984 ( .I(n31621), .Z(n59011) );
  INHSV2 U36985 ( .I(n59011), .ZN(n31536) );
  CLKNHSV1 U36986 ( .I(n31537), .ZN(n31538) );
  CLKNAND2HSV0 U36987 ( .A1(n31538), .A2(n31621), .ZN(n31680) );
  NAND3HSV4 U36988 ( .A1(n31676), .A2(n29668), .A3(n31680), .ZN(n31638) );
  NAND2HSV2 U36989 ( .A1(\pe6/ti_7t [7]), .A2(n48001), .ZN(n51439) );
  CLKNAND2HSV2 U36990 ( .A1(n31743), .A2(n51439), .ZN(n46123) );
  INHSV2 U36991 ( .I(n31903), .ZN(n31902) );
  CLKNAND2HSV2 U36992 ( .A1(n46123), .A2(n31902), .ZN(n31589) );
  BUFHSV2 U36993 ( .I(n29742), .Z(n35798) );
  CLKNAND2HSV3 U36994 ( .A1(n31621), .A2(n35798), .ZN(n48002) );
  INHSV2 U36995 ( .I(n48002), .ZN(n31539) );
  INHSV4 U36996 ( .I(n31625), .ZN(n48003) );
  CLKNAND2HSV2 U36997 ( .A1(n31539), .A2(n48003), .ZN(n31672) );
  NAND2HSV4 U36998 ( .A1(n31541), .A2(n31540), .ZN(n31683) );
  CLKNAND2HSV2 U36999 ( .A1(n31683), .A2(n35798), .ZN(n48004) );
  BUFHSV2 U37000 ( .I(n31625), .Z(n31670) );
  AOI21HSV2 U37001 ( .A1(n48004), .A2(n31670), .B(n36023), .ZN(n31542) );
  CLKNAND2HSV1 U37002 ( .A1(n31672), .A2(n31542), .ZN(n31543) );
  NAND2HSV2 U37003 ( .A1(\pe6/ti_7t [6]), .A2(n36050), .ZN(n31706) );
  CLKNAND2HSV3 U37004 ( .A1(n31543), .A2(n31706), .ZN(n31769) );
  NAND2HSV2 U37005 ( .A1(n31769), .A2(\pe6/got [28]), .ZN(n31587) );
  BUFHSV4 U37006 ( .I(n32697), .Z(n32384) );
  INHSV2 U37007 ( .I(n46750), .ZN(n31861) );
  NAND2HSV2 U37008 ( .A1(n59594), .A2(n31861), .ZN(n31583) );
  NAND2HSV2 U37009 ( .A1(n31990), .A2(n36153), .ZN(n31545) );
  CLKNHSV0 U37010 ( .I(n31908), .ZN(n31820) );
  CLKNAND2HSV0 U37011 ( .A1(n31820), .A2(n59061), .ZN(n31544) );
  XOR2HSV0 U37012 ( .A1(n31545), .A2(n31544), .Z(n31548) );
  INHSV2 U37013 ( .I(n49003), .ZN(n58714) );
  CLKNAND2HSV1 U37014 ( .A1(n33016), .A2(n58714), .ZN(n31546) );
  XNOR2HSV1 U37015 ( .A1(n31546), .A2(\pe6/phq [11]), .ZN(n31547) );
  XNOR2HSV1 U37016 ( .A1(n31548), .A2(n31547), .ZN(n31550) );
  NAND2HSV2 U37017 ( .A1(n31831), .A2(n59065), .ZN(n31793) );
  INHSV2 U37018 ( .I(n59194), .ZN(n31845) );
  INHSV2 U37019 ( .I(n32193), .ZN(n31910) );
  CLKNAND2HSV1 U37020 ( .A1(n31845), .A2(n31910), .ZN(n35734) );
  XOR2HSV0 U37021 ( .A1(n31793), .A2(n35734), .Z(n31549) );
  XOR2HSV0 U37022 ( .A1(n31550), .A2(n31549), .Z(n31552) );
  NOR2HSV0 U37023 ( .A1(n31366), .A2(n49315), .ZN(n31551) );
  XOR2HSV0 U37024 ( .A1(n31552), .A2(n31551), .Z(n31571) );
  INHSV2 U37025 ( .I(\pe6/bq[22] ), .ZN(n31979) );
  INHSV2 U37026 ( .I(n31979), .ZN(n31925) );
  NAND2HSV2 U37027 ( .A1(n31925), .A2(n59276), .ZN(n31554) );
  INHSV2 U37028 ( .I(\pe6/bq[23] ), .ZN(n32068) );
  INHSV2 U37029 ( .I(n32068), .ZN(n31830) );
  NAND2HSV0 U37030 ( .A1(n31830), .A2(n44446), .ZN(n31553) );
  XOR2HSV0 U37031 ( .A1(n31554), .A2(n31553), .Z(n31559) );
  CLKNHSV0 U37032 ( .I(n31425), .ZN(n35740) );
  NAND2HSV2 U37033 ( .A1(n35740), .A2(n59239), .ZN(n31557) );
  CLKNHSV0 U37034 ( .I(n31924), .ZN(n31555) );
  INHSV2 U37035 ( .I(n31555), .ZN(n35817) );
  CLKNAND2HSV0 U37036 ( .A1(n59206), .A2(n31829), .ZN(n31556) );
  XOR2HSV0 U37037 ( .A1(n31557), .A2(n31556), .Z(n31558) );
  XOR2HSV0 U37038 ( .A1(n31559), .A2(n31558), .Z(n31569) );
  CLKNAND2HSV1 U37039 ( .A1(n32576), .A2(n49831), .ZN(n31563) );
  INHSV2 U37040 ( .I(n31561), .ZN(n46135) );
  INHSV2 U37041 ( .I(n32079), .ZN(n31785) );
  NAND2HSV0 U37042 ( .A1(n46135), .A2(n31785), .ZN(n31562) );
  XOR2HSV0 U37043 ( .A1(n31563), .A2(n31562), .Z(n31567) );
  INHSV2 U37044 ( .I(n46663), .ZN(n32605) );
  CLKNAND2HSV0 U37045 ( .A1(n31718), .A2(n32605), .ZN(n31564) );
  XOR2HSV0 U37046 ( .A1(n31565), .A2(n31564), .Z(n31566) );
  XOR2HSV0 U37047 ( .A1(n31567), .A2(n31566), .Z(n31568) );
  XOR2HSV0 U37048 ( .A1(n31569), .A2(n31568), .Z(n31570) );
  XNOR2HSV1 U37049 ( .A1(n31571), .A2(n31570), .ZN(n31577) );
  XNOR2HSV4 U37050 ( .A1(n31573), .A2(n31572), .ZN(n52700) );
  NAND2HSV2 U37051 ( .A1(n52700), .A2(n31817), .ZN(n31574) );
  OAI21HSV4 U37052 ( .A1(n31575), .A2(n32685), .B(n31574), .ZN(n31944) );
  CLKNAND2HSV0 U37053 ( .A1(n31944), .A2(n31717), .ZN(n31576) );
  CLKXOR2HSV2 U37054 ( .A1(n31577), .A2(n31576), .Z(n31582) );
  NAND3HSV2 U37055 ( .A1(n31579), .A2(n31578), .A3(n32463), .ZN(n31580) );
  NAND2HSV2 U37056 ( .A1(\pe6/ti_7t [4]), .A2(n32949), .ZN(n48011) );
  NAND2HSV4 U37057 ( .A1(n31580), .A2(n48011), .ZN(n31949) );
  BUFHSV3 U37058 ( .I(n31949), .Z(n58940) );
  NAND2HSV2 U37059 ( .A1(n58940), .A2(n32242), .ZN(n31581) );
  XOR3HSV2 U37060 ( .A1(n31583), .A2(n31582), .A3(n31581), .Z(n31585) );
  CLKBUFHSV4 U37061 ( .I(n31683), .Z(n59595) );
  BUFHSV2 U37062 ( .I(\pe6/got [27]), .Z(n35789) );
  NAND2HSV2 U37063 ( .A1(n59595), .A2(n35789), .ZN(n31584) );
  XOR2HSV0 U37064 ( .A1(n31585), .A2(n31584), .Z(n31586) );
  XOR2HSV2 U37065 ( .A1(n31587), .A2(n31586), .Z(n31588) );
  XNOR2HSV4 U37066 ( .A1(n31589), .A2(n31588), .ZN(n31643) );
  CLKNAND2HSV1 U37067 ( .A1(n31592), .A2(n36101), .ZN(n31601) );
  NAND2HSV2 U37068 ( .A1(n31718), .A2(n46643), .ZN(n46645) );
  NAND2HSV0 U37069 ( .A1(n31593), .A2(\pe6/pvq [8]), .ZN(n31594) );
  XOR2HSV0 U37070 ( .A1(n46645), .A2(n31594), .Z(n31599) );
  CLKNAND2HSV1 U37071 ( .A1(n31595), .A2(n31829), .ZN(n31597) );
  CLKNAND2HSV1 U37072 ( .A1(n31990), .A2(n31785), .ZN(n31596) );
  XOR2HSV0 U37073 ( .A1(n31597), .A2(n31596), .Z(n31598) );
  XOR2HSV0 U37074 ( .A1(n31599), .A2(n31598), .Z(n31600) );
  XNOR2HSV4 U37075 ( .A1(n31601), .A2(n31600), .ZN(n31614) );
  CLKNAND2HSV1 U37076 ( .A1(n31644), .A2(n32991), .ZN(n31603) );
  CLKNAND2HSV1 U37077 ( .A1(n46624), .A2(n59276), .ZN(n31602) );
  XOR2HSV0 U37078 ( .A1(n31603), .A2(n31602), .Z(n31607) );
  INHSV2 U37079 ( .I(n31791), .ZN(n48035) );
  NAND2HSV2 U37080 ( .A1(n48035), .A2(n44446), .ZN(n31605) );
  INHSV2 U37081 ( .I(n46663), .ZN(n59087) );
  XOR2HSV0 U37082 ( .A1(n31605), .A2(n31604), .Z(n31606) );
  XOR2HSV0 U37083 ( .A1(n31607), .A2(n31606), .Z(n31612) );
  NAND2HSV2 U37084 ( .A1(n33016), .A2(n31710), .ZN(n31608) );
  XNOR2HSV1 U37085 ( .A1(n31608), .A2(\pe6/phq [8]), .ZN(n31610) );
  XNOR2HSV1 U37086 ( .A1(n31610), .A2(n31609), .ZN(n31611) );
  XNOR2HSV1 U37087 ( .A1(n31612), .A2(n31611), .ZN(n31613) );
  XNOR2HSV1 U37088 ( .A1(n31614), .A2(n31613), .ZN(n31615) );
  XNOR2HSV4 U37089 ( .A1(n31616), .A2(n31615), .ZN(n31618) );
  BUFHSV2 U37090 ( .I(\pe6/got [27]), .Z(n32815) );
  CLKAND2HSV1 U37091 ( .A1(n31944), .A2(n32815), .Z(n31617) );
  XNOR2HSV4 U37092 ( .A1(n31618), .A2(n31617), .ZN(n31620) );
  XNOR2HSV4 U37093 ( .A1(n31620), .A2(n31619), .ZN(n31623) );
  INHSV2 U37094 ( .I(n35710), .ZN(n32411) );
  CLKNAND2HSV1 U37095 ( .A1(n31621), .A2(n32411), .ZN(n31622) );
  XNOR2HSV4 U37096 ( .A1(n31623), .A2(n31622), .ZN(n31635) );
  CLKNAND2HSV2 U37097 ( .A1(n31683), .A2(n31624), .ZN(n31629) );
  INHSV2 U37098 ( .I(n31684), .ZN(n31626) );
  CLKNAND2HSV1 U37099 ( .A1(n31629), .A2(n31626), .ZN(n31633) );
  INHSV2 U37100 ( .I(n36050), .ZN(n36083) );
  NAND3HSV2 U37101 ( .A1(n31628), .A2(n31627), .A3(n36083), .ZN(n31681) );
  INHSV2 U37102 ( .I(n31630), .ZN(n31632) );
  AND2HSV2 U37103 ( .A1(n31673), .A2(n46574), .Z(n31631) );
  NAND3HSV4 U37104 ( .A1(n31633), .A2(n31632), .A3(n31631), .ZN(n31634) );
  XNOR2HSV4 U37105 ( .A1(n31635), .A2(n31634), .ZN(n51437) );
  NOR2HSV4 U37106 ( .A1(n51437), .A2(n31636), .ZN(n31748) );
  CLKAND2HSV2 U37107 ( .A1(n44369), .A2(\pe6/ti_7t [8]), .Z(n31637) );
  NOR2HSV4 U37108 ( .A1(n31748), .A2(n31637), .ZN(n31754) );
  INHSV3 U37109 ( .I(n31754), .ZN(n31641) );
  CLKNAND2HSV2 U37110 ( .A1(n51437), .A2(n31690), .ZN(n31640) );
  NOR2HSV2 U37111 ( .A1(n48000), .A2(n36066), .ZN(n31639) );
  NOR2HSV4 U37112 ( .A1(n31639), .A2(n31640), .ZN(n31753) );
  NOR2HSV4 U37113 ( .A1(n31641), .A2(n31753), .ZN(n31705) );
  INHSV4 U37114 ( .I(n31705), .ZN(n31768) );
  NAND2HSV2 U37115 ( .A1(n31768), .A2(n46155), .ZN(n31642) );
  XNOR2HSV4 U37116 ( .A1(n31643), .A2(n31642), .ZN(n31700) );
  CLKNAND2HSV1 U37117 ( .A1(n31949), .A2(n31590), .ZN(n31666) );
  INAND2HSV2 U37118 ( .A1(n35817), .B1(n31644), .ZN(n32372) );
  NAND2HSV2 U37119 ( .A1(n32198), .A2(\pe6/pvq [9]), .ZN(n31645) );
  XOR2HSV0 U37120 ( .A1(n32372), .A2(n31645), .Z(n31649) );
  NAND2HSV2 U37121 ( .A1(n48035), .A2(n31910), .ZN(n31647) );
  CLKNAND2HSV0 U37122 ( .A1(n46624), .A2(n59278), .ZN(n31646) );
  XOR2HSV0 U37123 ( .A1(n31647), .A2(n31646), .Z(n31648) );
  XOR2HSV0 U37124 ( .A1(n31649), .A2(n31648), .Z(n31662) );
  INHSV2 U37125 ( .I(n50837), .ZN(n59074) );
  NAND2HSV2 U37126 ( .A1(n59259), .A2(n59074), .ZN(n31651) );
  CLKNAND2HSV0 U37127 ( .A1(n31776), .A2(n31785), .ZN(n31650) );
  XOR2HSV0 U37128 ( .A1(n31651), .A2(n31650), .Z(n31655) );
  CLKNAND2HSV1 U37129 ( .A1(n46135), .A2(n46643), .ZN(n31653) );
  CLKNAND2HSV0 U37130 ( .A1(\pe6/bq[24] ), .A2(n59276), .ZN(n31652) );
  XOR2HSV0 U37131 ( .A1(n31653), .A2(n31652), .Z(n31654) );
  XOR2HSV0 U37132 ( .A1(n31655), .A2(n31654), .Z(n31661) );
  BUFHSV2 U37133 ( .I(n46620), .Z(n36124) );
  NOR2HSV2 U37134 ( .A1(n36124), .A2(n32589), .ZN(n31657) );
  INHSV2 U37135 ( .I(n46663), .ZN(n31932) );
  CLKNAND2HSV0 U37136 ( .A1(n59261), .A2(n31932), .ZN(n31656) );
  CLKNAND2HSV1 U37137 ( .A1(n59236), .A2(n31717), .ZN(n31658) );
  XOR2HSV0 U37138 ( .A1(n31658), .A2(\pe6/phq [9]), .Z(n31659) );
  CLKNAND2HSV1 U37139 ( .A1(n31944), .A2(n36101), .ZN(n31663) );
  XNOR2HSV1 U37140 ( .A1(n31664), .A2(n31663), .ZN(n31665) );
  XNOR2HSV4 U37141 ( .A1(n31666), .A2(n31665), .ZN(n31669) );
  NAND2HSV2 U37142 ( .A1(n48004), .A2(n31670), .ZN(n31671) );
  CLKNAND2HSV2 U37143 ( .A1(n31672), .A2(n31671), .ZN(n31675) );
  CLKNAND2HSV1 U37144 ( .A1(n31673), .A2(n35808), .ZN(n31674) );
  INHSV2 U37145 ( .I(n31676), .ZN(n31694) );
  CLKNHSV0 U37146 ( .I(n31681), .ZN(n31682) );
  NAND2HSV2 U37147 ( .A1(n31682), .A2(n59011), .ZN(n31689) );
  BUFHSV2 U37148 ( .I(n31683), .Z(n35668) );
  NOR2HSV2 U37149 ( .A1(n31684), .A2(n35668), .ZN(n31687) );
  OR2HSV1 U37150 ( .A1(n31685), .A2(n36050), .Z(n31686) );
  NOR2HSV2 U37151 ( .A1(n31687), .A2(n31686), .ZN(n31688) );
  INHSV1 U37152 ( .I(\pe6/ti_7t [7]), .ZN(n31691) );
  AOI21HSV2 U37153 ( .A1(n31691), .A2(n32057), .B(n32239), .ZN(n31692) );
  INHSV2 U37154 ( .I(n31757), .ZN(n31763) );
  NAND3HSV2 U37155 ( .A1(n31768), .A2(n31762), .A3(n33089), .ZN(n31697) );
  NOR2HSV2 U37156 ( .A1(n31817), .A2(\pe6/ti_7t [9]), .ZN(n31746) );
  INHSV1 U37157 ( .I(n31746), .ZN(n31695) );
  CLKAND2HSV2 U37158 ( .A1(n31695), .A2(n59339), .Z(n31696) );
  CLKNAND2HSV2 U37159 ( .A1(n31697), .A2(n31696), .ZN(n31698) );
  AOI21HSV4 U37160 ( .A1(n31699), .A2(n31765), .B(n31698), .ZN(n31701) );
  NAND2HSV2 U37161 ( .A1(n31700), .A2(n31701), .ZN(n31704) );
  INHSV2 U37162 ( .I(n31700), .ZN(n31703) );
  INHSV2 U37163 ( .I(n31701), .ZN(n31702) );
  CLKNHSV0 U37164 ( .I(n31706), .ZN(n31708) );
  AOI21HSV2 U37165 ( .A1(n31706), .A2(n32329), .B(n31373), .ZN(n31707) );
  NAND2HSV2 U37166 ( .A1(n59595), .A2(\pe6/got [28]), .ZN(n31742) );
  BUFHSV2 U37167 ( .I(n32697), .Z(n59594) );
  NAND2HSV2 U37168 ( .A1(n59594), .A2(n36101), .ZN(n31740) );
  CLKNAND2HSV1 U37169 ( .A1(n31944), .A2(n31710), .ZN(n31737) );
  NAND2HSV2 U37170 ( .A1(n32198), .A2(\pe6/pvq [10]), .ZN(n31716) );
  INHSV2 U37171 ( .I(n49315), .ZN(n49002) );
  NAND2HSV2 U37172 ( .A1(n33016), .A2(n49002), .ZN(n31711) );
  XNOR2HSV1 U37173 ( .A1(n31711), .A2(\pe6/phq [10]), .ZN(n31715) );
  CLKNAND2HSV1 U37174 ( .A1(n46135), .A2(n59061), .ZN(n31713) );
  INHSV2 U37175 ( .I(n50837), .ZN(n31909) );
  CLKNAND2HSV0 U37176 ( .A1(n32992), .A2(n31909), .ZN(n31712) );
  XOR2HSV0 U37177 ( .A1(n31713), .A2(n31712), .Z(n31714) );
  XOR3HSV2 U37178 ( .A1(n31716), .A2(n31715), .A3(n31714), .Z(n31735) );
  NAND2HSV2 U37179 ( .A1(n31454), .A2(n31717), .ZN(n31734) );
  NAND2HSV2 U37180 ( .A1(n35743), .A2(\pe6/aot [23]), .ZN(n31720) );
  CLKNAND2HSV0 U37181 ( .A1(n31718), .A2(n31785), .ZN(n31719) );
  XOR2HSV0 U37182 ( .A1(n31720), .A2(n31719), .Z(n31724) );
  CLKNAND2HSV0 U37183 ( .A1(n31820), .A2(n46643), .ZN(n31722) );
  CLKNAND2HSV0 U37184 ( .A1(n31831), .A2(n31829), .ZN(n31721) );
  XOR2HSV0 U37185 ( .A1(n31722), .A2(n31721), .Z(n31723) );
  XOR2HSV0 U37186 ( .A1(n31724), .A2(n31723), .Z(n31732) );
  CLKNAND2HSV1 U37187 ( .A1(n59206), .A2(n31910), .ZN(n31726) );
  INHSV2 U37188 ( .I(n59194), .ZN(n44453) );
  NAND2HSV0 U37189 ( .A1(n44453), .A2(n44446), .ZN(n31725) );
  XOR2HSV0 U37190 ( .A1(n31726), .A2(n31725), .Z(n31730) );
  CLKNAND2HSV0 U37191 ( .A1(n31830), .A2(n59276), .ZN(n31728) );
  CLKNAND2HSV1 U37192 ( .A1(n31776), .A2(n32605), .ZN(n31727) );
  XOR2HSV0 U37193 ( .A1(n31728), .A2(n31727), .Z(n31729) );
  XOR2HSV0 U37194 ( .A1(n31730), .A2(n31729), .Z(n31731) );
  XOR2HSV0 U37195 ( .A1(n31732), .A2(n31731), .Z(n31733) );
  XOR3HSV2 U37196 ( .A1(n31735), .A2(n31734), .A3(n31733), .Z(n31736) );
  XOR2HSV0 U37197 ( .A1(n31737), .A2(n31736), .Z(n31739) );
  CLKNAND2HSV1 U37198 ( .A1(n31949), .A2(n35789), .ZN(n31738) );
  XOR3HSV2 U37199 ( .A1(n31740), .A2(n31739), .A3(n31738), .Z(n31741) );
  NOR2HSV1 U37200 ( .A1(n31746), .A2(n46549), .ZN(n31747) );
  CLKNHSV0 U37201 ( .I(n31747), .ZN(n31749) );
  NOR3HSV2 U37202 ( .A1(n31753), .A2(n31749), .A3(n25868), .ZN(n31750) );
  INHSV2 U37203 ( .I(n31750), .ZN(n31751) );
  CLKNHSV0 U37204 ( .I(n31753), .ZN(n31756) );
  CLKAND2HSV2 U37205 ( .A1(n31754), .A2(n31461), .Z(n31755) );
  INHSV2 U37206 ( .I(n47996), .ZN(n31758) );
  OAI21HSV2 U37207 ( .A1(n52701), .A2(\pe6/ti_7t [11]), .B(n33063), .ZN(n31761) );
  CLKNHSV2 U37208 ( .I(n31761), .ZN(n31760) );
  NAND2HSV0 U37209 ( .A1(n31762), .A2(n31768), .ZN(n31875) );
  CLKNHSV2 U37210 ( .I(n31763), .ZN(n31764) );
  NAND2HSV2 U37211 ( .A1(\pe6/ti_7t [9]), .A2(n36023), .ZN(n31876) );
  CLKNHSV0 U37212 ( .I(n31876), .ZN(n31766) );
  OAI21HSV2 U37213 ( .A1(n31766), .A2(n52701), .B(n59168), .ZN(n31767) );
  BUFHSV8 U37214 ( .I(n31768), .Z(n31958) );
  NAND2HSV2 U37215 ( .A1(n46123), .A2(\pe6/got [28]), .ZN(n31811) );
  INHSV4 U37216 ( .I(n31769), .ZN(n31905) );
  CLKNAND2HSV2 U37217 ( .A1(n31769), .A2(n35789), .ZN(n31809) );
  CLKNAND2HSV1 U37218 ( .A1(n59594), .A2(n32970), .ZN(n31805) );
  CLKNAND2HSV0 U37219 ( .A1(n31454), .A2(n32009), .ZN(n31802) );
  CLKNAND2HSV1 U37220 ( .A1(n31990), .A2(\pe6/aot [22]), .ZN(n31771) );
  BUFHSV2 U37221 ( .I(n46620), .Z(n35653) );
  INHSV2 U37222 ( .I(n35653), .ZN(n32168) );
  CLKNAND2HSV0 U37223 ( .A1(n32168), .A2(n31909), .ZN(n31770) );
  XOR2HSV0 U37224 ( .A1(n31771), .A2(n31770), .Z(n31775) );
  BUFHSV2 U37225 ( .I(n31487), .Z(n32086) );
  NAND2HSV2 U37226 ( .A1(n32973), .A2(n31925), .ZN(n31773) );
  CLKNAND2HSV0 U37227 ( .A1(n31845), .A2(n31829), .ZN(n31772) );
  XOR2HSV0 U37228 ( .A1(n31773), .A2(n31772), .Z(n31774) );
  XOR2HSV0 U37229 ( .A1(n31775), .A2(n31774), .Z(n31784) );
  INHSV2 U37230 ( .I(\pe6/aot [21]), .ZN(n35864) );
  CLKNAND2HSV0 U37231 ( .A1(n59259), .A2(\pe6/aot [21]), .ZN(n31778) );
  NAND2HSV0 U37232 ( .A1(n31776), .A2(\pe6/aot [23]), .ZN(n31777) );
  XOR2HSV0 U37233 ( .A1(n31778), .A2(n31777), .Z(n31782) );
  CLKNAND2HSV0 U37234 ( .A1(n31830), .A2(n31910), .ZN(n31780) );
  INHSV2 U37235 ( .I(n59205), .ZN(n45813) );
  CLKNAND2HSV1 U37236 ( .A1(n45813), .A2(n59276), .ZN(n31779) );
  XOR2HSV0 U37237 ( .A1(n31780), .A2(n31779), .Z(n31781) );
  XOR2HSV0 U37238 ( .A1(n31782), .A2(n31781), .Z(n31783) );
  XOR2HSV0 U37239 ( .A1(n31784), .A2(n31783), .Z(n31799) );
  CLKNAND2HSV0 U37240 ( .A1(n31820), .A2(n31785), .ZN(n31787) );
  NAND2HSV0 U37241 ( .A1(n46135), .A2(n31932), .ZN(n31786) );
  XOR2HSV0 U37242 ( .A1(n31787), .A2(n31786), .Z(n31790) );
  XNOR2HSV1 U37243 ( .A1(n31788), .A2(\pe6/phq [12]), .ZN(n31789) );
  XNOR2HSV1 U37244 ( .A1(n31790), .A2(n31789), .ZN(n31797) );
  CLKNAND2HSV0 U37245 ( .A1(n59206), .A2(n59061), .ZN(n31828) );
  NAND2HSV2 U37246 ( .A1(n59206), .A2(n59065), .ZN(n32739) );
  OAI21HSV1 U37247 ( .A1(n46192), .A2(n32589), .B(n32739), .ZN(n31792) );
  OAI21HSV1 U37248 ( .A1(n31828), .A2(n31793), .B(n31792), .ZN(n31795) );
  CLKNAND2HSV1 U37249 ( .A1(n32198), .A2(\pe6/pvq [12]), .ZN(n31794) );
  XOR2HSV0 U37250 ( .A1(n31795), .A2(n31794), .Z(n31796) );
  XNOR2HSV1 U37251 ( .A1(n31797), .A2(n31796), .ZN(n31798) );
  XNOR2HSV1 U37252 ( .A1(n31799), .A2(n31798), .ZN(n31801) );
  NAND2HSV0 U37253 ( .A1(n31944), .A2(n59174), .ZN(n31800) );
  XOR3HSV2 U37254 ( .A1(n31802), .A2(n31801), .A3(n31800), .Z(n31804) );
  BUFHSV3 U37255 ( .I(n31949), .Z(n59121) );
  NAND2HSV2 U37256 ( .A1(n59121), .A2(n31861), .ZN(n31803) );
  XOR3HSV2 U37257 ( .A1(n31805), .A2(n31804), .A3(n31803), .Z(n31807) );
  NAND2HSV2 U37258 ( .A1(n59595), .A2(n36101), .ZN(n31806) );
  XNOR2HSV1 U37259 ( .A1(n31807), .A2(n31806), .ZN(n31808) );
  XNOR2HSV2 U37260 ( .A1(n31811), .A2(n31810), .ZN(n31812) );
  INHSV2 U37261 ( .I(n32463), .ZN(n32949) );
  NAND2HSV2 U37262 ( .A1(n32949), .A2(\pe6/ti_7t [10]), .ZN(n31901) );
  INHSV2 U37263 ( .I(n31901), .ZN(n31869) );
  CLKNHSV0 U37264 ( .I(\pe6/ti_7t [12]), .ZN(n31818) );
  NAND2HSV2 U37265 ( .A1(n46123), .A2(\pe6/got [27]), .ZN(n31867) );
  BUFHSV2 U37266 ( .I(\pe6/got [26]), .Z(n32354) );
  NAND2HSV0 U37267 ( .A1(n31769), .A2(n32354), .ZN(n31865) );
  NAND2HSV0 U37268 ( .A1(n31925), .A2(n31910), .ZN(n31822) );
  NAND2HSV0 U37269 ( .A1(n31820), .A2(n31932), .ZN(n31821) );
  XOR2HSV0 U37270 ( .A1(n31822), .A2(n31821), .Z(n31826) );
  CLKNAND2HSV1 U37271 ( .A1(n35740), .A2(n49831), .ZN(n31824) );
  INHSV2 U37272 ( .I(n35837), .ZN(n46137) );
  CLKNAND2HSV0 U37273 ( .A1(n46137), .A2(n59276), .ZN(n31823) );
  XOR2HSV0 U37274 ( .A1(n31824), .A2(n31823), .Z(n31825) );
  XOR2HSV0 U37275 ( .A1(n31826), .A2(n31825), .Z(n31837) );
  CLKNAND2HSV1 U37276 ( .A1(n31593), .A2(\pe6/pvq [13]), .ZN(n31827) );
  XOR2HSV0 U37277 ( .A1(n31828), .A2(n31827), .Z(n31835) );
  NAND2HSV0 U37278 ( .A1(n31830), .A2(n31829), .ZN(n31833) );
  CLKNHSV0 U37279 ( .I(n32079), .ZN(n31972) );
  NAND2HSV0 U37280 ( .A1(n31831), .A2(n31972), .ZN(n31832) );
  XOR2HSV0 U37281 ( .A1(n31833), .A2(n31832), .Z(n31834) );
  XOR2HSV0 U37282 ( .A1(n31835), .A2(n31834), .Z(n31836) );
  XOR2HSV0 U37283 ( .A1(n31837), .A2(n31836), .Z(n31854) );
  NAND2HSV2 U37284 ( .A1(n32172), .A2(n32973), .ZN(n31839) );
  NAND2HSV0 U37285 ( .A1(n46135), .A2(n31909), .ZN(n31838) );
  XOR2HSV0 U37286 ( .A1(n31839), .A2(n31838), .Z(n31843) );
  NAND2HSV2 U37287 ( .A1(n32168), .A2(\pe6/aot [23]), .ZN(n31841) );
  CLKNAND2HSV1 U37288 ( .A1(n31990), .A2(\pe6/aot [21]), .ZN(n31840) );
  XOR2HSV0 U37289 ( .A1(n31841), .A2(n31840), .Z(n31842) );
  XOR2HSV0 U37290 ( .A1(n31843), .A2(n31842), .Z(n31852) );
  NOR2HSV2 U37291 ( .A1(n31560), .A2(n35607), .ZN(n31847) );
  CLKNAND2HSV0 U37292 ( .A1(n31845), .A2(n32171), .ZN(n31846) );
  XOR2HSV0 U37293 ( .A1(n31847), .A2(n31846), .Z(n31850) );
  XOR2HSV0 U37294 ( .A1(n31848), .A2(\pe6/phq [13]), .Z(n31849) );
  XOR2HSV0 U37295 ( .A1(n31850), .A2(n31849), .Z(n31851) );
  XOR2HSV0 U37296 ( .A1(n31852), .A2(n31851), .Z(n31853) );
  XOR2HSV0 U37297 ( .A1(n31854), .A2(n31853), .Z(n31858) );
  CLKNAND2HSV0 U37298 ( .A1(n31944), .A2(n32009), .ZN(n31857) );
  CLKNAND2HSV0 U37299 ( .A1(n44426), .A2(n59328), .ZN(n31856) );
  CLKNAND2HSV1 U37300 ( .A1(n32384), .A2(n35812), .ZN(n31855) );
  XOR4HSV1 U37301 ( .A1(n31858), .A2(n31857), .A3(n31856), .A4(n31855), .Z(
        n31860) );
  CLKNAND2HSV1 U37302 ( .A1(n58940), .A2(n59165), .ZN(n31859) );
  XOR2HSV0 U37303 ( .A1(n31860), .A2(n31859), .Z(n31863) );
  NAND2HSV2 U37304 ( .A1(n35668), .A2(n31861), .ZN(n31862) );
  XNOR2HSV1 U37305 ( .A1(n31863), .A2(n31862), .ZN(n31864) );
  XNOR2HSV1 U37306 ( .A1(n31865), .A2(n31864), .ZN(n31866) );
  XNOR2HSV2 U37307 ( .A1(n31867), .A2(n31866), .ZN(n31868) );
  CLKNAND2HSV0 U37308 ( .A1(n32822), .A2(n32411), .ZN(n32444) );
  NAND2HSV0 U37309 ( .A1(n31869), .A2(n32647), .ZN(n31872) );
  NAND2HSV0 U37310 ( .A1(n31901), .A2(n47950), .ZN(n31884) );
  CLKNHSV0 U37311 ( .I(n31884), .ZN(n31870) );
  NOR2HSV0 U37312 ( .A1(n31870), .A2(n44376), .ZN(n31871) );
  NAND3HSV2 U37313 ( .A1(n31875), .A2(n31874), .A3(n32961), .ZN(n31877) );
  CLKNAND2HSV2 U37314 ( .A1(n31877), .A2(n31876), .ZN(n59673) );
  INHSV4 U37315 ( .I(n59673), .ZN(n31970) );
  NAND2HSV2 U37316 ( .A1(\pe6/ti_7t [11]), .A2(n32148), .ZN(n32133) );
  INOR2HSV1 U37317 ( .A1(n31884), .B1(n46159), .ZN(n31896) );
  NAND2HSV0 U37318 ( .A1(n31896), .A2(n32133), .ZN(n31885) );
  CLKNHSV0 U37319 ( .I(n31896), .ZN(n31886) );
  NAND2HSV0 U37320 ( .A1(n31886), .A2(n32133), .ZN(n31888) );
  INOR2HSV1 U37321 ( .A1(n32133), .B1(n32961), .ZN(n32024) );
  NOR2HSV0 U37322 ( .A1(n32024), .A2(n32530), .ZN(n31887) );
  AOI21HSV2 U37323 ( .A1(n31890), .A2(n31898), .B(n31889), .ZN(n31891) );
  CLKNHSV1 U37324 ( .I(n31893), .ZN(n35704) );
  BUFHSV2 U37325 ( .I(n47934), .Z(n32793) );
  INHSV2 U37326 ( .I(n46591), .ZN(n48018) );
  NAND2HSV2 U37327 ( .A1(\pe6/ti_7t [13]), .A2(n48018), .ZN(n32052) );
  BUFHSV2 U37328 ( .I(n32052), .Z(n32059) );
  INHSV2 U37329 ( .I(n51445), .ZN(n31894) );
  NAND2HSV2 U37330 ( .A1(\pe6/ti_7t [12]), .A2(n32148), .ZN(n32060) );
  CLKNHSV0 U37331 ( .I(n32060), .ZN(n32029) );
  CLKNHSV0 U37332 ( .I(n35917), .ZN(n46574) );
  CLKNAND2HSV1 U37333 ( .A1(n32029), .A2(n46574), .ZN(n31895) );
  NOR2HSV1 U37334 ( .A1(n32024), .A2(n44376), .ZN(n31899) );
  NAND2HSV2 U37335 ( .A1(n59596), .A2(n31902), .ZN(n31964) );
  INHSV1 U37336 ( .I(n31903), .ZN(n59166) );
  CLKNHSV0 U37337 ( .I(n31590), .ZN(n31904) );
  NAND2HSV2 U37338 ( .A1(n32218), .A2(n32354), .ZN(n31957) );
  INHSV3 U37339 ( .I(n31905), .ZN(n32167) );
  NAND2HSV2 U37340 ( .A1(n32167), .A2(\pe6/got [25]), .ZN(n31955) );
  CLKNHSV0 U37341 ( .I(n59194), .ZN(n32173) );
  NAND2HSV0 U37342 ( .A1(n32173), .A2(n46662), .ZN(n31907) );
  CLKNHSV0 U37343 ( .I(n32068), .ZN(n32276) );
  INHSV2 U37344 ( .I(n35816), .ZN(n32171) );
  CLKNAND2HSV1 U37345 ( .A1(n32276), .A2(n32171), .ZN(n31906) );
  XOR2HSV0 U37346 ( .A1(n31907), .A2(n31906), .Z(n31914) );
  CLKNHSV0 U37347 ( .I(n31908), .ZN(n45812) );
  NAND2HSV0 U37348 ( .A1(n45812), .A2(n31909), .ZN(n31912) );
  NAND2HSV0 U37349 ( .A1(n32172), .A2(n31910), .ZN(n31911) );
  XOR2HSV0 U37350 ( .A1(n31912), .A2(n31911), .Z(n31913) );
  XOR2HSV0 U37351 ( .A1(n31914), .A2(n31913), .Z(n31921) );
  NOR2HSV0 U37352 ( .A1(n44411), .A2(n35607), .ZN(n31916) );
  NAND2HSV0 U37353 ( .A1(n46135), .A2(\pe6/aot [23]), .ZN(n31915) );
  XOR2HSV0 U37354 ( .A1(n31916), .A2(n31915), .Z(n31919) );
  INHSV2 U37355 ( .I(\pe6/got [19]), .ZN(n44494) );
  INHSV2 U37356 ( .I(n44494), .ZN(n49096) );
  CLKNAND2HSV0 U37357 ( .A1(n59236), .A2(n49096), .ZN(n31917) );
  XOR2HSV0 U37358 ( .A1(n31917), .A2(\pe6/phq [14]), .Z(n31918) );
  XOR2HSV0 U37359 ( .A1(n31919), .A2(n31918), .Z(n31920) );
  XOR2HSV0 U37360 ( .A1(n31921), .A2(n31920), .Z(n31923) );
  INHSV2 U37361 ( .I(n32125), .ZN(n32563) );
  NAND2HSV0 U37362 ( .A1(n31454), .A2(n32563), .ZN(n31922) );
  XNOR2HSV1 U37363 ( .A1(n31923), .A2(n31922), .ZN(n31943) );
  BUFHSV2 U37364 ( .I(n31924), .Z(n32266) );
  INHSV2 U37365 ( .I(n32266), .ZN(n59234) );
  CLKNAND2HSV0 U37366 ( .A1(n31925), .A2(n59234), .ZN(n31927) );
  INHSV2 U37367 ( .I(n31560), .ZN(n59259) );
  NAND2HSV2 U37368 ( .A1(n59259), .A2(\pe6/aot [19]), .ZN(n31926) );
  XOR2HSV0 U37369 ( .A1(n31927), .A2(n31926), .Z(n31941) );
  INHSV2 U37370 ( .I(n44397), .ZN(n50829) );
  CLKNAND2HSV1 U37371 ( .A1(n50829), .A2(n33004), .ZN(n32744) );
  OAI22HSV0 U37372 ( .A1(n31253), .A2(n44397), .B1(n31928), .B2(n32373), .ZN(
        n31929) );
  OAI21HSV0 U37373 ( .A1(n33019), .A2(n32744), .B(n31929), .ZN(n31931) );
  CLKNAND2HSV0 U37374 ( .A1(n48036), .A2(\pe6/pvq [14]), .ZN(n31930) );
  XNOR2HSV1 U37375 ( .A1(n31931), .A2(n31930), .ZN(n31940) );
  NAND2HSV0 U37376 ( .A1(n48035), .A2(n31932), .ZN(n31934) );
  NAND2HSV0 U37377 ( .A1(n59206), .A2(n31972), .ZN(n31933) );
  XOR2HSV0 U37378 ( .A1(n31934), .A2(n31933), .Z(n31938) );
  CLKNHSV0 U37379 ( .I(n31425), .ZN(n59071) );
  CLKNAND2HSV1 U37380 ( .A1(n59071), .A2(\pe6/aot [21]), .ZN(n31936) );
  NAND2HSV0 U37381 ( .A1(n46137), .A2(n36114), .ZN(n31935) );
  XOR2HSV0 U37382 ( .A1(n31936), .A2(n31935), .Z(n31937) );
  XOR2HSV0 U37383 ( .A1(n31938), .A2(n31937), .Z(n31939) );
  XOR3HSV2 U37384 ( .A1(n31941), .A2(n31940), .A3(n31939), .Z(n31942) );
  XNOR2HSV1 U37385 ( .A1(n31943), .A2(n31942), .ZN(n31946) );
  BUFHSV2 U37386 ( .I(n31944), .Z(n32286) );
  CLKNAND2HSV1 U37387 ( .A1(n32286), .A2(n59328), .ZN(n31945) );
  XOR2HSV0 U37388 ( .A1(n31946), .A2(n31945), .Z(n31948) );
  NAND2HSV0 U37389 ( .A1(n59594), .A2(n32009), .ZN(n31947) );
  XNOR2HSV1 U37390 ( .A1(n31948), .A2(n31947), .ZN(n31951) );
  BUFHSV3 U37391 ( .I(n31949), .Z(n59670) );
  CLKNAND2HSV1 U37392 ( .A1(n59670), .A2(n35812), .ZN(n31950) );
  CLKNAND2HSV1 U37393 ( .A1(n32293), .A2(n31717), .ZN(n31952) );
  XNOR2HSV1 U37394 ( .A1(n31953), .A2(n31952), .ZN(n31954) );
  XNOR2HSV1 U37395 ( .A1(n31957), .A2(n31956), .ZN(n31960) );
  BUFHSV2 U37396 ( .I(\pe6/got [27]), .Z(n49665) );
  XNOR2HSV1 U37397 ( .A1(n31960), .A2(n31959), .ZN(n31961) );
  XNOR2HSV4 U37398 ( .A1(n31962), .A2(n31961), .ZN(n31963) );
  MUX2NHSV4 U37399 ( .I0(n31964), .I1(n29665), .S(n31963), .ZN(n31965) );
  XNOR2HSV4 U37400 ( .A1(n31966), .A2(n31965), .ZN(n32042) );
  XNOR2HSV4 U37401 ( .A1(n31967), .A2(n32042), .ZN(n32146) );
  INHSV2 U37402 ( .I(n32146), .ZN(n31968) );
  INHSV2 U37403 ( .I(n31968), .ZN(n31969) );
  CLKNAND2HSV1 U37404 ( .A1(n32218), .A2(\pe6/got [25]), .ZN(n32017) );
  CLKNAND2HSV1 U37405 ( .A1(n32167), .A2(n32970), .ZN(n32015) );
  NAND2HSV0 U37406 ( .A1(n46137), .A2(n32991), .ZN(n31974) );
  NAND2HSV0 U37407 ( .A1(n32173), .A2(n31972), .ZN(n31973) );
  XOR2HSV0 U37408 ( .A1(n31974), .A2(n31973), .Z(n31978) );
  CLKNAND2HSV1 U37409 ( .A1(n59259), .A2(n32573), .ZN(n31976) );
  NAND2HSV0 U37410 ( .A1(n59206), .A2(n32605), .ZN(n31975) );
  XOR2HSV0 U37411 ( .A1(n31976), .A2(n31975), .Z(n31977) );
  XOR2HSV0 U37412 ( .A1(n31978), .A2(n31977), .Z(n31987) );
  NAND2HSV0 U37413 ( .A1(n32276), .A2(n46662), .ZN(n31981) );
  CLKNHSV0 U37414 ( .I(n31979), .ZN(n44700) );
  CLKNAND2HSV0 U37415 ( .A1(n44700), .A2(n32171), .ZN(n31980) );
  XOR2HSV0 U37416 ( .A1(n31981), .A2(n31980), .Z(n31985) );
  CLKNAND2HSV0 U37417 ( .A1(n45812), .A2(\pe6/aot [23]), .ZN(n31983) );
  CLKNHSV0 U37418 ( .I(\pe6/bq[28] ), .ZN(n36123) );
  INHSV1 U37419 ( .I(n36123), .ZN(n32999) );
  NAND2HSV0 U37420 ( .A1(n32999), .A2(\pe6/aot [22]), .ZN(n31982) );
  XOR2HSV0 U37421 ( .A1(n31983), .A2(n31982), .Z(n31984) );
  XOR2HSV0 U37422 ( .A1(n31985), .A2(n31984), .Z(n31986) );
  XOR2HSV0 U37423 ( .A1(n31987), .A2(n31986), .Z(n31989) );
  CLKNHSV1 U37424 ( .I(n52706), .ZN(n35612) );
  INHSV2 U37425 ( .I(\pe6/got [19]), .ZN(n32696) );
  CLKNAND2HSV0 U37426 ( .A1(n35612), .A2(n49096), .ZN(n31988) );
  XNOR2HSV1 U37427 ( .A1(n31989), .A2(n31988), .ZN(n32004) );
  NAND2HSV0 U37428 ( .A1(n31990), .A2(\pe6/aot [19]), .ZN(n32271) );
  NAND2HSV0 U37429 ( .A1(\pe6/bq[18] ), .A2(n59276), .ZN(n32590) );
  XOR2HSV0 U37430 ( .A1(n32271), .A2(n32590), .Z(n32002) );
  NAND2HSV0 U37431 ( .A1(n32252), .A2(n59239), .ZN(n31992) );
  INHSV2 U37432 ( .I(n44397), .ZN(n32486) );
  NAND2HSV0 U37433 ( .A1(n32486), .A2(n32973), .ZN(n31991) );
  XOR2HSV0 U37434 ( .A1(n31992), .A2(n31991), .Z(n31995) );
  XNOR2HSV1 U37435 ( .A1(n31993), .A2(\pe6/phq [15]), .ZN(n31994) );
  XNOR2HSV1 U37436 ( .A1(n31995), .A2(n31994), .ZN(n32001) );
  NOR2HSV2 U37437 ( .A1(n32484), .A2(n35607), .ZN(n35609) );
  CLKNAND2HSV0 U37438 ( .A1(n32172), .A2(n59234), .ZN(n32268) );
  XOR2HSV0 U37439 ( .A1(n35609), .A2(n32268), .Z(n31999) );
  NAND2HSV0 U37440 ( .A1(n59201), .A2(\pe6/pvq [15]), .ZN(n31997) );
  NAND2HSV0 U37441 ( .A1(n32168), .A2(\pe6/aot [21]), .ZN(n31996) );
  XOR2HSV0 U37442 ( .A1(n31997), .A2(n31996), .Z(n31998) );
  XOR2HSV0 U37443 ( .A1(n31999), .A2(n31998), .Z(n32000) );
  XOR3HSV2 U37444 ( .A1(n32002), .A2(n32001), .A3(n32000), .Z(n32003) );
  XNOR2HSV1 U37445 ( .A1(n32004), .A2(n32003), .ZN(n32006) );
  CLKNAND2HSV0 U37446 ( .A1(n32286), .A2(n32563), .ZN(n32005) );
  XNOR2HSV1 U37447 ( .A1(n32006), .A2(n32005), .ZN(n32008) );
  NAND2HSV0 U37448 ( .A1(n32384), .A2(n59328), .ZN(n32007) );
  XNOR2HSV1 U37449 ( .A1(n32008), .A2(n32007), .ZN(n32011) );
  CLKNAND2HSV0 U37450 ( .A1(n59670), .A2(n32009), .ZN(n32010) );
  XOR2HSV0 U37451 ( .A1(n32011), .A2(n32010), .Z(n32013) );
  CLKNAND2HSV1 U37452 ( .A1(n32293), .A2(n59174), .ZN(n32012) );
  XNOR2HSV1 U37453 ( .A1(n32013), .A2(n32012), .ZN(n32014) );
  XNOR2HSV1 U37454 ( .A1(n32015), .A2(n32014), .ZN(n32016) );
  XNOR2HSV1 U37455 ( .A1(n32017), .A2(n32016), .ZN(n32019) );
  CLKNAND2HSV1 U37456 ( .A1(n44476), .A2(n32354), .ZN(n32018) );
  XNOR2HSV1 U37457 ( .A1(n32019), .A2(n32018), .ZN(n32020) );
  BUFHSV2 U37458 ( .I(n32466), .Z(n32640) );
  CLKNAND2HSV1 U37459 ( .A1(n59596), .A2(n33061), .ZN(n32022) );
  XOR2HSV2 U37460 ( .A1(n32023), .A2(n32022), .Z(n32028) );
  CLKNHSV0 U37461 ( .I(n32024), .ZN(n32025) );
  XNOR2HSV4 U37462 ( .A1(n32028), .A2(n32027), .ZN(n32032) );
  OAI21HSV1 U37463 ( .A1(n32029), .A2(n35797), .B(n32647), .ZN(n32030) );
  AOI21HSV1 U37464 ( .A1(n51445), .A2(n32060), .B(n32030), .ZN(n32031) );
  XNOR2HSV4 U37465 ( .A1(n32032), .A2(n32031), .ZN(n32050) );
  INHSV2 U37466 ( .I(n32033), .ZN(n32038) );
  OAI21HSV1 U37467 ( .A1(n47934), .A2(\pe6/ti_7t [13]), .B(n46567), .ZN(n32034) );
  AOI21HSV4 U37468 ( .A1(n29646), .A2(n32038), .B(n32034), .ZN(n32040) );
  CLKNHSV2 U37469 ( .I(n32035), .ZN(n32036) );
  CLKNAND2HSV4 U37470 ( .A1(n32040), .A2(n32039), .ZN(n32049) );
  XNOR2HSV4 U37471 ( .A1(n32042), .A2(n32041), .ZN(n32325) );
  NOR2HSV0 U37472 ( .A1(n35797), .A2(\pe6/ti_7t [14]), .ZN(n32043) );
  NOR2HSV2 U37473 ( .A1(n32043), .A2(n51438), .ZN(n32145) );
  INHSV2 U37474 ( .I(n32145), .ZN(n47973) );
  NOR2HSV2 U37475 ( .A1(n47973), .A2(n33079), .ZN(n32315) );
  CLKNHSV0 U37476 ( .I(n32315), .ZN(n32045) );
  NOR2HSV2 U37477 ( .A1(n32146), .A2(n47973), .ZN(n32046) );
  CLKNAND2HSV1 U37478 ( .A1(n32046), .A2(n32159), .ZN(n32048) );
  NAND2HSV0 U37479 ( .A1(n32145), .A2(n32157), .ZN(n32051) );
  NAND2HSV2 U37480 ( .A1(n31350), .A2(\pe6/ti_7t [15]), .ZN(n32152) );
  BUFHSV2 U37481 ( .I(n32152), .Z(n32513) );
  NAND3HSV2 U37482 ( .A1(n32155), .A2(n32512), .A3(n32513), .ZN(n32345) );
  BUFHSV2 U37483 ( .I(n32345), .Z(n35898) );
  NAND2HSV2 U37484 ( .A1(n35898), .A2(n49665), .ZN(n32144) );
  INHSV2 U37485 ( .I(n32052), .ZN(n32163) );
  CLKNAND2HSV0 U37486 ( .A1(n32052), .A2(n48018), .ZN(n32054) );
  AND2HSV2 U37487 ( .A1(n32054), .A2(n32783), .Z(n32055) );
  CLKNHSV2 U37488 ( .I(\pe6/ti_7t [14]), .ZN(n32058) );
  MUX2NHSV4 U37489 ( .I0(n52765), .I1(n32058), .S(n32057), .ZN(n59914) );
  NAND2HSV2 U37490 ( .A1(n32059), .A2(n32157), .ZN(n44391) );
  CLKNAND2HSV0 U37491 ( .A1(n44391), .A2(n31861), .ZN(n32140) );
  OAI21HSV2 U37492 ( .A1(n51445), .A2(n35704), .B(n32060), .ZN(n32353) );
  INHSV2 U37493 ( .I(n32353), .ZN(n32061) );
  CLKNAND2HSV1 U37494 ( .A1(n59034), .A2(n32970), .ZN(n32138) );
  BUFHSV2 U37495 ( .I(n26109), .Z(n58939) );
  CLKNAND2HSV0 U37496 ( .A1(n58939), .A2(n59328), .ZN(n32129) );
  NAND2HSV0 U37497 ( .A1(n32841), .A2(n49096), .ZN(n32124) );
  NAND2HSV0 U37498 ( .A1(n35813), .A2(\pe6/got [18]), .ZN(n32122) );
  CLKNAND2HSV0 U37499 ( .A1(n32286), .A2(n35991), .ZN(n32116) );
  BUFHSV2 U37500 ( .I(n32384), .Z(n36108) );
  CLKNAND2HSV0 U37501 ( .A1(n36108), .A2(\pe6/got [15]), .ZN(n32115) );
  NAND2HSV0 U37502 ( .A1(n46624), .A2(\pe6/aot [19]), .ZN(n32063) );
  NAND2HSV0 U37503 ( .A1(n46672), .A2(n58943), .ZN(n32062) );
  XOR2HSV0 U37504 ( .A1(n32063), .A2(n32062), .Z(n32067) );
  CLKNHSV0 U37505 ( .I(\pe6/bq[27] ), .ZN(n35647) );
  INHSV2 U37506 ( .I(\pe6/aot [17]), .ZN(n58851) );
  NAND2HSV0 U37507 ( .A1(n59267), .A2(\pe6/aot [17]), .ZN(n32065) );
  CLKNHSV0 U37508 ( .I(\pe6/bq[22] ), .ZN(n50822) );
  INHSV2 U37509 ( .I(n50822), .ZN(n32886) );
  NAND2HSV0 U37510 ( .A1(n32886), .A2(n33004), .ZN(n32064) );
  XOR2HSV0 U37511 ( .A1(n32065), .A2(n32064), .Z(n32066) );
  XOR2HSV0 U37512 ( .A1(n32067), .A2(n32066), .Z(n32076) );
  BUFHSV2 U37513 ( .I(n35631), .Z(n32269) );
  INHSV2 U37514 ( .I(\pe6/aot [13]), .ZN(n58983) );
  CLKNAND2HSV0 U37515 ( .A1(n32992), .A2(\pe6/aot [13]), .ZN(n32070) );
  CLKNHSV0 U37516 ( .I(n32068), .ZN(n44702) );
  NAND2HSV0 U37517 ( .A1(n44702), .A2(\pe6/aot [21]), .ZN(n32069) );
  XOR2HSV0 U37518 ( .A1(n32070), .A2(n32069), .Z(n32074) );
  CLKNAND2HSV1 U37519 ( .A1(n36161), .A2(\pe6/pvq [21]), .ZN(n32072) );
  CLKNHSV0 U37520 ( .I(n44397), .ZN(n35761) );
  CLKNHSV0 U37521 ( .I(n46663), .ZN(n59245) );
  NAND2HSV0 U37522 ( .A1(n35761), .A2(n59245), .ZN(n32071) );
  XOR2HSV0 U37523 ( .A1(n32072), .A2(n32071), .Z(n32073) );
  XOR2HSV0 U37524 ( .A1(n32074), .A2(n32073), .Z(n32075) );
  XOR2HSV0 U37525 ( .A1(n32076), .A2(n32075), .Z(n32078) );
  NAND2HSV0 U37526 ( .A1(n35612), .A2(n58654), .ZN(n32077) );
  XNOR2HSV1 U37527 ( .A1(n32078), .A2(n32077), .ZN(n32113) );
  INHSV2 U37528 ( .I(\pe6/bq[16] ), .ZN(n32732) );
  INHSV2 U37529 ( .I(n32732), .ZN(n32567) );
  NAND2HSV0 U37530 ( .A1(n32567), .A2(n58991), .ZN(n32081) );
  BUFHSV3 U37531 ( .I(n32079), .Z(n32976) );
  CLKNHSV1 U37532 ( .I(n32976), .ZN(n32876) );
  NAND2HSV0 U37533 ( .A1(n33023), .A2(n32876), .ZN(n32080) );
  XOR2HSV0 U37534 ( .A1(n32081), .A2(n32080), .Z(n32085) );
  NAND2HSV0 U37535 ( .A1(n33005), .A2(n33022), .ZN(n32083) );
  CLKNHSV0 U37536 ( .I(n32245), .ZN(n35726) );
  NAND2HSV0 U37537 ( .A1(n32252), .A2(n35726), .ZN(n32082) );
  XOR2HSV0 U37538 ( .A1(n32083), .A2(n32082), .Z(n32084) );
  XOR2HSV0 U37539 ( .A1(n32085), .A2(n32084), .Z(n32094) );
  NAND2HSV0 U37540 ( .A1(n32568), .A2(n36153), .ZN(n32088) );
  INHSV2 U37541 ( .I(n46853), .ZN(n33000) );
  NAND2HSV0 U37542 ( .A1(n33000), .A2(n36114), .ZN(n32087) );
  XOR2HSV0 U37543 ( .A1(n32088), .A2(n32087), .Z(n32092) );
  NAND2HSV0 U37544 ( .A1(\pe6/bq[14] ), .A2(n35925), .ZN(n32090) );
  INHSV2 U37545 ( .I(n44396), .ZN(n33024) );
  NAND2HSV0 U37546 ( .A1(n35768), .A2(n33024), .ZN(n32089) );
  XOR2HSV0 U37547 ( .A1(n32090), .A2(n32089), .Z(n32091) );
  XOR2HSV0 U37548 ( .A1(n32092), .A2(n32091), .Z(n32093) );
  XOR2HSV0 U37549 ( .A1(n32094), .A2(n32093), .Z(n32111) );
  NOR2HSV0 U37550 ( .A1(n59194), .A2(n35607), .ZN(n32096) );
  CLKNHSV0 U37551 ( .I(n32589), .ZN(n32981) );
  NAND2HSV0 U37552 ( .A1(n32982), .A2(n32981), .ZN(n32095) );
  XOR2HSV0 U37553 ( .A1(n32096), .A2(n32095), .Z(n32099) );
  NAND2HSV0 U37554 ( .A1(n33016), .A2(n33039), .ZN(n32097) );
  XOR2HSV0 U37555 ( .A1(n32097), .A2(\pe6/phq [21]), .Z(n32098) );
  XOR2HSV0 U37556 ( .A1(n32099), .A2(n32098), .Z(n32109) );
  OAI22HSV0 U37557 ( .A1(n31560), .A2(n49188), .B1(n48047), .B2(n35817), .ZN(
        n32103) );
  NAND2HSV0 U37558 ( .A1(n59045), .A2(\pe6/aot [12]), .ZN(n50846) );
  CLKNHSV1 U37559 ( .I(n50846), .ZN(n32100) );
  NAND2HSV0 U37560 ( .A1(n32101), .A2(n32100), .ZN(n32102) );
  CLKNAND2HSV1 U37561 ( .A1(n32103), .A2(n32102), .ZN(n32107) );
  INHSV2 U37562 ( .I(n46789), .ZN(n59044) );
  NAND2HSV0 U37563 ( .A1(n48051), .A2(n59044), .ZN(n58866) );
  INHSV2 U37564 ( .I(n46789), .ZN(n59189) );
  NAND2HSV0 U37565 ( .A1(n32999), .A2(n59189), .ZN(n46646) );
  OAI21HSV0 U37566 ( .A1(n31253), .A2(n59094), .B(n46646), .ZN(n32104) );
  OAI21HSV0 U37567 ( .A1(n32105), .A2(n58866), .B(n32104), .ZN(n32106) );
  XOR2HSV0 U37568 ( .A1(n32107), .A2(n32106), .Z(n32108) );
  XOR2HSV0 U37569 ( .A1(n32109), .A2(n32108), .Z(n32110) );
  XNOR2HSV1 U37570 ( .A1(n32111), .A2(n32110), .ZN(n32112) );
  XOR2HSV0 U37571 ( .A1(n32113), .A2(n32112), .Z(n32114) );
  XOR3HSV2 U37572 ( .A1(n32116), .A2(n32115), .A3(n32114), .Z(n32118) );
  BUFHSV2 U37573 ( .I(n59121), .Z(n32900) );
  NAND2HSV0 U37574 ( .A1(n32900), .A2(n46171), .ZN(n32117) );
  XNOR2HSV1 U37575 ( .A1(n32118), .A2(n32117), .ZN(n32120) );
  INHSV2 U37576 ( .I(n53103), .ZN(n32971) );
  NAND2HSV0 U37577 ( .A1(n36183), .A2(n32971), .ZN(n32119) );
  XNOR2HSV1 U37578 ( .A1(n32120), .A2(n32119), .ZN(n32121) );
  XNOR2HSV1 U37579 ( .A1(n32122), .A2(n32121), .ZN(n32123) );
  XNOR2HSV1 U37580 ( .A1(n32124), .A2(n32123), .ZN(n32127) );
  CLKBUFHSV4 U37581 ( .I(n44476), .Z(n36185) );
  CLKNAND2HSV0 U37582 ( .A1(n36185), .A2(\pe6/got [20]), .ZN(n32126) );
  XNOR2HSV1 U37583 ( .A1(n32127), .A2(n32126), .ZN(n32128) );
  CLKNHSV2 U37584 ( .I(n59596), .ZN(n32130) );
  CLKNAND2HSV0 U37585 ( .A1(n32165), .A2(\pe6/got [22]), .ZN(n32131) );
  XNOR2HSV1 U37586 ( .A1(n32132), .A2(n32131), .ZN(n32136) );
  BUFHSV2 U37587 ( .I(n32133), .Z(n32134) );
  INHSV2 U37588 ( .I(n32306), .ZN(n32506) );
  XNOR2HSV1 U37589 ( .A1(n32136), .A2(n32135), .ZN(n32137) );
  XOR2HSV0 U37590 ( .A1(n32138), .A2(n32137), .Z(n32139) );
  XNOR2HSV1 U37591 ( .A1(n32140), .A2(n32139), .ZN(n32141) );
  XOR2HSV0 U37592 ( .A1(n32142), .A2(n32141), .Z(n32143) );
  XOR2HSV2 U37593 ( .A1(n32144), .A2(n32143), .Z(n32237) );
  NAND2HSV2 U37594 ( .A1(n32145), .A2(n32152), .ZN(n32151) );
  NOR2HSV2 U37595 ( .A1(n32146), .A2(n32151), .ZN(n32147) );
  NAND2HSV2 U37596 ( .A1(n32147), .A2(n32407), .ZN(n32150) );
  CLKNAND2HSV0 U37597 ( .A1(n32152), .A2(n32148), .ZN(n32149) );
  AOI21HSV4 U37598 ( .A1(n52780), .A2(n32348), .B(n46584), .ZN(n32228) );
  INOR2HSV4 U37599 ( .A1(n32155), .B1(n32154), .ZN(n32350) );
  INHSV1 U37600 ( .I(n32162), .ZN(n47977) );
  NOR2HSV2 U37601 ( .A1(n36083), .A2(\pe6/ti_7t [14]), .ZN(n32467) );
  NOR2HSV0 U37602 ( .A1(n32467), .A2(n32530), .ZN(n32322) );
  AOI21HSV4 U37603 ( .A1(n29757), .A2(n46587), .B(n32158), .ZN(n32324) );
  NOR2HSV4 U37604 ( .A1(n32324), .A2(n32160), .ZN(n32227) );
  CLKNHSV0 U37605 ( .I(n32444), .ZN(n32161) );
  INHSV2 U37606 ( .I(n32651), .ZN(n46155) );
  CLKNAND2HSV0 U37607 ( .A1(n32163), .A2(n46155), .ZN(n32164) );
  CLKNAND2HSV1 U37608 ( .A1(n59166), .A2(n32353), .ZN(n32224) );
  CLKNHSV0 U37609 ( .I(\pe6/got [26]), .ZN(n32166) );
  CLKNAND2HSV1 U37610 ( .A1(n32167), .A2(n58808), .ZN(n32217) );
  INHSV2 U37611 ( .I(n35607), .ZN(n58856) );
  NAND2HSV0 U37612 ( .A1(n32168), .A2(n58856), .ZN(n32170) );
  NAND2HSV0 U37613 ( .A1(\pe6/bq[18] ), .A2(n32973), .ZN(n32169) );
  XOR2HSV0 U37614 ( .A1(n32170), .A2(n32169), .Z(n32177) );
  NAND2HSV0 U37615 ( .A1(n32172), .A2(n32171), .ZN(n32175) );
  NAND2HSV0 U37616 ( .A1(n32173), .A2(n32605), .ZN(n32174) );
  XOR2HSV0 U37617 ( .A1(n32175), .A2(n32174), .Z(n32176) );
  XOR2HSV0 U37618 ( .A1(n32177), .A2(n32176), .Z(n32185) );
  CLKNAND2HSV1 U37619 ( .A1(n32276), .A2(n31972), .ZN(n32179) );
  INHSV2 U37620 ( .I(n32269), .ZN(n59261) );
  INHSV2 U37621 ( .I(n32245), .ZN(n32573) );
  CLKNAND2HSV1 U37622 ( .A1(n59261), .A2(n32573), .ZN(n32178) );
  XOR2HSV0 U37623 ( .A1(n32179), .A2(n32178), .Z(n32183) );
  NAND2HSV0 U37624 ( .A1(n59206), .A2(n33022), .ZN(n32181) );
  CLKNAND2HSV1 U37625 ( .A1(n35760), .A2(\pe6/aot [21]), .ZN(n32180) );
  XOR2HSV0 U37626 ( .A1(n32181), .A2(n32180), .Z(n32182) );
  XOR2HSV0 U37627 ( .A1(n32183), .A2(n32182), .Z(n32184) );
  XOR2HSV0 U37628 ( .A1(n32185), .A2(n32184), .Z(n32187) );
  CLKNAND2HSV1 U37629 ( .A1(n35612), .A2(n53101), .ZN(n32186) );
  XNOR2HSV1 U37630 ( .A1(n32187), .A2(n32186), .ZN(n32207) );
  CLKNAND2HSV1 U37631 ( .A1(n59259), .A2(\pe6/aot [17]), .ZN(n32189) );
  NAND2HSV0 U37632 ( .A1(n44700), .A2(n46662), .ZN(n32188) );
  XOR2HSV0 U37633 ( .A1(n32189), .A2(n32188), .Z(n32192) );
  CLKNHSV2 U37634 ( .I(n53103), .ZN(n49174) );
  CLKNAND2HSV0 U37635 ( .A1(n59236), .A2(n49174), .ZN(n32190) );
  XNOR2HSV1 U37636 ( .A1(n32190), .A2(\pe6/phq [16]), .ZN(n32191) );
  XNOR2HSV1 U37637 ( .A1(n32192), .A2(n32191), .ZN(n32197) );
  CLKNAND2HSV1 U37638 ( .A1(n32486), .A2(\pe6/aot [19]), .ZN(n35928) );
  OAI22HSV1 U37639 ( .A1(n32484), .A2(n46637), .B1(n44397), .B2(n32714), .ZN(
        n32194) );
  OAI21HSV0 U37640 ( .A1(n46179), .A2(n35928), .B(n32194), .ZN(n32195) );
  NAND2HSV0 U37641 ( .A1(\pe6/bq[17] ), .A2(n59276), .ZN(n32880) );
  XNOR2HSV1 U37642 ( .A1(n32195), .A2(n32880), .ZN(n32196) );
  XNOR2HSV1 U37643 ( .A1(n32197), .A2(n32196), .ZN(n32205) );
  CLKNAND2HSV0 U37644 ( .A1(n32252), .A2(\pe6/aot [23]), .ZN(n32585) );
  CLKNAND2HSV1 U37645 ( .A1(n59201), .A2(\pe6/pvq [16]), .ZN(n32199) );
  XOR2HSV0 U37646 ( .A1(n32585), .A2(n32199), .Z(n32203) );
  CLKNAND2HSV1 U37647 ( .A1(n32606), .A2(n59234), .ZN(n32201) );
  NAND2HSV0 U37648 ( .A1(n45812), .A2(n33004), .ZN(n32200) );
  XOR2HSV0 U37649 ( .A1(n32201), .A2(n32200), .Z(n32202) );
  XOR2HSV0 U37650 ( .A1(n32203), .A2(n32202), .Z(n32204) );
  XNOR2HSV1 U37651 ( .A1(n32205), .A2(n32204), .ZN(n32206) );
  XNOR2HSV1 U37652 ( .A1(n32207), .A2(n32206), .ZN(n32209) );
  CLKNAND2HSV0 U37653 ( .A1(n32286), .A2(n49096), .ZN(n32208) );
  XNOR2HSV1 U37654 ( .A1(n32209), .A2(n32208), .ZN(n32211) );
  NAND2HSV0 U37655 ( .A1(n32384), .A2(n32563), .ZN(n32210) );
  XNOR2HSV1 U37656 ( .A1(n32211), .A2(n32210), .ZN(n32213) );
  CLKNAND2HSV0 U37657 ( .A1(n59670), .A2(n59328), .ZN(n32212) );
  XOR2HSV0 U37658 ( .A1(n32213), .A2(n32212), .Z(n32215) );
  CLKNAND2HSV1 U37659 ( .A1(n32293), .A2(n49825), .ZN(n32214) );
  XNOR2HSV1 U37660 ( .A1(n32215), .A2(n32214), .ZN(n32216) );
  XOR2HSV0 U37661 ( .A1(n32217), .A2(n32216), .Z(n32220) );
  CLKNAND2HSV0 U37662 ( .A1(n32218), .A2(n32970), .ZN(n32219) );
  XOR2HSV0 U37663 ( .A1(n32220), .A2(n32219), .Z(n32222) );
  CLKNAND2HSV1 U37664 ( .A1(n44476), .A2(n46283), .ZN(n32221) );
  XNOR2HSV4 U37665 ( .A1(n32224), .A2(n32223), .ZN(n32321) );
  XNOR2HSV4 U37666 ( .A1(n32225), .A2(n32321), .ZN(n32226) );
  XNOR2HSV4 U37667 ( .A1(n32227), .A2(n32226), .ZN(n52779) );
  OAI21HSV4 U37668 ( .A1(n32228), .A2(n32350), .B(n52779), .ZN(n32230) );
  INHSV2 U37669 ( .I(\pe6/ti_7t [16]), .ZN(n32330) );
  NOR2HSV2 U37670 ( .A1(n32330), .A2(n52710), .ZN(n32349) );
  INHSV2 U37671 ( .I(n32349), .ZN(n32229) );
  INHSV2 U37672 ( .I(n52780), .ZN(n32231) );
  NOR2HSV4 U37673 ( .A1(n29751), .A2(n32231), .ZN(n32524) );
  CLKNAND2HSV3 U37674 ( .A1(n32233), .A2(n32232), .ZN(n32426) );
  AND2HSV2 U37675 ( .A1(n32822), .A2(n36029), .Z(n32234) );
  CLKNAND2HSV4 U37676 ( .A1(n32524), .A2(n32235), .ZN(n32351) );
  NOR2HSV1 U37677 ( .A1(n32814), .A2(n32241), .ZN(n32236) );
  XOR2HSV2 U37678 ( .A1(n32237), .A2(n32236), .Z(n32347) );
  INHSV2 U37679 ( .I(n32238), .ZN(n32423) );
  NAND2HSV4 U37680 ( .A1(n52765), .A2(n47934), .ZN(n32469) );
  NOR2HSV2 U37681 ( .A1(n32467), .A2(n44376), .ZN(n32240) );
  CLKNAND2HSV1 U37682 ( .A1(n59596), .A2(n32242), .ZN(n32305) );
  CLKNAND2HSV1 U37683 ( .A1(n32841), .A2(n59027), .ZN(n32299) );
  NAND2HSV2 U37684 ( .A1(n59597), .A2(n32009), .ZN(n32297) );
  CLKNAND2HSV1 U37685 ( .A1(n36150), .A2(n35925), .ZN(n32244) );
  CLKNAND2HSV0 U37686 ( .A1(n44700), .A2(n32876), .ZN(n32243) );
  XOR2HSV0 U37687 ( .A1(n32244), .A2(n32243), .Z(n32249) );
  CLKNHSV0 U37688 ( .I(n31425), .ZN(n46672) );
  INHSV2 U37689 ( .I(n32245), .ZN(n49760) );
  NAND2HSV2 U37690 ( .A1(n46672), .A2(n49760), .ZN(n32247) );
  NAND2HSV0 U37691 ( .A1(\pe6/bq[17] ), .A2(n36114), .ZN(n32246) );
  XOR2HSV0 U37692 ( .A1(n32247), .A2(n32246), .Z(n32248) );
  XOR2HSV0 U37693 ( .A1(n32249), .A2(n32248), .Z(n32258) );
  INHSV2 U37694 ( .I(n35607), .ZN(n32564) );
  NAND2HSV2 U37695 ( .A1(n59251), .A2(n32564), .ZN(n32251) );
  NAND2HSV0 U37696 ( .A1(\pe6/bq[16] ), .A2(n59276), .ZN(n32250) );
  XOR2HSV0 U37697 ( .A1(n32251), .A2(n32250), .Z(n32256) );
  NAND2HSV0 U37698 ( .A1(n59206), .A2(n36153), .ZN(n32254) );
  NAND2HSV0 U37699 ( .A1(n32252), .A2(\pe6/aot [22]), .ZN(n32253) );
  XOR2HSV0 U37700 ( .A1(n32254), .A2(n32253), .Z(n32255) );
  XOR2HSV0 U37701 ( .A1(n32256), .A2(n32255), .Z(n32257) );
  XOR2HSV0 U37702 ( .A1(n32258), .A2(n32257), .Z(n32260) );
  INHSV2 U37703 ( .I(n53103), .ZN(n35723) );
  NAND2HSV0 U37704 ( .A1(n35612), .A2(n35723), .ZN(n32259) );
  XNOR2HSV1 U37705 ( .A1(n32260), .A2(n32259), .ZN(n32285) );
  NOR2HSV2 U37706 ( .A1(n35647), .A2(n35864), .ZN(n32262) );
  CLKNHSV0 U37707 ( .I(n59194), .ZN(n33003) );
  NAND2HSV0 U37708 ( .A1(n33003), .A2(n33022), .ZN(n32261) );
  XOR2HSV0 U37709 ( .A1(n32262), .A2(n32261), .Z(n32265) );
  INHSV4 U37710 ( .I(\pe6/got [16]), .ZN(n49666) );
  INHSV2 U37711 ( .I(n49666), .ZN(n59031) );
  NAND2HSV0 U37712 ( .A1(n59236), .A2(n59031), .ZN(n32263) );
  XOR2HSV0 U37713 ( .A1(n32263), .A2(\pe6/phq [17]), .Z(n32264) );
  XOR2HSV0 U37714 ( .A1(n32265), .A2(n32264), .Z(n32275) );
  INHSV2 U37715 ( .I(n32589), .ZN(n32588) );
  CLKNAND2HSV1 U37716 ( .A1(n32486), .A2(n32588), .ZN(n32487) );
  OAI22HSV0 U37717 ( .A1(n32266), .A2(n44397), .B1(n59205), .B2(n32589), .ZN(
        n32267) );
  OAI21HSV2 U37718 ( .A1(n32268), .A2(n32487), .B(n32267), .ZN(n32273) );
  CLKNAND2HSV1 U37719 ( .A1(n59247), .A2(\pe6/aot [17]), .ZN(n32490) );
  OAI22HSV0 U37720 ( .A1(n32269), .A2(n58851), .B1(n36124), .B2(n46637), .ZN(
        n32270) );
  OAI21HSV1 U37721 ( .A1(n32271), .A2(n32490), .B(n32270), .ZN(n32272) );
  XOR2HSV0 U37722 ( .A1(n32273), .A2(n32272), .Z(n32274) );
  XOR2HSV0 U37723 ( .A1(n32275), .A2(n32274), .Z(n32283) );
  NAND2HSV0 U37724 ( .A1(n32276), .A2(n32605), .ZN(n36120) );
  CLKNAND2HSV1 U37725 ( .A1(n36161), .A2(\pe6/pvq [17]), .ZN(n32277) );
  XOR2HSV0 U37726 ( .A1(n36120), .A2(n32277), .Z(n32281) );
  INHSV2 U37727 ( .I(n46789), .ZN(n46217) );
  CLKNAND2HSV1 U37728 ( .A1(n32576), .A2(n46217), .ZN(n32279) );
  INHSV1 U37729 ( .I(n35816), .ZN(n58991) );
  CLKNAND2HSV0 U37730 ( .A1(n32606), .A2(n58991), .ZN(n32278) );
  XOR2HSV0 U37731 ( .A1(n32279), .A2(n32278), .Z(n32280) );
  XOR2HSV0 U37732 ( .A1(n32281), .A2(n32280), .Z(n32282) );
  XNOR2HSV1 U37733 ( .A1(n32283), .A2(n32282), .ZN(n32284) );
  XNOR2HSV1 U37734 ( .A1(n32285), .A2(n32284), .ZN(n32288) );
  CLKNAND2HSV1 U37735 ( .A1(n32286), .A2(n36104), .ZN(n32287) );
  XNOR2HSV1 U37736 ( .A1(n32288), .A2(n32287), .ZN(n32290) );
  NAND2HSV0 U37737 ( .A1(n32384), .A2(n49096), .ZN(n32289) );
  XNOR2HSV1 U37738 ( .A1(n32290), .A2(n32289), .ZN(n32292) );
  CLKNAND2HSV1 U37739 ( .A1(n59670), .A2(n32563), .ZN(n32291) );
  XOR2HSV0 U37740 ( .A1(n32292), .A2(n32291), .Z(n32295) );
  CLKNAND2HSV0 U37741 ( .A1(n32293), .A2(n59328), .ZN(n32294) );
  XNOR2HSV1 U37742 ( .A1(n32295), .A2(n32294), .ZN(n32296) );
  XNOR2HSV1 U37743 ( .A1(n32297), .A2(n32296), .ZN(n32298) );
  XOR2HSV0 U37744 ( .A1(n32299), .A2(n32298), .Z(n32301) );
  CLKNAND2HSV0 U37745 ( .A1(n36185), .A2(n32970), .ZN(n32300) );
  XNOR2HSV1 U37746 ( .A1(n32301), .A2(n32300), .ZN(n32302) );
  XOR2HSV0 U37747 ( .A1(n32303), .A2(n32302), .Z(n32304) );
  XNOR2HSV1 U37748 ( .A1(n32305), .A2(n32304), .ZN(n32308) );
  CLKAND2HSV1 U37749 ( .A1(n32306), .A2(n49665), .Z(n32307) );
  XNOR2HSV4 U37750 ( .A1(n32313), .A2(n32429), .ZN(n32531) );
  INHSV2 U37751 ( .I(n32531), .ZN(n32341) );
  CLKNAND2HSV0 U37752 ( .A1(n32514), .A2(n32333), .ZN(n32319) );
  CLKNHSV0 U37753 ( .I(n32335), .ZN(n32317) );
  CLKNAND2HSV0 U37754 ( .A1(n32514), .A2(n32317), .ZN(n32318) );
  NAND2HSV2 U37755 ( .A1(n32319), .A2(n32318), .ZN(n32435) );
  XNOR2HSV4 U37756 ( .A1(n32321), .A2(n32320), .ZN(n32343) );
  CLKNHSV1 U37757 ( .I(n32322), .ZN(n32323) );
  NOR2HSV4 U37758 ( .A1(n32324), .A2(n32323), .ZN(n32328) );
  CLKNHSV0 U37759 ( .I(n32325), .ZN(n32326) );
  NAND2HSV2 U37760 ( .A1(n32326), .A2(n32159), .ZN(n32327) );
  AOI21HSV0 U37761 ( .A1(n32330), .A2(n32329), .B(n46549), .ZN(n32344) );
  INHSV2 U37762 ( .I(n47970), .ZN(n32332) );
  CLKNAND2HSV3 U37763 ( .A1(n32337), .A2(n32332), .ZN(n32331) );
  NAND2HSV4 U37764 ( .A1(n32331), .A2(n46591), .ZN(n32434) );
  NOR2HSV0 U37765 ( .A1(n32333), .A2(n47970), .ZN(n32334) );
  CLKNAND2HSV0 U37766 ( .A1(n32335), .A2(n32334), .ZN(n32339) );
  CLKNAND2HSV0 U37767 ( .A1(n29647), .A2(n32336), .ZN(n32338) );
  AOI21HSV2 U37768 ( .A1(n32339), .A2(n32338), .B(n32337), .ZN(n32436) );
  AOI21HSV4 U37769 ( .A1(n32435), .A2(n32434), .B(n32436), .ZN(n32642) );
  NAND2HSV4 U37770 ( .A1(n32341), .A2(n32642), .ZN(n32812) );
  NAND3HSV2 U37771 ( .A1(n32514), .A2(n32513), .A3(n32512), .ZN(n32838) );
  XNOR2HSV4 U37772 ( .A1(n32343), .A2(n32342), .ZN(n32418) );
  NAND2HSV2 U37773 ( .A1(n32344), .A2(n32793), .ZN(n32417) );
  CLKBUFHSV4 U37774 ( .I(n32345), .Z(n49381) );
  NAND3HSV4 U37775 ( .A1(n32531), .A2(n32648), .A3(n32644), .ZN(n32813) );
  INHSV2 U37776 ( .I(n32533), .ZN(n32652) );
  BUFHSV2 U37777 ( .I(n32652), .Z(n32811) );
  NAND3HSV4 U37778 ( .A1(n32812), .A2(n32813), .A3(n32811), .ZN(n32692) );
  CLKXOR2HSV4 U37779 ( .A1(n32347), .A2(n32346), .Z(n32446) );
  CLKNAND2HSV2 U37780 ( .A1(n32521), .A2(n52779), .ZN(n32352) );
  AOI21HSV4 U37781 ( .A1(n29751), .A2(n32350), .B(n32349), .ZN(n32519) );
  BUFHSV2 U37782 ( .I(n32353), .Z(n59420) );
  INHSV2 U37783 ( .I(n32506), .ZN(n59036) );
  NAND2HSV2 U37784 ( .A1(n59036), .A2(n32354), .ZN(n32402) );
  NAND2HSV2 U37785 ( .A1(n32165), .A2(n46283), .ZN(n32400) );
  CLKNAND2HSV1 U37786 ( .A1(n32841), .A2(n32009), .ZN(n32394) );
  CLKNAND2HSV1 U37787 ( .A1(n59597), .A2(n59328), .ZN(n32392) );
  CLKNAND2HSV1 U37788 ( .A1(n32576), .A2(\pe6/aot [15]), .ZN(n32356) );
  CLKNAND2HSV0 U37789 ( .A1(n59247), .A2(n32573), .ZN(n32355) );
  XOR2HSV0 U37790 ( .A1(n32356), .A2(n32355), .Z(n32360) );
  CLKNAND2HSV1 U37791 ( .A1(n59251), .A2(\pe6/aot [19]), .ZN(n32358) );
  CLKNAND2HSV0 U37792 ( .A1(\pe6/bq[17] ), .A2(n59040), .ZN(n32357) );
  XOR2HSV0 U37793 ( .A1(n32358), .A2(n32357), .Z(n32359) );
  XOR2HSV0 U37794 ( .A1(n32360), .A2(n32359), .Z(n32368) );
  NAND2HSV2 U37795 ( .A1(n32567), .A2(n36114), .ZN(n32362) );
  CLKNAND2HSV1 U37796 ( .A1(n32568), .A2(n31972), .ZN(n32361) );
  XOR2HSV0 U37797 ( .A1(n32362), .A2(n32361), .Z(n32366) );
  NAND2HSV0 U37798 ( .A1(n44700), .A2(n32605), .ZN(n32364) );
  CLKNAND2HSV0 U37799 ( .A1(n33003), .A2(\pe6/aot [23]), .ZN(n32363) );
  XOR2HSV0 U37800 ( .A1(n32364), .A2(n32363), .Z(n32365) );
  XOR2HSV0 U37801 ( .A1(n32366), .A2(n32365), .Z(n32367) );
  XOR2HSV0 U37802 ( .A1(n32368), .A2(n32367), .Z(n32370) );
  NAND2HSV0 U37803 ( .A1(n35612), .A2(n59316), .ZN(n32369) );
  XNOR2HSV1 U37804 ( .A1(n32370), .A2(n32369), .ZN(n32381) );
  CLKNAND2HSV1 U37805 ( .A1(n32606), .A2(n32588), .ZN(n32489) );
  CLKNAND2HSV1 U37806 ( .A1(n46626), .A2(\pe6/pvq [18]), .ZN(n32371) );
  XOR2HSV0 U37807 ( .A1(n32489), .A2(n32371), .Z(n32379) );
  CLKNAND2HSV0 U37808 ( .A1(n33023), .A2(n32564), .ZN(n35929) );
  NAND2HSV0 U37809 ( .A1(n45812), .A2(n32564), .ZN(n49682) );
  NAND2HSV2 U37810 ( .A1(n59261), .A2(n59044), .ZN(n35839) );
  INHSV2 U37811 ( .I(n31253), .ZN(n32740) );
  XOR2HSV0 U37812 ( .A1(n32375), .A2(n32374), .Z(n32376) );
  XOR4HSV1 U37813 ( .A1(n32379), .A2(n32378), .A3(n32377), .A4(n32376), .Z(
        n32380) );
  XNOR2HSV1 U37814 ( .A1(n32381), .A2(n32380), .ZN(n32383) );
  CLKNAND2HSV1 U37815 ( .A1(n32286), .A2(n35723), .ZN(n32382) );
  XNOR2HSV1 U37816 ( .A1(n32383), .A2(n32382), .ZN(n32386) );
  NAND2HSV0 U37817 ( .A1(n32384), .A2(\pe6/got [18]), .ZN(n32385) );
  XNOR2HSV1 U37818 ( .A1(n32386), .A2(n32385), .ZN(n32388) );
  CLKNAND2HSV1 U37819 ( .A1(n58940), .A2(n35922), .ZN(n32387) );
  XOR2HSV0 U37820 ( .A1(n32388), .A2(n32387), .Z(n32390) );
  CLKNAND2HSV1 U37821 ( .A1(n59295), .A2(n32563), .ZN(n32389) );
  XNOR2HSV1 U37822 ( .A1(n32390), .A2(n32389), .ZN(n32391) );
  XNOR2HSV1 U37823 ( .A1(n32392), .A2(n32391), .ZN(n32393) );
  XNOR2HSV1 U37824 ( .A1(n32394), .A2(n32393), .ZN(n32396) );
  CLKNAND2HSV1 U37825 ( .A1(n59917), .A2(n58808), .ZN(n32395) );
  XNOR2HSV1 U37826 ( .A1(n32396), .A2(n32395), .ZN(n32397) );
  XOR2HSV0 U37827 ( .A1(n32398), .A2(n32397), .Z(n32399) );
  XNOR2HSV1 U37828 ( .A1(n32400), .A2(n32399), .ZN(n32401) );
  XNOR2HSV1 U37829 ( .A1(n32402), .A2(n32401), .ZN(n32404) );
  AOI21HSV2 U37830 ( .A1(n59420), .A2(n49665), .B(n32404), .ZN(n32403) );
  INHSV2 U37831 ( .I(n32403), .ZN(n32406) );
  NAND3HSV2 U37832 ( .A1(n32404), .A2(n59420), .A3(n35789), .ZN(n32405) );
  NAND2HSV2 U37833 ( .A1(n32406), .A2(n32405), .ZN(n32409) );
  CLKNAND2HSV0 U37834 ( .A1(n32407), .A2(n33061), .ZN(n32408) );
  CLKNHSV1 U37835 ( .I(\pe6/got [29]), .ZN(n35777) );
  NOR2HSV1 U37836 ( .A1(n32467), .A2(n35777), .ZN(n32410) );
  INHSV2 U37837 ( .I(n32412), .ZN(n32413) );
  NAND2HSV2 U37838 ( .A1(n32413), .A2(n32458), .ZN(n32414) );
  NOR2HSV0 U37839 ( .A1(n32838), .A2(n32533), .ZN(n32415) );
  AO22HSV1 U37840 ( .A1(n32417), .A2(n32652), .B1(n32416), .B2(n32415), .Z(
        n32432) );
  CLKNAND2HSV0 U37841 ( .A1(n32418), .A2(n32652), .ZN(n32419) );
  INAND2HSV2 U37842 ( .A1(n32419), .B1(n35898), .ZN(n32420) );
  INHSV2 U37843 ( .I(n32420), .ZN(n32431) );
  CLKNAND2HSV0 U37844 ( .A1(n32422), .A2(n32421), .ZN(n32425) );
  CLKNAND2HSV1 U37845 ( .A1(n32423), .A2(n32422), .ZN(n32424) );
  NAND2HSV2 U37846 ( .A1(n32425), .A2(n32424), .ZN(n32427) );
  INHSV2 U37847 ( .I(n32646), .ZN(n32430) );
  OAI21HSV2 U37848 ( .A1(n32432), .A2(n32431), .B(n32430), .ZN(n32442) );
  INHSV2 U37849 ( .I(n32433), .ZN(n32643) );
  INHSV2 U37850 ( .I(n32434), .ZN(n32438) );
  CLKNHSV2 U37851 ( .I(n33063), .ZN(n32439) );
  NAND2HSV2 U37852 ( .A1(n32558), .A2(n32557), .ZN(n32691) );
  INHSV4 U37853 ( .I(n32558), .ZN(n32560) );
  CLKNAND2HSV2 U37854 ( .A1(n32691), .A2(n32690), .ZN(n32445) );
  INHSV2 U37855 ( .I(\pe6/ti_7t [18]), .ZN(n32460) );
  NOR2HSV1 U37856 ( .A1(n32460), .A2(n52701), .ZN(n32824) );
  INHSV2 U37857 ( .I(n32824), .ZN(n32925) );
  OAI22HSV4 U37858 ( .A1(n32445), .A2(n32444), .B1(n32443), .B2(n32925), .ZN(
        n32447) );
  CLKNAND2HSV1 U37859 ( .A1(n32446), .A2(n32447), .ZN(n32451) );
  NAND2HSV2 U37860 ( .A1(n32451), .A2(n32450), .ZN(n32556) );
  NOR2HSV4 U37861 ( .A1(n32692), .A2(n44380), .ZN(n32543) );
  NAND2HSV2 U37862 ( .A1(n32453), .A2(n36229), .ZN(n32455) );
  NAND2HSV2 U37863 ( .A1(n32453), .A2(n32814), .ZN(n32454) );
  NAND3HSV4 U37864 ( .A1(n32456), .A2(n32455), .A3(n32454), .ZN(n32542) );
  NAND2HSV2 U37865 ( .A1(n32813), .A2(n32812), .ZN(n32545) );
  AO21HSV0 U37866 ( .A1(n32460), .A2(n31350), .B(n46159), .Z(n32546) );
  CLKNHSV2 U37867 ( .I(n32546), .ZN(n32461) );
  CLKNHSV2 U37868 ( .I(n32463), .ZN(n35806) );
  INHSV2 U37869 ( .I(n32465), .ZN(n32541) );
  NOR2HSV0 U37870 ( .A1(n32467), .A2(n35907), .ZN(n32468) );
  CLKNAND2HSV1 U37871 ( .A1(n32469), .A2(n32468), .ZN(n32518) );
  CLKNAND2HSV1 U37872 ( .A1(n44391), .A2(n49665), .ZN(n32511) );
  CLKNAND2HSV1 U37873 ( .A1(n32165), .A2(n32970), .ZN(n32505) );
  NAND2HSV2 U37874 ( .A1(n58939), .A2(n59174), .ZN(n32503) );
  CLKNAND2HSV1 U37875 ( .A1(n32841), .A2(n59328), .ZN(n32499) );
  CLKNAND2HSV1 U37876 ( .A1(n59597), .A2(n32563), .ZN(n32497) );
  CLKNAND2HSV1 U37877 ( .A1(n36108), .A2(n35723), .ZN(n32493) );
  NAND2HSV0 U37878 ( .A1(n44702), .A2(\pe6/aot [23]), .ZN(n32470) );
  NAND2HSV0 U37879 ( .A1(n33003), .A2(\pe6/aot [22]), .ZN(n32472) );
  NAND2HSV0 U37880 ( .A1(n32982), .A2(n59234), .ZN(n32471) );
  CLKNAND2HSV0 U37881 ( .A1(n32576), .A2(\pe6/aot [14]), .ZN(n32474) );
  NAND2HSV0 U37882 ( .A1(n46624), .A2(\pe6/aot [21]), .ZN(n32473) );
  CLKNAND2HSV0 U37883 ( .A1(n36161), .A2(\pe6/pvq [19]), .ZN(n32476) );
  NAND2HSV0 U37884 ( .A1(n32886), .A2(n33022), .ZN(n32475) );
  NOR2HSV1 U37885 ( .A1(n31791), .A2(n35607), .ZN(n32478) );
  NAND2HSV0 U37886 ( .A1(n32568), .A2(n32605), .ZN(n32477) );
  CLKNAND2HSV0 U37887 ( .A1(n33023), .A2(n58991), .ZN(n32480) );
  CLKNAND2HSV0 U37888 ( .A1(n32567), .A2(n35925), .ZN(n32479) );
  NOR2HSV2 U37889 ( .A1(n48047), .A2(n32086), .ZN(n32482) );
  CLKNAND2HSV0 U37890 ( .A1(n35760), .A2(n32573), .ZN(n32481) );
  NAND2HSV0 U37891 ( .A1(n59236), .A2(n35991), .ZN(n32483) );
  NAND2HSV2 U37892 ( .A1(n59071), .A2(n33024), .ZN(n32591) );
  OAI22HSV0 U37893 ( .A1(n32484), .A2(n46789), .B1(n44411), .B2(n44396), .ZN(
        n32485) );
  CLKNAND2HSV0 U37894 ( .A1(n32486), .A2(n32876), .ZN(n32604) );
  OAI21HSV1 U37895 ( .A1(n35837), .A2(n32877), .B(n32487), .ZN(n32488) );
  CLKNAND2HSV1 U37896 ( .A1(n59267), .A2(\pe6/aot [19]), .ZN(n46636) );
  INHSV2 U37897 ( .I(n49666), .ZN(n36106) );
  CLKNAND2HSV0 U37898 ( .A1(n58940), .A2(n53101), .ZN(n32491) );
  XOR3HSV2 U37899 ( .A1(n32493), .A2(n32492), .A3(n32491), .Z(n32495) );
  CLKNAND2HSV1 U37900 ( .A1(n36183), .A2(n58807), .ZN(n32494) );
  XNOR2HSV1 U37901 ( .A1(n32495), .A2(n32494), .ZN(n32496) );
  XNOR2HSV1 U37902 ( .A1(n32497), .A2(n32496), .ZN(n32498) );
  XNOR2HSV1 U37903 ( .A1(n32499), .A2(n32498), .ZN(n32501) );
  CLKNAND2HSV0 U37904 ( .A1(n29737), .A2(n49825), .ZN(n32500) );
  XNOR2HSV1 U37905 ( .A1(n32501), .A2(n32500), .ZN(n32502) );
  XOR2HSV0 U37906 ( .A1(n32503), .A2(n32502), .Z(n32504) );
  XNOR2HSV1 U37907 ( .A1(n32505), .A2(n32504), .ZN(n32509) );
  INAND2HSV2 U37908 ( .A1(n44507), .B1(n49743), .ZN(n32508) );
  NAND2HSV2 U37909 ( .A1(n59034), .A2(\pe6/got [26]), .ZN(n32507) );
  XOR3HSV2 U37910 ( .A1(n32509), .A2(n32508), .A3(n32507), .Z(n32510) );
  XNOR2HSV1 U37911 ( .A1(n32511), .A2(n32510), .ZN(n32517) );
  NAND3HSV2 U37912 ( .A1(n32514), .A2(n32513), .A3(n32512), .ZN(n32515) );
  NAND2HSV2 U37913 ( .A1(n32515), .A2(n31902), .ZN(n32516) );
  XOR3HSV2 U37914 ( .A1(n32518), .A2(n32517), .A3(n32516), .Z(n32529) );
  NAND3HSV2 U37915 ( .A1(n32521), .A2(n52779), .A3(n35808), .ZN(n32526) );
  NOR2HSV1 U37916 ( .A1(n32522), .A2(n35710), .ZN(n32523) );
  XNOR2HSV4 U37917 ( .A1(n32529), .A2(n32528), .ZN(n32539) );
  NOR2HSV3 U37918 ( .A1(n32531), .A2(n32530), .ZN(n32532) );
  XNOR2HSV4 U37919 ( .A1(n32539), .A2(n32538), .ZN(n32664) );
  INHSV4 U37920 ( .I(n32664), .ZN(n32673) );
  INHSV2 U37921 ( .I(n32673), .ZN(n32540) );
  CLKNAND2HSV2 U37922 ( .A1(n32541), .A2(n32540), .ZN(n32554) );
  CLKNHSV0 U37923 ( .I(n32544), .ZN(n32549) );
  CLKNHSV0 U37924 ( .I(n32545), .ZN(n32548) );
  INHSV2 U37925 ( .I(n32551), .ZN(n32782) );
  NOR2HSV1 U37926 ( .A1(n32546), .A2(n32782), .ZN(n32547) );
  NAND2HSV0 U37927 ( .A1(n32551), .A2(n36050), .ZN(n32784) );
  NAND2HSV2 U37928 ( .A1(n32784), .A2(n46163), .ZN(n32552) );
  CLKNAND2HSV2 U37929 ( .A1(n32553), .A2(n32554), .ZN(n32555) );
  XNOR2HSV4 U37930 ( .A1(n32556), .A2(n32555), .ZN(n32684) );
  INHSV3 U37931 ( .I(n32684), .ZN(n32682) );
  NAND2HSV2 U37932 ( .A1(n32558), .A2(n32557), .ZN(n32561) );
  CLKNHSV2 U37933 ( .I(n36065), .ZN(n32562) );
  NOR2HSV8 U37934 ( .A1(n32820), .A2(n32562), .ZN(n32796) );
  NAND2HSV2 U37935 ( .A1(n59034), .A2(\pe6/got [25]), .ZN(n32636) );
  CLKNAND2HSV0 U37936 ( .A1(n32165), .A2(n35812), .ZN(n32634) );
  CLKNAND2HSV1 U37937 ( .A1(n58939), .A2(n32009), .ZN(n32630) );
  NAND2HSV0 U37938 ( .A1(n32841), .A2(n32563), .ZN(n32626) );
  CLKNAND2HSV0 U37939 ( .A1(n35813), .A2(n58807), .ZN(n32624) );
  NAND2HSV0 U37940 ( .A1(n59247), .A2(n59044), .ZN(n32566) );
  CLKNAND2HSV0 U37941 ( .A1(n46624), .A2(n32564), .ZN(n32565) );
  XOR2HSV0 U37942 ( .A1(n32566), .A2(n32565), .Z(n32572) );
  NAND2HSV0 U37943 ( .A1(n32567), .A2(n59234), .ZN(n32570) );
  NAND2HSV0 U37944 ( .A1(n32568), .A2(n33022), .ZN(n32569) );
  XOR2HSV0 U37945 ( .A1(n32570), .A2(n32569), .Z(n32571) );
  XOR2HSV0 U37946 ( .A1(n32572), .A2(n32571), .Z(n32582) );
  CLKNAND2HSV0 U37947 ( .A1(n59267), .A2(n32573), .ZN(n32575) );
  CLKNAND2HSV0 U37948 ( .A1(n58668), .A2(n36114), .ZN(n32574) );
  XOR2HSV0 U37949 ( .A1(n32575), .A2(n32574), .Z(n32580) );
  CLKNAND2HSV0 U37950 ( .A1(n32576), .A2(\pe6/aot [13]), .ZN(n32578) );
  NAND2HSV0 U37951 ( .A1(n32982), .A2(n46643), .ZN(n32577) );
  XOR2HSV0 U37952 ( .A1(n32578), .A2(n32577), .Z(n32579) );
  XOR2HSV0 U37953 ( .A1(n32580), .A2(n32579), .Z(n32581) );
  XOR2HSV0 U37954 ( .A1(n32582), .A2(n32581), .Z(n32595) );
  NAND2HSV0 U37955 ( .A1(n59236), .A2(\pe6/got [13]), .ZN(n32583) );
  XOR2HSV0 U37956 ( .A1(n32583), .A2(\pe6/phq [20]), .Z(n32587) );
  CLKNAND2HSV0 U37957 ( .A1(n32886), .A2(\pe6/aot [19]), .ZN(n49011) );
  OAI22HSV0 U37958 ( .A1(n31791), .A2(n46637), .B1(n50822), .B2(n49699), .ZN(
        n32584) );
  OAI21HSV0 U37959 ( .A1(n32585), .A2(n49011), .B(n32584), .ZN(n32586) );
  XNOR2HSV1 U37960 ( .A1(n32587), .A2(n32586), .ZN(n32593) );
  NAND2HSV0 U37961 ( .A1(n33000), .A2(n32588), .ZN(n35739) );
  BUFHSV2 U37962 ( .I(n31253), .Z(n32878) );
  XNOR2HSV1 U37963 ( .A1(n32593), .A2(n32592), .ZN(n32594) );
  XNOR2HSV1 U37964 ( .A1(n32595), .A2(n32594), .ZN(n32618) );
  CLKNAND2HSV1 U37965 ( .A1(n32286), .A2(n32596), .ZN(n32617) );
  NAND2HSV0 U37966 ( .A1(n44702), .A2(\pe6/aot [22]), .ZN(n32598) );
  NAND2HSV0 U37967 ( .A1(n33003), .A2(\pe6/aot [21]), .ZN(n32597) );
  XOR2HSV0 U37968 ( .A1(n32598), .A2(n32597), .Z(n32602) );
  CLKNAND2HSV0 U37969 ( .A1(n35760), .A2(\pe6/aot [17]), .ZN(n32600) );
  NAND2HSV0 U37970 ( .A1(n59261), .A2(n49208), .ZN(n32599) );
  XOR2HSV0 U37971 ( .A1(n32600), .A2(n32599), .Z(n32601) );
  XOR2HSV0 U37972 ( .A1(n32602), .A2(n32601), .Z(n32612) );
  NAND2HSV2 U37973 ( .A1(n36161), .A2(\pe6/pvq [20]), .ZN(n32603) );
  XOR2HSV0 U37974 ( .A1(n32604), .A2(n32603), .Z(n32610) );
  NAND2HSV0 U37975 ( .A1(n32606), .A2(n32605), .ZN(n32608) );
  CLKNAND2HSV0 U37976 ( .A1(n59045), .A2(n35925), .ZN(n32607) );
  XOR2HSV0 U37977 ( .A1(n32608), .A2(n32607), .Z(n32609) );
  XOR2HSV0 U37978 ( .A1(n32610), .A2(n32609), .Z(n32611) );
  XOR2HSV0 U37979 ( .A1(n32612), .A2(n32611), .Z(n32614) );
  NAND2HSV0 U37980 ( .A1(n35612), .A2(n35991), .ZN(n32613) );
  XNOR2HSV1 U37981 ( .A1(n32614), .A2(n32613), .ZN(n32616) );
  CLKNAND2HSV1 U37982 ( .A1(n36108), .A2(n46171), .ZN(n32615) );
  XOR4HSV1 U37983 ( .A1(n32618), .A2(n32617), .A3(n32616), .A4(n32615), .Z(
        n32620) );
  CLKNAND2HSV0 U37984 ( .A1(n32900), .A2(n35723), .ZN(n32619) );
  XOR2HSV0 U37985 ( .A1(n32620), .A2(n32619), .Z(n32622) );
  CLKNAND2HSV0 U37986 ( .A1(n36183), .A2(\pe6/got [18]), .ZN(n32621) );
  XNOR2HSV1 U37987 ( .A1(n32622), .A2(n32621), .ZN(n32623) );
  XNOR2HSV1 U37988 ( .A1(n32624), .A2(n32623), .ZN(n32625) );
  XNOR2HSV1 U37989 ( .A1(n32626), .A2(n32625), .ZN(n32628) );
  NAND2HSV0 U37990 ( .A1(n58886), .A2(n59328), .ZN(n32627) );
  XNOR2HSV1 U37991 ( .A1(n32628), .A2(n32627), .ZN(n32629) );
  XOR2HSV0 U37992 ( .A1(n32630), .A2(n32629), .Z(n32633) );
  CLKNAND2HSV1 U37993 ( .A1(n49743), .A2(n31717), .ZN(n32632) );
  XOR3HSV2 U37994 ( .A1(n32634), .A2(n32633), .A3(n32632), .Z(n32635) );
  XNOR2HSV1 U37995 ( .A1(n32636), .A2(n32635), .ZN(n32638) );
  CLKNAND2HSV0 U37996 ( .A1(n44391), .A2(n32242), .ZN(n32637) );
  XNOR2HSV1 U37997 ( .A1(n32638), .A2(n32637), .ZN(n32639) );
  INHSV2 U37998 ( .I(n32640), .ZN(n59171) );
  NAND2HSV2 U37999 ( .A1(n49381), .A2(n59171), .ZN(n32641) );
  CLKAND2HSV2 U38000 ( .A1(n32642), .A2(n32647), .Z(n32656) );
  CLKBUFHSV4 U38001 ( .I(n32643), .Z(n47971) );
  CLKNHSV0 U38002 ( .I(n32644), .ZN(n32645) );
  NOR2HSV2 U38003 ( .A1(n32646), .A2(n32645), .ZN(n32650) );
  CLKAND2HSV1 U38004 ( .A1(n32648), .A2(n32647), .Z(n32649) );
  OR2HSV1 U38005 ( .A1(n32652), .A2(n32651), .Z(n32653) );
  CLKNAND2HSV2 U38006 ( .A1(n32654), .A2(n32653), .ZN(n32655) );
  AOI21HSV4 U38007 ( .A1(n32656), .A2(n47971), .B(n32655), .ZN(n32657) );
  XNOR2HSV4 U38008 ( .A1(n32658), .A2(n32657), .ZN(n32672) );
  MUX2NHSV1 U38009 ( .I0(n32820), .I1(n32796), .S(n32672), .ZN(n32661) );
  XNOR2HSV4 U38010 ( .A1(n32658), .A2(n32657), .ZN(n32667) );
  INHSV2 U38011 ( .I(n32659), .ZN(n32660) );
  INHSV4 U38012 ( .I(n32662), .ZN(n32790) );
  CLKNAND2HSV3 U38013 ( .A1(n32664), .A2(n32663), .ZN(n32688) );
  CLKNHSV0 U38014 ( .I(n32686), .ZN(n32665) );
  OAI21HSV4 U38015 ( .A1(n32686), .A2(n32674), .B(n32673), .ZN(n32942) );
  CLKNAND2HSV2 U38016 ( .A1(n32786), .A2(n32942), .ZN(n47961) );
  NOR2HSV4 U38017 ( .A1(n47961), .A2(n33079), .ZN(n32680) );
  INHSV4 U38018 ( .I(n32667), .ZN(n32948) );
  NOR2HSV3 U38019 ( .A1(n32796), .A2(n32148), .ZN(n32671) );
  CLKNHSV0 U38020 ( .I(\pe6/ti_7t [20]), .ZN(n32668) );
  NAND2HSV0 U38021 ( .A1(n32668), .A2(n36050), .ZN(n32952) );
  CLKNHSV2 U38022 ( .I(n32952), .ZN(n32669) );
  NOR2HSV2 U38023 ( .A1(n32669), .A2(n36066), .ZN(n32675) );
  INHSV2 U38024 ( .I(n32675), .ZN(n32670) );
  AOI21HSV4 U38025 ( .A1(n32948), .A2(n32671), .B(n32670), .ZN(n32678) );
  NAND2HSV2 U38026 ( .A1(n32672), .A2(n32796), .ZN(n32794) );
  INHSV2 U38027 ( .I(n32676), .ZN(n32677) );
  AOI21HSV4 U38028 ( .A1(n32790), .A2(n32680), .B(n32679), .ZN(n32683) );
  INHSV3 U38029 ( .I(n32683), .ZN(n32681) );
  CLKNAND2HSV1 U38030 ( .A1(n47950), .A2(\pe6/ti_7t [21]), .ZN(n35778) );
  INHSV2 U38031 ( .I(n32941), .ZN(n32685) );
  NOR2HSV2 U38032 ( .A1(n32688), .A2(n32687), .ZN(n32689) );
  NOR2HSV4 U38033 ( .A1(n32689), .A2(n32782), .ZN(n32940) );
  OAI21HSV4 U38034 ( .A1(n32942), .A2(n32941), .B(n32940), .ZN(n46170) );
  CLKNAND2HSV1 U38035 ( .A1(n46170), .A2(n46289), .ZN(n32781) );
  CLKNAND2HSV1 U38036 ( .A1(n46592), .A2(n49665), .ZN(n32779) );
  AND2HSV2 U38037 ( .A1(n32692), .A2(n59025), .Z(n32694) );
  BUFHSV2 U38038 ( .I(n32814), .Z(n50805) );
  INHSV2 U38039 ( .I(n50805), .ZN(n35775) );
  CLKNAND2HSV1 U38040 ( .A1(n35775), .A2(n31710), .ZN(n32693) );
  XNOR2HSV1 U38041 ( .A1(n32694), .A2(n32693), .ZN(n32778) );
  BUFHSV2 U38042 ( .I(n32833), .Z(n59032) );
  BUFHSV2 U38043 ( .I(n44391), .Z(n46172) );
  CLKNAND2HSV0 U38044 ( .A1(n46172), .A2(n49825), .ZN(n32774) );
  CLKNHSV0 U38045 ( .I(n59328), .ZN(n32695) );
  INAND2HSV0 U38046 ( .A1(n32695), .B1(n59034), .ZN(n32772) );
  BUFHSV2 U38047 ( .I(n49743), .Z(n35722) );
  NAND2HSV2 U38048 ( .A1(n35722), .A2(n46818), .ZN(n32770) );
  BUFHSV2 U38049 ( .I(n32165), .Z(n58815) );
  NAND2HSV2 U38050 ( .A1(n58815), .A2(\pe6/got [19]), .ZN(n32768) );
  NAND2HSV0 U38051 ( .A1(n26109), .A2(n58715), .ZN(n32766) );
  CLKNAND2HSV1 U38052 ( .A1(n32218), .A2(n36106), .ZN(n32762) );
  NAND2HSV2 U38053 ( .A1(n59597), .A2(\pe6/got [15]), .ZN(n32760) );
  BUFHSV2 U38054 ( .I(n32697), .Z(n35724) );
  BUFHSV2 U38055 ( .I(\pe6/got [12]), .Z(n58719) );
  NAND2HSV0 U38056 ( .A1(n35724), .A2(n58719), .ZN(n32699) );
  CLKNHSV0 U38057 ( .I(n53110), .ZN(n33034) );
  NAND2HSV0 U38058 ( .A1(n32286), .A2(n33034), .ZN(n32698) );
  XOR2HSV0 U38059 ( .A1(n32699), .A2(n32698), .Z(n32754) );
  NAND2HSV2 U38060 ( .A1(n32982), .A2(n59239), .ZN(n32701) );
  CLKNHSV0 U38061 ( .I(\pe6/bq[23] ), .ZN(n44403) );
  INHSV2 U38062 ( .I(n44403), .ZN(n59202) );
  NAND2HSV0 U38063 ( .A1(n59202), .A2(n35726), .ZN(n32700) );
  XOR2HSV0 U38064 ( .A1(n32701), .A2(n32700), .Z(n32705) );
  NAND2HSV0 U38065 ( .A1(n58976), .A2(n46677), .ZN(n32703) );
  NAND2HSV0 U38066 ( .A1(n35768), .A2(n58631), .ZN(n32702) );
  XOR2HSV0 U38067 ( .A1(n32703), .A2(n32702), .Z(n32704) );
  XOR2HSV0 U38068 ( .A1(n32705), .A2(n32704), .Z(n32713) );
  CLKNHSV1 U38069 ( .I(n35607), .ZN(n44439) );
  NAND2HSV0 U38070 ( .A1(n32568), .A2(n44439), .ZN(n32707) );
  NAND2HSV0 U38071 ( .A1(n59267), .A2(n49208), .ZN(n32706) );
  XOR2HSV0 U38072 ( .A1(n32707), .A2(n32706), .Z(n32711) );
  NAND2HSV0 U38073 ( .A1(n44453), .A2(\pe6/aot [17]), .ZN(n32709) );
  CLKNHSV0 U38074 ( .I(n31560), .ZN(n35743) );
  NAND2HSV0 U38075 ( .A1(n35743), .A2(n58999), .ZN(n32708) );
  XOR2HSV0 U38076 ( .A1(n32709), .A2(n32708), .Z(n32710) );
  XOR2HSV0 U38077 ( .A1(n32711), .A2(n32710), .Z(n32712) );
  XOR2HSV0 U38078 ( .A1(n32713), .A2(n32712), .Z(n32731) );
  NAND2HSV0 U38079 ( .A1(n35750), .A2(n32991), .ZN(n32716) );
  NAND2HSV0 U38080 ( .A1(n35740), .A2(\pe6/aot [11]), .ZN(n32715) );
  XOR2HSV0 U38081 ( .A1(n32716), .A2(n32715), .Z(n32720) );
  NAND2HSV0 U38082 ( .A1(n33023), .A2(n36153), .ZN(n32718) );
  NAND2HSV0 U38083 ( .A1(n59217), .A2(n33024), .ZN(n32717) );
  XOR2HSV0 U38084 ( .A1(n32718), .A2(n32717), .Z(n32719) );
  XOR2HSV0 U38085 ( .A1(n32720), .A2(n32719), .Z(n32729) );
  NOR2HSV2 U38086 ( .A1(n48047), .A2(n32877), .ZN(n32722) );
  NAND2HSV0 U38087 ( .A1(n33005), .A2(\pe6/aot [21]), .ZN(n32721) );
  XOR2HSV0 U38088 ( .A1(n32722), .A2(n32721), .Z(n32727) );
  CLKNAND2HSV1 U38089 ( .A1(n36161), .A2(\pe6/pvq [24]), .ZN(n32725) );
  NAND2HSV0 U38090 ( .A1(n44336), .A2(n32973), .ZN(n32724) );
  XOR2HSV0 U38091 ( .A1(n32725), .A2(n32724), .Z(n32726) );
  XOR2HSV0 U38092 ( .A1(n32727), .A2(n32726), .Z(n32728) );
  XOR2HSV0 U38093 ( .A1(n32729), .A2(n32728), .Z(n32730) );
  XOR2HSV0 U38094 ( .A1(n32731), .A2(n32730), .Z(n32752) );
  NAND2HSV0 U38095 ( .A1(n35760), .A2(\pe6/aot [13]), .ZN(n32734) );
  INHSV2 U38096 ( .I(n32732), .ZN(n36168) );
  NAND2HSV0 U38097 ( .A1(n36168), .A2(n59245), .ZN(n32733) );
  XOR2HSV0 U38098 ( .A1(n32734), .A2(n32733), .Z(n32737) );
  BUFHSV2 U38099 ( .I(\pe6/got [9]), .Z(n46633) );
  NAND2HSV0 U38100 ( .A1(n33016), .A2(n46633), .ZN(n32735) );
  XNOR2HSV1 U38101 ( .A1(n32735), .A2(\pe6/phq [24]), .ZN(n32736) );
  XNOR2HSV1 U38102 ( .A1(n32737), .A2(n32736), .ZN(n32743) );
  CLKNAND2HSV1 U38103 ( .A1(n36143), .A2(n35732), .ZN(n58982) );
  OAI22HSV0 U38104 ( .A1(n35816), .A2(n46853), .B1(n36132), .B2(n46789), .ZN(
        n32738) );
  OAI21HSV0 U38105 ( .A1(n32739), .A2(n58982), .B(n32738), .ZN(n32741) );
  INHSV2 U38106 ( .I(\pe6/bq[9] ), .ZN(n44436) );
  INHSV2 U38107 ( .I(n44436), .ZN(n48044) );
  NAND2HSV0 U38108 ( .A1(n48044), .A2(n32740), .ZN(n35736) );
  XNOR2HSV1 U38109 ( .A1(n32741), .A2(n35736), .ZN(n32742) );
  XNOR2HSV1 U38110 ( .A1(n32743), .A2(n32742), .ZN(n32748) );
  XOR2HSV0 U38111 ( .A1(n32744), .A2(n49011), .Z(n32746) );
  INHSV2 U38112 ( .I(\pe6/aot [10]), .ZN(n58463) );
  CLKNAND2HSV0 U38113 ( .A1(n32992), .A2(n58488), .ZN(n46657) );
  CLKNAND2HSV0 U38114 ( .A1(n58668), .A2(n32981), .ZN(n46661) );
  XOR2HSV0 U38115 ( .A1(n46657), .A2(n46661), .Z(n32745) );
  XOR2HSV0 U38116 ( .A1(n32746), .A2(n32745), .Z(n32747) );
  XNOR2HSV1 U38117 ( .A1(n32748), .A2(n32747), .ZN(n32750) );
  NAND2HSV0 U38118 ( .A1(n35725), .A2(n44393), .ZN(n32749) );
  XNOR2HSV1 U38119 ( .A1(n32750), .A2(n32749), .ZN(n32751) );
  XNOR2HSV1 U38120 ( .A1(n32752), .A2(n32751), .ZN(n32753) );
  XNOR2HSV1 U38121 ( .A1(n32754), .A2(n32753), .ZN(n32756) );
  NAND2HSV0 U38122 ( .A1(n59121), .A2(n58811), .ZN(n32755) );
  XOR2HSV0 U38123 ( .A1(n32756), .A2(n32755), .Z(n32758) );
  NAND2HSV0 U38124 ( .A1(n59295), .A2(n58713), .ZN(n32757) );
  XNOR2HSV1 U38125 ( .A1(n32758), .A2(n32757), .ZN(n32759) );
  XNOR2HSV1 U38126 ( .A1(n32760), .A2(n32759), .ZN(n32761) );
  XNOR2HSV1 U38127 ( .A1(n32762), .A2(n32761), .ZN(n32764) );
  CLKNAND2HSV1 U38128 ( .A1(n44476), .A2(n35723), .ZN(n32763) );
  XNOR2HSV1 U38129 ( .A1(n32764), .A2(n32763), .ZN(n32765) );
  XOR2HSV0 U38130 ( .A1(n32766), .A2(n32765), .Z(n32767) );
  XOR2HSV0 U38131 ( .A1(n32768), .A2(n32767), .Z(n32769) );
  XOR2HSV0 U38132 ( .A1(n32770), .A2(n32769), .Z(n32771) );
  XOR2HSV0 U38133 ( .A1(n32772), .A2(n32771), .Z(n32773) );
  XNOR2HSV1 U38134 ( .A1(n32774), .A2(n32773), .ZN(n32775) );
  XNOR2HSV1 U38135 ( .A1(n32776), .A2(n32775), .ZN(n32777) );
  XNOR2HSV1 U38136 ( .A1(n32781), .A2(n32780), .ZN(n32808) );
  NAND2HSV0 U38137 ( .A1(n32784), .A2(n32783), .ZN(n32950) );
  INHSV2 U38138 ( .I(n32950), .ZN(n32946) );
  CLKNAND2HSV1 U38139 ( .A1(n32801), .A2(n32946), .ZN(n32785) );
  INHSV2 U38140 ( .I(n32785), .ZN(n32789) );
  CLKNAND2HSV0 U38141 ( .A1(n29725), .A2(n31350), .ZN(n32787) );
  AOI21HSV2 U38142 ( .A1(n32789), .A2(n29725), .B(n32788), .ZN(n32792) );
  CLKNAND2HSV1 U38143 ( .A1(n32792), .A2(n32791), .ZN(n32806) );
  CLKNAND2HSV1 U38144 ( .A1(n32794), .A2(n32793), .ZN(n32799) );
  AND2HSV2 U38145 ( .A1(n32824), .A2(n46163), .Z(n32795) );
  NOR2HSV4 U38146 ( .A1(n32796), .A2(n32795), .ZN(n32947) );
  NAND2HSV0 U38147 ( .A1(n32947), .A2(n32948), .ZN(n32797) );
  CLKNAND2HSV1 U38148 ( .A1(n32797), .A2(n32946), .ZN(n32798) );
  NOR2HSV2 U38149 ( .A1(n32799), .A2(n32798), .ZN(n32804) );
  INHSV2 U38150 ( .I(n32800), .ZN(n32803) );
  INHSV2 U38151 ( .I(n32801), .ZN(n32802) );
  CLKNAND2HSV0 U38152 ( .A1(n35788), .A2(n35705), .ZN(n32807) );
  XNOR2HSV1 U38153 ( .A1(n32808), .A2(n32807), .ZN(n32809) );
  INHSV2 U38154 ( .I(n32825), .ZN(n32816) );
  NAND2HSV2 U38155 ( .A1(n35721), .A2(n33061), .ZN(n32818) );
  INHSV2 U38156 ( .I(n32816), .ZN(n32817) );
  AOI22HSV4 U38157 ( .A1(n35721), .A2(n32819), .B1(n32818), .B2(n32817), .ZN(
        n32927) );
  CLKNHSV0 U38158 ( .I(n32820), .ZN(n32821) );
  NAND2HSV0 U38159 ( .A1(n32822), .A2(n35705), .ZN(n32930) );
  CLKNHSV0 U38160 ( .I(n32930), .ZN(n32823) );
  CLKNAND2HSV1 U38161 ( .A1(n29677), .A2(n32823), .ZN(n32929) );
  NAND2HSV0 U38162 ( .A1(n32824), .A2(n35705), .ZN(n32826) );
  AOI21HSV0 U38163 ( .A1(n32925), .A2(n44380), .B(n35777), .ZN(n32827) );
  MUX2NHSV1 U38164 ( .I0(n32826), .I1(n32827), .S(n32825), .ZN(n32831) );
  MUX2NHSV1 U38165 ( .I0(n32827), .I1(n32826), .S(n32825), .ZN(n32828) );
  INHSV2 U38166 ( .I(n32828), .ZN(n32829) );
  CLKNAND2HSV2 U38167 ( .A1(n32829), .A2(n59171), .ZN(n32830) );
  OAI22HSV4 U38168 ( .A1(n32832), .A2(n32831), .B1(n32830), .B2(n26472), .ZN(
        n32932) );
  INAND2HSV2 U38169 ( .A1(n44507), .B1(n32833), .ZN(n32835) );
  XNOR2HSV1 U38170 ( .A1(n32835), .A2(n32834), .ZN(n32837) );
  NAND2HSV2 U38171 ( .A1(n46172), .A2(n32970), .ZN(n32836) );
  INAND2HSV2 U38172 ( .A1(n59025), .B1(n32839), .ZN(n32918) );
  CLKNHSV1 U38173 ( .I(n32918), .ZN(n32915) );
  NAND2HSV0 U38174 ( .A1(n32838), .A2(\pe6/got [26]), .ZN(n32840) );
  CLKNAND2HSV1 U38175 ( .A1(n59034), .A2(n35812), .ZN(n32914) );
  INAND2HSV2 U38176 ( .A1(n49003), .B1(n49743), .ZN(n32912) );
  CLKNAND2HSV0 U38177 ( .A1(n32165), .A2(n59328), .ZN(n32910) );
  CLKNAND2HSV0 U38178 ( .A1(n26109), .A2(n46818), .ZN(n32908) );
  CLKNAND2HSV0 U38179 ( .A1(n32841), .A2(\pe6/got [18]), .ZN(n32906) );
  NAND2HSV2 U38180 ( .A1(n35724), .A2(n58713), .ZN(n32843) );
  CLKNAND2HSV1 U38181 ( .A1(n59038), .A2(n58711), .ZN(n32842) );
  XOR2HSV0 U38182 ( .A1(n32843), .A2(n32842), .Z(n32899) );
  CLKNAND2HSV1 U38183 ( .A1(n59206), .A2(n35726), .ZN(n32845) );
  NAND2HSV2 U38184 ( .A1(n31820), .A2(n59189), .ZN(n32844) );
  XOR2HSV0 U38185 ( .A1(n32845), .A2(n32844), .Z(n32849) );
  NAND2HSV2 U38186 ( .A1(n59217), .A2(\pe6/aot [17]), .ZN(n32847) );
  CLKNAND2HSV1 U38187 ( .A1(n33000), .A2(n35925), .ZN(n32846) );
  XOR2HSV0 U38188 ( .A1(n32847), .A2(n32846), .Z(n32848) );
  XOR2HSV0 U38189 ( .A1(n32849), .A2(n32848), .Z(n32857) );
  NAND2HSV2 U38190 ( .A1(n35751), .A2(n32171), .ZN(n32851) );
  NAND2HSV0 U38191 ( .A1(n58668), .A2(n46677), .ZN(n32850) );
  XOR2HSV0 U38192 ( .A1(n32851), .A2(n32850), .Z(n32855) );
  CLKNAND2HSV0 U38193 ( .A1(n32999), .A2(n33024), .ZN(n32853) );
  NAND2HSV2 U38194 ( .A1(n59202), .A2(n44439), .ZN(n32852) );
  XOR2HSV0 U38195 ( .A1(n32853), .A2(n32852), .Z(n32854) );
  XOR2HSV0 U38196 ( .A1(n32855), .A2(n32854), .Z(n32856) );
  XOR2HSV0 U38197 ( .A1(n32857), .A2(n32856), .Z(n32873) );
  NAND2HSV2 U38198 ( .A1(n35768), .A2(n49208), .ZN(n32860) );
  CLKNAND2HSV1 U38199 ( .A1(n32568), .A2(n33004), .ZN(n32859) );
  XOR2HSV0 U38200 ( .A1(n32860), .A2(n32859), .Z(n32864) );
  NAND2HSV2 U38201 ( .A1(n59240), .A2(n32973), .ZN(n32862) );
  CLKNAND2HSV1 U38202 ( .A1(n35743), .A2(\pe6/aot [11]), .ZN(n32861) );
  XOR2HSV0 U38203 ( .A1(n32862), .A2(n32861), .Z(n32863) );
  XOR2HSV0 U38204 ( .A1(n32864), .A2(n32863), .Z(n32871) );
  NOR2HSV2 U38205 ( .A1(n32484), .A2(n58983), .ZN(n32866) );
  CLKNAND2HSV1 U38206 ( .A1(n33023), .A2(n59245), .ZN(n32865) );
  XOR2HSV0 U38207 ( .A1(n32866), .A2(n32865), .Z(n32869) );
  NAND2HSV0 U38208 ( .A1(n33016), .A2(n33034), .ZN(n32867) );
  XOR2HSV0 U38209 ( .A1(n32867), .A2(\pe6/phq [22]), .Z(n32868) );
  XOR2HSV0 U38210 ( .A1(n32869), .A2(n32868), .Z(n32870) );
  XOR2HSV0 U38211 ( .A1(n32871), .A2(n32870), .Z(n32872) );
  XOR2HSV0 U38212 ( .A1(n32873), .A2(n32872), .Z(n32897) );
  NAND2HSV2 U38213 ( .A1(n32992), .A2(n32972), .ZN(n32875) );
  CLKNAND2HSV1 U38214 ( .A1(n35761), .A2(n33022), .ZN(n32874) );
  XOR2HSV0 U38215 ( .A1(n32875), .A2(n32874), .Z(n32893) );
  CLKNAND2HSV1 U38216 ( .A1(n35750), .A2(n32876), .ZN(n36163) );
  OAI22HSV1 U38217 ( .A1(n32878), .A2(n46850), .B1(n46688), .B2(n32877), .ZN(
        n32879) );
  OAI21HSV0 U38218 ( .A1(n36163), .A2(n32880), .B(n32879), .ZN(n32883) );
  BUFHSV2 U38219 ( .I(n26513), .Z(n59201) );
  NAND2HSV2 U38220 ( .A1(n59902), .A2(\pe6/pvq [22]), .ZN(n32882) );
  XNOR2HSV1 U38221 ( .A1(n32883), .A2(n32882), .ZN(n32892) );
  NAND2HSV0 U38222 ( .A1(n33003), .A2(\pe6/aot [19]), .ZN(n32885) );
  CLKNAND2HSV1 U38223 ( .A1(n36168), .A2(n32981), .ZN(n32884) );
  XOR2HSV0 U38224 ( .A1(n32885), .A2(n32884), .Z(n32890) );
  NAND2HSV2 U38225 ( .A1(n33005), .A2(\pe6/aot [23]), .ZN(n32888) );
  NAND2HSV0 U38226 ( .A1(n32886), .A2(\pe6/aot [21]), .ZN(n32887) );
  XOR2HSV0 U38227 ( .A1(n32888), .A2(n32887), .Z(n32889) );
  XOR2HSV0 U38228 ( .A1(n32890), .A2(n32889), .Z(n32891) );
  XOR3HSV2 U38229 ( .A1(n32893), .A2(n32892), .A3(n32891), .Z(n32895) );
  NAND2HSV0 U38230 ( .A1(n35725), .A2(n33039), .ZN(n32894) );
  XNOR2HSV1 U38231 ( .A1(n32895), .A2(n32894), .ZN(n32896) );
  XOR2HSV0 U38232 ( .A1(n32897), .A2(n32896), .Z(n32898) );
  XNOR2HSV1 U38233 ( .A1(n32899), .A2(n32898), .ZN(n32902) );
  CLKNAND2HSV1 U38234 ( .A1(n32900), .A2(\pe6/got [15]), .ZN(n32901) );
  XNOR2HSV1 U38235 ( .A1(n32902), .A2(n32901), .ZN(n32904) );
  NAND2HSV2 U38236 ( .A1(n32293), .A2(n46171), .ZN(n32903) );
  XNOR2HSV1 U38237 ( .A1(n32904), .A2(n32903), .ZN(n32905) );
  XNOR2HSV1 U38238 ( .A1(n32906), .A2(n32905), .ZN(n32907) );
  XOR2HSV0 U38239 ( .A1(n32908), .A2(n32907), .Z(n32909) );
  XNOR2HSV1 U38240 ( .A1(n32910), .A2(n32909), .ZN(n32911) );
  XOR2HSV0 U38241 ( .A1(n32912), .A2(n32911), .Z(n32913) );
  XNOR2HSV1 U38242 ( .A1(n32914), .A2(n32913), .ZN(n32916) );
  OAI21HSV2 U38243 ( .A1(n32915), .A2(n32919), .B(n32916), .ZN(n32923) );
  CLKNHSV0 U38244 ( .I(n32916), .ZN(n32917) );
  CLKAND2HSV2 U38245 ( .A1(n32918), .A2(n32917), .Z(n32921) );
  INHSV1 U38246 ( .I(n32919), .ZN(n32920) );
  CLKNAND2HSV1 U38247 ( .A1(n32921), .A2(n32920), .ZN(n32922) );
  NAND2HSV2 U38248 ( .A1(n32923), .A2(n32922), .ZN(n32934) );
  CLKNAND2HSV2 U38249 ( .A1(n32932), .A2(n32934), .ZN(n32924) );
  INHSV2 U38250 ( .I(n32924), .ZN(n32928) );
  INAND2HSV4 U38251 ( .A1(n32927), .B1(n32926), .ZN(n32933) );
  NAND3HSV2 U38252 ( .A1(n32929), .A2(n32928), .A3(n32933), .ZN(n32939) );
  NOR2HSV1 U38253 ( .A1(n32934), .A2(n32930), .ZN(n32931) );
  NAND2HSV2 U38254 ( .A1(n29677), .A2(n32931), .ZN(n32938) );
  CLKNAND2HSV2 U38255 ( .A1(n32933), .A2(n32932), .ZN(n32936) );
  INHSV2 U38256 ( .I(n32934), .ZN(n32935) );
  CLKNAND2HSV3 U38257 ( .A1(n32936), .A2(n32935), .ZN(n32937) );
  NAND3HSV4 U38258 ( .A1(n32939), .A2(n32938), .A3(n32937), .ZN(n32945) );
  XNOR2HSV4 U38259 ( .A1(n32945), .A2(n32944), .ZN(n32957) );
  XNOR2HSV4 U38260 ( .A1(n32948), .A2(n32947), .ZN(n47953) );
  NOR2HSV0 U38261 ( .A1(n32950), .A2(n33079), .ZN(n32951) );
  AND2HSV2 U38262 ( .A1(n32952), .A2(n36095), .Z(n32953) );
  AOI21HSV4 U38263 ( .A1(n29637), .A2(n47952), .B(n32955), .ZN(n32956) );
  XNOR2HSV4 U38264 ( .A1(n32957), .A2(n32956), .ZN(n33069) );
  INHSV2 U38265 ( .I(n35778), .ZN(n35782) );
  CLKNHSV2 U38266 ( .I(n35782), .ZN(n32958) );
  INOR2HSV0 U38267 ( .A1(n35778), .B1(n32961), .ZN(n32968) );
  NAND2HSV2 U38268 ( .A1(n44369), .A2(\pe6/ti_7t [22]), .ZN(n35703) );
  NAND2HSV0 U38269 ( .A1(n35703), .A2(n36023), .ZN(n32963) );
  NAND2HSV2 U38270 ( .A1(n32963), .A2(n59339), .ZN(n32964) );
  AOI21HSV2 U38271 ( .A1(n51451), .A2(n35703), .B(n32964), .ZN(n32965) );
  XNOR2HSV4 U38272 ( .A1(n32966), .A2(n32965), .ZN(n35717) );
  NOR2HSV2 U38273 ( .A1(n35717), .A2(n32941), .ZN(n33087) );
  CLKNHSV0 U38274 ( .I(n32443), .ZN(n32967) );
  INHSV2 U38275 ( .I(n32968), .ZN(n35919) );
  NAND2HSV2 U38276 ( .A1(n35919), .A2(n59339), .ZN(n32969) );
  NOR2HSV4 U38277 ( .A1(n35921), .A2(n32969), .ZN(n33078) );
  INAND2HSV0 U38278 ( .A1(n49003), .B1(n59034), .ZN(n33060) );
  CLKNAND2HSV1 U38279 ( .A1(n35722), .A2(n59328), .ZN(n33058) );
  NAND2HSV0 U38280 ( .A1(n59596), .A2(\pe6/got [20]), .ZN(n33056) );
  NAND2HSV0 U38281 ( .A1(n26109), .A2(n58807), .ZN(n33054) );
  CLKNAND2HSV0 U38282 ( .A1(n32841), .A2(n32971), .ZN(n33050) );
  NAND2HSV0 U38283 ( .A1(n35813), .A2(n36106), .ZN(n33048) );
  NAND2HSV0 U38284 ( .A1(n59071), .A2(n32972), .ZN(n32975) );
  NAND2HSV0 U38285 ( .A1(n35750), .A2(n32973), .ZN(n32974) );
  XOR2HSV0 U38286 ( .A1(n32975), .A2(n32974), .Z(n32980) );
  NAND2HSV0 U38287 ( .A1(n32568), .A2(\pe6/aot [21]), .ZN(n32978) );
  CLKNHSV0 U38288 ( .I(n32976), .ZN(n59272) );
  NAND2HSV0 U38289 ( .A1(n36168), .A2(n59272), .ZN(n32977) );
  XOR2HSV0 U38290 ( .A1(n32978), .A2(n32977), .Z(n32979) );
  XOR2HSV0 U38291 ( .A1(n32980), .A2(n32979), .Z(n32990) );
  NAND2HSV0 U38292 ( .A1(n35751), .A2(n32981), .ZN(n32984) );
  NAND2HSV0 U38293 ( .A1(n32982), .A2(n59245), .ZN(n32983) );
  XOR2HSV0 U38294 ( .A1(n32984), .A2(n32983), .Z(n32988) );
  NAND2HSV0 U38295 ( .A1(n59202), .A2(\pe6/aot [19]), .ZN(n32986) );
  NAND2HSV0 U38296 ( .A1(n35743), .A2(\pe6/aot [10]), .ZN(n32985) );
  XOR2HSV0 U38297 ( .A1(n32986), .A2(n32985), .Z(n32987) );
  XOR2HSV0 U38298 ( .A1(n32988), .A2(n32987), .Z(n32989) );
  XOR2HSV0 U38299 ( .A1(n32990), .A2(n32989), .Z(n33013) );
  NAND2HSV0 U38300 ( .A1(n59240), .A2(n32991), .ZN(n32994) );
  NAND2HSV0 U38301 ( .A1(n32992), .A2(\pe6/aot [11]), .ZN(n32993) );
  XOR2HSV0 U38302 ( .A1(n32994), .A2(n32993), .Z(n32998) );
  NAND2HSV0 U38303 ( .A1(n35761), .A2(n36153), .ZN(n32996) );
  NAND2HSV0 U38304 ( .A1(n59206), .A2(\pe6/aot [17]), .ZN(n32995) );
  XOR2HSV0 U38305 ( .A1(n32996), .A2(n32995), .Z(n32997) );
  XOR2HSV0 U38306 ( .A1(n32998), .A2(n32997), .Z(n33011) );
  NAND2HSV0 U38307 ( .A1(n32999), .A2(n49208), .ZN(n33002) );
  NAND2HSV0 U38308 ( .A1(n33000), .A2(n46677), .ZN(n33001) );
  XOR2HSV0 U38309 ( .A1(n33002), .A2(n33001), .Z(n33009) );
  NAND2HSV0 U38310 ( .A1(n33003), .A2(n35726), .ZN(n33007) );
  NAND2HSV0 U38311 ( .A1(n33005), .A2(n33004), .ZN(n33006) );
  XOR2HSV0 U38312 ( .A1(n33007), .A2(n33006), .Z(n33008) );
  XOR2HSV0 U38313 ( .A1(n33009), .A2(n33008), .Z(n33010) );
  XOR2HSV0 U38314 ( .A1(n33011), .A2(n33010), .Z(n33012) );
  XOR2HSV0 U38315 ( .A1(n33013), .A2(n33012), .Z(n33038) );
  NAND2HSV0 U38316 ( .A1(n59201), .A2(\pe6/pvq [23]), .ZN(n33015) );
  NAND2HSV0 U38317 ( .A1(n59217), .A2(n59189), .ZN(n33014) );
  XOR2HSV0 U38318 ( .A1(n33015), .A2(n33014), .Z(n33033) );
  NAND2HSV0 U38319 ( .A1(n33016), .A2(n44393), .ZN(n33017) );
  XOR2HSV0 U38320 ( .A1(n33017), .A2(\pe6/phq [23]), .Z(n33021) );
  NAND2HSV0 U38321 ( .A1(n44336), .A2(\pe6/aot [13]), .ZN(n49853) );
  OAI22HSV0 U38322 ( .A1(n31253), .A2(n49680), .B1(n36124), .B2(n58983), .ZN(
        n33018) );
  OAI21HSV0 U38323 ( .A1(n33019), .A2(n49853), .B(n33018), .ZN(n33020) );
  XNOR2HSV1 U38324 ( .A1(n33021), .A2(n33020), .ZN(n33032) );
  NAND2HSV0 U38325 ( .A1(n33023), .A2(n33022), .ZN(n33026) );
  NAND2HSV0 U38326 ( .A1(n59267), .A2(n33024), .ZN(n33025) );
  XOR2HSV0 U38327 ( .A1(n33026), .A2(n33025), .Z(n33030) );
  NAND2HSV0 U38328 ( .A1(n58668), .A2(n58991), .ZN(n33028) );
  NAND2HSV0 U38329 ( .A1(n59100), .A2(n44439), .ZN(n33027) );
  XOR2HSV0 U38330 ( .A1(n33028), .A2(n33027), .Z(n33029) );
  XOR2HSV0 U38331 ( .A1(n33030), .A2(n33029), .Z(n33031) );
  XOR3HSV2 U38332 ( .A1(n33033), .A2(n33032), .A3(n33031), .Z(n33036) );
  NAND2HSV0 U38333 ( .A1(n35725), .A2(n33034), .ZN(n33035) );
  XNOR2HSV1 U38334 ( .A1(n33036), .A2(n33035), .ZN(n33037) );
  XOR2HSV0 U38335 ( .A1(n33038), .A2(n33037), .Z(n33044) );
  NAND2HSV0 U38336 ( .A1(n35724), .A2(n58654), .ZN(n33041) );
  NAND2HSV0 U38337 ( .A1(n32286), .A2(n33039), .ZN(n33040) );
  XOR2HSV0 U38338 ( .A1(n33041), .A2(n33040), .Z(n33043) );
  NAND2HSV0 U38339 ( .A1(n59121), .A2(n35991), .ZN(n33042) );
  XOR3HSV2 U38340 ( .A1(n33044), .A2(n33043), .A3(n33042), .Z(n33046) );
  NAND2HSV0 U38341 ( .A1(n59295), .A2(\pe6/got [15]), .ZN(n33045) );
  XNOR2HSV1 U38342 ( .A1(n33046), .A2(n33045), .ZN(n33047) );
  XNOR2HSV1 U38343 ( .A1(n33048), .A2(n33047), .ZN(n33049) );
  XNOR2HSV1 U38344 ( .A1(n33050), .A2(n33049), .ZN(n33052) );
  NAND2HSV0 U38345 ( .A1(n36185), .A2(n58715), .ZN(n33051) );
  XNOR2HSV1 U38346 ( .A1(n33052), .A2(n33051), .ZN(n33053) );
  XOR2HSV0 U38347 ( .A1(n33054), .A2(n33053), .Z(n33055) );
  XNOR2HSV1 U38348 ( .A1(n33056), .A2(n33055), .ZN(n33057) );
  XOR2HSV0 U38349 ( .A1(n33058), .A2(n33057), .Z(n33059) );
  CLKBUFHSV4 U38350 ( .I(n46592), .Z(n36102) );
  CLKNAND2HSV1 U38351 ( .A1(n46589), .A2(n44519), .ZN(n33062) );
  AOI21HSV2 U38352 ( .A1(n33078), .A2(n33076), .B(n33062), .ZN(n33065) );
  INHSV2 U38353 ( .I(n33078), .ZN(n46590) );
  CLKAND2HSV2 U38354 ( .A1(n46588), .A2(n51438), .Z(n33077) );
  CLKNAND2HSV1 U38355 ( .A1(n46590), .A2(n33077), .ZN(n33064) );
  CLKNAND2HSV1 U38356 ( .A1(n33065), .A2(n33064), .ZN(n33066) );
  AOI21HSV2 U38357 ( .A1(n51451), .A2(n33067), .B(n33066), .ZN(n33074) );
  XNOR2HSV4 U38358 ( .A1(n33069), .A2(n33068), .ZN(n33085) );
  CLKNAND2HSV3 U38359 ( .A1(n33074), .A2(n33073), .ZN(n35904) );
  NOR2HSV4 U38360 ( .A1(n33084), .A2(n36066), .ZN(n33075) );
  INAND2HSV2 U38361 ( .A1(n33078), .B1(n33076), .ZN(n33082) );
  NAND2HSV2 U38362 ( .A1(n33078), .A2(n33077), .ZN(n33081) );
  NOR2HSV2 U38363 ( .A1(n46589), .A2(n33079), .ZN(n33080) );
  AOI21HSV4 U38364 ( .A1(n33085), .A2(n25855), .B(n33083), .ZN(n35708) );
  NAND2HSV2 U38365 ( .A1(n44369), .A2(\pe6/ti_7t [23]), .ZN(n35903) );
  NAND3HSV4 U38366 ( .A1(n35904), .A2(n35709), .A3(n35903), .ZN(n33086) );
  CLKNAND2HSV4 U38367 ( .A1(n33086), .A2(n31624), .ZN(n33088) );
  CLKNAND2HSV1 U38368 ( .A1(n32941), .A2(\pe6/ti_7t [24]), .ZN(n36024) );
  INHSV2 U38369 ( .I(n36024), .ZN(n36030) );
  AOI21HSV4 U38370 ( .A1(n33087), .A2(n35719), .B(n36030), .ZN(n36206) );
  INHSV4 U38371 ( .I(\pe2/aot [28]), .ZN(n44212) );
  INHSV2 U38372 ( .I(n44212), .ZN(n59759) );
  INHSV2 U38373 ( .I(n33687), .ZN(n33093) );
  CLKNHSV2 U38374 ( .I(n33779), .ZN(n33339) );
  CLKNHSV0 U38375 ( .I(\pe4/ti_7t [9]), .ZN(n33340) );
  INHSV2 U38376 ( .I(n33785), .ZN(n59997) );
  INHSV4 U38377 ( .I(\pe4/ctrq ), .ZN(n33090) );
  CLKNHSV2 U38378 ( .I(n33095), .ZN(n34983) );
  CLKBUFHSV4 U38379 ( .I(\pe4/bq[32] ), .Z(n33249) );
  INHSV4 U38380 ( .I(\pe4/aot [31]), .ZN(n33114) );
  INHSV2 U38381 ( .I(\pe4/aot [32]), .ZN(n33893) );
  BUFHSV2 U38382 ( .I(n33184), .Z(n33457) );
  INHSV2 U38383 ( .I(n33457), .ZN(n34203) );
  INHSV2 U38384 ( .I(n33785), .ZN(n33849) );
  NOR2HSV4 U38385 ( .A1(n33118), .A2(n33098), .ZN(n33100) );
  NAND2HSV2 U38386 ( .A1(\pe4/aot [32]), .A2(\pe4/bq[30] ), .ZN(n33099) );
  XNOR2HSV4 U38387 ( .A1(n33100), .A2(n33099), .ZN(n33102) );
  INHSV2 U38388 ( .I(n34631), .ZN(n57106) );
  CLKBUFHSV4 U38389 ( .I(\pe4/bq[32] ), .Z(n35075) );
  NAND2HSV2 U38390 ( .A1(n57106), .A2(n35075), .ZN(n33105) );
  NAND2HSV2 U38391 ( .A1(n57242), .A2(n33103), .ZN(n33104) );
  XOR2HSV0 U38392 ( .A1(n33105), .A2(n33104), .Z(n33106) );
  CLKBUFHSV4 U38393 ( .I(n33189), .Z(n34328) );
  CLKNHSV2 U38394 ( .I(n33779), .ZN(n33403) );
  NOR2HSV4 U38395 ( .A1(n34226), .A2(n33403), .ZN(n33997) );
  INHSV2 U38396 ( .I(n33696), .ZN(n35283) );
  NAND2HSV2 U38397 ( .A1(n29766), .A2(n35283), .ZN(n33107) );
  BUFHSV2 U38398 ( .I(n33687), .Z(n35311) );
  INHSV2 U38399 ( .I(n33184), .ZN(n47778) );
  OAI21HSV2 U38400 ( .A1(n35311), .A2(\pe4/ti_7t [3]), .B(n47778), .ZN(n33109)
         );
  INHSV2 U38401 ( .I(n34631), .ZN(n33624) );
  INHSV2 U38402 ( .I(n33112), .ZN(n33110) );
  NAND2HSV4 U38403 ( .A1(n33624), .A2(n33110), .ZN(n33203) );
  INHSV2 U38404 ( .I(n33103), .ZN(n33113) );
  CLKBUFHSV4 U38405 ( .I(n33112), .Z(n34117) );
  INHSV4 U38406 ( .I(\pe4/aot [32]), .ZN(n33355) );
  XNOR2HSV1 U38407 ( .A1(n33117), .A2(n33116), .ZN(n33124) );
  INHSV4 U38408 ( .I(\pe4/got [29]), .ZN(n57199) );
  BUFHSV8 U38409 ( .I(n57199), .Z(n34187) );
  INHSV2 U38410 ( .I(n34187), .ZN(n33215) );
  INHSV2 U38411 ( .I(n34479), .ZN(n59834) );
  NAND2HSV2 U38412 ( .A1(n59834), .A2(n35075), .ZN(n33119) );
  XNOR2HSV4 U38413 ( .A1(n33120), .A2(n33119), .ZN(n33122) );
  CLKBUFHSV4 U38414 ( .I(n48082), .Z(n34138) );
  NAND2HSV2 U38415 ( .A1(n34138), .A2(\pe4/pvq [4]), .ZN(n33121) );
  XNOR2HSV4 U38416 ( .A1(n33122), .A2(n33121), .ZN(n33123) );
  XNOR2HSV4 U38417 ( .A1(n33124), .A2(n33123), .ZN(n33126) );
  INHSV2 U38418 ( .I(\pe4/ti_7t [1]), .ZN(n33151) );
  NOR2HSV4 U38419 ( .A1(n33785), .A2(n33151), .ZN(n33175) );
  INHSV2 U38420 ( .I(\pe4/got [30]), .ZN(n34851) );
  INHSV2 U38421 ( .I(n34851), .ZN(n59955) );
  CLKBUFHSV4 U38422 ( .I(n33153), .Z(n59577) );
  INHSV2 U38423 ( .I(\pe4/got [30]), .ZN(n34108) );
  BUFHSV4 U38424 ( .I(n33097), .Z(n33522) );
  INHSV2 U38425 ( .I(n33522), .ZN(n33852) );
  NOR2HSV2 U38426 ( .A1(n34851), .A2(n33852), .ZN(n33982) );
  AOI22HSV4 U38427 ( .A1(n33175), .A2(n34017), .B1(n59577), .B2(n33982), .ZN(
        n33125) );
  XNOR2HSV4 U38428 ( .A1(n33126), .A2(n33125), .ZN(n33127) );
  INHSV2 U38429 ( .I(\pe4/got [31]), .ZN(n33282) );
  CLKNHSV1 U38430 ( .I(n33779), .ZN(n35316) );
  INHSV2 U38431 ( .I(n35316), .ZN(n34220) );
  INHSV2 U38432 ( .I(n33785), .ZN(n33774) );
  NAND2HSV2 U38433 ( .A1(\pe4/ti_7t [4]), .A2(n33774), .ZN(n33201) );
  INHSV2 U38434 ( .I(n57199), .ZN(n57208) );
  NAND2HSV2 U38435 ( .A1(n46611), .A2(n57208), .ZN(n33166) );
  CLKBUFHSV4 U38436 ( .I(n26218), .Z(n33307) );
  BUFHSV2 U38437 ( .I(n33175), .Z(n33130) );
  AOI21HSV4 U38438 ( .A1(n59577), .A2(n33687), .B(n33130), .ZN(n33308) );
  INHSV2 U38439 ( .I(n33308), .ZN(n33247) );
  INHSV4 U38440 ( .I(\pe4/got [26]), .ZN(n34456) );
  INHSV2 U38441 ( .I(n34456), .ZN(n33306) );
  CLKNAND2HSV1 U38442 ( .A1(n33247), .A2(n33306), .ZN(n33131) );
  INHSV2 U38443 ( .I(\pe4/bq[25] ), .ZN(n33325) );
  INHSV2 U38444 ( .I(n33325), .ZN(n33615) );
  NAND2HSV0 U38445 ( .A1(n33415), .A2(n33615), .ZN(n33133) );
  INHSV2 U38446 ( .I(n34631), .ZN(n59383) );
  CLKNAND2HSV1 U38447 ( .A1(n59383), .A2(n33427), .ZN(n33132) );
  XOR2HSV0 U38448 ( .A1(n33133), .A2(n33132), .Z(n33137) );
  INHSV2 U38449 ( .I(n57026), .ZN(n59838) );
  BUFHSV2 U38450 ( .I(n33249), .Z(n48074) );
  NAND2HSV2 U38451 ( .A1(n59838), .A2(n48074), .ZN(n33135) );
  INHSV2 U38452 ( .I(n33350), .ZN(n48071) );
  NAND2HSV0 U38453 ( .A1(n57242), .A2(n48071), .ZN(n33134) );
  XOR2HSV0 U38454 ( .A1(n33135), .A2(n33134), .Z(n33136) );
  XOR2HSV0 U38455 ( .A1(n33137), .A2(n33136), .Z(n33141) );
  INHSV2 U38456 ( .I(n34479), .ZN(n33420) );
  CLKNAND2HSV1 U38457 ( .A1(n33420), .A2(n48069), .ZN(n33138) );
  XNOR2HSV1 U38458 ( .A1(n33139), .A2(n33138), .ZN(n33140) );
  XNOR2HSV1 U38459 ( .A1(n33141), .A2(n33140), .ZN(n33149) );
  INHSV2 U38460 ( .I(n33250), .ZN(n59598) );
  NAND2HSV2 U38461 ( .A1(n59598), .A2(n33326), .ZN(n33143) );
  INHSV2 U38462 ( .I(n47661), .ZN(n59390) );
  BUFHSV2 U38463 ( .I(n33112), .Z(n33414) );
  INHSV2 U38464 ( .I(n33414), .ZN(n33313) );
  CLKNAND2HSV1 U38465 ( .A1(n59390), .A2(n33313), .ZN(n33142) );
  XOR2HSV0 U38466 ( .A1(n33143), .A2(n33142), .Z(n33147) );
  INHSV4 U38467 ( .I(\pe4/aot [26]), .ZN(n57509) );
  INHSV2 U38468 ( .I(n57509), .ZN(n33614) );
  INHSV2 U38469 ( .I(n33113), .ZN(n33423) );
  NAND2HSV2 U38470 ( .A1(n33614), .A2(n33423), .ZN(n33145) );
  NAND2HSV0 U38471 ( .A1(n57190), .A2(n35370), .ZN(n33144) );
  XOR2HSV0 U38472 ( .A1(n33145), .A2(n33144), .Z(n33146) );
  XOR2HSV0 U38473 ( .A1(n33147), .A2(n33146), .Z(n33148) );
  XNOR2HSV1 U38474 ( .A1(n33149), .A2(n33148), .ZN(n33150) );
  AOI21HSV2 U38475 ( .A1(n33151), .A2(n33156), .B(n34328), .ZN(n33152) );
  NAND2HSV2 U38476 ( .A1(n33155), .A2(n33154), .ZN(n33160) );
  INHSV4 U38477 ( .I(n26218), .ZN(n33463) );
  INHSV4 U38478 ( .I(n33463), .ZN(n33181) );
  BUFHSV2 U38479 ( .I(n33687), .Z(n35604) );
  NOR2HSV2 U38480 ( .A1(n47778), .A2(n59997), .ZN(n35013) );
  INHSV2 U38481 ( .I(n35013), .ZN(n33387) );
  OAI21HSV4 U38482 ( .A1(n33159), .A2(n33158), .B(n33387), .ZN(n33162) );
  CLKNAND2HSV3 U38483 ( .A1(n33162), .A2(n52699), .ZN(n33164) );
  INHSV2 U38484 ( .I(n33779), .ZN(n34566) );
  NAND2HSV2 U38485 ( .A1(n34566), .A2(\pe4/ti_7t [3]), .ZN(n33163) );
  XOR2HSV2 U38486 ( .A1(n33166), .A2(n33165), .Z(n33197) );
  CLKNHSV0 U38487 ( .I(n34220), .ZN(n33167) );
  NOR2HSV4 U38488 ( .A1(n59578), .A2(n33167), .ZN(n33196) );
  NAND2HSV2 U38489 ( .A1(n29650), .A2(n33181), .ZN(n33168) );
  BUFHSV2 U38490 ( .I(n33189), .Z(n34712) );
  INHSV2 U38491 ( .I(n34712), .ZN(n33169) );
  INHSV2 U38492 ( .I(n33785), .ZN(n35294) );
  CLKNHSV2 U38493 ( .I(n33170), .ZN(n33171) );
  INHSV4 U38494 ( .I(n33114), .ZN(n59523) );
  INHSV2 U38495 ( .I(n34117), .ZN(n57254) );
  NAND2HSV2 U38496 ( .A1(n34138), .A2(\pe4/pvq [5]), .ZN(n33174) );
  INHSV2 U38497 ( .I(n33538), .ZN(n33248) );
  INHSV2 U38498 ( .I(n33355), .ZN(n59485) );
  NOR2HSV2 U38499 ( .A1(n59577), .A2(n33175), .ZN(n33177) );
  BUFHSV2 U38500 ( .I(n33785), .Z(n34834) );
  OAI21HSV2 U38501 ( .A1(n33175), .A2(n34834), .B(n57208), .ZN(n33176) );
  AOI21HSV4 U38502 ( .A1(n33181), .A2(n29650), .B(n33180), .ZN(n33218) );
  NAND2HSV0 U38503 ( .A1(n33218), .A2(n33170), .ZN(n33183) );
  CLKNAND2HSV1 U38504 ( .A1(n33170), .A2(n34718), .ZN(n33182) );
  INHSV2 U38505 ( .I(n33774), .ZN(n35021) );
  INHSV2 U38506 ( .I(n33184), .ZN(n33676) );
  OAI21HSV2 U38507 ( .A1(n35311), .A2(\pe4/ti_7t [4]), .B(n33676), .ZN(n33185)
         );
  INHSV2 U38508 ( .I(n33185), .ZN(n33188) );
  OR2HSV1 U38509 ( .A1(n33188), .A2(n33171), .Z(n33186) );
  OA21HSV2 U38510 ( .A1(n33171), .A2(n35021), .B(n33186), .Z(n33187) );
  INHSV2 U38511 ( .I(n33188), .ZN(n33290) );
  BUFHSV2 U38512 ( .I(n33189), .Z(n35286) );
  CLKNHSV2 U38513 ( .I(n35286), .ZN(n33190) );
  INHSV2 U38514 ( .I(n33292), .ZN(n33191) );
  NAND2HSV2 U38515 ( .A1(n33191), .A2(n29740), .ZN(n33193) );
  INHSV2 U38516 ( .I(n34571), .ZN(n33695) );
  CLKNHSV2 U38517 ( .I(n33695), .ZN(n33192) );
  INHSV2 U38518 ( .I(n25856), .ZN(n33498) );
  INHSV2 U38519 ( .I(n34108), .ZN(n33507) );
  INHSV4 U38520 ( .I(n33198), .ZN(n33200) );
  NOR2HSV4 U38521 ( .A1(n33200), .A2(n33199), .ZN(n33246) );
  CLKNAND2HSV1 U38522 ( .A1(n33201), .A2(n33774), .ZN(n33245) );
  INHSV2 U38523 ( .I(n33282), .ZN(n35274) );
  NAND2HSV2 U38524 ( .A1(n33245), .A2(n35274), .ZN(n33202) );
  NOR2HSV4 U38525 ( .A1(n33246), .A2(n33202), .ZN(n33237) );
  INHSV2 U38526 ( .I(n47661), .ZN(n33474) );
  XNOR2HSV4 U38527 ( .A1(n33203), .A2(\pe4/phq [6]), .ZN(n33205) );
  CLKBUFHSV4 U38528 ( .I(\pe4/ctrq ), .Z(n34496) );
  CLKBUFHSV4 U38529 ( .I(n34496), .Z(n34770) );
  NAND2HSV2 U38530 ( .A1(n34770), .A2(\pe4/pvq [6]), .ZN(n33204) );
  XNOR2HSV4 U38531 ( .A1(n33205), .A2(n33204), .ZN(n33206) );
  XNOR2HSV4 U38532 ( .A1(n33207), .A2(n33206), .ZN(n33212) );
  INHSV2 U38533 ( .I(n33250), .ZN(n57510) );
  NAND2HSV0 U38534 ( .A1(n59834), .A2(n33816), .ZN(n33209) );
  CLKNAND2HSV1 U38535 ( .A1(n59485), .A2(n33427), .ZN(n33208) );
  XNOR2HSV4 U38536 ( .A1(n33212), .A2(n33211), .ZN(n33214) );
  CLKNAND2HSV1 U38537 ( .A1(n33247), .A2(n33263), .ZN(n33213) );
  XOR2HSV2 U38538 ( .A1(n33214), .A2(n33213), .Z(n33217) );
  CLKNAND2HSV3 U38539 ( .A1(n33307), .A2(n33215), .ZN(n33216) );
  XNOR2HSV4 U38540 ( .A1(n33217), .A2(n33216), .ZN(n33219) );
  CLKNAND2HSV3 U38541 ( .A1(n57166), .A2(n33507), .ZN(n33220) );
  INHSV2 U38542 ( .I(n33220), .ZN(n33221) );
  XNOR2HSV4 U38543 ( .A1(n33237), .A2(n33238), .ZN(n33344) );
  AND2HSV2 U38544 ( .A1(n33344), .A2(n34983), .Z(n33230) );
  NOR2HSV4 U38545 ( .A1(n33344), .A2(n33852), .ZN(n33225) );
  NAND2HSV4 U38546 ( .A1(n33240), .A2(n33225), .ZN(n33243) );
  INHSV2 U38547 ( .I(n35274), .ZN(n35303) );
  INHSV2 U38548 ( .I(n35303), .ZN(n34428) );
  NAND2HSV2 U38549 ( .A1(n33226), .A2(n34428), .ZN(n33227) );
  IAO21HSV4 U38550 ( .A1(n33344), .A2(n33387), .B(n33227), .ZN(n33228) );
  CLKNAND2HSV2 U38551 ( .A1(n33243), .A2(n33228), .ZN(n33229) );
  AOI21HSV2 U38552 ( .A1(n33498), .A2(n33230), .B(n33229), .ZN(n33232) );
  CLKNAND2HSV1 U38553 ( .A1(n33231), .A2(n33232), .ZN(n33236) );
  INHSV2 U38554 ( .I(n33232), .ZN(n33233) );
  CLKNAND2HSV4 U38555 ( .A1(n33236), .A2(n33235), .ZN(n33391) );
  CLKBUFHSV3 U38556 ( .I(n33391), .Z(n46607) );
  XNOR2HSV4 U38557 ( .A1(n33239), .A2(n33238), .ZN(n52725) );
  NOR2HSV4 U38558 ( .A1(n52725), .A2(n34565), .ZN(n33242) );
  CLKNAND2HSV2 U38559 ( .A1(n33226), .A2(n52723), .ZN(n33241) );
  AOI21HSV4 U38560 ( .A1(n33242), .A2(n33224), .B(n33241), .ZN(n33244) );
  CLKNHSV4 U38561 ( .I(n52731), .ZN(n33284) );
  CLKNAND2HSV1 U38562 ( .A1(n33247), .A2(n33748), .ZN(n33266) );
  NAND2HSV2 U38563 ( .A1(n33313), .A2(n33631), .ZN(n34355) );
  CLKNAND2HSV1 U38564 ( .A1(n59383), .A2(n33248), .ZN(n57343) );
  XOR2HSV0 U38565 ( .A1(n34355), .A2(n57343), .Z(n33255) );
  INHSV2 U38566 ( .I(n57509), .ZN(n57327) );
  INHSV2 U38567 ( .I(n35084), .ZN(n33621) );
  NAND2HSV2 U38568 ( .A1(n34054), .A2(\pe4/pvq [7]), .ZN(n33256) );
  XNOR2HSV1 U38569 ( .A1(n33256), .A2(\pe4/phq [7]), .ZN(n33260) );
  NAND2HSV2 U38570 ( .A1(n59390), .A2(n33326), .ZN(n33258) );
  NAND2HSV0 U38571 ( .A1(n33415), .A2(n48071), .ZN(n33257) );
  XOR2HSV0 U38572 ( .A1(n33258), .A2(n33257), .Z(n33259) );
  XNOR2HSV1 U38573 ( .A1(n33260), .A2(n33259), .ZN(n33261) );
  CLKXOR2HSV4 U38574 ( .A1(n33262), .A2(n33261), .Z(n33265) );
  XOR3HSV2 U38575 ( .A1(n33266), .A2(n33265), .A3(n33264), .Z(n33268) );
  XNOR2HSV4 U38576 ( .A1(n33268), .A2(n33267), .ZN(n33269) );
  XNOR2HSV4 U38577 ( .A1(n33270), .A2(n33269), .ZN(n52729) );
  MUX2NHSV2 U38578 ( .I0(n52730), .I1(n33694), .S(n52729), .ZN(n33272) );
  CLKXOR2HSV4 U38579 ( .A1(n33270), .A2(n33269), .Z(n33273) );
  OAI21HSV2 U38580 ( .A1(n33273), .A2(n29780), .B(n33588), .ZN(n33271) );
  NOR2HSV4 U38581 ( .A1(n33272), .A2(n33271), .ZN(n33283) );
  CLKNHSV0 U38582 ( .I(n33282), .ZN(n34436) );
  MUX2NHSV2 U38583 ( .I0(n52730), .I1(n34436), .S(n33273), .ZN(n33275) );
  OAI21HSV2 U38584 ( .A1(n52729), .A2(n29780), .B(n33588), .ZN(n33274) );
  NOR2HSV4 U38585 ( .A1(n33275), .A2(n33274), .ZN(n33279) );
  NAND2HSV2 U38586 ( .A1(n35294), .A2(\pe4/ti_7t [8]), .ZN(n33389) );
  CLKNAND2HSV3 U38587 ( .A1(n46607), .A2(n29676), .ZN(n33276) );
  CLKNHSV1 U38588 ( .I(n33527), .ZN(n33278) );
  INHSV4 U38589 ( .I(n33391), .ZN(n33394) );
  NAND3HSV3 U38590 ( .A1(n33394), .A2(n33389), .A3(n33393), .ZN(n33516) );
  CLKNAND2HSV1 U38591 ( .A1(n33278), .A2(n33516), .ZN(n33338) );
  INHSV2 U38592 ( .I(n33279), .ZN(n33280) );
  INHSV2 U38593 ( .I(n33280), .ZN(n33289) );
  NAND2HSV0 U38594 ( .A1(n52731), .A2(n33796), .ZN(n33281) );
  INHSV2 U38595 ( .I(n33281), .ZN(n33288) );
  CLKNHSV1 U38596 ( .I(n33282), .ZN(n33796) );
  NAND3HSV4 U38597 ( .A1(n33284), .A2(n33283), .A3(n33796), .ZN(n33286) );
  NAND2HSV2 U38598 ( .A1(n47788), .A2(\pe4/ti_7t [7]), .ZN(n33382) );
  INHSV2 U38599 ( .I(n33382), .ZN(n33411) );
  CLKNAND2HSV1 U38600 ( .A1(n33411), .A2(n47773), .ZN(n33285) );
  CLKNAND2HSV3 U38601 ( .A1(n33286), .A2(n33285), .ZN(n33287) );
  AOI21HSV4 U38602 ( .A1(n33289), .A2(n33288), .B(n33287), .ZN(n33337) );
  NOR2HSV4 U38603 ( .A1(n33291), .A2(n33290), .ZN(n33293) );
  INHSV2 U38604 ( .I(n33097), .ZN(n34423) );
  AOI21HSV2 U38605 ( .A1(n60082), .A2(n25420), .B(n34423), .ZN(n33345) );
  INHSV1 U38606 ( .I(n33345), .ZN(n33295) );
  CLKNHSV2 U38607 ( .I(n52725), .ZN(n33341) );
  CLKNAND2HSV2 U38608 ( .A1(n33341), .A2(n35445), .ZN(n33294) );
  NOR2HSV2 U38609 ( .A1(n33295), .A2(n33294), .ZN(n33305) );
  INHSV1 U38610 ( .I(n33305), .ZN(n33299) );
  NAND2HSV2 U38611 ( .A1(n60082), .A2(n33277), .ZN(n33342) );
  CLKNHSV0 U38612 ( .I(n34108), .ZN(n33801) );
  INAND2HSV2 U38613 ( .A1(n33342), .B1(n33801), .ZN(n33303) );
  INHSV1 U38614 ( .I(n33303), .ZN(n33296) );
  CLKBUFHSV2 U38615 ( .I(n52725), .Z(n33300) );
  CLKNAND2HSV0 U38616 ( .A1(\pe4/ti_7t [6]), .A2(n33774), .ZN(n33346) );
  CLKNHSV0 U38617 ( .I(n33346), .ZN(n33297) );
  NAND2HSV2 U38618 ( .A1(n33297), .A2(n33507), .ZN(n33301) );
  CLKNHSV1 U38619 ( .I(n52725), .ZN(n33302) );
  OAI21HSV2 U38620 ( .A1(n33303), .A2(n33302), .B(n33301), .ZN(n33304) );
  NOR2HSV2 U38621 ( .A1(n33305), .A2(n33304), .ZN(n33334) );
  BUFHSV2 U38622 ( .I(n59956), .Z(n35598) );
  CLKNAND2HSV1 U38623 ( .A1(n29781), .A2(n35598), .ZN(n33332) );
  INHSV2 U38624 ( .I(n33564), .ZN(n33461) );
  NAND2HSV2 U38625 ( .A1(n33307), .A2(n33306), .ZN(n33310) );
  BUFHSV2 U38626 ( .I(n33308), .Z(n33464) );
  BUFHSV2 U38627 ( .I(n33859), .Z(n50314) );
  NOR2HSV2 U38628 ( .A1(n33464), .A2(n50314), .ZN(n33309) );
  CLKNAND2HSV1 U38629 ( .A1(n57727), .A2(n48074), .ZN(n33312) );
  INHSV2 U38630 ( .I(n33350), .ZN(n33713) );
  CLKNAND2HSV0 U38631 ( .A1(n59383), .A2(n33713), .ZN(n33311) );
  XOR2HSV0 U38632 ( .A1(n33312), .A2(n33311), .Z(n33317) );
  NAND2HSV0 U38633 ( .A1(n33420), .A2(n33427), .ZN(n33315) );
  CLKNAND2HSV0 U38634 ( .A1(n59598), .A2(n33313), .ZN(n33314) );
  XOR2HSV0 U38635 ( .A1(n33315), .A2(n33314), .Z(n33316) );
  XOR2HSV0 U38636 ( .A1(n33317), .A2(n33316), .Z(n33324) );
  NAND2HSV0 U38637 ( .A1(n33415), .A2(\pe4/bq[24] ), .ZN(n33319) );
  NAND2HSV0 U38638 ( .A1(n33474), .A2(n48069), .ZN(n33318) );
  XOR2HSV0 U38639 ( .A1(n33319), .A2(n33318), .Z(n33322) );
  CLKNAND2HSV1 U38640 ( .A1(n33808), .A2(\pe4/pvq [9]), .ZN(n33320) );
  XOR2HSV0 U38641 ( .A1(n33320), .A2(\pe4/phq [9]), .Z(n33321) );
  XOR2HSV0 U38642 ( .A1(n33322), .A2(n33321), .Z(n33323) );
  XOR2HSV0 U38643 ( .A1(n33324), .A2(n33323), .Z(n33328) );
  INHSV2 U38644 ( .I(n33325), .ZN(n34030) );
  INHSV2 U38645 ( .I(n57026), .ZN(n57499) );
  NAND2HSV2 U38646 ( .A1(n57499), .A2(n33423), .ZN(n34145) );
  INHSV2 U38647 ( .I(n57509), .ZN(n59661) );
  XNOR2HSV1 U38648 ( .A1(n33328), .A2(n33327), .ZN(n33329) );
  CLKNAND2HSV1 U38649 ( .A1(n34043), .A2(n59350), .ZN(n33330) );
  XNOR2HSV4 U38650 ( .A1(n33332), .A2(n33331), .ZN(n33333) );
  NOR2HSV4 U38651 ( .A1(n33337), .A2(n25880), .ZN(n33405) );
  XNOR2HSV1 U38652 ( .A1(n33338), .A2(n33518), .ZN(n60038) );
  NOR2HSV2 U38653 ( .A1(n33342), .A2(n33341), .ZN(n33343) );
  BUFHSV2 U38654 ( .I(n33413), .Z(n50266) );
  CLKNAND2HSV0 U38655 ( .A1(n50266), .A2(\pe4/got [24]), .ZN(n33381) );
  BUFHSV2 U38656 ( .I(n46611), .Z(n57325) );
  BUFHSV2 U38657 ( .I(n57325), .Z(n34109) );
  CLKNAND2HSV0 U38658 ( .A1(n34109), .A2(n59601), .ZN(n33377) );
  INHSV4 U38659 ( .I(\pe4/bq[23] ), .ZN(n50248) );
  BUFHSV2 U38660 ( .I(n50248), .Z(n48056) );
  CLKNAND2HSV0 U38661 ( .A1(n35377), .A2(n57368), .ZN(n34148) );
  NAND2HSV0 U38662 ( .A1(n33808), .A2(\pe4/pvq [15]), .ZN(n33347) );
  CLKNHSV0 U38663 ( .I(n34117), .ZN(n57377) );
  CLKNAND2HSV1 U38664 ( .A1(n59839), .A2(n57377), .ZN(n33813) );
  INHSV2 U38665 ( .I(n34485), .ZN(n33816) );
  NAND2HSV2 U38666 ( .A1(n59951), .A2(n33816), .ZN(n33710) );
  BUFHSV2 U38667 ( .I(n34117), .Z(n35043) );
  OAI22HSV0 U38668 ( .A1(n34485), .A2(n49982), .B1(n50008), .B2(n35043), .ZN(
        n33348) );
  OAI21HSV0 U38669 ( .A1(n33813), .A2(n33710), .B(n33348), .ZN(n33349) );
  NAND2HSV0 U38670 ( .A1(n59390), .A2(n33711), .ZN(n33352) );
  INHSV2 U38671 ( .I(\pe4/aot [24]), .ZN(n33467) );
  INHSV2 U38672 ( .I(n33350), .ZN(n34629) );
  NAND2HSV0 U38673 ( .A1(n33726), .A2(n34629), .ZN(n33351) );
  BUFHSV2 U38674 ( .I(n35084), .Z(n57260) );
  NAND2HSV0 U38675 ( .A1(n33716), .A2(n34598), .ZN(n33354) );
  INHSV2 U38676 ( .I(n33830), .ZN(n59372) );
  CLKNHSV0 U38677 ( .I(n46618), .ZN(n57157) );
  NAND2HSV0 U38678 ( .A1(n59372), .A2(n57157), .ZN(n33353) );
  BUFHSV4 U38679 ( .I(n34285), .Z(n57359) );
  INHSV2 U38680 ( .I(n33860), .ZN(n33831) );
  NAND2HSV0 U38681 ( .A1(n33965), .A2(n33966), .ZN(n33357) );
  BUFHSV2 U38682 ( .I(n33355), .Z(n34501) );
  INHSV2 U38683 ( .I(n48026), .ZN(n34359) );
  CLKNAND2HSV0 U38684 ( .A1(n35201), .A2(n34359), .ZN(n33356) );
  XOR2HSV0 U38685 ( .A1(n33357), .A2(n33356), .Z(n33361) );
  NAND2HSV0 U38686 ( .A1(n34240), .A2(n34030), .ZN(n33359) );
  INHSV2 U38687 ( .I(n57605), .ZN(n34047) );
  NAND2HSV0 U38688 ( .A1(n34047), .A2(n33611), .ZN(n33358) );
  XOR2HSV0 U38689 ( .A1(n33359), .A2(n33358), .Z(n33360) );
  XOR2HSV0 U38690 ( .A1(n33361), .A2(n33360), .Z(n33369) );
  CLKNHSV0 U38691 ( .I(\pe4/aot [26]), .ZN(n34249) );
  INHSV2 U38692 ( .I(n34249), .ZN(n33947) );
  CLKNAND2HSV0 U38693 ( .A1(n33947), .A2(n34120), .ZN(n33363) );
  CLKNHSV0 U38694 ( .I(n34631), .ZN(n33960) );
  INHSV2 U38695 ( .I(n48023), .ZN(n34243) );
  NAND2HSV0 U38696 ( .A1(n33960), .A2(n34243), .ZN(n33362) );
  XOR2HSV0 U38697 ( .A1(n33363), .A2(n33362), .Z(n33367) );
  CLKNHSV1 U38698 ( .I(n34479), .ZN(n33631) );
  NAND2HSV0 U38699 ( .A1(n33631), .A2(n33969), .ZN(n33365) );
  BUFHSV2 U38700 ( .I(n35075), .Z(n34888) );
  CLKNAND2HSV0 U38701 ( .A1(\pe4/aot [18]), .A2(n33934), .ZN(n33364) );
  XOR2HSV0 U38702 ( .A1(n33365), .A2(n33364), .Z(n33366) );
  XOR2HSV0 U38703 ( .A1(n33367), .A2(n33366), .Z(n33368) );
  XOR2HSV0 U38704 ( .A1(n33369), .A2(n33368), .Z(n33371) );
  CLKNHSV0 U38705 ( .I(n33464), .ZN(n33976) );
  CLKNAND2HSV0 U38706 ( .A1(n33976), .A2(n59602), .ZN(n33370) );
  XNOR2HSV1 U38707 ( .A1(n33371), .A2(n33370), .ZN(n33372) );
  XNOR2HSV1 U38708 ( .A1(n33373), .A2(n33372), .ZN(n33375) );
  CLKNHSV0 U38709 ( .I(n35501), .ZN(n35340) );
  CLKNAND2HSV1 U38710 ( .A1(n35340), .A2(n34948), .ZN(n33374) );
  XNOR2HSV1 U38711 ( .A1(n33375), .A2(n33374), .ZN(n33376) );
  XNOR2HSV1 U38712 ( .A1(n33377), .A2(n33376), .ZN(n33379) );
  CLKNAND2HSV0 U38713 ( .A1(n59662), .A2(n59369), .ZN(n33378) );
  XNOR2HSV1 U38714 ( .A1(n33379), .A2(n33378), .ZN(n33380) );
  XNOR2HSV1 U38715 ( .A1(n33381), .A2(n33380), .ZN(n33386) );
  BUFHSV2 U38716 ( .I(n45806), .Z(n34595) );
  INHSV2 U38717 ( .I(n33859), .ZN(n34672) );
  CLKNAND2HSV1 U38718 ( .A1(n34595), .A2(n34672), .ZN(n33385) );
  XNOR2HSV1 U38719 ( .A1(n33386), .A2(n33385), .ZN(n33397) );
  INHSV2 U38720 ( .I(n33389), .ZN(n33390) );
  AOI21HSV4 U38721 ( .A1(n33392), .A2(n33391), .B(n33390), .ZN(n33505) );
  CLKNAND2HSV4 U38722 ( .A1(n33395), .A2(n33394), .ZN(n33506) );
  CLKNAND2HSV3 U38723 ( .A1(n33505), .A2(n33506), .ZN(n33565) );
  INHSV3 U38724 ( .I(n33565), .ZN(n44697) );
  CLKBUFHSV2 U38725 ( .I(n44697), .Z(n33750) );
  CLKNHSV0 U38726 ( .I(n33708), .ZN(n35587) );
  OR2HSV1 U38727 ( .A1(n33750), .A2(n35587), .Z(n33396) );
  XOR2HSV0 U38728 ( .A1(n33397), .A2(n33396), .Z(n33398) );
  XNOR2HSV1 U38729 ( .A1(n33399), .A2(n33398), .ZN(n33455) );
  NOR2HSV4 U38730 ( .A1(n33400), .A2(n35295), .ZN(n33402) );
  NOR2HSV2 U38731 ( .A1(n33588), .A2(\pe4/ti_7t [9]), .ZN(n33660) );
  AOI21HSV4 U38732 ( .A1(n33402), .A2(n33565), .B(n33401), .ZN(n33408) );
  CLKNAND2HSV3 U38733 ( .A1(n33505), .A2(n33506), .ZN(n33444) );
  INHSV3 U38734 ( .I(n33444), .ZN(n33909) );
  NOR2HSV4 U38735 ( .A1(n33406), .A2(n33405), .ZN(n33513) );
  CLKNAND2HSV1 U38736 ( .A1(n33909), .A2(n33513), .ZN(n33407) );
  CLKNHSV2 U38737 ( .I(n33573), .ZN(n33409) );
  INHSV4 U38738 ( .I(n33410), .ZN(n45802) );
  NOR2HSV4 U38739 ( .A1(n33412), .A2(n33411), .ZN(n33655) );
  NOR2HSV4 U38740 ( .A1(n33655), .A2(n34416), .ZN(n33443) );
  CLKNHSV0 U38741 ( .I(n33414), .ZN(n33533) );
  CLKNAND2HSV1 U38742 ( .A1(n59661), .A2(n33533), .ZN(n33417) );
  INHSV4 U38743 ( .I(n50248), .ZN(n57592) );
  NAND2HSV0 U38744 ( .A1(n33415), .A2(n57592), .ZN(n33416) );
  INHSV2 U38745 ( .I(n46143), .ZN(n33546) );
  CLKNAND2HSV1 U38746 ( .A1(n33546), .A2(n48074), .ZN(n33419) );
  INHSV2 U38747 ( .I(n34463), .ZN(n33620) );
  CLKNAND2HSV1 U38748 ( .A1(n33620), .A2(n34120), .ZN(n33418) );
  CLKNAND2HSV0 U38749 ( .A1(n59598), .A2(n48069), .ZN(n33422) );
  NAND2HSV0 U38750 ( .A1(n33420), .A2(n33713), .ZN(n33421) );
  NAND2HSV2 U38751 ( .A1(\pe4/aot [25]), .A2(n46617), .ZN(n33425) );
  CLKNAND2HSV0 U38752 ( .A1(n33726), .A2(n33423), .ZN(n33424) );
  CLKNAND2HSV1 U38753 ( .A1(n59383), .A2(n34030), .ZN(n33432) );
  NAND2HSV2 U38754 ( .A1(n47659), .A2(\pe4/pvq [10]), .ZN(n33426) );
  XNOR2HSV1 U38755 ( .A1(n33426), .A2(\pe4/phq [10]), .ZN(n33431) );
  NAND2HSV0 U38756 ( .A1(n33474), .A2(n33427), .ZN(n33429) );
  CLKNAND2HSV1 U38757 ( .A1(n59369), .A2(n33897), .ZN(n33428) );
  XOR2HSV0 U38758 ( .A1(n33429), .A2(n33428), .Z(n33430) );
  XOR3HSV2 U38759 ( .A1(n33432), .A2(n33431), .A3(n33430), .Z(n33433) );
  XNOR2HSV1 U38760 ( .A1(n33434), .A2(n33433), .ZN(n33440) );
  INHSV2 U38761 ( .I(n33859), .ZN(n59600) );
  CLKBUFHSV4 U38762 ( .I(n33464), .Z(n35099) );
  INHSV2 U38763 ( .I(n35099), .ZN(n33735) );
  NAND2HSV2 U38764 ( .A1(n33735), .A2(n33556), .ZN(n33435) );
  XNOR2HSV4 U38765 ( .A1(n33436), .A2(n33435), .ZN(n33439) );
  INHSV2 U38766 ( .I(n33858), .ZN(n59599) );
  NAND2HSV2 U38767 ( .A1(n59501), .A2(n59599), .ZN(n33438) );
  XNOR2HSV4 U38768 ( .A1(n33443), .A2(n33442), .ZN(n33449) );
  INHSV4 U38769 ( .I(n33449), .ZN(n45803) );
  NAND2HSV4 U38770 ( .A1(n45802), .A2(n45803), .ZN(n33447) );
  CLKNAND2HSV1 U38771 ( .A1(n33450), .A2(n33444), .ZN(n33445) );
  NAND2HSV2 U38772 ( .A1(n33445), .A2(n33449), .ZN(n33446) );
  NAND2HSV2 U38773 ( .A1(n33993), .A2(\pe4/ti_7t [10]), .ZN(n33574) );
  INHSV2 U38774 ( .I(n33574), .ZN(n33456) );
  AOI21HSV4 U38775 ( .A1(n45804), .A2(n33448), .B(n33456), .ZN(n33453) );
  AOI21HSV4 U38776 ( .A1(n45802), .A2(n33449), .B(n33695), .ZN(n33570) );
  CLKNAND2HSV2 U38777 ( .A1(n33570), .A2(n33569), .ZN(n33459) );
  INHSV2 U38778 ( .I(n33459), .ZN(n33451) );
  INHSV2 U38779 ( .I(n33573), .ZN(n33578) );
  CLKNAND2HSV2 U38780 ( .A1(n33451), .A2(n33578), .ZN(n33452) );
  CLKNAND2HSV3 U38781 ( .A1(n33453), .A2(n33452), .ZN(n33594) );
  NAND2HSV2 U38782 ( .A1(n59928), .A2(n33707), .ZN(n33454) );
  XNOR2HSV4 U38783 ( .A1(n33455), .A2(n33454), .ZN(n33525) );
  INHSV2 U38784 ( .I(n33456), .ZN(n33458) );
  CLKNAND2HSV2 U38785 ( .A1(n33667), .A2(n33460), .ZN(n33521) );
  NAND2HSV2 U38786 ( .A1(n45806), .A2(n35598), .ZN(n33504) );
  NAND2HSV2 U38787 ( .A1(n33413), .A2(n33461), .ZN(n33502) );
  CLKNHSV2 U38788 ( .I(n33556), .ZN(n33462) );
  NOR2HSV1 U38789 ( .A1(n33464), .A2(n35488), .ZN(n33465) );
  XOR2HSV2 U38790 ( .A1(n33466), .A2(n33465), .Z(n33493) );
  CLKNAND2HSV0 U38791 ( .A1(\pe4/aot [22]), .A2(n48074), .ZN(n33469) );
  INHSV2 U38792 ( .I(n33467), .ZN(n59388) );
  CLKNAND2HSV0 U38793 ( .A1(n59388), .A2(n46617), .ZN(n33468) );
  XOR2HSV0 U38794 ( .A1(n33469), .A2(n33468), .Z(n33473) );
  NAND2HSV0 U38795 ( .A1(n59598), .A2(n33621), .ZN(n33471) );
  CLKNAND2HSV0 U38796 ( .A1(n33614), .A2(n33966), .ZN(n33470) );
  XOR2HSV0 U38797 ( .A1(n33471), .A2(n33470), .Z(n33472) );
  XOR2HSV0 U38798 ( .A1(n33473), .A2(n33472), .Z(n33482) );
  NAND2HSV0 U38799 ( .A1(n33474), .A2(n33713), .ZN(n33476) );
  CLKNAND2HSV1 U38800 ( .A1(n33546), .A2(n33611), .ZN(n33475) );
  XOR2HSV0 U38801 ( .A1(n33476), .A2(n33475), .Z(n33480) );
  CLKNAND2HSV1 U38802 ( .A1(n35370), .A2(\pe4/got [22]), .ZN(n33478) );
  AND2HSV2 U38803 ( .A1(n33624), .A2(n50007), .Z(n33477) );
  XNOR2HSV1 U38804 ( .A1(n33478), .A2(n33477), .ZN(n33479) );
  XOR2HSV0 U38805 ( .A1(n33480), .A2(n33479), .Z(n33481) );
  XOR2HSV0 U38806 ( .A1(n33482), .A2(n33481), .Z(n33491) );
  CLKNAND2HSV1 U38807 ( .A1(n33620), .A2(n57592), .ZN(n33484) );
  INHSV2 U38808 ( .I(n34501), .ZN(n33727) );
  CLKNAND2HSV1 U38809 ( .A1(n33727), .A2(\pe4/bq[22] ), .ZN(n33483) );
  XOR2HSV0 U38810 ( .A1(n33484), .A2(n33483), .Z(n33487) );
  CLKNAND2HSV0 U38811 ( .A1(n34054), .A2(\pe4/pvq [11]), .ZN(n33485) );
  XNOR2HSV1 U38812 ( .A1(n33485), .A2(\pe4/phq [11]), .ZN(n33486) );
  XNOR2HSV1 U38813 ( .A1(n33487), .A2(n33486), .ZN(n33489) );
  INHSV2 U38814 ( .I(n57026), .ZN(n34240) );
  XNOR2HSV1 U38815 ( .A1(n33489), .A2(n33488), .ZN(n33490) );
  XNOR2HSV1 U38816 ( .A1(n33491), .A2(n33490), .ZN(n33492) );
  XOR2HSV0 U38817 ( .A1(n33493), .A2(n33492), .Z(n33495) );
  CLKNAND2HSV0 U38818 ( .A1(n34043), .A2(n34672), .ZN(n33494) );
  XNOR2HSV1 U38819 ( .A1(n33495), .A2(n33494), .ZN(n33496) );
  XNOR2HSV1 U38820 ( .A1(n33497), .A2(n33496), .ZN(n33500) );
  CLKNAND2HSV0 U38821 ( .A1(n29781), .A2(\pe4/got [27]), .ZN(n33499) );
  XNOR2HSV1 U38822 ( .A1(n33500), .A2(n33499), .ZN(n33501) );
  XNOR2HSV4 U38823 ( .A1(n33504), .A2(n33503), .ZN(n33510) );
  NAND2HSV0 U38824 ( .A1(n33506), .A2(n33505), .ZN(n33508) );
  XNOR2HSV4 U38825 ( .A1(n33510), .A2(n33509), .ZN(n33592) );
  CLKNAND2HSV3 U38826 ( .A1(n33527), .A2(n33513), .ZN(n33663) );
  NOR2HSV0 U38827 ( .A1(n33660), .A2(n34712), .ZN(n33511) );
  CLKNAND2HSV2 U38828 ( .A1(n33663), .A2(n33511), .ZN(n33515) );
  INHSV2 U38829 ( .I(n33516), .ZN(n33512) );
  CLKNAND2HSV3 U38830 ( .A1(n33513), .A2(n33512), .ZN(n33662) );
  NOR2HSV4 U38831 ( .A1(n33515), .A2(n33514), .ZN(n33520) );
  CLKNAND2HSV1 U38832 ( .A1(n33516), .A2(n35021), .ZN(n33517) );
  INHSV2 U38833 ( .I(n33400), .ZN(n33518) );
  NAND2HSV4 U38834 ( .A1(n33520), .A2(n33661), .ZN(n33591) );
  XNOR2HSV4 U38835 ( .A1(n33592), .A2(n33591), .ZN(n33587) );
  XNOR2HSV4 U38836 ( .A1(n33521), .A2(n33587), .ZN(n60031) );
  CLKNAND2HSV1 U38837 ( .A1(n60031), .A2(n33848), .ZN(n33524) );
  NAND2HSV2 U38838 ( .A1(\pe4/ti_7t [11]), .A2(n35483), .ZN(n33523) );
  INHSV2 U38839 ( .I(n34187), .ZN(n33805) );
  NOR2HSV0 U38840 ( .A1(n33660), .A2(n34851), .ZN(n33526) );
  NAND2HSV2 U38841 ( .A1(n33662), .A2(n33526), .ZN(n33530) );
  NAND3HSV1 U38842 ( .A1(n33400), .A2(n35011), .A3(n33527), .ZN(n33528) );
  NAND2HSV2 U38843 ( .A1(n33661), .A2(n33528), .ZN(n33529) );
  NAND2HSV2 U38844 ( .A1(n33413), .A2(n33748), .ZN(n33563) );
  NAND2HSV2 U38845 ( .A1(n57325), .A2(n59600), .ZN(n33559) );
  INHSV2 U38846 ( .I(n50207), .ZN(n59370) );
  CLKNAND2HSV0 U38847 ( .A1(n59370), .A2(n33897), .ZN(n33532) );
  CLKNAND2HSV0 U38848 ( .A1(n33965), .A2(n33611), .ZN(n33531) );
  XOR2HSV0 U38849 ( .A1(n33532), .A2(n33531), .Z(n33537) );
  CLKNAND2HSV0 U38850 ( .A1(n59388), .A2(n33533), .ZN(n33535) );
  NAND2HSV0 U38851 ( .A1(n33624), .A2(n57592), .ZN(n33534) );
  XOR2HSV0 U38852 ( .A1(n33535), .A2(n33534), .Z(n33536) );
  XOR2HSV0 U38853 ( .A1(n33537), .A2(n33536), .Z(n33544) );
  NOR2HSV1 U38854 ( .A1(n57026), .A2(n35092), .ZN(n57232) );
  NAND2HSV0 U38855 ( .A1(n59598), .A2(n33713), .ZN(n57012) );
  XOR2HSV0 U38856 ( .A1(n57232), .A2(n57012), .Z(n33542) );
  NAND2HSV0 U38857 ( .A1(n33614), .A2(n33621), .ZN(n33540) );
  CLKNAND2HSV0 U38858 ( .A1(n33631), .A2(n33712), .ZN(n33539) );
  XOR2HSV0 U38859 ( .A1(n33540), .A2(n33539), .Z(n33541) );
  XOR2HSV0 U38860 ( .A1(n33542), .A2(n33541), .Z(n33543) );
  XOR2HSV0 U38861 ( .A1(n33544), .A2(n33543), .Z(n33545) );
  CLKNAND2HSV0 U38862 ( .A1(n33546), .A2(n46617), .ZN(n33548) );
  CLKNAND2HSV1 U38863 ( .A1(n33727), .A2(n34254), .ZN(n33547) );
  XOR2HSV0 U38864 ( .A1(n33548), .A2(n33547), .Z(n33552) );
  NAND2HSV0 U38865 ( .A1(n59390), .A2(n33615), .ZN(n33550) );
  CLKNAND2HSV1 U38866 ( .A1(\pe4/aot [21]), .A2(n34888), .ZN(n33549) );
  XOR2HSV0 U38867 ( .A1(n33550), .A2(n33549), .Z(n33551) );
  XOR2HSV0 U38868 ( .A1(n33552), .A2(n33551), .Z(n33554) );
  CLKNAND2HSV1 U38869 ( .A1(n33620), .A2(n34044), .ZN(n33950) );
  XNOR2HSV1 U38870 ( .A1(n33554), .A2(n33553), .ZN(n33555) );
  CLKNAND2HSV1 U38871 ( .A1(n59501), .A2(n33556), .ZN(n33557) );
  XNOR2HSV1 U38872 ( .A1(n33559), .A2(n33558), .ZN(n33561) );
  XNOR2HSV1 U38873 ( .A1(n33561), .A2(n33560), .ZN(n33562) );
  INHSV2 U38874 ( .I(n33564), .ZN(n33707) );
  NAND2HSV2 U38875 ( .A1(n45806), .A2(n33707), .ZN(n33567) );
  NAND2HSV2 U38876 ( .A1(n35598), .A2(n33565), .ZN(n33566) );
  CLKNAND2HSV0 U38877 ( .A1(n33569), .A2(n33796), .ZN(n33572) );
  CLKNHSV0 U38878 ( .I(n33570), .ZN(n33571) );
  NOR2HSV2 U38879 ( .A1(n33572), .A2(n33571), .ZN(n33579) );
  CLKNAND2HSV2 U38880 ( .A1(n33573), .A2(n33986), .ZN(n33576) );
  OAI22HSV2 U38881 ( .A1(n33576), .A2(n33575), .B1(n34727), .B2(n33574), .ZN(
        n33577) );
  AOI21HSV2 U38882 ( .A1(n33579), .A2(n33578), .B(n33577), .ZN(n33581) );
  NAND2HSV2 U38883 ( .A1(n33580), .A2(n33581), .ZN(n33585) );
  INHSV2 U38884 ( .I(n33580), .ZN(n33583) );
  INHSV2 U38885 ( .I(n33581), .ZN(n33582) );
  CLKNAND2HSV3 U38886 ( .A1(n33582), .A2(n33583), .ZN(n33584) );
  CLKNAND2HSV4 U38887 ( .A1(n33584), .A2(n33585), .ZN(n33678) );
  BUFHSV2 U38888 ( .I(n33678), .Z(n52757) );
  CLKNAND2HSV0 U38889 ( .A1(\pe4/ti_7t [12]), .A2(n33849), .ZN(n33700) );
  INHSV2 U38890 ( .I(n33700), .ZN(n33597) );
  OAI21HSV0 U38891 ( .A1(n35604), .A2(\pe4/ti_7t [11]), .B(n33676), .ZN(n33598) );
  INHSV1 U38892 ( .I(n33598), .ZN(n46603) );
  INHSV2 U38893 ( .I(n46603), .ZN(n33586) );
  NOR2HSV4 U38894 ( .A1(n33603), .A2(n33586), .ZN(n33590) );
  CLKNHSV2 U38895 ( .I(n33587), .ZN(n33589) );
  NAND2HSV4 U38896 ( .A1(n33589), .A2(n33588), .ZN(n33600) );
  CLKNAND2HSV2 U38897 ( .A1(n33590), .A2(n33600), .ZN(n33699) );
  XNOR2HSV4 U38898 ( .A1(n33592), .A2(n33591), .ZN(n33593) );
  CLKAND2HSV1 U38899 ( .A1(n33697), .A2(n33700), .Z(n33595) );
  CLKNAND2HSV1 U38900 ( .A1(n33595), .A2(n29674), .ZN(n33596) );
  NOR2HSV2 U38901 ( .A1(n33598), .A2(n34565), .ZN(n33702) );
  CLKNHSV1 U38902 ( .I(n33702), .ZN(n33599) );
  NOR2HSV1 U38903 ( .A1(n33678), .A2(n33599), .ZN(n33604) );
  INHSV4 U38904 ( .I(n33600), .ZN(n33601) );
  CLKNAND2HSV4 U38905 ( .A1(n33602), .A2(n33601), .ZN(n46604) );
  NAND2HSV4 U38906 ( .A1(n46604), .A2(n46602), .ZN(n33705) );
  INHSV4 U38907 ( .I(n33705), .ZN(n52758) );
  CLKNAND2HSV1 U38908 ( .A1(n33604), .A2(n52758), .ZN(n33605) );
  CLKNHSV0 U38909 ( .I(n34108), .ZN(n34017) );
  NAND2HSV2 U38910 ( .A1(n34458), .A2(n34017), .ZN(n33606) );
  XNOR2HSV4 U38911 ( .A1(n33607), .A2(n33606), .ZN(n33789) );
  INHSV2 U38912 ( .I(n44697), .ZN(n33608) );
  CLKNAND2HSV2 U38913 ( .A1(n33608), .A2(n33707), .ZN(n33659) );
  CLKNAND2HSV0 U38914 ( .A1(n57325), .A2(n57574), .ZN(n33652) );
  INHSV2 U38915 ( .I(n49965), .ZN(n34351) );
  CLKNAND2HSV0 U38916 ( .A1(n34285), .A2(n34351), .ZN(n33610) );
  NOR2HSV1 U38917 ( .A1(n35099), .A2(n50207), .ZN(n33609) );
  XNOR2HSV1 U38918 ( .A1(n33610), .A2(n33609), .ZN(n33648) );
  NAND2HSV2 U38919 ( .A1(n33965), .A2(n33816), .ZN(n33613) );
  INHSV2 U38920 ( .I(n50008), .ZN(n34637) );
  CLKNAND2HSV0 U38921 ( .A1(n34637), .A2(n33611), .ZN(n33612) );
  XOR2HSV0 U38922 ( .A1(n33613), .A2(n33612), .Z(n33619) );
  NAND2HSV0 U38923 ( .A1(n33614), .A2(n33713), .ZN(n33617) );
  NAND2HSV0 U38924 ( .A1(n34110), .A2(n33615), .ZN(n33616) );
  XOR2HSV0 U38925 ( .A1(n33617), .A2(n33616), .Z(n33618) );
  XOR2HSV0 U38926 ( .A1(n33619), .A2(n33618), .Z(n33630) );
  NAND2HSV0 U38927 ( .A1(n33620), .A2(n34254), .ZN(n33623) );
  NAND2HSV0 U38928 ( .A1(n57499), .A2(n33621), .ZN(n33622) );
  XOR2HSV0 U38929 ( .A1(n33623), .A2(n33622), .Z(n33628) );
  NAND2HSV0 U38930 ( .A1(n59390), .A2(n33712), .ZN(n33626) );
  NAND2HSV0 U38931 ( .A1(n33624), .A2(n33711), .ZN(n33625) );
  XOR2HSV0 U38932 ( .A1(n33626), .A2(n33625), .Z(n33627) );
  XOR2HSV0 U38933 ( .A1(n33628), .A2(n33627), .Z(n33629) );
  XOR2HSV0 U38934 ( .A1(n33630), .A2(n33629), .Z(n33646) );
  CLKNAND2HSV0 U38935 ( .A1(n33631), .A2(n57592), .ZN(n33633) );
  CLKNAND2HSV1 U38936 ( .A1(n33716), .A2(n57377), .ZN(n33632) );
  XOR2HSV0 U38937 ( .A1(n33633), .A2(n33632), .Z(n33637) );
  NAND2HSV0 U38938 ( .A1(n33726), .A2(n33966), .ZN(n33635) );
  CLKNAND2HSV0 U38939 ( .A1(n59386), .A2(n57157), .ZN(n33634) );
  XOR2HSV0 U38940 ( .A1(n33635), .A2(n33634), .Z(n33636) );
  XOR2HSV0 U38941 ( .A1(n33637), .A2(n33636), .Z(n33644) );
  CLKNAND2HSV1 U38942 ( .A1(\pe4/aot [20]), .A2(n34888), .ZN(n33639) );
  CLKNAND2HSV0 U38943 ( .A1(n33727), .A2(\pe4/bq[20] ), .ZN(n33638) );
  XOR2HSV0 U38944 ( .A1(n33639), .A2(n33638), .Z(n33642) );
  NAND2HSV0 U38945 ( .A1(n34770), .A2(\pe4/pvq [13]), .ZN(n33640) );
  XOR2HSV0 U38946 ( .A1(n33640), .A2(\pe4/phq [13]), .Z(n33641) );
  XOR2HSV0 U38947 ( .A1(n33642), .A2(n33641), .Z(n33643) );
  XOR2HSV0 U38948 ( .A1(n33644), .A2(n33643), .Z(n33645) );
  XOR2HSV0 U38949 ( .A1(n33646), .A2(n33645), .Z(n33647) );
  XOR2HSV0 U38950 ( .A1(n33648), .A2(n33647), .Z(n33650) );
  INHSV4 U38951 ( .I(n35488), .ZN(n57672) );
  CLKNAND2HSV0 U38952 ( .A1(n59501), .A2(n57672), .ZN(n33649) );
  XNOR2HSV1 U38953 ( .A1(n33650), .A2(n33649), .ZN(n33651) );
  XNOR2HSV1 U38954 ( .A1(n33652), .A2(n33651), .ZN(n33654) );
  NAND2HSV2 U38955 ( .A1(n50266), .A2(n33708), .ZN(n33656) );
  XOR3HSV2 U38956 ( .A1(n33657), .A2(n33656), .A3(n29658), .Z(n33658) );
  XNOR2HSV4 U38957 ( .A1(n33659), .A2(n33658), .ZN(n33665) );
  XNOR2HSV4 U38958 ( .A1(n33665), .A2(n33664), .ZN(n33669) );
  XNOR2HSV4 U38959 ( .A1(n33669), .A2(n33668), .ZN(n52756) );
  INHSV2 U38960 ( .I(n52756), .ZN(n33670) );
  INHSV2 U38961 ( .I(\pe4/ti_7t [13]), .ZN(n33674) );
  OR2HSV1 U38962 ( .A1(n34834), .A2(n33674), .Z(n33677) );
  CLKNAND2HSV1 U38963 ( .A1(n29718), .A2(n33677), .ZN(n33680) );
  NOR2HSV2 U38964 ( .A1(n33678), .A2(n33680), .ZN(n33682) );
  INHSV4 U38965 ( .I(n33678), .ZN(n33704) );
  AOI21HSV4 U38966 ( .A1(n33679), .A2(n46604), .B(n33704), .ZN(n52759) );
  CLKNHSV0 U38967 ( .I(n33680), .ZN(n33681) );
  AOI22HSV2 U38968 ( .A1(n52758), .A2(n33682), .B1(n52759), .B2(n33681), .ZN(
        n33683) );
  CLKNAND2HSV2 U38969 ( .A1(n33684), .A2(n33683), .ZN(n33693) );
  INHSV2 U38970 ( .I(n52759), .ZN(n33686) );
  NAND2HSV2 U38971 ( .A1(n52758), .A2(n33704), .ZN(n33685) );
  NAND2HSV2 U38972 ( .A1(n33686), .A2(n33685), .ZN(n33691) );
  NAND2HSV2 U38973 ( .A1(n29718), .A2(n33848), .ZN(n33688) );
  NOR2HSV2 U38974 ( .A1(n33689), .A2(n33688), .ZN(n33690) );
  CLKNAND2HSV3 U38975 ( .A1(n33691), .A2(n33690), .ZN(n33692) );
  CLKNHSV4 U38976 ( .I(n33802), .ZN(n48892) );
  INHSV2 U38977 ( .I(n34718), .ZN(n33986) );
  XNOR2HSV4 U38978 ( .A1(n33789), .A2(n33788), .ZN(n46599) );
  CLKNAND2HSV0 U38979 ( .A1(n33695), .A2(\pe4/ti_7t [15]), .ZN(n33775) );
  INHSV2 U38980 ( .I(n33775), .ZN(n33783) );
  NAND2HSV2 U38981 ( .A1(n33699), .A2(n33698), .ZN(n33701) );
  AND2HSV2 U38982 ( .A1(n33702), .A2(n33986), .Z(n33703) );
  NOR2HSV3 U38983 ( .A1(n33706), .A2(n33705), .ZN(n33762) );
  NOR2HSV2 U38984 ( .A1(n33763), .A2(n33762), .ZN(n33760) );
  CLKBUFHSV4 U38985 ( .I(n35560), .Z(n34537) );
  CLKNAND2HSV0 U38986 ( .A1(n45806), .A2(n33708), .ZN(n33754) );
  NAND2HSV2 U38987 ( .A1(n50266), .A2(n59600), .ZN(n33747) );
  NAND2HSV2 U38988 ( .A1(n34109), .A2(n57672), .ZN(n33743) );
  NAND2HSV2 U38989 ( .A1(n57359), .A2(n59370), .ZN(n33725) );
  NAND2HSV0 U38990 ( .A1(n33947), .A2(n34030), .ZN(n33709) );
  XOR2HSV0 U38991 ( .A1(n33710), .A2(n33709), .Z(n33723) );
  CLKNAND2HSV1 U38992 ( .A1(n33965), .A2(n33711), .ZN(n34248) );
  NAND2HSV0 U38993 ( .A1(n34110), .A2(n33712), .ZN(n50339) );
  NAND2HSV0 U38994 ( .A1(n34240), .A2(n33713), .ZN(n33715) );
  CLKNAND2HSV0 U38995 ( .A1(n50404), .A2(n57157), .ZN(n33714) );
  XOR2HSV0 U38996 ( .A1(n33715), .A2(n33714), .Z(n33720) );
  NAND2HSV0 U38997 ( .A1(n59390), .A2(\pe4/bq[23] ), .ZN(n33718) );
  NAND2HSV0 U38998 ( .A1(n33716), .A2(n33966), .ZN(n33717) );
  XOR2HSV0 U38999 ( .A1(n33718), .A2(n33717), .Z(n33719) );
  XOR2HSV0 U39000 ( .A1(n33720), .A2(n33719), .Z(n33721) );
  XOR3HSV2 U39001 ( .A1(n33723), .A2(n33722), .A3(n33721), .Z(n33724) );
  XOR2HSV0 U39002 ( .A1(n33725), .A2(n33724), .Z(n33739) );
  INHSV2 U39003 ( .I(n57605), .ZN(n57859) );
  NAND2HSV2 U39004 ( .A1(n35377), .A2(\pe4/bq[20] ), .ZN(n33729) );
  CLKNAND2HSV0 U39005 ( .A1(n33727), .A2(\pe4/bq[19] ), .ZN(n33728) );
  XOR2HSV0 U39006 ( .A1(n33729), .A2(n33728), .Z(n33732) );
  NAND2HSV0 U39007 ( .A1(n33808), .A2(\pe4/pvq [14]), .ZN(n33730) );
  XOR2HSV0 U39008 ( .A1(n33730), .A2(\pe4/phq [14]), .Z(n33731) );
  XOR2HSV0 U39009 ( .A1(n33732), .A2(n33731), .Z(n33733) );
  XOR2HSV0 U39010 ( .A1(n33734), .A2(n33733), .Z(n33737) );
  CLKNAND2HSV0 U39011 ( .A1(n33735), .A2(n33831), .ZN(n33736) );
  XNOR2HSV1 U39012 ( .A1(n33737), .A2(n33736), .ZN(n33738) );
  XNOR2HSV1 U39013 ( .A1(n33739), .A2(n33738), .ZN(n33741) );
  NAND2HSV0 U39014 ( .A1(n34043), .A2(n59601), .ZN(n33740) );
  XNOR2HSV1 U39015 ( .A1(n33741), .A2(n33740), .ZN(n33742) );
  XNOR2HSV1 U39016 ( .A1(n33743), .A2(n33742), .ZN(n33745) );
  CLKNAND2HSV1 U39017 ( .A1(n29738), .A2(\pe4/got [24]), .ZN(n33744) );
  XOR2HSV0 U39018 ( .A1(n33745), .A2(n33744), .Z(n33746) );
  XOR2HSV0 U39019 ( .A1(n33747), .A2(n33746), .Z(n33753) );
  NOR2HSV2 U39020 ( .A1(n44697), .A2(n33749), .ZN(n33751) );
  INHSV2 U39021 ( .I(n33751), .ZN(n33752) );
  XOR3HSV2 U39022 ( .A1(n33754), .A2(n33753), .A3(n33752), .Z(n33755) );
  XNOR2HSV4 U39023 ( .A1(n33756), .A2(n33755), .ZN(n33757) );
  XNOR2HSV4 U39024 ( .A1(n33758), .A2(n33757), .ZN(n33761) );
  INHSV2 U39025 ( .I(n33761), .ZN(n33759) );
  CLKNAND2HSV2 U39026 ( .A1(n33760), .A2(n33759), .ZN(n33769) );
  OAI21HSV2 U39027 ( .A1(n33763), .A2(n33762), .B(n33761), .ZN(n33768) );
  CLKNAND2HSV1 U39028 ( .A1(n33769), .A2(n33768), .ZN(n33766) );
  INHSV2 U39029 ( .I(n45801), .ZN(n33764) );
  NOR2HSV2 U39030 ( .A1(n33764), .A2(n34416), .ZN(n33767) );
  INHSV1 U39031 ( .I(n33767), .ZN(n33765) );
  NAND2HSV2 U39032 ( .A1(n33766), .A2(n33765), .ZN(n33771) );
  NAND3HSV2 U39033 ( .A1(n33769), .A2(n33768), .A3(n33767), .ZN(n33770) );
  NOR2HSV2 U39034 ( .A1(n33850), .A2(n34565), .ZN(n33784) );
  INHSV2 U39035 ( .I(\pe4/ti_7t [14]), .ZN(n33794) );
  AOI21HSV1 U39036 ( .A1(n33794), .A2(n47788), .B(n52696), .ZN(n46597) );
  INHSV1 U39037 ( .I(n46597), .ZN(n33772) );
  NOR2HSV2 U39038 ( .A1(n33772), .A2(n33783), .ZN(n33778) );
  INHSV4 U39039 ( .I(n33802), .ZN(n33795) );
  NAND2HSV0 U39040 ( .A1(n33778), .A2(n48892), .ZN(n33773) );
  NOR2HSV2 U39041 ( .A1(n33784), .A2(n33773), .ZN(n33777) );
  AND2HSV2 U39042 ( .A1(n33775), .A2(n33774), .Z(n33776) );
  NOR2HSV4 U39043 ( .A1(n33777), .A2(n33776), .ZN(n33781) );
  CLKAND2HSV4 U39044 ( .A1(n33781), .A2(n33780), .Z(n33782) );
  OAI21HSV4 U39045 ( .A1(n46599), .A2(n33783), .B(n33782), .ZN(n33793) );
  CLKNAND2HSV1 U39046 ( .A1(n33784), .A2(n25326), .ZN(n46596) );
  AND2HSV2 U39047 ( .A1(n46597), .A2(n33785), .Z(n33786) );
  CLKNAND2HSV1 U39048 ( .A1(n46596), .A2(n33786), .ZN(n33787) );
  NOR2HSV2 U39049 ( .A1(n33857), .A2(n25326), .ZN(n46595) );
  NOR2HSV2 U39050 ( .A1(n33787), .A2(n46595), .ZN(n33791) );
  XOR2HSV0 U39051 ( .A1(n33789), .A2(n33788), .Z(n33790) );
  CLKNAND2HSV2 U39052 ( .A1(n34408), .A2(n25420), .ZN(n33847) );
  NOR2HSV2 U39053 ( .A1(n34419), .A2(n33794), .ZN(n33983) );
  INHSV2 U39054 ( .I(n33850), .ZN(n33854) );
  INHSV2 U39055 ( .I(n47777), .ZN(n35153) );
  AOI22HSV4 U39056 ( .A1(n33796), .A2(n33983), .B1(n60042), .B2(n33997), .ZN(
        n33927) );
  INHSV2 U39057 ( .I(n33564), .ZN(n57195) );
  CLKNAND2HSV1 U39058 ( .A1(n45801), .A2(n57195), .ZN(n33798) );
  CLKAND2HSV2 U39059 ( .A1(n59928), .A2(n33748), .Z(n33797) );
  XNOR2HSV1 U39060 ( .A1(n33798), .A2(n33797), .ZN(n33800) );
  CLKNHSV0 U39061 ( .I(n33800), .ZN(n33799) );
  NOR2HSV2 U39062 ( .A1(n33799), .A2(n34851), .ZN(n33804) );
  AOI21HSV0 U39063 ( .A1(n33802), .A2(n33801), .B(n33800), .ZN(n33803) );
  CLKNAND2HSV1 U39064 ( .A1(n34458), .A2(n33805), .ZN(n33845) );
  BUFHSV2 U39065 ( .I(n34456), .Z(n33858) );
  INHSV2 U39066 ( .I(n33858), .ZN(n34020) );
  NAND2HSV2 U39067 ( .A1(n25616), .A2(n34020), .ZN(n33843) );
  BUFHSV2 U39068 ( .I(n33413), .Z(n35036) );
  NAND2HSV2 U39069 ( .A1(n57530), .A2(n57672), .ZN(n33837) );
  CLKNAND2HSV1 U39070 ( .A1(n34109), .A2(n57567), .ZN(n33833) );
  NAND2HSV0 U39071 ( .A1(n59388), .A2(n34030), .ZN(n33807) );
  CLKNAND2HSV1 U39072 ( .A1(n59605), .A2(n34738), .ZN(n33806) );
  XOR2HSV0 U39073 ( .A1(n33807), .A2(n33806), .Z(n33811) );
  NAND2HSV0 U39074 ( .A1(n33808), .A2(\pe4/pvq [16]), .ZN(n33809) );
  XNOR2HSV1 U39075 ( .A1(n33809), .A2(\pe4/phq [16]), .ZN(n33810) );
  XNOR2HSV1 U39076 ( .A1(n33811), .A2(n33810), .ZN(n33815) );
  CLKNAND2HSV1 U39077 ( .A1(n33947), .A2(n34044), .ZN(n33948) );
  CLKNAND2HSV1 U39078 ( .A1(n33965), .A2(n34598), .ZN(n33818) );
  CLKNAND2HSV0 U39079 ( .A1(n34047), .A2(n33816), .ZN(n33817) );
  XOR2HSV0 U39080 ( .A1(n33818), .A2(n33817), .Z(n33821) );
  NAND2HSV2 U39081 ( .A1(n35201), .A2(n57850), .ZN(n34062) );
  INHSV2 U39082 ( .I(n46143), .ZN(n34022) );
  CLKNAND2HSV1 U39083 ( .A1(n34022), .A2(n34629), .ZN(n33819) );
  XOR2HSV0 U39084 ( .A1(n34062), .A2(n33819), .Z(n33820) );
  INHSV2 U39085 ( .I(n50052), .ZN(n35321) );
  CLKNAND2HSV1 U39086 ( .A1(n35377), .A2(n34359), .ZN(n33823) );
  NAND2HSV0 U39087 ( .A1(n59951), .A2(n33966), .ZN(n33822) );
  CLKNAND2HSV1 U39088 ( .A1(n33960), .A2(n57368), .ZN(n33825) );
  INHSV2 U39089 ( .I(n47861), .ZN(n59353) );
  CLKNAND2HSV0 U39090 ( .A1(n59353), .A2(n57157), .ZN(n33824) );
  CLKNHSV0 U39091 ( .I(n47661), .ZN(n34033) );
  CLKNAND2HSV1 U39092 ( .A1(n34033), .A2(n33969), .ZN(n33827) );
  CLKNAND2HSV1 U39093 ( .A1(n57014), .A2(n33934), .ZN(n33826) );
  CLKNHSV0 U39094 ( .I(n34479), .ZN(n34029) );
  CLKNAND2HSV1 U39095 ( .A1(n34029), .A2(n34243), .ZN(n33829) );
  NAND2HSV0 U39096 ( .A1(n57499), .A2(n34120), .ZN(n33828) );
  INHSV2 U39097 ( .I(n33830), .ZN(n34042) );
  CLKNHSV0 U39098 ( .I(n35501), .ZN(n57285) );
  XNOR2HSV1 U39099 ( .A1(n33833), .A2(n33832), .ZN(n33835) );
  CLKNAND2HSV1 U39100 ( .A1(n57526), .A2(n59601), .ZN(n33834) );
  XNOR2HSV1 U39101 ( .A1(n33835), .A2(n33834), .ZN(n33836) );
  XNOR2HSV1 U39102 ( .A1(n33837), .A2(n33836), .ZN(n33839) );
  CLKNAND2HSV1 U39103 ( .A1(n34595), .A2(n33556), .ZN(n33838) );
  XNOR2HSV1 U39104 ( .A1(n33839), .A2(n33838), .ZN(n33841) );
  NAND2HSV2 U39105 ( .A1(n47742), .A2(n34672), .ZN(n33840) );
  XOR2HSV0 U39106 ( .A1(n33841), .A2(n33840), .Z(n33842) );
  XNOR2HSV1 U39107 ( .A1(n33843), .A2(n33842), .ZN(n33844) );
  XNOR2HSV4 U39108 ( .A1(n33927), .A2(n33926), .ZN(n33994) );
  XNOR2HSV4 U39109 ( .A1(n33847), .A2(n33994), .ZN(pov4[16]) );
  NAND2HSV2 U39110 ( .A1(\pe4/ti_7t [16]), .A2(n33849), .ZN(n34015) );
  INHSV4 U39111 ( .I(n34408), .ZN(n47972) );
  CLKNHSV1 U39112 ( .I(n34187), .ZN(n34019) );
  NAND2HSV2 U39113 ( .A1(n34955), .A2(n34019), .ZN(n33925) );
  INAND2HSV2 U39114 ( .A1(n33852), .B1(n33850), .ZN(n33857) );
  INHSV2 U39115 ( .I(n33851), .ZN(n33856) );
  NOR2HSV0 U39116 ( .A1(n33852), .A2(n46581), .ZN(n33853) );
  AOI31HSV2 U39117 ( .A1(n33854), .A2(n57188), .A3(n33853), .B(n33983), .ZN(
        n33855) );
  CLKBUFHSV4 U39118 ( .I(n35569), .Z(n34593) );
  NAND2HSV2 U39119 ( .A1(n34593), .A2(n57195), .ZN(n33923) );
  BUFHSV4 U39120 ( .I(n34458), .Z(n46601) );
  INHSV2 U39121 ( .I(n33858), .ZN(n47771) );
  CLKNAND2HSV1 U39122 ( .A1(n46601), .A2(n47771), .ZN(n33921) );
  CLKNAND2HSV1 U39123 ( .A1(n34459), .A2(\pe4/got [25]), .ZN(n33917) );
  BUFHSV2 U39124 ( .I(n34867), .Z(n35322) );
  CLKNAND2HSV1 U39125 ( .A1(n35322), .A2(n34239), .ZN(n33913) );
  BUFHSV2 U39126 ( .I(n34109), .Z(n47733) );
  NAND2HSV0 U39127 ( .A1(n47658), .A2(n34243), .ZN(n33862) );
  NAND2HSV0 U39128 ( .A1(n34029), .A2(\pe4/bq[17] ), .ZN(n33861) );
  XOR2HSV0 U39129 ( .A1(n33862), .A2(n33861), .Z(n33866) );
  NAND2HSV0 U39130 ( .A1(n34033), .A2(n34359), .ZN(n33864) );
  NAND2HSV0 U39131 ( .A1(n34110), .A2(n57929), .ZN(n33863) );
  XOR2HSV0 U39132 ( .A1(n33864), .A2(n33863), .Z(n33865) );
  XOR2HSV0 U39133 ( .A1(n33866), .A2(n33865), .Z(n33875) );
  CLKNHSV0 U39134 ( .I(n34631), .ZN(n35091) );
  CLKNAND2HSV1 U39135 ( .A1(n35091), .A2(n49943), .ZN(n33869) );
  CLKNAND2HSV0 U39136 ( .A1(n33867), .A2(n48069), .ZN(n33868) );
  XOR2HSV0 U39137 ( .A1(n33869), .A2(n33868), .Z(n33873) );
  NAND2HSV0 U39138 ( .A1(n34743), .A2(n34629), .ZN(n33871) );
  CLKNAND2HSV1 U39139 ( .A1(\pe4/aot [14]), .A2(n57098), .ZN(n33870) );
  XOR2HSV0 U39140 ( .A1(n33871), .A2(n33870), .Z(n33872) );
  XOR2HSV0 U39141 ( .A1(n33873), .A2(n33872), .Z(n33874) );
  XOR2HSV0 U39142 ( .A1(n33875), .A2(n33874), .Z(n33877) );
  CLKNHSV0 U39143 ( .I(n35099), .ZN(n34127) );
  INHSV2 U39144 ( .I(n50212), .ZN(n57307) );
  NAND2HSV0 U39145 ( .A1(n34127), .A2(n57307), .ZN(n33876) );
  XNOR2HSV1 U39146 ( .A1(n33877), .A2(n33876), .ZN(n33908) );
  NAND2HSV0 U39147 ( .A1(n34043), .A2(n59353), .ZN(n33907) );
  BUFHSV2 U39148 ( .I(n34254), .Z(n34636) );
  NAND2HSV0 U39149 ( .A1(n34240), .A2(n34636), .ZN(n33879) );
  NAND2HSV0 U39150 ( .A1(\pe4/aot [17]), .A2(n57377), .ZN(n33878) );
  XOR2HSV0 U39151 ( .A1(n33879), .A2(n33878), .Z(n33883) );
  NAND2HSV0 U39152 ( .A1(\pe4/aot [22]), .A2(n34120), .ZN(n33881) );
  NAND2HSV0 U39153 ( .A1(n34637), .A2(n34030), .ZN(n33880) );
  XOR2HSV0 U39154 ( .A1(n33881), .A2(n33880), .Z(n33882) );
  XOR2HSV0 U39155 ( .A1(n33883), .A2(n33882), .Z(n33891) );
  CLKNHSV0 U39156 ( .I(n57605), .ZN(n34874) );
  INHSV2 U39157 ( .I(n57260), .ZN(n35207) );
  NAND2HSV0 U39158 ( .A1(n34874), .A2(n35207), .ZN(n33885) );
  NAND2HSV0 U39159 ( .A1(n57852), .A2(n34738), .ZN(n33884) );
  XOR2HSV0 U39160 ( .A1(n33885), .A2(n33884), .Z(n33889) );
  NAND2HSV0 U39161 ( .A1(n59388), .A2(n34044), .ZN(n33887) );
  CLKNAND2HSV0 U39162 ( .A1(n34022), .A2(n57476), .ZN(n33886) );
  XOR2HSV0 U39163 ( .A1(n33887), .A2(n33886), .Z(n33888) );
  XOR2HSV0 U39164 ( .A1(n33889), .A2(n33888), .Z(n33890) );
  XOR2HSV0 U39165 ( .A1(n33891), .A2(n33890), .Z(n33903) );
  CLKNHSV0 U39166 ( .I(n33808), .ZN(n35493) );
  NAND2HSV2 U39167 ( .A1(\pe4/pvq [19]), .A2(n47659), .ZN(n33892) );
  XOR2HSV0 U39168 ( .A1(n33892), .A2(\pe4/phq [19]), .Z(n33896) );
  INHSV2 U39169 ( .I(n47818), .ZN(n57348) );
  NAND2HSV2 U39170 ( .A1(n35201), .A2(n57348), .ZN(n34060) );
  CLKNHSV0 U39171 ( .I(n34463), .ZN(n34387) );
  CLKNAND2HSV0 U39172 ( .A1(n34387), .A2(n57139), .ZN(n34146) );
  BUFHSV2 U39173 ( .I(n33355), .Z(n35058) );
  OAI22HSV0 U39174 ( .A1(n33114), .A2(n47818), .B1(n35058), .B2(n57387), .ZN(
        n33894) );
  OAI21HSV1 U39175 ( .A1(n34060), .A2(n34146), .B(n33894), .ZN(n33895) );
  XNOR2HSV1 U39176 ( .A1(n33896), .A2(n33895), .ZN(n33901) );
  NAND2HSV0 U39177 ( .A1(n59952), .A2(n34021), .ZN(n33899) );
  INHSV2 U39178 ( .I(n50042), .ZN(n57424) );
  NAND2HSV0 U39179 ( .A1(n57424), .A2(n47679), .ZN(n33898) );
  XOR2HSV0 U39180 ( .A1(n33899), .A2(n33898), .Z(n33900) );
  XNOR2HSV1 U39181 ( .A1(n33901), .A2(n33900), .ZN(n33902) );
  XNOR2HSV1 U39182 ( .A1(n33903), .A2(n33902), .ZN(n33905) );
  CLKNAND2HSV0 U39183 ( .A1(n59382), .A2(n57189), .ZN(n33904) );
  XNOR2HSV1 U39184 ( .A1(n33905), .A2(n33904), .ZN(n33906) );
  CLKNHSV0 U39185 ( .I(n33909), .ZN(n35401) );
  NAND2HSV0 U39186 ( .A1(n35401), .A2(n34351), .ZN(n33910) );
  XOR2HSV0 U39187 ( .A1(n33911), .A2(n33910), .Z(n33912) );
  XNOR2HSV1 U39188 ( .A1(n33913), .A2(n33912), .ZN(n33915) );
  NAND2HSV0 U39189 ( .A1(n59928), .A2(n59603), .ZN(n33914) );
  XNOR2HSV1 U39190 ( .A1(n33915), .A2(n33914), .ZN(n33916) );
  XNOR2HSV1 U39191 ( .A1(n33917), .A2(n33916), .ZN(n33920) );
  CLKNAND2HSV1 U39192 ( .A1(n33918), .A2(n59350), .ZN(n33919) );
  XOR3HSV2 U39193 ( .A1(n33921), .A2(n33920), .A3(n33919), .Z(n33922) );
  XNOR2HSV1 U39194 ( .A1(n33923), .A2(n33922), .ZN(n33924) );
  XNOR2HSV4 U39195 ( .A1(n33925), .A2(n33924), .ZN(n34105) );
  XNOR2HSV4 U39196 ( .A1(n34106), .A2(n34105), .ZN(n34230) );
  XNOR2HSV4 U39197 ( .A1(n33927), .A2(n33926), .ZN(n33989) );
  CLKNHSV0 U39198 ( .I(n35032), .ZN(n33929) );
  NOR2HSV2 U39199 ( .A1(n33795), .A2(n33929), .ZN(n33933) );
  NAND2HSV2 U39200 ( .A1(n34459), .A2(n59350), .ZN(n33931) );
  CLKNAND2HSV0 U39201 ( .A1(n59928), .A2(n34020), .ZN(n33930) );
  INHSV2 U39202 ( .I(n33564), .ZN(n34410) );
  CLKNAND2HSV1 U39203 ( .A1(n25616), .A2(n34672), .ZN(n33979) );
  CLKNAND2HSV0 U39204 ( .A1(n59952), .A2(n33934), .ZN(n33936) );
  CLKNAND2HSV0 U39205 ( .A1(n34033), .A2(n34243), .ZN(n33935) );
  XOR2HSV0 U39206 ( .A1(n33936), .A2(n33935), .Z(n33939) );
  NAND2HSV0 U39207 ( .A1(n34022), .A2(n34030), .ZN(n34914) );
  NAND2HSV0 U39208 ( .A1(n59388), .A2(n50007), .ZN(n33937) );
  XOR2HSV0 U39209 ( .A1(n34914), .A2(n33937), .Z(n33938) );
  XOR2HSV0 U39210 ( .A1(n33939), .A2(n33938), .Z(n33957) );
  CLKNAND2HSV1 U39211 ( .A1(n34637), .A2(n35207), .ZN(n33941) );
  NAND2HSV0 U39212 ( .A1(n47656), .A2(n57157), .ZN(n33940) );
  XOR2HSV0 U39213 ( .A1(n33941), .A2(n33940), .Z(n33944) );
  NAND2HSV0 U39214 ( .A1(n34138), .A2(\pe4/pvq [17]), .ZN(n33942) );
  XOR2HSV0 U39215 ( .A1(n33942), .A2(\pe4/phq [17]), .Z(n33943) );
  XOR2HSV0 U39216 ( .A1(n33944), .A2(n33943), .Z(n33954) );
  NAND2HSV2 U39217 ( .A1(\pe4/aot [17]), .A2(n49943), .ZN(n57131) );
  CLKNAND2HSV0 U39218 ( .A1(n35201), .A2(\pe4/bq[16] ), .ZN(n34152) );
  OAI21HSV2 U39219 ( .A1(n35175), .A2(n35068), .B(n34152), .ZN(n33945) );
  NAND2HSV0 U39220 ( .A1(n33947), .A2(n57850), .ZN(n34353) );
  OAI21HSV0 U39221 ( .A1(n47809), .A2(n34463), .B(n33948), .ZN(n33949) );
  OAI21HSV0 U39222 ( .A1(n33950), .A2(n34353), .B(n33949), .ZN(n33951) );
  XOR2HSV0 U39223 ( .A1(n33952), .A2(n33951), .Z(n33953) );
  XNOR2HSV1 U39224 ( .A1(n33954), .A2(n33953), .ZN(n33956) );
  CLKNAND2HSV1 U39225 ( .A1(n57359), .A2(n34042), .ZN(n33955) );
  NAND2HSV0 U39226 ( .A1(n57218), .A2(n34021), .ZN(n33959) );
  CLKNAND2HSV0 U39227 ( .A1(n34029), .A2(\pe4/bq[19] ), .ZN(n33958) );
  XOR2HSV0 U39228 ( .A1(n33959), .A2(n33958), .Z(n33964) );
  NAND2HSV0 U39229 ( .A1(n34240), .A2(n57476), .ZN(n33962) );
  NAND2HSV0 U39230 ( .A1(n33960), .A2(n34359), .ZN(n33961) );
  XOR2HSV0 U39231 ( .A1(n33962), .A2(n33961), .Z(n33963) );
  XOR2HSV0 U39232 ( .A1(n33964), .A2(n33963), .Z(n33975) );
  NAND2HSV0 U39233 ( .A1(n33965), .A2(n34629), .ZN(n33968) );
  NAND2HSV0 U39234 ( .A1(n59839), .A2(n33966), .ZN(n33967) );
  XOR2HSV0 U39235 ( .A1(n33968), .A2(n33967), .Z(n33973) );
  NAND2HSV0 U39236 ( .A1(n34047), .A2(n57377), .ZN(n33971) );
  NAND2HSV0 U39237 ( .A1(n34110), .A2(n33969), .ZN(n33970) );
  XOR2HSV0 U39238 ( .A1(n33971), .A2(n33970), .Z(n33972) );
  XOR2HSV0 U39239 ( .A1(n33973), .A2(n33972), .Z(n33974) );
  INHSV2 U39240 ( .I(n47861), .ZN(n57753) );
  CLKNAND2HSV1 U39241 ( .A1(n35401), .A2(n33556), .ZN(n33977) );
  XNOR2HSV4 U39242 ( .A1(n33981), .A2(n33980), .ZN(n33985) );
  AOI22HSV2 U39243 ( .A1(n33983), .A2(n47655), .B1(n60042), .B2(n33982), .ZN(
        n33984) );
  XNOR2HSV4 U39244 ( .A1(n33985), .A2(n33984), .ZN(n34010) );
  INHSV2 U39245 ( .I(n34010), .ZN(n33987) );
  CLKNAND2HSV2 U39246 ( .A1(n34408), .A2(n33986), .ZN(n34011) );
  XNOR2HSV4 U39247 ( .A1(n33987), .A2(n34011), .ZN(n52797) );
  CLKNAND2HSV0 U39248 ( .A1(n52796), .A2(n52797), .ZN(n33988) );
  INHSV2 U39249 ( .I(n33988), .ZN(n33992) );
  CLKNHSV0 U39250 ( .I(n33989), .ZN(n33998) );
  OAI21HSV2 U39251 ( .A1(n33848), .A2(\pe4/ti_7t [16]), .B(n47778), .ZN(n52793) );
  NOR2HSV2 U39252 ( .A1(n52793), .A2(n34221), .ZN(n34009) );
  CLKNAND2HSV1 U39253 ( .A1(n34009), .A2(n34843), .ZN(n33990) );
  AOI21HSV2 U39254 ( .A1(n33998), .A2(n57816), .B(n33990), .ZN(n33991) );
  NAND2HSV4 U39255 ( .A1(n33992), .A2(n33991), .ZN(n34001) );
  CLKNAND2HSV1 U39256 ( .A1(n47788), .A2(\pe4/ti_7t [17]), .ZN(n34005) );
  OR2HSV1 U39257 ( .A1(n34005), .A2(n57204), .Z(n34000) );
  INHSV2 U39258 ( .I(n34008), .ZN(n33996) );
  NOR2HSV0 U39259 ( .A1(n34408), .A2(n52793), .ZN(n33995) );
  NAND2HSV2 U39260 ( .A1(n33996), .A2(n33995), .ZN(n34196) );
  NOR2HSV2 U39261 ( .A1(n47972), .A2(n52793), .ZN(n34003) );
  CLKNHSV2 U39262 ( .I(n34349), .ZN(n34101) );
  NOR2HSV4 U39263 ( .A1(n34004), .A2(n52797), .ZN(n34006) );
  INHSV2 U39264 ( .I(n34005), .ZN(n34204) );
  NOR2HSV4 U39265 ( .A1(n34006), .A2(n34204), .ZN(n34014) );
  CLKNHSV0 U39266 ( .I(n47972), .ZN(n34007) );
  NAND3HSV4 U39267 ( .A1(n52796), .A2(n52795), .A3(n34009), .ZN(n34012) );
  XNOR2HSV4 U39268 ( .A1(n34011), .A2(n34010), .ZN(n34197) );
  NOR2HSV4 U39269 ( .A1(n34012), .A2(n34197), .ZN(n34207) );
  NAND2HSV4 U39270 ( .A1(n34014), .A2(n34013), .ZN(n34447) );
  NOR2HSV4 U39271 ( .A1(n34099), .A2(n33993), .ZN(n34103) );
  NOR2HSV0 U39272 ( .A1(n47972), .A2(n34416), .ZN(n34018) );
  INHSV2 U39273 ( .I(n34018), .ZN(n34092) );
  CLKNAND2HSV1 U39274 ( .A1(n35569), .A2(n34019), .ZN(n34089) );
  NAND2HSV2 U39275 ( .A1(n46601), .A2(n59350), .ZN(n34087) );
  NAND2HSV2 U39276 ( .A1(n34459), .A2(n34020), .ZN(n34084) );
  NAND2HSV2 U39277 ( .A1(n35322), .A2(n59603), .ZN(n34080) );
  BUFHSV2 U39278 ( .I(n34109), .Z(n34868) );
  CLKNAND2HSV0 U39279 ( .A1(\pe4/aot [17]), .A2(n34021), .ZN(n34024) );
  NAND2HSV0 U39280 ( .A1(n34022), .A2(n34120), .ZN(n34023) );
  XOR2HSV0 U39281 ( .A1(n34024), .A2(n34023), .Z(n34028) );
  NAND2HSV2 U39282 ( .A1(n34387), .A2(\pe4/bq[16] ), .ZN(n34026) );
  NAND2HSV2 U39283 ( .A1(n57852), .A2(n57098), .ZN(n34025) );
  XOR2HSV0 U39284 ( .A1(n34026), .A2(n34025), .Z(n34027) );
  XOR2HSV0 U39285 ( .A1(n34028), .A2(n34027), .Z(n34039) );
  NAND2HSV0 U39286 ( .A1(n34029), .A2(n34359), .ZN(n34032) );
  NAND2HSV0 U39287 ( .A1(n33965), .A2(n34030), .ZN(n34031) );
  XOR2HSV0 U39288 ( .A1(n34032), .A2(n34031), .Z(n34037) );
  NAND2HSV0 U39289 ( .A1(n34637), .A2(n34629), .ZN(n34035) );
  NAND2HSV0 U39290 ( .A1(n34033), .A2(n50250), .ZN(n34034) );
  XOR2HSV0 U39291 ( .A1(n34035), .A2(n34034), .Z(n34036) );
  XOR2HSV0 U39292 ( .A1(n34037), .A2(n34036), .Z(n34038) );
  XOR2HSV0 U39293 ( .A1(n34039), .A2(n34038), .Z(n34041) );
  CLKNAND2HSV1 U39294 ( .A1(n34127), .A2(n57189), .ZN(n34040) );
  XNOR2HSV1 U39295 ( .A1(n34041), .A2(n34040), .ZN(n34074) );
  NAND2HSV0 U39296 ( .A1(n34043), .A2(n34042), .ZN(n34073) );
  NAND2HSV0 U39297 ( .A1(n34240), .A2(n34044), .ZN(n34046) );
  NAND2HSV0 U39298 ( .A1(\pe4/aot [16]), .A2(n34738), .ZN(n34045) );
  XOR2HSV0 U39299 ( .A1(n34046), .A2(n34045), .Z(n34051) );
  NAND2HSV2 U39300 ( .A1(n47658), .A2(n34636), .ZN(n34049) );
  NAND2HSV0 U39301 ( .A1(n34047), .A2(n33966), .ZN(n34048) );
  XOR2HSV0 U39302 ( .A1(n34049), .A2(n34048), .Z(n34050) );
  XOR2HSV0 U39303 ( .A1(n34051), .A2(n34050), .Z(n34059) );
  NAND2HSV0 U39304 ( .A1(n59388), .A2(n57476), .ZN(n34053) );
  NAND2HSV0 U39305 ( .A1(\pe4/aot [18]), .A2(n57377), .ZN(n34052) );
  XOR2HSV0 U39306 ( .A1(n34053), .A2(n34052), .Z(n34057) );
  NAND2HSV0 U39307 ( .A1(n34054), .A2(\pe4/pvq [18]), .ZN(n34055) );
  XOR2HSV0 U39308 ( .A1(n34055), .A2(\pe4/phq [18]), .Z(n34056) );
  XOR2HSV0 U39309 ( .A1(n34057), .A2(n34056), .Z(n34058) );
  XOR2HSV0 U39310 ( .A1(n34059), .A2(n34058), .Z(n34069) );
  INHSV2 U39311 ( .I(n47818), .ZN(n58084) );
  CLKNAND2HSV1 U39312 ( .A1(n35091), .A2(n58084), .ZN(n34153) );
  OAI21HSV0 U39313 ( .A1(n47809), .A2(n34631), .B(n34060), .ZN(n34061) );
  OAI21HSV0 U39314 ( .A1(n34062), .A2(n34153), .B(n34061), .ZN(n34063) );
  CLKNAND2HSV0 U39315 ( .A1(n34743), .A2(n35207), .ZN(n34278) );
  XNOR2HSV1 U39316 ( .A1(n34063), .A2(n34278), .ZN(n34067) );
  NAND2HSV0 U39317 ( .A1(n34110), .A2(n34243), .ZN(n34065) );
  CLKNAND2HSV0 U39318 ( .A1(\pe4/got [15]), .A2(n47679), .ZN(n34064) );
  XOR2HSV0 U39319 ( .A1(n34065), .A2(n34064), .Z(n34066) );
  XNOR2HSV1 U39320 ( .A1(n34067), .A2(n34066), .ZN(n34068) );
  XNOR2HSV1 U39321 ( .A1(n34069), .A2(n34068), .ZN(n34071) );
  INHSV2 U39322 ( .I(n47861), .ZN(n35167) );
  NAND2HSV2 U39323 ( .A1(n57359), .A2(n35167), .ZN(n34070) );
  XNOR2HSV1 U39324 ( .A1(n34071), .A2(n34070), .ZN(n34072) );
  CLKNAND2HSV1 U39325 ( .A1(n59681), .A2(n34351), .ZN(n34075) );
  XNOR2HSV1 U39326 ( .A1(n34076), .A2(n34075), .ZN(n34078) );
  NAND2HSV0 U39327 ( .A1(n47742), .A2(n59369), .ZN(n34077) );
  XOR2HSV0 U39328 ( .A1(n34078), .A2(n34077), .Z(n34079) );
  XNOR2HSV1 U39329 ( .A1(n34080), .A2(n34079), .ZN(n34082) );
  CLKNAND2HSV1 U39330 ( .A1(n34405), .A2(\pe4/got [25]), .ZN(n34081) );
  XNOR2HSV1 U39331 ( .A1(n34082), .A2(n34081), .ZN(n34083) );
  XNOR2HSV1 U39332 ( .A1(n34084), .A2(n34083), .ZN(n34086) );
  NAND2HSV2 U39333 ( .A1(n50384), .A2(n57195), .ZN(n34085) );
  XOR3HSV2 U39334 ( .A1(n34087), .A2(n34086), .A3(n34085), .Z(n34088) );
  XOR2HSV0 U39335 ( .A1(n34089), .A2(n34088), .Z(n34090) );
  CLKNHSV2 U39336 ( .I(n34090), .ZN(n34091) );
  XNOR2HSV4 U39337 ( .A1(n34092), .A2(n34091), .ZN(n34210) );
  INHSV2 U39338 ( .I(n34210), .ZN(n34205) );
  CLKNAND2HSV1 U39339 ( .A1(n34097), .A2(n34205), .ZN(n34095) );
  AND2HSV1 U39340 ( .A1(n34210), .A2(n34843), .Z(n34093) );
  OAI21HSV2 U39341 ( .A1(n33848), .A2(\pe4/ti_7t [18]), .B(n25420), .ZN(n34317) );
  NOR2HSV1 U39342 ( .A1(n34210), .A2(n34712), .ZN(n34096) );
  NAND3HSV4 U39343 ( .A1(n34100), .A2(n34099), .A3(n35011), .ZN(n34320) );
  NAND3HSV4 U39344 ( .A1(n34101), .A2(n52820), .A3(n35011), .ZN(n47962) );
  CLKNAND2HSV4 U39345 ( .A1(n34103), .A2(n34102), .ZN(n34343) );
  NOR2HSV1 U39346 ( .A1(n34317), .A2(n47788), .ZN(n34323) );
  INHSV2 U39347 ( .I(\pe4/ti_7t [19]), .ZN(n34327) );
  XNOR2HSV4 U39348 ( .A1(n34106), .A2(n34105), .ZN(n34107) );
  XNOR2HSV4 U39349 ( .A1(n34107), .A2(n25879), .ZN(n34345) );
  INHSV1 U39350 ( .I(n34108), .ZN(n47655) );
  CLKNAND2HSV4 U39351 ( .A1(n29759), .A2(n47655), .ZN(n34192) );
  NAND2HSV2 U39352 ( .A1(n34593), .A2(n59350), .ZN(n34184) );
  NAND2HSV2 U39353 ( .A1(n46601), .A2(n57190), .ZN(n34182) );
  CLKNAND2HSV1 U39354 ( .A1(n34459), .A2(n59603), .ZN(n34179) );
  BUFHSV2 U39355 ( .I(n25616), .Z(n34352) );
  NAND2HSV2 U39356 ( .A1(n34352), .A2(n34351), .ZN(n34175) );
  NAND2HSV0 U39357 ( .A1(n35036), .A2(n35321), .ZN(n34169) );
  NAND2HSV0 U39358 ( .A1(n34109), .A2(n59353), .ZN(n34165) );
  CLKNAND2HSV1 U39359 ( .A1(n34022), .A2(n34044), .ZN(n34112) );
  NAND2HSV0 U39360 ( .A1(n34110), .A2(n34359), .ZN(n34111) );
  XOR2HSV0 U39361 ( .A1(n34112), .A2(n34111), .Z(n34116) );
  CLKNAND2HSV1 U39362 ( .A1(n35533), .A2(n57926), .ZN(n34114) );
  CLKNAND2HSV1 U39363 ( .A1(n59953), .A2(n57134), .ZN(n34113) );
  XOR2HSV0 U39364 ( .A1(n34114), .A2(n34113), .Z(n34115) );
  XOR2HSV0 U39365 ( .A1(n34116), .A2(n34115), .Z(n34126) );
  CLKNAND2HSV1 U39366 ( .A1(\pe4/aot [16]), .A2(n33313), .ZN(n34119) );
  CLKNHSV0 U39367 ( .I(\pe4/bq[25] ), .ZN(n48070) );
  INHSV2 U39368 ( .I(n48070), .ZN(n57459) );
  NAND2HSV0 U39369 ( .A1(n59839), .A2(n57459), .ZN(n34118) );
  XOR2HSV0 U39370 ( .A1(n34119), .A2(n34118), .Z(n34124) );
  NAND2HSV0 U39371 ( .A1(n59605), .A2(n35207), .ZN(n34122) );
  NAND2HSV0 U39372 ( .A1(n34637), .A2(n34120), .ZN(n34121) );
  XOR2HSV0 U39373 ( .A1(n34122), .A2(n34121), .Z(n34123) );
  XOR2HSV0 U39374 ( .A1(n34124), .A2(n34123), .Z(n34125) );
  XOR2HSV0 U39375 ( .A1(n34126), .A2(n34125), .Z(n34129) );
  NAND2HSV0 U39376 ( .A1(n34127), .A2(n57424), .ZN(n34128) );
  XNOR2HSV1 U39377 ( .A1(n34129), .A2(n34128), .ZN(n34163) );
  INHSV1 U39378 ( .I(n47793), .ZN(n59604) );
  NAND2HSV0 U39379 ( .A1(n57285), .A2(n59604), .ZN(n34162) );
  CLKNAND2HSV1 U39380 ( .A1(n33726), .A2(n34636), .ZN(n34131) );
  INHSV2 U39381 ( .I(n44338), .ZN(n58163) );
  CLKNAND2HSV0 U39382 ( .A1(n58163), .A2(n33934), .ZN(n34130) );
  XOR2HSV0 U39383 ( .A1(n34131), .A2(n34130), .Z(n34135) );
  NAND2HSV0 U39384 ( .A1(\pe4/aot [22]), .A2(n57592), .ZN(n34133) );
  CLKNHSV0 U39385 ( .I(n58189), .ZN(n57820) );
  NAND2HSV0 U39386 ( .A1(n57820), .A2(n47679), .ZN(n34132) );
  XOR2HSV0 U39387 ( .A1(n34133), .A2(n34132), .Z(n34134) );
  XOR2HSV0 U39388 ( .A1(n34135), .A2(n34134), .Z(n34143) );
  NOR2HSV0 U39389 ( .A1(n35175), .A2(n35092), .ZN(n34137) );
  NAND2HSV0 U39390 ( .A1(n34874), .A2(n34629), .ZN(n34136) );
  XOR2HSV0 U39391 ( .A1(n34137), .A2(n34136), .Z(n34141) );
  NAND2HSV0 U39392 ( .A1(n34138), .A2(\pe4/pvq [20]), .ZN(n34139) );
  XOR2HSV0 U39393 ( .A1(n34139), .A2(\pe4/phq [20]), .Z(n34140) );
  XOR2HSV0 U39394 ( .A1(n34141), .A2(n34140), .Z(n34142) );
  XOR2HSV0 U39395 ( .A1(n34143), .A2(n34142), .Z(n34158) );
  NAND2HSV0 U39396 ( .A1(\pe4/aot [14]), .A2(n34243), .ZN(n47669) );
  OAI22HSV0 U39397 ( .A1(n35068), .A2(n34470), .B1(n57026), .B2(n48023), .ZN(
        n34144) );
  OAI21HSV0 U39398 ( .A1(n34145), .A2(n47669), .B(n34144), .ZN(n34150) );
  CLKNAND2HSV0 U39399 ( .A1(n47658), .A2(n57139), .ZN(n34920) );
  OAI21HSV0 U39400 ( .A1(n48022), .A2(n57509), .B(n34146), .ZN(n34147) );
  OAI21HSV0 U39401 ( .A1(n34920), .A2(n34148), .B(n34147), .ZN(n34149) );
  XOR2HSV0 U39402 ( .A1(n34150), .A2(n34149), .Z(n34156) );
  CLKNHSV0 U39403 ( .I(n34479), .ZN(n35491) );
  CLKNAND2HSV1 U39404 ( .A1(n35491), .A2(n34480), .ZN(n34641) );
  OAI22HSV0 U39405 ( .A1(n35058), .A2(n53219), .B1(n34479), .B2(n48024), .ZN(
        n34151) );
  OAI21HSV0 U39406 ( .A1(n34152), .A2(n34641), .B(n34151), .ZN(n34154) );
  XNOR2HSV1 U39407 ( .A1(n34154), .A2(n34153), .ZN(n34155) );
  XNOR2HSV1 U39408 ( .A1(n34156), .A2(n34155), .ZN(n34157) );
  XNOR2HSV1 U39409 ( .A1(n34158), .A2(n34157), .ZN(n34160) );
  CLKNHSV1 U39410 ( .I(n50212), .ZN(n34937) );
  CLKNAND2HSV0 U39411 ( .A1(n34285), .A2(n34937), .ZN(n34159) );
  XNOR2HSV1 U39412 ( .A1(n34160), .A2(n34159), .ZN(n34161) );
  XOR3HSV2 U39413 ( .A1(n34163), .A2(n34162), .A3(n34161), .Z(n34164) );
  XNOR2HSV1 U39414 ( .A1(n34165), .A2(n34164), .ZN(n34167) );
  CLKNAND2HSV0 U39415 ( .A1(n57526), .A2(n59372), .ZN(n34166) );
  XNOR2HSV1 U39416 ( .A1(n34167), .A2(n34166), .ZN(n34168) );
  XNOR2HSV1 U39417 ( .A1(n34169), .A2(n34168), .ZN(n34171) );
  CLKNAND2HSV0 U39418 ( .A1(n57405), .A2(n59386), .ZN(n34170) );
  XNOR2HSV1 U39419 ( .A1(n34171), .A2(n34170), .ZN(n34173) );
  CLKNHSV1 U39420 ( .I(n33750), .ZN(n57679) );
  CLKNAND2HSV1 U39421 ( .A1(n57679), .A2(n59370), .ZN(n34172) );
  XOR2HSV0 U39422 ( .A1(n34173), .A2(n34172), .Z(n34174) );
  XNOR2HSV1 U39423 ( .A1(n34175), .A2(n34174), .ZN(n34177) );
  CLKNAND2HSV0 U39424 ( .A1(n34405), .A2(n34239), .ZN(n34176) );
  XNOR2HSV1 U39425 ( .A1(n34177), .A2(n34176), .ZN(n34178) );
  XNOR2HSV1 U39426 ( .A1(n34179), .A2(n34178), .ZN(n34181) );
  NAND2HSV2 U39427 ( .A1(n25894), .A2(n47771), .ZN(n34180) );
  XOR3HSV2 U39428 ( .A1(n34182), .A2(n34181), .A3(n34180), .Z(n34183) );
  XNOR2HSV1 U39429 ( .A1(n34184), .A2(n34183), .ZN(n34186) );
  NAND2HSV2 U39430 ( .A1(n34007), .A2(n34410), .ZN(n34185) );
  XNOR2HSV1 U39431 ( .A1(n34186), .A2(n34185), .ZN(n34189) );
  INHSV2 U39432 ( .I(n34187), .ZN(n35032) );
  CLKNHSV2 U39433 ( .I(n34227), .ZN(n47965) );
  CLKNAND2HSV2 U39434 ( .A1(n34190), .A2(n47965), .ZN(n34195) );
  NAND3HSV2 U39435 ( .A1(n34193), .A2(n47962), .A3(n34235), .ZN(n34194) );
  NAND2HSV4 U39436 ( .A1(n34195), .A2(n34194), .ZN(n34700) );
  NAND2HSV2 U39437 ( .A1(n34197), .A2(n34196), .ZN(n34198) );
  CLKNHSV2 U39438 ( .I(n34198), .ZN(n34202) );
  INHSV1 U39439 ( .I(n34199), .ZN(n34200) );
  NOR2HSV2 U39440 ( .A1(n34200), .A2(n33095), .ZN(n34201) );
  CLKNAND2HSV2 U39441 ( .A1(n34202), .A2(n34201), .ZN(n34212) );
  AND2HSV2 U39442 ( .A1(n34204), .A2(n34203), .Z(n34208) );
  INHSV2 U39443 ( .I(n34208), .ZN(n34209) );
  NAND4HSV4 U39444 ( .A1(n34212), .A2(n34211), .A3(n34210), .A4(n34209), .ZN(
        n34213) );
  NAND2HSV4 U39445 ( .A1(n34214), .A2(n34213), .ZN(n46594) );
  INHSV2 U39446 ( .I(n46594), .ZN(n34217) );
  AND2HSV2 U39447 ( .A1(n34220), .A2(n59345), .Z(n34215) );
  CLKAND2HSV2 U39448 ( .A1(n34865), .A2(n34215), .Z(n34216) );
  CLKNAND2HSV2 U39449 ( .A1(n34217), .A2(n34216), .ZN(n34225) );
  CLKNHSV1 U39450 ( .I(n34218), .ZN(n34219) );
  NOR2HSV4 U39451 ( .A1(n34219), .A2(n34727), .ZN(n46593) );
  NOR2HSV2 U39452 ( .A1(n46593), .A2(n34221), .ZN(n34223) );
  CLKAND2HSV2 U39453 ( .A1(n47788), .A2(\pe4/ti_7t [18]), .Z(n34222) );
  AOI21HSV4 U39454 ( .A1(n46594), .A2(n34223), .B(n34222), .ZN(n34224) );
  CLKNAND2HSV4 U39455 ( .A1(n34225), .A2(n34224), .ZN(n34446) );
  INHSV2 U39456 ( .I(n34226), .ZN(n47773) );
  CLKNAND2HSV1 U39457 ( .A1(n47967), .A2(n35021), .ZN(n34580) );
  INHSV4 U39458 ( .I(n34580), .ZN(n34701) );
  NOR2HSV1 U39459 ( .A1(n34834), .A2(\pe4/ti_7t [21]), .ZN(n34970) );
  CLKNAND2HSV3 U39460 ( .A1(n34227), .A2(n47963), .ZN(n34228) );
  INHSV3 U39461 ( .I(n34228), .ZN(n34336) );
  XNOR2HSV4 U39462 ( .A1(n34230), .A2(n25879), .ZN(n52821) );
  CLKNAND2HSV2 U39463 ( .A1(n34336), .A2(n47964), .ZN(n34577) );
  CLKNHSV2 U39464 ( .I(n34233), .ZN(n34234) );
  NOR2HSV3 U39465 ( .A1(n34235), .A2(n34234), .ZN(n34238) );
  AND2HSV2 U39466 ( .A1(n33094), .A2(n47773), .Z(n34236) );
  CLKNAND2HSV2 U39467 ( .A1(n34446), .A2(n34236), .ZN(n34237) );
  NOR2HSV4 U39468 ( .A1(n34238), .A2(n34237), .ZN(n34337) );
  NAND2HSV2 U39469 ( .A1(n34446), .A2(n47655), .ZN(n34315) );
  CLKNAND2HSV1 U39470 ( .A1(n57324), .A2(\pe4/got [24]), .ZN(n34309) );
  NAND2HSV0 U39471 ( .A1(n34459), .A2(n34239), .ZN(n34306) );
  INHSV2 U39472 ( .I(n50207), .ZN(n34594) );
  CLKNAND2HSV1 U39473 ( .A1(n34352), .A2(n34594), .ZN(n34302) );
  NAND2HSV0 U39474 ( .A1(n35036), .A2(n59372), .ZN(n34296) );
  CLKNAND2HSV0 U39475 ( .A1(n34868), .A2(n59604), .ZN(n34292) );
  CLKNHSV0 U39476 ( .I(n33250), .ZN(n35508) );
  NAND2HSV2 U39477 ( .A1(n35508), .A2(n57926), .ZN(n34242) );
  NAND2HSV0 U39478 ( .A1(n34240), .A2(n57368), .ZN(n34241) );
  XOR2HSV0 U39479 ( .A1(n34242), .A2(n34241), .Z(n34247) );
  NAND2HSV0 U39480 ( .A1(n33726), .A2(n34243), .ZN(n34245) );
  NAND2HSV0 U39481 ( .A1(n34637), .A2(\pe4/bq[23] ), .ZN(n34244) );
  XOR2HSV0 U39482 ( .A1(n34245), .A2(n34244), .Z(n34246) );
  XOR2HSV0 U39483 ( .A1(n34247), .A2(n34246), .Z(n34251) );
  CLKNAND2HSV0 U39484 ( .A1(n35091), .A2(n58069), .ZN(n34633) );
  INHSV2 U39485 ( .I(n47818), .ZN(n57846) );
  XOR2HSV0 U39486 ( .A1(n34251), .A2(n34250), .Z(n34253) );
  CLKNHSV0 U39487 ( .I(n35099), .ZN(n35227) );
  CLKNAND2HSV0 U39488 ( .A1(n35227), .A2(n57820), .ZN(n34252) );
  XNOR2HSV1 U39489 ( .A1(n34253), .A2(n34252), .ZN(n34290) );
  NAND2HSV0 U39490 ( .A1(n57285), .A2(n57752), .ZN(n34289) );
  NAND2HSV0 U39491 ( .A1(n57384), .A2(n34254), .ZN(n34256) );
  NAND2HSV0 U39492 ( .A1(n34387), .A2(n34480), .ZN(n34255) );
  XOR2HSV0 U39493 ( .A1(n34256), .A2(n34255), .Z(n34260) );
  CLKNAND2HSV0 U39494 ( .A1(\pe4/aot [14]), .A2(n57134), .ZN(n34258) );
  INHSV2 U39495 ( .I(n49954), .ZN(n57888) );
  NAND2HSV0 U39496 ( .A1(n57888), .A2(n57157), .ZN(n34257) );
  XOR2HSV0 U39497 ( .A1(n34258), .A2(n34257), .Z(n34259) );
  XOR2HSV0 U39498 ( .A1(n34260), .A2(n34259), .Z(n34268) );
  NAND2HSV0 U39499 ( .A1(\pe4/aot [16]), .A2(n48069), .ZN(n34262) );
  INHSV1 U39500 ( .I(n48070), .ZN(n57691) );
  CLKNAND2HSV0 U39501 ( .A1(n34874), .A2(n57691), .ZN(n34261) );
  XOR2HSV0 U39502 ( .A1(n34262), .A2(n34261), .Z(n34266) );
  CLKNAND2HSV0 U39503 ( .A1(n59343), .A2(n34888), .ZN(n34264) );
  NAND2HSV0 U39504 ( .A1(n35533), .A2(\pe4/bq[16] ), .ZN(n34263) );
  XOR2HSV0 U39505 ( .A1(n34264), .A2(n34263), .Z(n34265) );
  XOR2HSV0 U39506 ( .A1(n34266), .A2(n34265), .Z(n34267) );
  XOR2HSV0 U39507 ( .A1(n34268), .A2(n34267), .Z(n34284) );
  NOR2HSV0 U39508 ( .A1(n44338), .A2(n35068), .ZN(n34270) );
  NAND2HSV0 U39509 ( .A1(n33727), .A2(\pe4/bq[12] ), .ZN(n34269) );
  XOR2HSV0 U39510 ( .A1(n34270), .A2(n34269), .Z(n34274) );
  NAND2HSV0 U39511 ( .A1(n59605), .A2(n34629), .ZN(n34272) );
  CLKNAND2HSV0 U39512 ( .A1(n59953), .A2(n33313), .ZN(n34271) );
  XOR2HSV0 U39513 ( .A1(n34272), .A2(n34271), .Z(n34273) );
  XOR2HSV0 U39514 ( .A1(n34274), .A2(n34273), .Z(n34282) );
  NAND2HSV0 U39515 ( .A1(n34770), .A2(\pe4/pvq [21]), .ZN(n34275) );
  XOR2HSV0 U39516 ( .A1(n34275), .A2(\pe4/phq [21]), .Z(n34280) );
  NAND2HSV0 U39517 ( .A1(\pe4/aot [17]), .A2(n50007), .ZN(n34779) );
  OAI22HSV0 U39518 ( .A1(n34276), .A2(n49982), .B1(n35175), .B2(n57260), .ZN(
        n34277) );
  OAI21HSV0 U39519 ( .A1(n34779), .A2(n34278), .B(n34277), .ZN(n34279) );
  XOR2HSV0 U39520 ( .A1(n34280), .A2(n34279), .Z(n34281) );
  XNOR2HSV1 U39521 ( .A1(n34282), .A2(n34281), .ZN(n34283) );
  XNOR2HSV1 U39522 ( .A1(n34284), .A2(n34283), .ZN(n34287) );
  CLKNHSV0 U39523 ( .I(n50042), .ZN(n35490) );
  CLKNAND2HSV1 U39524 ( .A1(n59382), .A2(n35490), .ZN(n34286) );
  XNOR2HSV1 U39525 ( .A1(n34287), .A2(n34286), .ZN(n34288) );
  XOR3HSV2 U39526 ( .A1(n34290), .A2(n34289), .A3(n34288), .Z(n34291) );
  XNOR2HSV1 U39527 ( .A1(n34292), .A2(n34291), .ZN(n34294) );
  CLKNAND2HSV0 U39528 ( .A1(n57526), .A2(n59353), .ZN(n34293) );
  XNOR2HSV1 U39529 ( .A1(n34294), .A2(n34293), .ZN(n34295) );
  XNOR2HSV1 U39530 ( .A1(n34296), .A2(n34295), .ZN(n34298) );
  NAND2HSV0 U39531 ( .A1(n34595), .A2(n35321), .ZN(n34297) );
  XNOR2HSV1 U39532 ( .A1(n34298), .A2(n34297), .ZN(n34300) );
  NAND2HSV0 U39533 ( .A1(n35401), .A2(n59386), .ZN(n34299) );
  XOR2HSV0 U39534 ( .A1(n34300), .A2(n34299), .Z(n34301) );
  XNOR2HSV1 U39535 ( .A1(n34302), .A2(n34301), .ZN(n34304) );
  NAND2HSV0 U39536 ( .A1(n34405), .A2(n34351), .ZN(n34303) );
  XNOR2HSV1 U39537 ( .A1(n34304), .A2(n34303), .ZN(n34305) );
  XNOR2HSV1 U39538 ( .A1(n34306), .A2(n34305), .ZN(n34308) );
  CLKNAND2HSV1 U39539 ( .A1(n25894), .A2(n57190), .ZN(n34307) );
  XOR3HSV2 U39540 ( .A1(n34309), .A2(n34308), .A3(n34307), .Z(n34310) );
  INHSV2 U39541 ( .I(n34592), .ZN(n34457) );
  NAND2HSV2 U39542 ( .A1(n34409), .A2(n34410), .ZN(n34312) );
  CLKNAND2HSV2 U39543 ( .A1(n29758), .A2(n35032), .ZN(n34311) );
  XOR3HSV2 U39544 ( .A1(n34313), .A2(n34312), .A3(n34311), .Z(n34314) );
  CLKNAND2HSV0 U39545 ( .A1(n34317), .A2(n33522), .ZN(n34318) );
  CLKNAND2HSV2 U39546 ( .A1(n34321), .A2(n34350), .ZN(n34332) );
  INHSV4 U39547 ( .I(n35286), .ZN(n59345) );
  NAND2HSV0 U39548 ( .A1(n34343), .A2(n59345), .ZN(n34322) );
  NOR2HSV2 U39549 ( .A1(n34345), .A2(n34322), .ZN(n34326) );
  CLKNHSV0 U39550 ( .I(n34323), .ZN(n34324) );
  CLKNAND2HSV1 U39551 ( .A1(n34326), .A2(n34347), .ZN(n34331) );
  NOR2HSV2 U39552 ( .A1(n34220), .A2(n34327), .ZN(n34346) );
  CLKNHSV0 U39553 ( .I(n34346), .ZN(n34329) );
  OR2HSV1 U39554 ( .A1(n34329), .A2(n34328), .Z(n34330) );
  NAND3HSV4 U39555 ( .A1(n34332), .A2(n34331), .A3(n34330), .ZN(n34433) );
  XNOR2HSV4 U39556 ( .A1(n34434), .A2(n34433), .ZN(n34587) );
  CLKNHSV0 U39557 ( .I(n34696), .ZN(n34422) );
  MUX2NHSV2 U39558 ( .I0(n47965), .I1(n34336), .S(n47964), .ZN(n34338) );
  NAND2HSV2 U39559 ( .A1(n34338), .A2(n34337), .ZN(n34424) );
  CLKNHSV0 U39560 ( .I(n34424), .ZN(n34339) );
  INHSV4 U39561 ( .I(n34451), .ZN(n34341) );
  CLKNAND2HSV2 U39562 ( .A1(n34575), .A2(n34587), .ZN(n34697) );
  INHSV2 U39563 ( .I(n34860), .ZN(n34717) );
  CLKNAND2HSV1 U39564 ( .A1(n34697), .A2(n34717), .ZN(n34421) );
  CLKNHSV2 U39565 ( .I(n34343), .ZN(n34344) );
  AOI21HSV4 U39566 ( .A1(n34348), .A2(n34347), .B(n34346), .ZN(n34686) );
  INHSV1 U39567 ( .I(n34108), .ZN(n35487) );
  NAND2HSV2 U39568 ( .A1(n34446), .A2(n35032), .ZN(n34415) );
  CLKNAND2HSV1 U39569 ( .A1(n34352), .A2(n59386), .ZN(n34404) );
  INHSV2 U39570 ( .I(n47861), .ZN(n34797) );
  NAND2HSV2 U39571 ( .A1(n57404), .A2(n34797), .ZN(n34398) );
  NAND2HSV0 U39572 ( .A1(n59605), .A2(n57459), .ZN(n50342) );
  XOR2HSV0 U39573 ( .A1(n34353), .A2(n50342), .Z(n34366) );
  CLKNHSV1 U39574 ( .I(n53217), .ZN(n57139) );
  NAND2HSV2 U39575 ( .A1(\pe4/aot [14]), .A2(n57139), .ZN(n50363) );
  CLKNHSV1 U39576 ( .I(\pe4/bq[14] ), .ZN(n57387) );
  OAI22HSV0 U39577 ( .A1(n34479), .A2(n57387), .B1(n34470), .B2(n35043), .ZN(
        n34354) );
  OAI21HSV0 U39578 ( .A1(n34355), .A2(n50363), .B(n34354), .ZN(n34356) );
  NAND2HSV0 U39579 ( .A1(\pe4/aot [22]), .A2(\pe4/bq[21] ), .ZN(n50350) );
  XNOR2HSV1 U39580 ( .A1(n34356), .A2(n50350), .ZN(n34365) );
  CLKNAND2HSV0 U39581 ( .A1(n58163), .A2(n57134), .ZN(n34358) );
  NAND2HSV0 U39582 ( .A1(\pe4/got [11]), .A2(n57157), .ZN(n34357) );
  XOR2HSV0 U39583 ( .A1(n34358), .A2(n34357), .Z(n34363) );
  NAND2HSV0 U39584 ( .A1(n34240), .A2(n34359), .ZN(n34361) );
  NAND2HSV0 U39585 ( .A1(\pe4/aot [17]), .A2(n34629), .ZN(n34360) );
  XOR2HSV0 U39586 ( .A1(n34361), .A2(n34360), .Z(n34362) );
  XOR2HSV0 U39587 ( .A1(n34363), .A2(n34362), .Z(n34364) );
  CLKNHSV0 U39588 ( .I(n50042), .ZN(n59630) );
  CLKNAND2HSV1 U39589 ( .A1(n57384), .A2(n57785), .ZN(n34368) );
  CLKNAND2HSV0 U39590 ( .A1(n35508), .A2(n49943), .ZN(n34367) );
  XOR2HSV0 U39591 ( .A1(n34368), .A2(n34367), .Z(n34372) );
  NAND2HSV0 U39592 ( .A1(n59683), .A2(n33934), .ZN(n34370) );
  NAND2HSV0 U39593 ( .A1(\pe4/aot [24]), .A2(n57368), .ZN(n34369) );
  XOR2HSV0 U39594 ( .A1(n34370), .A2(n34369), .Z(n34371) );
  XOR2HSV0 U39595 ( .A1(n34372), .A2(n34371), .Z(n34380) );
  CLKNHSV0 U39596 ( .I(n34631), .ZN(n47709) );
  CLKNAND2HSV1 U39597 ( .A1(n47709), .A2(n34480), .ZN(n34374) );
  NAND2HSV0 U39598 ( .A1(n34874), .A2(n50007), .ZN(n34373) );
  XOR2HSV0 U39599 ( .A1(n34374), .A2(n34373), .Z(n34378) );
  NAND2HSV0 U39600 ( .A1(n34637), .A2(n34044), .ZN(n34376) );
  NAND2HSV0 U39601 ( .A1(\pe4/aot [16]), .A2(n35207), .ZN(n34375) );
  XOR2HSV0 U39602 ( .A1(n34376), .A2(n34375), .Z(n34377) );
  XOR2HSV0 U39603 ( .A1(n34378), .A2(n34377), .Z(n34379) );
  XOR2HSV0 U39604 ( .A1(n34380), .A2(n34379), .Z(n34395) );
  NAND2HSV0 U39605 ( .A1(n57852), .A2(n48069), .ZN(n34382) );
  NAND2HSV0 U39606 ( .A1(n35533), .A2(n57846), .ZN(n34381) );
  XOR2HSV0 U39607 ( .A1(n34382), .A2(n34381), .Z(n34386) );
  NAND2HSV0 U39608 ( .A1(n34743), .A2(\pe4/bq[23] ), .ZN(n34384) );
  NAND2HSV0 U39609 ( .A1(n34873), .A2(n34738), .ZN(n34383) );
  XOR2HSV0 U39610 ( .A1(n34384), .A2(n34383), .Z(n34385) );
  XOR2HSV0 U39611 ( .A1(n34386), .A2(n34385), .Z(n34394) );
  NAND2HSV0 U39612 ( .A1(n34387), .A2(\pe4/bq[12] ), .ZN(n34389) );
  NAND2HSV0 U39613 ( .A1(n35201), .A2(\pe4/bq[11] ), .ZN(n34388) );
  XOR2HSV0 U39614 ( .A1(n34389), .A2(n34388), .Z(n34392) );
  NAND2HSV0 U39615 ( .A1(n34770), .A2(\pe4/pvq [22]), .ZN(n34390) );
  XOR2HSV0 U39616 ( .A1(n34390), .A2(\pe4/phq [22]), .Z(n34391) );
  XOR2HSV0 U39617 ( .A1(n34392), .A2(n34391), .Z(n34393) );
  INHSV2 U39618 ( .I(n58189), .ZN(n47657) );
  XNOR2HSV1 U39619 ( .A1(n34398), .A2(n34397), .ZN(n34400) );
  NAND2HSV0 U39620 ( .A1(n34595), .A2(n59372), .ZN(n34399) );
  XNOR2HSV1 U39621 ( .A1(n34400), .A2(n34399), .ZN(n34402) );
  CLKNAND2HSV0 U39622 ( .A1(n57679), .A2(n35321), .ZN(n34401) );
  XOR2HSV0 U39623 ( .A1(n34402), .A2(n34401), .Z(n34403) );
  XNOR2HSV1 U39624 ( .A1(n34404), .A2(n34403), .ZN(n34406) );
  CLKNHSV0 U39625 ( .I(n34408), .ZN(n35570) );
  CLKNAND2HSV3 U39626 ( .A1(n29759), .A2(n34410), .ZN(n34411) );
  XOR3HSV2 U39627 ( .A1(n34413), .A2(n34412), .A3(n34411), .Z(n34414) );
  XNOR2HSV4 U39628 ( .A1(n34415), .A2(n34414), .ZN(n34417) );
  IOA21HSV4 U39629 ( .A1(n34733), .A2(n35487), .B(n34417), .ZN(n34427) );
  NOR2HSV4 U39630 ( .A1(n34417), .A2(n34416), .ZN(n34418) );
  CLKNAND2HSV2 U39631 ( .A1(n34418), .A2(n34733), .ZN(n34426) );
  CLKNAND2HSV1 U39632 ( .A1(n34721), .A2(n34717), .ZN(n34420) );
  OAI21HSV2 U39633 ( .A1(n34422), .A2(n34421), .B(n34420), .ZN(n34559) );
  INAND2HSV2 U39634 ( .A1(n34559), .B1(n34019), .ZN(n34445) );
  NAND2HSV2 U39635 ( .A1(n34423), .A2(\pe4/ti_7t [20]), .ZN(n34699) );
  CLKNAND2HSV2 U39636 ( .A1(n34424), .A2(n34699), .ZN(n34425) );
  INHSV4 U39637 ( .I(n34425), .ZN(n34450) );
  NAND2HSV4 U39638 ( .A1(n34340), .A2(n34450), .ZN(n34429) );
  BUFHSV8 U39639 ( .I(n34429), .Z(n34967) );
  CLKNAND2HSV4 U39640 ( .A1(n34426), .A2(n34427), .ZN(n34702) );
  INHSV4 U39641 ( .I(n34702), .ZN(n34726) );
  AND2HSV2 U39642 ( .A1(n34967), .A2(n34726), .Z(n34432) );
  BUFHSV2 U39643 ( .I(n34702), .Z(n34441) );
  CLKNAND2HSV2 U39644 ( .A1(n34429), .A2(n34428), .ZN(n34724) );
  NAND2HSV2 U39645 ( .A1(n34441), .A2(n34724), .ZN(n34430) );
  CLKNAND2HSV2 U39646 ( .A1(n34430), .A2(n34717), .ZN(n34431) );
  NOR2HSV4 U39647 ( .A1(n34432), .A2(n34431), .ZN(n34560) );
  XNOR2HSV4 U39648 ( .A1(n34434), .A2(n34433), .ZN(n34581) );
  INAND2HSV2 U39649 ( .A1(n34436), .B1(n34702), .ZN(n34437) );
  CLKNAND2HSV1 U39650 ( .A1(n34437), .A2(n34571), .ZN(n34438) );
  INHSV2 U39651 ( .I(n34438), .ZN(n34716) );
  INHSV2 U39652 ( .I(n34716), .ZN(n34439) );
  NOR2HSV8 U39653 ( .A1(n34440), .A2(n34439), .ZN(n34858) );
  CLKNAND2HSV0 U39654 ( .A1(n34724), .A2(n34726), .ZN(n34442) );
  CLKNAND2HSV3 U39655 ( .A1(n34443), .A2(n34442), .ZN(n34557) );
  NAND2HSV2 U39656 ( .A1(n34858), .A2(n34557), .ZN(n34444) );
  BUFHSV4 U39657 ( .I(n34446), .Z(n35320) );
  CLKNAND2HSV1 U39658 ( .A1(n35320), .A2(n35318), .ZN(n34449) );
  BUFHSV2 U39659 ( .I(n34447), .Z(n58060) );
  BUFHSV2 U39660 ( .I(n58060), .Z(n49951) );
  CLKAND2HSV2 U39661 ( .A1(n49951), .A2(n59603), .Z(n34448) );
  XNOR2HSV1 U39662 ( .A1(n34449), .A2(n34448), .ZN(n34453) );
  AOI21HSV1 U39663 ( .A1(n34967), .A2(n59350), .B(n34453), .ZN(n34454) );
  AOI21HSV2 U39664 ( .A1(n34455), .A2(n50065), .B(n34454), .ZN(n34554) );
  BUFHSV2 U39665 ( .I(n34456), .Z(n35035) );
  CLKNHSV2 U39666 ( .I(n34457), .ZN(n59526) );
  INHSV2 U39667 ( .I(n35488), .ZN(n57309) );
  NAND2HSV0 U39668 ( .A1(n59526), .A2(n57309), .ZN(n34550) );
  BUFHSV3 U39669 ( .I(n34593), .Z(n44695) );
  BUFHSV2 U39670 ( .I(n44695), .Z(n34866) );
  INHSV2 U39671 ( .I(n50207), .ZN(n34948) );
  NAND2HSV2 U39672 ( .A1(n34866), .A2(n34948), .ZN(n34546) );
  BUFHSV2 U39673 ( .I(n34458), .Z(n35489) );
  CLKNAND2HSV1 U39674 ( .A1(n35489), .A2(\pe4/got [19]), .ZN(n34544) );
  NAND2HSV2 U39675 ( .A1(n57209), .A2(n57754), .ZN(n34541) );
  NAND2HSV2 U39676 ( .A1(n34352), .A2(\pe4/got [16]), .ZN(n34536) );
  NAND2HSV2 U39677 ( .A1(n57530), .A2(n35400), .ZN(n34530) );
  NAND2HSV0 U39678 ( .A1(n47733), .A2(n58153), .ZN(n34526) );
  BUFHSV2 U39679 ( .I(n59382), .Z(n57251) );
  INHSV1 U39680 ( .I(\pe4/got [9]), .ZN(n59628) );
  CLKNAND2HSV1 U39681 ( .A1(n57251), .A2(n58041), .ZN(n34462) );
  INHSV2 U39682 ( .I(\pe4/got [8]), .ZN(n58253) );
  NOR2HSV0 U39683 ( .A1(n35099), .A2(n58253), .ZN(n34461) );
  XNOR2HSV1 U39684 ( .A1(n34462), .A2(n34461), .ZN(n34524) );
  NAND2HSV0 U39685 ( .A1(n57166), .A2(n59663), .ZN(n34523) );
  CLKNAND2HSV0 U39686 ( .A1(n35377), .A2(n35184), .ZN(n34465) );
  INHSV2 U39687 ( .I(n48026), .ZN(n57089) );
  CLKNAND2HSV1 U39688 ( .A1(n59951), .A2(n57089), .ZN(n34464) );
  XOR2HSV0 U39689 ( .A1(n34465), .A2(n34464), .Z(n34469) );
  NAND2HSV0 U39690 ( .A1(n57499), .A2(n57139), .ZN(n34467) );
  CLKNAND2HSV0 U39691 ( .A1(\pe4/aot [20]), .A2(n57929), .ZN(n34466) );
  XOR2HSV0 U39692 ( .A1(n34467), .A2(n34466), .Z(n34468) );
  XOR2HSV0 U39693 ( .A1(n34469), .A2(n34468), .Z(n34476) );
  CLKNHSV0 U39694 ( .I(n47661), .ZN(n57210) );
  CLKNAND2HSV0 U39695 ( .A1(n57210), .A2(\pe4/bq[11] ), .ZN(n34472) );
  NAND2HSV0 U39696 ( .A1(n59952), .A2(n57476), .ZN(n34471) );
  XOR2HSV0 U39697 ( .A1(n34472), .A2(n34471), .Z(n34473) );
  XOR2HSV0 U39698 ( .A1(n34474), .A2(n34473), .Z(n34475) );
  XOR2HSV0 U39699 ( .A1(n34476), .A2(n34475), .Z(n34495) );
  NAND2HSV0 U39700 ( .A1(n57014), .A2(n33711), .ZN(n34478) );
  NAND2HSV0 U39701 ( .A1(n34874), .A2(\pe4/bq[20] ), .ZN(n34477) );
  XOR2HSV0 U39702 ( .A1(n34478), .A2(n34477), .Z(n34484) );
  CLKNHSV0 U39703 ( .I(n34479), .ZN(n57138) );
  CLKNAND2HSV1 U39704 ( .A1(n57138), .A2(n58116), .ZN(n34482) );
  NAND2HSV0 U39705 ( .A1(n33947), .A2(n34480), .ZN(n34481) );
  XOR2HSV0 U39706 ( .A1(n34482), .A2(n34481), .Z(n34483) );
  XOR2HSV0 U39707 ( .A1(n34484), .A2(n34483), .Z(n34493) );
  NOR2HSV0 U39708 ( .A1(n46143), .A2(n48024), .ZN(n34487) );
  INHSV2 U39709 ( .I(\pe4/aot [9]), .ZN(n34897) );
  CLKNAND2HSV1 U39710 ( .A1(\pe4/aot [9]), .A2(n34021), .ZN(n34486) );
  XOR2HSV0 U39711 ( .A1(n34487), .A2(n34486), .Z(n34491) );
  CLKNHSV0 U39712 ( .I(n50064), .ZN(n59957) );
  NAND2HSV0 U39713 ( .A1(n59957), .A2(n47679), .ZN(n34489) );
  INHSV2 U39714 ( .I(n57775), .ZN(n57506) );
  NAND2HSV0 U39715 ( .A1(n57506), .A2(n33611), .ZN(n34488) );
  XOR2HSV0 U39716 ( .A1(n34489), .A2(n34488), .Z(n34490) );
  XOR2HSV0 U39717 ( .A1(n34491), .A2(n34490), .Z(n34492) );
  XOR2HSV0 U39718 ( .A1(n34493), .A2(n34492), .Z(n34494) );
  XOR2HSV0 U39719 ( .A1(n34495), .A2(n34494), .Z(n34521) );
  BUFHSV2 U39720 ( .I(n34496), .Z(n53218) );
  NAND2HSV2 U39721 ( .A1(n48058), .A2(\pe4/pvq [26]), .ZN(n34497) );
  XNOR2HSV1 U39722 ( .A1(n34497), .A2(\pe4/phq [26]), .ZN(n34500) );
  NAND2HSV0 U39723 ( .A1(n59343), .A2(n35207), .ZN(n34499) );
  XNOR2HSV1 U39724 ( .A1(n34500), .A2(n34499), .ZN(n34519) );
  BUFHSV2 U39725 ( .I(\pe4/bq[9] ), .Z(n35220) );
  CLKNAND2HSV0 U39726 ( .A1(n47709), .A2(n35220), .ZN(n34503) );
  INHSV2 U39727 ( .I(n50114), .ZN(n35323) );
  CLKNAND2HSV1 U39728 ( .A1(n47692), .A2(n35323), .ZN(n34502) );
  XOR2HSV0 U39729 ( .A1(n34503), .A2(n34502), .Z(n34507) );
  CLKNHSV0 U39730 ( .I(n33250), .ZN(n35326) );
  CLKNAND2HSV0 U39731 ( .A1(n35326), .A2(n57986), .ZN(n34505) );
  NAND2HSV0 U39732 ( .A1(n47718), .A2(n33110), .ZN(n34504) );
  XOR2HSV0 U39733 ( .A1(n34505), .A2(n34504), .Z(n34506) );
  XOR2HSV0 U39734 ( .A1(n34507), .A2(n34506), .Z(n34518) );
  NAND2HSV2 U39735 ( .A1(\pe4/aot [11]), .A2(n35194), .ZN(n34509) );
  INHSV2 U39736 ( .I(n44338), .ZN(n35191) );
  NAND2HSV0 U39737 ( .A1(n35191), .A2(n33713), .ZN(n34508) );
  XOR2HSV0 U39738 ( .A1(n34509), .A2(n34508), .Z(n34517) );
  INHSV2 U39739 ( .I(n57918), .ZN(n35347) );
  NAND2HSV0 U39740 ( .A1(n35347), .A2(n50007), .ZN(n34511) );
  NAND2HSV0 U39741 ( .A1(n57218), .A2(\pe4/bq[21] ), .ZN(n34510) );
  XOR2HSV0 U39742 ( .A1(n34511), .A2(n34510), .Z(n34515) );
  NAND2HSV2 U39743 ( .A1(n33965), .A2(n57926), .ZN(n34513) );
  INHSV2 U39744 ( .I(\pe4/aot [7]), .ZN(n35042) );
  NAND2HSV0 U39745 ( .A1(n58198), .A2(n34888), .ZN(n34512) );
  XOR2HSV0 U39746 ( .A1(n34513), .A2(n34512), .Z(n34514) );
  XOR2HSV0 U39747 ( .A1(n34515), .A2(n34514), .Z(n34516) );
  XOR4HSV1 U39748 ( .A1(n34519), .A2(n34518), .A3(n34517), .A4(n34516), .Z(
        n34520) );
  XNOR2HSV1 U39749 ( .A1(n34521), .A2(n34520), .ZN(n34522) );
  XOR3HSV2 U39750 ( .A1(n34524), .A2(n34523), .A3(n34522), .Z(n34525) );
  XNOR2HSV1 U39751 ( .A1(n34526), .A2(n34525), .ZN(n34528) );
  CLKNHSV0 U39752 ( .I(n49954), .ZN(n59631) );
  CLKNAND2HSV1 U39753 ( .A1(n33498), .A2(n59631), .ZN(n34527) );
  XNOR2HSV1 U39754 ( .A1(n34528), .A2(n34527), .ZN(n34529) );
  XNOR2HSV1 U39755 ( .A1(n34530), .A2(n34529), .ZN(n34532) );
  BUFHSV2 U39756 ( .I(n34595), .Z(n35555) );
  CLKNHSV0 U39757 ( .I(n50042), .ZN(n35243) );
  CLKNAND2HSV1 U39758 ( .A1(n35555), .A2(n35243), .ZN(n34531) );
  XNOR2HSV1 U39759 ( .A1(n34532), .A2(n34531), .ZN(n34534) );
  NAND2HSV0 U39760 ( .A1(n57679), .A2(n34937), .ZN(n34533) );
  XOR2HSV0 U39761 ( .A1(n34534), .A2(n34533), .Z(n34535) );
  XNOR2HSV1 U39762 ( .A1(n34536), .A2(n34535), .ZN(n34539) );
  CLKNHSV0 U39763 ( .I(n34537), .ZN(n57414) );
  CLKNAND2HSV0 U39764 ( .A1(n57414), .A2(n35167), .ZN(n34538) );
  XNOR2HSV1 U39765 ( .A1(n34539), .A2(n34538), .ZN(n34540) );
  XNOR2HSV1 U39766 ( .A1(n34541), .A2(n34540), .ZN(n34543) );
  INHSV2 U39767 ( .I(\pe4/got [20]), .ZN(n57830) );
  CLKNAND2HSV1 U39768 ( .A1(n33918), .A2(n57564), .ZN(n34542) );
  XOR3HSV2 U39769 ( .A1(n34544), .A2(n34543), .A3(n34542), .Z(n34545) );
  XNOR2HSV1 U39770 ( .A1(n34546), .A2(n34545), .ZN(n34548) );
  XNOR2HSV1 U39771 ( .A1(n34548), .A2(n34547), .ZN(n34549) );
  XNOR2HSV1 U39772 ( .A1(n34550), .A2(n34549), .ZN(n34551) );
  CLKXOR2HSV4 U39773 ( .A1(n34554), .A2(n34553), .Z(n34561) );
  INHSV2 U39774 ( .I(n34561), .ZN(n34555) );
  CLKNAND2HSV2 U39775 ( .A1(n34556), .A2(n34555), .ZN(n34564) );
  CLKNAND2HSV4 U39776 ( .A1(n34858), .A2(n34557), .ZN(n34558) );
  OAI21HSV4 U39777 ( .A1(n34560), .A2(n34559), .B(n34558), .ZN(n35428) );
  CLKNAND2HSV3 U39778 ( .A1(n34564), .A2(n34563), .ZN(n34574) );
  INHSV2 U39779 ( .I(n34581), .ZN(n51449) );
  IOA21HSV2 U39780 ( .A1(n34819), .A2(n47778), .B(n51449), .ZN(n51448) );
  INHSV2 U39781 ( .I(n51448), .ZN(n34572) );
  NAND2HSV0 U39782 ( .A1(n47778), .A2(n34819), .ZN(n51450) );
  INHSV1 U39783 ( .I(n51450), .ZN(n34569) );
  NOR2HSV2 U39784 ( .A1(n51449), .A2(n34565), .ZN(n34568) );
  AND2HSV2 U39785 ( .A1(n34566), .A2(\pe4/ti_7t [21]), .Z(n34567) );
  AOI21HSV2 U39786 ( .A1(n34569), .A2(n34568), .B(n34567), .ZN(n34570) );
  IOA21HSV4 U39787 ( .A1(n34572), .A2(n34571), .B(n34570), .ZN(n47842) );
  CLKAND2HSV2 U39788 ( .A1(n47842), .A2(n34410), .Z(n34573) );
  XNOR2HSV4 U39789 ( .A1(n34574), .A2(n34573), .ZN(n35006) );
  NAND2HSV2 U39790 ( .A1(n34575), .A2(n34581), .ZN(n34823) );
  NOR2HSV0 U39791 ( .A1(n34970), .A2(n34712), .ZN(n34576) );
  AND2HSV4 U39792 ( .A1(n34823), .A2(n34576), .Z(n34694) );
  CLKNHSV1 U39793 ( .I(n33095), .ZN(n34837) );
  CLKNHSV0 U39794 ( .I(n34700), .ZN(n34584) );
  NAND2HSV2 U39795 ( .A1(n34584), .A2(n34583), .ZN(n34585) );
  INHSV3 U39796 ( .I(n34969), .ZN(n34590) );
  CLKNHSV2 U39797 ( .I(n35013), .ZN(n34588) );
  INHSV2 U39798 ( .I(n25875), .ZN(n34589) );
  NOR2HSV4 U39799 ( .A1(n34590), .A2(n34589), .ZN(n34693) );
  CLKNAND2HSV2 U39800 ( .A1(n34694), .A2(n34693), .ZN(n34710) );
  CLKNHSV0 U39801 ( .I(n34686), .ZN(n34683) );
  CLKNAND2HSV2 U39802 ( .A1(n29758), .A2(n59350), .ZN(n34678) );
  CLKNAND2HSV1 U39803 ( .A1(n34592), .A2(n47771), .ZN(n34676) );
  CLKNAND2HSV0 U39804 ( .A1(n34593), .A2(n59603), .ZN(n34671) );
  NAND2HSV0 U39805 ( .A1(n46601), .A2(n59601), .ZN(n34669) );
  NAND2HSV2 U39806 ( .A1(n34459), .A2(n34594), .ZN(n34666) );
  BUFHSV2 U39807 ( .I(n25616), .Z(n59682) );
  NAND2HSV2 U39808 ( .A1(n59682), .A2(n59602), .ZN(n34662) );
  NAND2HSV0 U39809 ( .A1(n34595), .A2(n34797), .ZN(n34660) );
  NAND2HSV0 U39810 ( .A1(n35036), .A2(n59604), .ZN(n34657) );
  NAND2HSV0 U39811 ( .A1(n34868), .A2(n59630), .ZN(n34653) );
  CLKNHSV0 U39812 ( .I(n49954), .ZN(n35397) );
  CLKNAND2HSV0 U39813 ( .A1(n59382), .A2(n35397), .ZN(n34597) );
  NAND2HSV0 U39814 ( .A1(n35227), .A2(n58153), .ZN(n34596) );
  XNOR2HSV1 U39815 ( .A1(n34597), .A2(n34596), .ZN(n34651) );
  NAND2HSV0 U39816 ( .A1(n59501), .A2(n59629), .ZN(n34650) );
  NAND2HSV0 U39817 ( .A1(n34873), .A2(n57134), .ZN(n34600) );
  NAND2HSV0 U39818 ( .A1(n57852), .A2(n34598), .ZN(n34599) );
  XOR2HSV0 U39819 ( .A1(n34600), .A2(n34599), .Z(n34604) );
  NAND2HSV0 U39820 ( .A1(\pe4/aot [17]), .A2(n57459), .ZN(n34602) );
  CLKNAND2HSV0 U39821 ( .A1(n34387), .A2(\pe4/bq[11] ), .ZN(n34601) );
  XOR2HSV0 U39822 ( .A1(n34602), .A2(n34601), .Z(n34603) );
  XOR2HSV0 U39823 ( .A1(n34604), .A2(n34603), .Z(n34612) );
  NAND2HSV0 U39824 ( .A1(n58163), .A2(n33313), .ZN(n34606) );
  NAND2HSV0 U39825 ( .A1(\pe4/got [10]), .A2(n57157), .ZN(n34605) );
  XOR2HSV0 U39826 ( .A1(n34606), .A2(n34605), .Z(n34610) );
  NAND2HSV0 U39827 ( .A1(\pe4/aot [14]), .A2(n33966), .ZN(n34608) );
  NAND2HSV0 U39828 ( .A1(n57384), .A2(n57368), .ZN(n34607) );
  XOR2HSV0 U39829 ( .A1(n34608), .A2(n34607), .Z(n34609) );
  XOR2HSV0 U39830 ( .A1(n34610), .A2(n34609), .Z(n34611) );
  XOR2HSV0 U39831 ( .A1(n34612), .A2(n34611), .Z(n34628) );
  NAND2HSV0 U39832 ( .A1(n34874), .A2(n57476), .ZN(n34614) );
  NAND2HSV0 U39833 ( .A1(n35201), .A2(\pe4/bq[10] ), .ZN(n34613) );
  XOR2HSV0 U39834 ( .A1(n34614), .A2(n34613), .Z(n34618) );
  NAND2HSV0 U39835 ( .A1(\pe4/aot [24]), .A2(n57906), .ZN(n34616) );
  NAND2HSV0 U39836 ( .A1(n35508), .A2(n57846), .ZN(n34615) );
  XOR2HSV0 U39837 ( .A1(n34616), .A2(n34615), .Z(n34617) );
  XOR2HSV0 U39838 ( .A1(n34618), .A2(n34617), .Z(n34626) );
  CLKNAND2HSV0 U39839 ( .A1(n47658), .A2(n49943), .ZN(n34620) );
  NAND2HSV0 U39840 ( .A1(\pe4/aot [10]), .A2(n33934), .ZN(n34619) );
  XOR2HSV0 U39841 ( .A1(n34620), .A2(n34619), .Z(n34624) );
  NAND2HSV0 U39842 ( .A1(n34743), .A2(n34044), .ZN(n34622) );
  NAND2HSV0 U39843 ( .A1(\pe4/aot [11]), .A2(n34738), .ZN(n34621) );
  XOR2HSV0 U39844 ( .A1(n34622), .A2(n34621), .Z(n34623) );
  XOR2HSV0 U39845 ( .A1(n34624), .A2(n34623), .Z(n34625) );
  XOR2HSV0 U39846 ( .A1(n34626), .A2(n34625), .Z(n34627) );
  XOR2HSV0 U39847 ( .A1(n34628), .A2(n34627), .Z(n34648) );
  NAND2HSV0 U39848 ( .A1(n57234), .A2(n34629), .ZN(n34912) );
  NAND2HSV0 U39849 ( .A1(n57499), .A2(n57926), .ZN(n57708) );
  XOR2HSV0 U39850 ( .A1(n34912), .A2(n57708), .Z(n34646) );
  NAND2HSV0 U39851 ( .A1(n48082), .A2(\pe4/pvq [23]), .ZN(n34630) );
  XOR2HSV0 U39852 ( .A1(n34630), .A2(\pe4/phq [23]), .Z(n34635) );
  CLKNAND2HSV1 U39853 ( .A1(n57210), .A2(\pe4/bq[12] ), .ZN(n34921) );
  OAI22HSV0 U39854 ( .A1(n34631), .A2(n57841), .B1(n47661), .B2(n57387), .ZN(
        n34632) );
  OAI21HSV1 U39855 ( .A1(n34633), .A2(n34921), .B(n34632), .ZN(n34634) );
  XNOR2HSV1 U39856 ( .A1(n34635), .A2(n34634), .ZN(n34645) );
  NAND2HSV0 U39857 ( .A1(n57218), .A2(n50007), .ZN(n34639) );
  NAND2HSV0 U39858 ( .A1(n34637), .A2(n34636), .ZN(n34638) );
  XOR2HSV0 U39859 ( .A1(n34639), .A2(n34638), .Z(n34643) );
  NAND2HSV0 U39860 ( .A1(n33965), .A2(n34243), .ZN(n34640) );
  XOR2HSV0 U39861 ( .A1(n34641), .A2(n34640), .Z(n34642) );
  XOR2HSV0 U39862 ( .A1(n34643), .A2(n34642), .Z(n34644) );
  XOR3HSV2 U39863 ( .A1(n34646), .A2(n34645), .A3(n34644), .Z(n34647) );
  XNOR2HSV1 U39864 ( .A1(n34648), .A2(n34647), .ZN(n34649) );
  XOR3HSV2 U39865 ( .A1(n34651), .A2(n34650), .A3(n34649), .Z(n34652) );
  XOR2HSV0 U39866 ( .A1(n34653), .A2(n34652), .Z(n34655) );
  CLKNAND2HSV0 U39867 ( .A1(n34396), .A2(n34937), .ZN(n34654) );
  XNOR2HSV1 U39868 ( .A1(n34655), .A2(n34654), .ZN(n34656) );
  XOR2HSV0 U39869 ( .A1(n34657), .A2(n34656), .Z(n34659) );
  NAND2HSV0 U39870 ( .A1(n57679), .A2(n59372), .ZN(n34658) );
  XOR3HSV2 U39871 ( .A1(n34660), .A2(n34659), .A3(n34658), .Z(n34661) );
  XNOR2HSV1 U39872 ( .A1(n34662), .A2(n34661), .ZN(n34664) );
  CLKNAND2HSV0 U39873 ( .A1(n57414), .A2(n57564), .ZN(n34663) );
  XNOR2HSV1 U39874 ( .A1(n34664), .A2(n34663), .ZN(n34665) );
  XNOR2HSV1 U39875 ( .A1(n34666), .A2(n34665), .ZN(n34668) );
  NAND2HSV2 U39876 ( .A1(n33918), .A2(n34239), .ZN(n34667) );
  XOR3HSV2 U39877 ( .A1(n34669), .A2(n34668), .A3(n34667), .Z(n34670) );
  XNOR2HSV1 U39878 ( .A1(n34671), .A2(n34670), .ZN(n34674) );
  CLKNAND2HSV0 U39879 ( .A1(n59932), .A2(n34672), .ZN(n34673) );
  XNOR2HSV1 U39880 ( .A1(n34674), .A2(n34673), .ZN(n34675) );
  XNOR2HSV1 U39881 ( .A1(n34676), .A2(n34675), .ZN(n34677) );
  BUFHSV2 U39882 ( .I(n57199), .Z(n57453) );
  CLKNHSV0 U39883 ( .I(n34684), .ZN(n34679) );
  AOI21HSV2 U39884 ( .A1(n34683), .A2(n34682), .B(n34681), .ZN(n34688) );
  NAND3HSV0 U39885 ( .A1(n34686), .A2(n34685), .A3(n34684), .ZN(n34687) );
  NAND2HSV2 U39886 ( .A1(n34688), .A2(n34687), .ZN(n34690) );
  INHSV2 U39887 ( .I(n33564), .ZN(n34966) );
  CLKAND2HSV2 U39888 ( .A1(n35320), .A2(n34966), .Z(n34689) );
  CLKXOR2HSV2 U39889 ( .A1(n34690), .A2(n34689), .Z(n34692) );
  CLKNAND2HSV2 U39890 ( .A1(n34819), .A2(n35487), .ZN(n34691) );
  XNOR2HSV4 U39891 ( .A1(n34692), .A2(n34691), .ZN(n34695) );
  INHSV2 U39892 ( .I(n34695), .ZN(n34709) );
  NAND2HSV2 U39893 ( .A1(n34710), .A2(n34709), .ZN(n34984) );
  NAND2HSV2 U39894 ( .A1(n35483), .A2(\pe4/ti_7t [23]), .ZN(n34991) );
  CLKNAND2HSV2 U39895 ( .A1(n34984), .A2(n34991), .ZN(n34708) );
  NAND3HSV4 U39896 ( .A1(n34695), .A2(n34693), .A3(n34694), .ZN(n34711) );
  INHSV4 U39897 ( .I(n34844), .ZN(n34986) );
  XNOR2HSV4 U39898 ( .A1(n34703), .A2(n34702), .ZN(n34704) );
  XNOR2HSV4 U39899 ( .A1(n34723), .A2(n34704), .ZN(n60045) );
  INHSV2 U39900 ( .I(n34705), .ZN(n34706) );
  CLKNAND2HSV3 U39901 ( .A1(n60045), .A2(n34706), .ZN(n34989) );
  CLKNAND2HSV3 U39902 ( .A1(n34989), .A2(n34991), .ZN(n34707) );
  OAI21HSV4 U39903 ( .A1(n34708), .A2(n34986), .B(n34707), .ZN(n34831) );
  NAND2HSV4 U39904 ( .A1(n60045), .A2(n47772), .ZN(n34987) );
  NAND3HSV4 U39905 ( .A1(n34987), .A2(n34842), .A3(n29636), .ZN(n34829) );
  NOR2HSV2 U39906 ( .A1(n34856), .A2(n34712), .ZN(n34714) );
  NAND2HSV2 U39907 ( .A1(n34714), .A2(n34713), .ZN(n34720) );
  CLKNHSV0 U39908 ( .I(n34724), .ZN(n34715) );
  NAND2HSV2 U39909 ( .A1(n34715), .A2(n34726), .ZN(n34855) );
  NAND2HSV2 U39910 ( .A1(n34855), .A2(n34716), .ZN(n34719) );
  OAI22HSV4 U39911 ( .A1(n34720), .A2(n34719), .B1(n34718), .B2(n34717), .ZN(
        n34732) );
  INHSV1 U39912 ( .I(n34721), .ZN(n34722) );
  NAND2HSV2 U39913 ( .A1(n34723), .A2(n34722), .ZN(n34854) );
  NOR2HSV0 U39914 ( .A1(n34726), .A2(n34724), .ZN(n34725) );
  INHSV2 U39915 ( .I(n34725), .ZN(n34850) );
  NAND2HSV2 U39916 ( .A1(n35317), .A2(n34726), .ZN(n34849) );
  CLKNAND2HSV1 U39917 ( .A1(n34849), .A2(n52755), .ZN(n34728) );
  INHSV2 U39918 ( .I(n34728), .ZN(n34729) );
  CLKNAND2HSV1 U39919 ( .A1(n34850), .A2(n34729), .ZN(n34730) );
  NOR2HSV2 U39920 ( .A1(n34854), .A2(n34730), .ZN(n34731) );
  NOR2HSV4 U39921 ( .A1(n34732), .A2(n34731), .ZN(n34826) );
  CLKBUFHSV4 U39922 ( .I(n34733), .Z(n59665) );
  CLKNAND2HSV1 U39923 ( .A1(n35320), .A2(n59350), .ZN(n34816) );
  NAND2HSV2 U39924 ( .A1(n34866), .A2(n34239), .ZN(n34810) );
  CLKNAND2HSV1 U39925 ( .A1(n35489), .A2(n34948), .ZN(n34808) );
  CLKNAND2HSV1 U39926 ( .A1(n34459), .A2(n57564), .ZN(n34805) );
  NAND2HSV0 U39927 ( .A1(n35322), .A2(n59372), .ZN(n34801) );
  CLKNAND2HSV1 U39928 ( .A1(n57404), .A2(n34937), .ZN(n34794) );
  NAND2HSV0 U39929 ( .A1(n34868), .A2(n59629), .ZN(n34790) );
  NAND2HSV0 U39930 ( .A1(n59382), .A2(n58153), .ZN(n34735) );
  NAND2HSV0 U39931 ( .A1(n35227), .A2(n57646), .ZN(n34734) );
  XNOR2HSV1 U39932 ( .A1(n34735), .A2(n34734), .ZN(n34788) );
  NAND2HSV0 U39933 ( .A1(n35340), .A2(n59631), .ZN(n34787) );
  NAND2HSV0 U39934 ( .A1(n57218), .A2(n57476), .ZN(n34737) );
  NAND2HSV0 U39935 ( .A1(\pe4/aot [14]), .A2(n35207), .ZN(n34736) );
  XOR2HSV0 U39936 ( .A1(n34737), .A2(n34736), .Z(n34742) );
  NAND2HSV0 U39937 ( .A1(n34873), .A2(n33533), .ZN(n34740) );
  NAND2HSV0 U39938 ( .A1(n47718), .A2(n34738), .ZN(n34739) );
  XOR2HSV0 U39939 ( .A1(n34740), .A2(n34739), .Z(n34741) );
  XOR2HSV0 U39940 ( .A1(n34742), .A2(n34741), .Z(n34751) );
  NAND2HSV0 U39941 ( .A1(n57384), .A2(n57906), .ZN(n34745) );
  NAND2HSV0 U39942 ( .A1(n34743), .A2(n33969), .ZN(n34744) );
  XOR2HSV0 U39943 ( .A1(n34745), .A2(n34744), .Z(n34749) );
  NAND2HSV0 U39944 ( .A1(n35191), .A2(n48069), .ZN(n34747) );
  NAND2HSV0 U39945 ( .A1(n57852), .A2(n33713), .ZN(n34746) );
  XOR2HSV0 U39946 ( .A1(n34747), .A2(n34746), .Z(n34748) );
  XOR2HSV0 U39947 ( .A1(n34749), .A2(n34748), .Z(n34750) );
  XOR2HSV0 U39948 ( .A1(n34751), .A2(n34750), .Z(n34767) );
  NAND2HSV0 U39949 ( .A1(n33965), .A2(n57929), .ZN(n34753) );
  NAND2HSV0 U39950 ( .A1(n47709), .A2(\pe4/bq[11] ), .ZN(n34752) );
  XOR2HSV0 U39951 ( .A1(n34753), .A2(n34752), .Z(n34757) );
  NAND2HSV0 U39952 ( .A1(n35491), .A2(n58077), .ZN(n34755) );
  NAND2HSV0 U39953 ( .A1(n47658), .A2(n34879), .ZN(n34754) );
  XOR2HSV0 U39954 ( .A1(n34755), .A2(n34754), .Z(n34756) );
  XOR2HSV0 U39955 ( .A1(n34757), .A2(n34756), .Z(n34765) );
  NAND2HSV0 U39956 ( .A1(\pe4/aot [11]), .A2(n57134), .ZN(n34759) );
  NAND2HSV0 U39957 ( .A1(n59951), .A2(\pe4/bq[20] ), .ZN(n34758) );
  XOR2HSV0 U39958 ( .A1(n34759), .A2(n34758), .Z(n34763) );
  INHSV2 U39959 ( .I(\pe4/aot [9]), .ZN(n57707) );
  NAND2HSV0 U39960 ( .A1(\pe4/aot [9]), .A2(n34888), .ZN(n34761) );
  NAND2HSV0 U39961 ( .A1(\pe4/got [9]), .A2(n47679), .ZN(n34760) );
  XOR2HSV0 U39962 ( .A1(n34761), .A2(n34760), .Z(n34762) );
  XOR2HSV0 U39963 ( .A1(n34763), .A2(n34762), .Z(n34764) );
  XOR2HSV0 U39964 ( .A1(n34765), .A2(n34764), .Z(n34766) );
  XOR2HSV0 U39965 ( .A1(n34767), .A2(n34766), .Z(n34785) );
  NAND2HSV0 U39966 ( .A1(n59952), .A2(n57459), .ZN(n34769) );
  CLKNAND2HSV0 U39967 ( .A1(n47692), .A2(n35220), .ZN(n34768) );
  XOR2HSV0 U39968 ( .A1(n34769), .A2(n34768), .Z(n34773) );
  NAND2HSV0 U39969 ( .A1(n34770), .A2(\pe4/pvq [24]), .ZN(n34771) );
  XNOR2HSV1 U39970 ( .A1(n34771), .A2(\pe4/phq [24]), .ZN(n34772) );
  XNOR2HSV1 U39971 ( .A1(n34773), .A2(n34772), .ZN(n34775) );
  NAND2HSV0 U39972 ( .A1(n33726), .A2(n49943), .ZN(n34919) );
  NOR2HSV0 U39973 ( .A1(n47661), .A2(n53219), .ZN(n57112) );
  XNOR2HSV1 U39974 ( .A1(n34775), .A2(n34774), .ZN(n34783) );
  CLKNAND2HSV0 U39975 ( .A1(n35326), .A2(n57139), .ZN(n34777) );
  CLKNAND2HSV0 U39976 ( .A1(n34387), .A2(n58116), .ZN(n34776) );
  XOR2HSV0 U39977 ( .A1(n34777), .A2(n34776), .Z(n34781) );
  NAND2HSV0 U39978 ( .A1(n34874), .A2(\pe4/bq[22] ), .ZN(n34778) );
  XOR2HSV0 U39979 ( .A1(n34779), .A2(n34778), .Z(n34780) );
  XOR2HSV0 U39980 ( .A1(n34781), .A2(n34780), .Z(n34782) );
  XNOR2HSV1 U39981 ( .A1(n34783), .A2(n34782), .ZN(n34784) );
  XNOR2HSV1 U39982 ( .A1(n34785), .A2(n34784), .ZN(n34786) );
  XOR3HSV2 U39983 ( .A1(n34788), .A2(n34787), .A3(n34786), .Z(n34789) );
  XNOR2HSV1 U39984 ( .A1(n34790), .A2(n34789), .ZN(n34792) );
  NAND2HSV0 U39985 ( .A1(n34396), .A2(n59630), .ZN(n34791) );
  XNOR2HSV1 U39986 ( .A1(n34792), .A2(n34791), .ZN(n34793) );
  XNOR2HSV1 U39987 ( .A1(n34794), .A2(n34793), .ZN(n34796) );
  CLKNAND2HSV1 U39988 ( .A1(n35555), .A2(n59604), .ZN(n34795) );
  XNOR2HSV1 U39989 ( .A1(n34796), .A2(n34795), .ZN(n34799) );
  NAND2HSV0 U39990 ( .A1(n35401), .A2(n34797), .ZN(n34798) );
  XOR2HSV0 U39991 ( .A1(n34799), .A2(n34798), .Z(n34800) );
  XNOR2HSV1 U39992 ( .A1(n34801), .A2(n34800), .ZN(n34803) );
  NAND2HSV0 U39993 ( .A1(n57414), .A2(n35321), .ZN(n34802) );
  XNOR2HSV1 U39994 ( .A1(n34803), .A2(n34802), .ZN(n34804) );
  XNOR2HSV1 U39995 ( .A1(n34805), .A2(n34804), .ZN(n34807) );
  CLKNAND2HSV1 U39996 ( .A1(n57188), .A2(n59601), .ZN(n34806) );
  XOR3HSV2 U39997 ( .A1(n34808), .A2(n34807), .A3(n34806), .Z(n34809) );
  XNOR2HSV1 U39998 ( .A1(n34810), .A2(n34809), .ZN(n34812) );
  NAND2HSV0 U39999 ( .A1(n57985), .A2(n59603), .ZN(n34811) );
  XNOR2HSV1 U40000 ( .A1(n34812), .A2(n34811), .ZN(n34813) );
  XOR2HSV0 U40001 ( .A1(n34816), .A2(n34815), .Z(n34817) );
  XOR2HSV2 U40002 ( .A1(n34818), .A2(n34817), .Z(n34821) );
  NAND2HSV2 U40003 ( .A1(n34819), .A2(n34019), .ZN(n34820) );
  XNOR2HSV4 U40004 ( .A1(n34821), .A2(n34820), .ZN(n34825) );
  NOR2HSV0 U40005 ( .A1(n34970), .A2(n34851), .ZN(n34822) );
  NAND3HSV2 U40006 ( .A1(n34969), .A2(n29709), .A3(n34823), .ZN(n34824) );
  XNOR2HSV4 U40007 ( .A1(n34825), .A2(n34824), .ZN(n35275) );
  XNOR2HSV4 U40008 ( .A1(n34826), .A2(n35275), .ZN(n34994) );
  INHSV4 U40009 ( .I(n34999), .ZN(n34833) );
  INHSV4 U40010 ( .I(n34833), .ZN(n52826) );
  INHSV4 U40011 ( .I(n34827), .ZN(n34828) );
  NAND2HSV4 U40012 ( .A1(n52826), .A2(n34828), .ZN(n35024) );
  CLKNAND2HSV1 U40013 ( .A1(n34829), .A2(n33192), .ZN(n34830) );
  NAND2HSV4 U40014 ( .A1(n34833), .A2(n34832), .ZN(n35022) );
  NOR2HSV0 U40015 ( .A1(n34834), .A2(\pe4/ti_7t [24]), .ZN(n35278) );
  NOR2HSV2 U40016 ( .A1(n35278), .A2(n46581), .ZN(n35028) );
  CLKNHSV0 U40017 ( .I(n35028), .ZN(n34835) );
  CLKNHSV2 U40018 ( .I(n34835), .ZN(n34836) );
  NAND3HSV4 U40019 ( .A1(n35024), .A2(n35022), .A3(n34836), .ZN(n34982) );
  INHSV2 U40020 ( .I(n60045), .ZN(n34839) );
  NAND2HSV2 U40021 ( .A1(n34837), .A2(n34843), .ZN(n34838) );
  NAND2HSV4 U40022 ( .A1(n34844), .A2(n34842), .ZN(n47943) );
  NOR2HSV2 U40023 ( .A1(n34991), .A2(n57204), .ZN(n34840) );
  CLKNAND2HSV1 U40024 ( .A1(n34842), .A2(n34419), .ZN(n34846) );
  NOR2HSV2 U40025 ( .A1(n34846), .A2(n34845), .ZN(n34847) );
  NAND2HSV2 U40026 ( .A1(n34850), .A2(n34849), .ZN(n34852) );
  NOR2HSV2 U40027 ( .A1(n34857), .A2(n34108), .ZN(n34859) );
  NAND2HSV2 U40028 ( .A1(n34859), .A2(n34858), .ZN(n34862) );
  CLKNAND2HSV0 U40029 ( .A1(n34860), .A2(n59955), .ZN(n34861) );
  NAND3HSV3 U40030 ( .A1(n34863), .A2(n34862), .A3(n34861), .ZN(n34978) );
  NAND2HSV2 U40031 ( .A1(n47835), .A2(n59350), .ZN(n34965) );
  CLKNAND2HSV1 U40032 ( .A1(n35320), .A2(n34864), .ZN(n34963) );
  NAND2HSV0 U40033 ( .A1(n34865), .A2(n59603), .ZN(n34959) );
  CLKNAND2HSV1 U40034 ( .A1(n34866), .A2(n59601), .ZN(n34954) );
  CLKNAND2HSV0 U40035 ( .A1(n35489), .A2(\pe4/got [20]), .ZN(n34952) );
  CLKNAND2HSV0 U40036 ( .A1(n34459), .A2(n59602), .ZN(n34947) );
  BUFHSV2 U40037 ( .I(n34867), .Z(n57458) );
  NAND2HSV2 U40038 ( .A1(n57458), .A2(n35167), .ZN(n34943) );
  CLKNAND2HSV1 U40039 ( .A1(n57404), .A2(n35243), .ZN(n34936) );
  NAND2HSV0 U40040 ( .A1(n34868), .A2(n59631), .ZN(n34932) );
  CLKNAND2HSV1 U40041 ( .A1(n57251), .A2(n59663), .ZN(n34870) );
  INHSV2 U40042 ( .I(n59628), .ZN(n57180) );
  NAND2HSV0 U40043 ( .A1(n35227), .A2(n57180), .ZN(n34869) );
  XNOR2HSV1 U40044 ( .A1(n34870), .A2(n34869), .ZN(n34930) );
  NAND2HSV0 U40045 ( .A1(n35340), .A2(n58153), .ZN(n34929) );
  NAND2HSV0 U40046 ( .A1(n47709), .A2(n58116), .ZN(n34872) );
  NAND2HSV0 U40047 ( .A1(\pe4/aot [11]), .A2(n33313), .ZN(n34871) );
  XOR2HSV0 U40048 ( .A1(n34872), .A2(n34871), .Z(n34878) );
  NAND2HSV0 U40049 ( .A1(n34873), .A2(n35194), .ZN(n34876) );
  NAND2HSV0 U40050 ( .A1(n34874), .A2(n57505), .ZN(n34875) );
  XOR2HSV0 U40051 ( .A1(n34876), .A2(n34875), .Z(n34877) );
  XOR2HSV0 U40052 ( .A1(n34878), .A2(n34877), .Z(n34887) );
  NOR2HSV0 U40053 ( .A1(n44338), .A2(n57260), .ZN(n34881) );
  NAND2HSV0 U40054 ( .A1(n59838), .A2(n34879), .ZN(n34880) );
  XOR2HSV0 U40055 ( .A1(n34881), .A2(n34880), .Z(n34885) );
  NAND2HSV0 U40056 ( .A1(n59839), .A2(\pe4/bq[20] ), .ZN(n34883) );
  NAND2HSV0 U40057 ( .A1(n34387), .A2(n35220), .ZN(n34882) );
  XOR2HSV0 U40058 ( .A1(n34883), .A2(n34882), .Z(n34884) );
  XOR2HSV0 U40059 ( .A1(n34885), .A2(n34884), .Z(n34886) );
  XOR2HSV0 U40060 ( .A1(n34887), .A2(n34886), .Z(n34905) );
  INHSV1 U40061 ( .I(n57775), .ZN(n50251) );
  NAND2HSV0 U40062 ( .A1(n50251), .A2(n34888), .ZN(n34890) );
  NAND2HSV0 U40063 ( .A1(\pe4/got [8]), .A2(n35370), .ZN(n34889) );
  XOR2HSV0 U40064 ( .A1(n34890), .A2(n34889), .Z(n34894) );
  NAND2HSV0 U40065 ( .A1(\pe4/aot [22]), .A2(n57906), .ZN(n34892) );
  NAND2HSV0 U40066 ( .A1(n47718), .A2(n57134), .ZN(n34891) );
  XOR2HSV0 U40067 ( .A1(n34892), .A2(n34891), .Z(n34893) );
  XOR2HSV0 U40068 ( .A1(n34894), .A2(n34893), .Z(n34903) );
  NOR2HSV0 U40069 ( .A1(n33250), .A2(n53219), .ZN(n34896) );
  CLKNAND2HSV0 U40070 ( .A1(\pe4/aot [21]), .A2(n57929), .ZN(n34895) );
  XOR2HSV0 U40071 ( .A1(n34896), .A2(n34895), .Z(n34901) );
  NAND2HSV0 U40072 ( .A1(n57138), .A2(\pe4/bq[11] ), .ZN(n34899) );
  INHSV2 U40073 ( .I(n34897), .ZN(n57504) );
  NAND2HSV0 U40074 ( .A1(n57504), .A2(n33611), .ZN(n34898) );
  XOR2HSV0 U40075 ( .A1(n34899), .A2(n34898), .Z(n34900) );
  XOR2HSV0 U40076 ( .A1(n34901), .A2(n34900), .Z(n34902) );
  XOR2HSV0 U40077 ( .A1(n34903), .A2(n34902), .Z(n34904) );
  XOR2HSV0 U40078 ( .A1(n34905), .A2(n34904), .Z(n34927) );
  NOR2HSV0 U40079 ( .A1(n35175), .A2(n50248), .ZN(n34907) );
  CLKNAND2HSV0 U40080 ( .A1(n47692), .A2(n35184), .ZN(n34906) );
  XOR2HSV0 U40081 ( .A1(n34907), .A2(n34906), .Z(n34910) );
  CLKNAND2HSV1 U40082 ( .A1(n53218), .A2(\pe4/pvq [25]), .ZN(n34908) );
  XOR2HSV0 U40083 ( .A1(n34908), .A2(\pe4/phq [25]), .Z(n34909) );
  XOR2HSV0 U40084 ( .A1(n34910), .A2(n34909), .Z(n34918) );
  NAND2HSV0 U40085 ( .A1(\pe4/aot [14]), .A2(n33712), .ZN(n35168) );
  OAI22HSV0 U40086 ( .A1(n34276), .A2(n57030), .B1(n34470), .B2(n33350), .ZN(
        n34911) );
  OAI21HSV1 U40087 ( .A1(n35168), .A2(n34912), .B(n34911), .ZN(n34916) );
  NAND2HSV0 U40088 ( .A1(n35347), .A2(n57850), .ZN(n57849) );
  OAI22HSV0 U40089 ( .A1(n48070), .A2(n57918), .B1(n46143), .B2(n47809), .ZN(
        n34913) );
  OAI21HSV0 U40090 ( .A1(n34914), .A2(n57849), .B(n34913), .ZN(n34915) );
  XOR2HSV0 U40091 ( .A1(n34916), .A2(n34915), .Z(n34917) );
  XOR2HSV0 U40092 ( .A1(n34918), .A2(n34917), .Z(n34925) );
  XOR2HSV0 U40093 ( .A1(n34920), .A2(n34919), .Z(n34923) );
  NAND2HSV0 U40094 ( .A1(n34044), .A2(n57218), .ZN(n50131) );
  XOR2HSV0 U40095 ( .A1(n34921), .A2(n50131), .Z(n34922) );
  XOR2HSV0 U40096 ( .A1(n34923), .A2(n34922), .Z(n34924) );
  XNOR2HSV1 U40097 ( .A1(n34925), .A2(n34924), .ZN(n34926) );
  XNOR2HSV1 U40098 ( .A1(n34927), .A2(n34926), .ZN(n34928) );
  XOR3HSV2 U40099 ( .A1(n34930), .A2(n34929), .A3(n34928), .Z(n34931) );
  XNOR2HSV1 U40100 ( .A1(n34932), .A2(n34931), .ZN(n34934) );
  CLKNAND2HSV1 U40101 ( .A1(n33498), .A2(n59629), .ZN(n34933) );
  XNOR2HSV1 U40102 ( .A1(n34934), .A2(n34933), .ZN(n34935) );
  XNOR2HSV1 U40103 ( .A1(n34936), .A2(n34935), .ZN(n34939) );
  CLKNAND2HSV0 U40104 ( .A1(n35555), .A2(n34937), .ZN(n34938) );
  XNOR2HSV1 U40105 ( .A1(n34939), .A2(n34938), .ZN(n34941) );
  NAND2HSV0 U40106 ( .A1(n35401), .A2(n57189), .ZN(n34940) );
  XOR2HSV0 U40107 ( .A1(n34941), .A2(n34940), .Z(n34942) );
  XNOR2HSV1 U40108 ( .A1(n34943), .A2(n34942), .ZN(n34945) );
  NAND2HSV0 U40109 ( .A1(n57414), .A2(n57834), .ZN(n34944) );
  XNOR2HSV1 U40110 ( .A1(n34945), .A2(n34944), .ZN(n34946) );
  XNOR2HSV1 U40111 ( .A1(n34947), .A2(n34946), .ZN(n34951) );
  CLKNAND2HSV0 U40112 ( .A1(n25243), .A2(n34948), .ZN(n34950) );
  XOR3HSV2 U40113 ( .A1(n34952), .A2(n34951), .A3(n34950), .Z(n34953) );
  NAND2HSV0 U40114 ( .A1(n57985), .A2(n57309), .ZN(n34956) );
  XNOR2HSV1 U40115 ( .A1(n34957), .A2(n34956), .ZN(n34958) );
  XNOR2HSV1 U40116 ( .A1(n34959), .A2(n34958), .ZN(n34961) );
  CLKNAND2HSV1 U40117 ( .A1(n58060), .A2(n57190), .ZN(n34960) );
  XNOR2HSV1 U40118 ( .A1(n34961), .A2(n34960), .ZN(n34962) );
  XNOR2HSV1 U40119 ( .A1(n34963), .A2(n34962), .ZN(n34964) );
  XNOR2HSV1 U40120 ( .A1(n34965), .A2(n34964), .ZN(n34976) );
  NAND2HSV2 U40121 ( .A1(n34967), .A2(n34966), .ZN(n34975) );
  NOR2HSV0 U40122 ( .A1(n34970), .A2(n57453), .ZN(n34971) );
  CLKNAND2HSV1 U40123 ( .A1(n25875), .A2(n34971), .ZN(n34972) );
  NOR2HSV4 U40124 ( .A1(n34973), .A2(n34972), .ZN(n34974) );
  XOR3HSV2 U40125 ( .A1(n34976), .A2(n34975), .A3(n34974), .Z(n34977) );
  XNOR2HSV4 U40126 ( .A1(n34978), .A2(n34977), .ZN(n35025) );
  INHSV4 U40127 ( .I(n35026), .ZN(n34980) );
  CLKNHSV2 U40128 ( .I(n35025), .ZN(n34979) );
  CLKNAND2HSV3 U40129 ( .A1(n34980), .A2(n34979), .ZN(n34981) );
  CLKNAND2HSV1 U40130 ( .A1(n34984), .A2(n34983), .ZN(n34985) );
  NOR2HSV4 U40131 ( .A1(n34985), .A2(n34986), .ZN(n34988) );
  NAND2HSV4 U40132 ( .A1(n34988), .A2(n34987), .ZN(n34996) );
  CLKNHSV0 U40133 ( .I(n34989), .ZN(n34990) );
  NAND2HSV2 U40134 ( .A1(n47943), .A2(n34990), .ZN(n34995) );
  CLKNHSV2 U40135 ( .I(n34991), .ZN(n34992) );
  CLKNAND2HSV0 U40136 ( .A1(n34992), .A2(n33676), .ZN(n34993) );
  CLKNHSV2 U40137 ( .I(n35029), .ZN(n35437) );
  CLKNAND2HSV0 U40138 ( .A1(n34995), .A2(n33779), .ZN(n34998) );
  CLKNHSV0 U40139 ( .I(n34996), .ZN(n34997) );
  NOR2HSV2 U40140 ( .A1(n34998), .A2(n34997), .ZN(n35001) );
  INHSV2 U40141 ( .I(n34999), .ZN(n35027) );
  INHSV2 U40142 ( .I(n35027), .ZN(n35000) );
  AOI22HSV2 U40143 ( .A1(\pe4/ti_7t [24]), .A2(n35295), .B1(n35001), .B2(
        n35000), .ZN(n35002) );
  INHSV2 U40144 ( .I(n35014), .ZN(n46582) );
  CLKNHSV0 U40145 ( .I(n33097), .ZN(n35482) );
  OAI21HSV2 U40146 ( .A1(\pe4/ti_7t [26]), .A2(n35011), .B(n33696), .ZN(n35012) );
  NOR2HSV1 U40147 ( .A1(n35016), .A2(n35007), .ZN(n35015) );
  INHSV2 U40148 ( .I(n35016), .ZN(n35287) );
  NOR2HSV2 U40149 ( .A1(n33696), .A2(n47777), .ZN(n35017) );
  NAND2HSV2 U40150 ( .A1(n35287), .A2(n35017), .ZN(n35018) );
  NAND2HSV2 U40151 ( .A1(n35020), .A2(n35463), .ZN(n35457) );
  AND2HSV2 U40152 ( .A1(n35028), .A2(n35021), .Z(n35023) );
  NAND2HSV2 U40153 ( .A1(n35482), .A2(\pe4/ti_7t [25]), .ZN(n35449) );
  INHSV2 U40154 ( .I(n35143), .ZN(n47846) );
  NOR2HSV4 U40155 ( .A1(n35027), .A2(n35483), .ZN(n35440) );
  INHSV2 U40156 ( .I(n35451), .ZN(n35030) );
  CLKNAND2HSV2 U40157 ( .A1(n35446), .A2(n35030), .ZN(n35031) );
  NAND2HSV4 U40158 ( .A1(n29635), .A2(n35031), .ZN(n47865) );
  CLKBUFHSV4 U40159 ( .I(n47865), .Z(n49921) );
  CLKNAND2HSV3 U40160 ( .A1(n47865), .A2(n35032), .ZN(n35150) );
  CLKNAND2HSV1 U40161 ( .A1(n59950), .A2(n33707), .ZN(n35148) );
  CLKNHSV0 U40162 ( .I(n34966), .ZN(n35034) );
  NOR2HSV1 U40163 ( .A1(n50301), .A2(n35034), .ZN(n35147) );
  INHSV2 U40164 ( .I(n35428), .ZN(n35583) );
  CLKNAND2HSV0 U40165 ( .A1(n50065), .A2(n59603), .ZN(n35138) );
  CLKNAND2HSV1 U40166 ( .A1(n59833), .A2(n59664), .ZN(n35123) );
  NAND2HSV0 U40167 ( .A1(n57458), .A2(n47657), .ZN(n35119) );
  BUFHSV2 U40168 ( .I(n35036), .Z(n59667) );
  CLKNAND2HSV0 U40169 ( .A1(n59667), .A2(n59663), .ZN(n35113) );
  NAND2HSV0 U40170 ( .A1(n47733), .A2(n57177), .ZN(n35109) );
  NAND2HSV0 U40171 ( .A1(n57251), .A2(n58184), .ZN(n35051) );
  CLKNAND2HSV1 U40172 ( .A1(n35347), .A2(n57505), .ZN(n49971) );
  NAND2HSV0 U40173 ( .A1(n59343), .A2(n50007), .ZN(n57126) );
  XOR2HSV0 U40174 ( .A1(n49971), .A2(n57126), .Z(n35039) );
  NAND2HSV0 U40175 ( .A1(n57234), .A2(n57785), .ZN(n57349) );
  NAND2HSV0 U40176 ( .A1(\pe4/aot [20]), .A2(\pe4/bq[16] ), .ZN(n35037) );
  XOR2HSV0 U40177 ( .A1(n57349), .A2(n35037), .Z(n35038) );
  XOR2HSV0 U40178 ( .A1(n35039), .A2(n35038), .Z(n35049) );
  NAND2HSV0 U40179 ( .A1(n57218), .A2(n57089), .ZN(n35041) );
  NAND2HSV0 U40180 ( .A1(\pe4/aot [14]), .A2(n34044), .ZN(n35040) );
  XOR2HSV0 U40181 ( .A1(n35041), .A2(n35040), .Z(n35047) );
  NOR2HSV0 U40182 ( .A1(n35175), .A2(n48022), .ZN(n35045) );
  NAND2HSV0 U40183 ( .A1(n58198), .A2(n57377), .ZN(n35044) );
  XOR2HSV0 U40184 ( .A1(n35045), .A2(n35044), .Z(n35046) );
  XOR2HSV0 U40185 ( .A1(n35047), .A2(n35046), .Z(n35048) );
  XOR2HSV0 U40186 ( .A1(n35049), .A2(n35048), .Z(n35050) );
  XOR2HSV0 U40187 ( .A1(n35051), .A2(n35050), .Z(n35107) );
  NOR2HSV0 U40188 ( .A1(n35501), .A2(n50064), .ZN(n35106) );
  NAND2HSV0 U40189 ( .A1(n47658), .A2(\pe4/bq[11] ), .ZN(n50355) );
  NAND2HSV0 U40190 ( .A1(\pe4/aot [25]), .A2(\pe4/bq[10] ), .ZN(n35492) );
  NOR2HSV0 U40191 ( .A1(n50355), .A2(n35492), .ZN(n35053) );
  AOI22HSV0 U40192 ( .A1(n57499), .A2(\pe4/bq[11] ), .B1(n59661), .B2(n58116), 
        .ZN(n35052) );
  NOR2HSV2 U40193 ( .A1(n35053), .A2(n35052), .ZN(n35065) );
  NAND2HSV0 U40194 ( .A1(n47659), .A2(\pe4/pvq [29]), .ZN(n35054) );
  XOR2HSV0 U40195 ( .A1(n35054), .A2(\pe4/phq [29]), .Z(n35064) );
  NOR2HSV0 U40196 ( .A1(n46143), .A2(n53219), .ZN(n35057) );
  NOR2HSV0 U40197 ( .A1(n50134), .A2(n57387), .ZN(n35056) );
  CLKNAND2HSV0 U40198 ( .A1(n33965), .A2(n34480), .ZN(n35494) );
  NOR2HSV0 U40199 ( .A1(n46143), .A2(n57387), .ZN(n35331) );
  CLKNHSV0 U40200 ( .I(n35331), .ZN(n35055) );
  OAI22HSV2 U40201 ( .A1(n35057), .A2(n35056), .B1(n35494), .B2(n35055), .ZN(
        n35062) );
  NAND2HSV0 U40202 ( .A1(n47692), .A2(\pe4/bq[5] ), .ZN(n35333) );
  NAND2HSV0 U40203 ( .A1(n59523), .A2(n57595), .ZN(n35495) );
  NOR2HSV0 U40204 ( .A1(n35333), .A2(n35495), .ZN(n35060) );
  AOI22HSV0 U40205 ( .A1(n35377), .A2(n57837), .B1(n47692), .B2(n57498), .ZN(
        n35059) );
  NOR2HSV1 U40206 ( .A1(n35060), .A2(n35059), .ZN(n35061) );
  XOR2HSV0 U40207 ( .A1(n35062), .A2(n35061), .Z(n35063) );
  XOR3HSV2 U40208 ( .A1(n35065), .A2(n35064), .A3(n35063), .Z(n35104) );
  CLKNHSV1 U40209 ( .I(n33350), .ZN(n57460) );
  CLKNAND2HSV0 U40210 ( .A1(n47718), .A2(n57460), .ZN(n35067) );
  CLKNHSV0 U40211 ( .I(n44338), .ZN(n57463) );
  NAND2HSV0 U40212 ( .A1(n57463), .A2(n57476), .ZN(n35066) );
  XOR2HSV0 U40213 ( .A1(n35067), .A2(n35066), .Z(n35072) );
  INHSV1 U40214 ( .I(n49929), .ZN(n58223) );
  NAND2HSV0 U40215 ( .A1(n58223), .A2(n34738), .ZN(n35070) );
  NAND2HSV0 U40216 ( .A1(n57338), .A2(n34021), .ZN(n35069) );
  XOR2HSV0 U40217 ( .A1(n35070), .A2(n35069), .Z(n35071) );
  XOR2HSV0 U40218 ( .A1(n35072), .A2(n35071), .Z(n35081) );
  BUFHSV2 U40219 ( .I(\pe4/bq[9] ), .Z(n57135) );
  NAND2HSV0 U40220 ( .A1(n57510), .A2(n57135), .ZN(n35074) );
  NAND2HSV0 U40221 ( .A1(n57138), .A2(n58003), .ZN(n35073) );
  XOR2HSV0 U40222 ( .A1(n35074), .A2(n35073), .Z(n35079) );
  INHSV2 U40223 ( .I(n57011), .ZN(n58307) );
  BUFHSV2 U40224 ( .I(n34888), .Z(n57098) );
  CLKNAND2HSV0 U40225 ( .A1(n58307), .A2(n57098), .ZN(n35077) );
  NAND2HSV0 U40226 ( .A1(n59683), .A2(n57691), .ZN(n35076) );
  XOR2HSV0 U40227 ( .A1(n35077), .A2(n35076), .Z(n35078) );
  XOR2HSV0 U40228 ( .A1(n35079), .A2(n35078), .Z(n35080) );
  XOR2HSV0 U40229 ( .A1(n35081), .A2(n35080), .Z(n35103) );
  NAND2HSV0 U40230 ( .A1(n57210), .A2(n58130), .ZN(n35083) );
  NAND2HSV0 U40231 ( .A1(n59951), .A2(n58084), .ZN(n35082) );
  XOR2HSV0 U40232 ( .A1(n35083), .A2(n35082), .Z(n35088) );
  NAND2HSV0 U40233 ( .A1(n57504), .A2(n34598), .ZN(n35086) );
  INHSV2 U40234 ( .I(n50091), .ZN(n58206) );
  NAND2HSV0 U40235 ( .A1(n58206), .A2(n47679), .ZN(n35085) );
  XOR2HSV0 U40236 ( .A1(n35086), .A2(n35085), .Z(n35087) );
  XOR2HSV0 U40237 ( .A1(n35088), .A2(n35087), .Z(n35098) );
  CLKNAND2HSV0 U40238 ( .A1(n57727), .A2(\pe4/bq[12] ), .ZN(n35090) );
  NAND2HSV0 U40239 ( .A1(n50215), .A2(n57926), .ZN(n35089) );
  XOR2HSV0 U40240 ( .A1(n35090), .A2(n35089), .Z(n35096) );
  INHSV2 U40241 ( .I(n50351), .ZN(n57851) );
  NAND2HSV0 U40242 ( .A1(n35091), .A2(n57851), .ZN(n35094) );
  INHSV2 U40243 ( .I(n57775), .ZN(n59668) );
  NAND2HSV0 U40244 ( .A1(n59668), .A2(n35194), .ZN(n35093) );
  XOR2HSV0 U40245 ( .A1(n35094), .A2(n35093), .Z(n35095) );
  XOR2HSV0 U40246 ( .A1(n35096), .A2(n35095), .Z(n35097) );
  XOR2HSV0 U40247 ( .A1(n35098), .A2(n35097), .Z(n35101) );
  NAND2HSV0 U40248 ( .A1(n35227), .A2(\pe4/got [5]), .ZN(n35100) );
  XNOR2HSV1 U40249 ( .A1(n35101), .A2(n35100), .ZN(n35102) );
  XOR3HSV2 U40250 ( .A1(n35104), .A2(n35103), .A3(n35102), .Z(n35105) );
  XOR3HSV2 U40251 ( .A1(n35107), .A2(n35106), .A3(n35105), .Z(n35108) );
  XNOR2HSV1 U40252 ( .A1(n35109), .A2(n35108), .ZN(n35111) );
  NAND2HSV0 U40253 ( .A1(n57526), .A2(n57180), .ZN(n35110) );
  XNOR2HSV1 U40254 ( .A1(n35111), .A2(n35110), .ZN(n35112) );
  XNOR2HSV1 U40255 ( .A1(n35113), .A2(n35112), .ZN(n35115) );
  NAND2HSV0 U40256 ( .A1(n35555), .A2(n58153), .ZN(n35114) );
  XNOR2HSV1 U40257 ( .A1(n35115), .A2(n35114), .ZN(n35117) );
  NAND2HSV0 U40258 ( .A1(n47742), .A2(n35397), .ZN(n35116) );
  XOR2HSV0 U40259 ( .A1(n35117), .A2(n35116), .Z(n35118) );
  XNOR2HSV1 U40260 ( .A1(n35119), .A2(n35118), .ZN(n35121) );
  NAND2HSV0 U40261 ( .A1(n57414), .A2(n35490), .ZN(n35120) );
  XNOR2HSV1 U40262 ( .A1(n35121), .A2(n35120), .ZN(n35122) );
  XNOR2HSV1 U40263 ( .A1(n35123), .A2(n35122), .ZN(n35125) );
  NAND2HSV0 U40264 ( .A1(n35489), .A2(n47656), .ZN(n35124) );
  XOR2HSV0 U40265 ( .A1(n35125), .A2(n35124), .Z(n35127) );
  CLKNHSV0 U40266 ( .I(n48892), .ZN(n50384) );
  NAND2HSV0 U40267 ( .A1(n25243), .A2(n59353), .ZN(n35126) );
  XOR2HSV0 U40268 ( .A1(n35127), .A2(n35126), .Z(n35130) );
  NAND2HSV0 U40269 ( .A1(n44695), .A2(n34042), .ZN(n35129) );
  NAND2HSV0 U40270 ( .A1(n57985), .A2(n50404), .ZN(n35128) );
  XOR3HSV2 U40271 ( .A1(n35130), .A2(n35129), .A3(n35128), .Z(n35133) );
  NAND2HSV2 U40272 ( .A1(n57550), .A2(n57564), .ZN(n35132) );
  INHSV2 U40273 ( .I(n50207), .ZN(n57567) );
  CLKNAND2HSV1 U40274 ( .A1(n57817), .A2(n57567), .ZN(n35131) );
  XNOR3HSV1 U40275 ( .A1(n35133), .A2(n35132), .A3(n35131), .ZN(n35136) );
  CLKNAND2HSV1 U40276 ( .A1(n35577), .A2(n57309), .ZN(n35135) );
  BUFHSV2 U40277 ( .I(n35320), .Z(n50288) );
  CLKNAND2HSV1 U40278 ( .A1(n50288), .A2(n59601), .ZN(n35134) );
  XOR3HSV2 U40279 ( .A1(n35136), .A2(n35135), .A3(n35134), .Z(n35137) );
  XOR2HSV0 U40280 ( .A1(n35138), .A2(n35137), .Z(n35139) );
  BUFHSV2 U40281 ( .I(n47842), .Z(n57560) );
  CLKAND2HSV2 U40282 ( .A1(n59672), .A2(n34672), .Z(n35141) );
  XOR2HSV0 U40283 ( .A1(n35142), .A2(n35141), .Z(n35145) );
  INHSV2 U40284 ( .I(n35143), .ZN(n47770) );
  CLKNAND2HSV1 U40285 ( .A1(n58103), .A2(n59350), .ZN(n35144) );
  XNOR2HSV1 U40286 ( .A1(n35145), .A2(n35144), .ZN(n35146) );
  MUX2NHSV1 U40287 ( .I0(n35148), .I1(n35147), .S(n35146), .ZN(n35149) );
  XNOR2HSV4 U40288 ( .A1(n35150), .A2(n35149), .ZN(n35151) );
  CLKXOR2HSV4 U40289 ( .A1(n35152), .A2(n35151), .Z(n46564) );
  INHSV2 U40290 ( .I(n35157), .ZN(n35158) );
  NAND2HSV4 U40291 ( .A1(n35159), .A2(n35158), .ZN(n35298) );
  AND2HSV2 U40292 ( .A1(n34571), .A2(n47772), .Z(n35162) );
  CLKNAND2HSV1 U40293 ( .A1(n46582), .A2(n35162), .ZN(n35164) );
  NAND2HSV0 U40294 ( .A1(n35162), .A2(n60030), .ZN(n35163) );
  IOA21HSV4 U40295 ( .A1(n35164), .A2(n35163), .B(n35454), .ZN(n35299) );
  INHSV4 U40296 ( .I(n35299), .ZN(n35165) );
  NAND2HSV2 U40297 ( .A1(n59574), .A2(n33805), .ZN(n35273) );
  CLKNAND2HSV0 U40298 ( .A1(n59526), .A2(\pe4/got [22]), .ZN(n35260) );
  NAND2HSV0 U40299 ( .A1(n44695), .A2(n57564), .ZN(n35256) );
  NAND2HSV0 U40300 ( .A1(n35489), .A2(n57834), .ZN(n35254) );
  CLKNAND2HSV0 U40301 ( .A1(n57209), .A2(n35167), .ZN(n35251) );
  NAND2HSV0 U40302 ( .A1(n35322), .A2(n59664), .ZN(n35247) );
  NAND2HSV0 U40303 ( .A1(n57404), .A2(n35397), .ZN(n35240) );
  NAND2HSV0 U40304 ( .A1(n47733), .A2(n59663), .ZN(n35236) );
  NAND2HSV0 U40305 ( .A1(n33173), .A2(n57177), .ZN(n35183) );
  CLKNAND2HSV0 U40306 ( .A1(n50215), .A2(n57929), .ZN(n49986) );
  XOR2HSV0 U40307 ( .A1(n35168), .A2(n49986), .Z(n35172) );
  NAND2HSV0 U40308 ( .A1(n59668), .A2(n34021), .ZN(n35170) );
  NAND2HSV0 U40309 ( .A1(n59632), .A2(n33611), .ZN(n35169) );
  XOR2HSV0 U40310 ( .A1(n35170), .A2(n35169), .Z(n35171) );
  XOR2HSV0 U40311 ( .A1(n35172), .A2(n35171), .Z(n35181) );
  NOR2HSV0 U40312 ( .A1(n50134), .A2(n48024), .ZN(n35174) );
  NAND2HSV0 U40313 ( .A1(n33947), .A2(n57986), .ZN(n35173) );
  XOR2HSV0 U40314 ( .A1(n35174), .A2(n35173), .Z(n35179) );
  CLKNAND2HSV0 U40315 ( .A1(n59839), .A2(n57089), .ZN(n35177) );
  CLKNAND2HSV0 U40316 ( .A1(n57014), .A2(\pe4/bq[21] ), .ZN(n35176) );
  XOR2HSV0 U40317 ( .A1(n35177), .A2(n35176), .Z(n35178) );
  XOR2HSV0 U40318 ( .A1(n35179), .A2(n35178), .Z(n35180) );
  XOR2HSV0 U40319 ( .A1(n35181), .A2(n35180), .Z(n35182) );
  XOR2HSV0 U40320 ( .A1(n35183), .A2(n35182), .Z(n35234) );
  NAND2HSV0 U40321 ( .A1(n59501), .A2(n57180), .ZN(n35233) );
  INHSV3 U40322 ( .I(\pe4/aot [6]), .ZN(n58174) );
  NAND2HSV0 U40323 ( .A1(n59352), .A2(n57098), .ZN(n35186) );
  NAND2HSV0 U40324 ( .A1(n47709), .A2(n35184), .ZN(n35185) );
  XOR2HSV0 U40325 ( .A1(n35186), .A2(n35185), .Z(n35190) );
  NAND2HSV0 U40326 ( .A1(n35326), .A2(\pe4/bq[11] ), .ZN(n35188) );
  NAND2HSV0 U40327 ( .A1(n33726), .A2(n57139), .ZN(n35187) );
  XOR2HSV0 U40328 ( .A1(n35188), .A2(n35187), .Z(n35189) );
  XOR2HSV0 U40329 ( .A1(n35190), .A2(n35189), .Z(n35200) );
  NAND2HSV0 U40330 ( .A1(n35191), .A2(n57691), .ZN(n35193) );
  NAND2HSV0 U40331 ( .A1(n59952), .A2(n34044), .ZN(n35192) );
  XOR2HSV0 U40332 ( .A1(n35193), .A2(n35192), .Z(n35198) );
  NAND2HSV0 U40333 ( .A1(n47718), .A2(n35194), .ZN(n35196) );
  NAND2HSV0 U40334 ( .A1(n59838), .A2(n34480), .ZN(n35195) );
  XOR2HSV0 U40335 ( .A1(n35196), .A2(n35195), .Z(n35197) );
  XOR2HSV0 U40336 ( .A1(n35198), .A2(n35197), .Z(n35199) );
  XOR2HSV0 U40337 ( .A1(n35200), .A2(n35199), .Z(n35211) );
  NAND2HSV0 U40338 ( .A1(n59523), .A2(n35323), .ZN(n35203) );
  CLKNHSV0 U40339 ( .I(n50351), .ZN(n58014) );
  NAND2HSV0 U40340 ( .A1(n35201), .A2(n58014), .ZN(n35202) );
  XOR2HSV0 U40341 ( .A1(n35203), .A2(n35202), .Z(n35206) );
  CLKNAND2HSV0 U40342 ( .A1(n48068), .A2(\pe4/pvq [27]), .ZN(n35204) );
  XNOR2HSV1 U40343 ( .A1(n35204), .A2(\pe4/phq [27]), .ZN(n35205) );
  XNOR2HSV1 U40344 ( .A1(n35206), .A2(n35205), .ZN(n35209) );
  NAND2HSV0 U40345 ( .A1(n57210), .A2(\pe4/bq[10] ), .ZN(n57330) );
  NAND2HSV0 U40346 ( .A1(n59683), .A2(n35207), .ZN(n50360) );
  XOR2HSV0 U40347 ( .A1(n57330), .A2(n50360), .Z(n35208) );
  XNOR2HSV1 U40348 ( .A1(n35209), .A2(n35208), .ZN(n35210) );
  XNOR2HSV1 U40349 ( .A1(n35211), .A2(n35210), .ZN(n35231) );
  NAND2HSV0 U40350 ( .A1(n33716), .A2(n57348), .ZN(n35213) );
  NAND2HSV0 U40351 ( .A1(\pe4/got [6]), .A2(n47679), .ZN(n35212) );
  XOR2HSV0 U40352 ( .A1(n35213), .A2(n35212), .Z(n35217) );
  NAND2HSV0 U40353 ( .A1(\pe4/aot [9]), .A2(n33110), .ZN(n35215) );
  NAND2HSV0 U40354 ( .A1(n59951), .A2(n57926), .ZN(n35214) );
  XOR2HSV0 U40355 ( .A1(n35215), .A2(n35214), .Z(n35216) );
  XOR2HSV0 U40356 ( .A1(n35217), .A2(n35216), .Z(n35226) );
  NOR2HSV0 U40357 ( .A1(n57918), .A2(n50248), .ZN(n35219) );
  NAND2HSV0 U40358 ( .A1(n59343), .A2(n33713), .ZN(n35218) );
  XOR2HSV0 U40359 ( .A1(n35219), .A2(n35218), .Z(n35224) );
  NAND2HSV0 U40360 ( .A1(n57218), .A2(n57785), .ZN(n35222) );
  NAND2HSV0 U40361 ( .A1(n57138), .A2(n35220), .ZN(n35221) );
  XOR2HSV0 U40362 ( .A1(n35222), .A2(n35221), .Z(n35223) );
  XOR2HSV0 U40363 ( .A1(n35224), .A2(n35223), .Z(n35225) );
  XOR2HSV0 U40364 ( .A1(n35226), .A2(n35225), .Z(n35229) );
  NAND2HSV0 U40365 ( .A1(n35227), .A2(n58036), .ZN(n35228) );
  XNOR2HSV1 U40366 ( .A1(n35229), .A2(n35228), .ZN(n35230) );
  XOR2HSV0 U40367 ( .A1(n35231), .A2(n35230), .Z(n35232) );
  XOR3HSV2 U40368 ( .A1(n35234), .A2(n35233), .A3(n35232), .Z(n35235) );
  XOR2HSV0 U40369 ( .A1(n35236), .A2(n35235), .Z(n35238) );
  NAND2HSV0 U40370 ( .A1(n34396), .A2(n58153), .ZN(n35237) );
  XNOR2HSV1 U40371 ( .A1(n35238), .A2(n35237), .ZN(n35239) );
  XNOR2HSV1 U40372 ( .A1(n35240), .A2(n35239), .ZN(n35242) );
  NAND2HSV0 U40373 ( .A1(n35555), .A2(n35400), .ZN(n35241) );
  XNOR2HSV1 U40374 ( .A1(n35242), .A2(n35241), .ZN(n35245) );
  NAND2HSV0 U40375 ( .A1(n47742), .A2(n35243), .ZN(n35244) );
  XOR2HSV0 U40376 ( .A1(n35245), .A2(n35244), .Z(n35246) );
  XNOR2HSV1 U40377 ( .A1(n35247), .A2(n35246), .ZN(n35249) );
  NAND2HSV0 U40378 ( .A1(n57414), .A2(\pe4/got [16]), .ZN(n35248) );
  XNOR2HSV1 U40379 ( .A1(n35249), .A2(n35248), .ZN(n35250) );
  XNOR2HSV1 U40380 ( .A1(n35251), .A2(n35250), .ZN(n35253) );
  CLKNAND2HSV1 U40381 ( .A1(n57188), .A2(n50404), .ZN(n35252) );
  XOR3HSV2 U40382 ( .A1(n35254), .A2(n35253), .A3(n35252), .Z(n35255) );
  XNOR2HSV1 U40383 ( .A1(n35256), .A2(n35255), .ZN(n35258) );
  NAND2HSV0 U40384 ( .A1(n57985), .A2(n57567), .ZN(n35257) );
  XNOR2HSV1 U40385 ( .A1(n35258), .A2(n35257), .ZN(n35259) );
  XNOR2HSV1 U40386 ( .A1(n35260), .A2(n35259), .ZN(n35262) );
  CLKNAND2HSV0 U40387 ( .A1(n49951), .A2(n57309), .ZN(n35261) );
  XNOR2HSV1 U40388 ( .A1(n35262), .A2(n35261), .ZN(n35264) );
  NAND2HSV0 U40389 ( .A1(n35320), .A2(n59603), .ZN(n35263) );
  NAND2HSV2 U40390 ( .A1(n50213), .A2(n34864), .ZN(n35265) );
  XNOR2HSV1 U40391 ( .A1(n35266), .A2(n35265), .ZN(n35268) );
  CLKNAND2HSV1 U40392 ( .A1(n47842), .A2(n59350), .ZN(n35267) );
  NAND2HSV0 U40393 ( .A1(n34966), .A2(n35428), .ZN(n35269) );
  CLKNHSV1 U40394 ( .I(n35269), .ZN(n35270) );
  XOR2HSV0 U40395 ( .A1(n35271), .A2(n35270), .Z(n35272) );
  XOR2HSV2 U40396 ( .A1(n35273), .A2(n35272), .Z(n35282) );
  NAND2HSV2 U40397 ( .A1(n35428), .A2(n35274), .ZN(n35276) );
  XOR2HSV2 U40398 ( .A1(n35276), .A2(n35275), .Z(n35277) );
  XNOR2HSV4 U40399 ( .A1(n35277), .A2(n35434), .ZN(n35280) );
  INHSV2 U40400 ( .I(n35278), .ZN(n35435) );
  CLKNAND2HSV1 U40401 ( .A1(n35435), .A2(n59955), .ZN(n35279) );
  AOI21HSV4 U40402 ( .A1(n35280), .A2(n33848), .B(n35279), .ZN(n35281) );
  XNOR2HSV4 U40403 ( .A1(n35282), .A2(n35281), .ZN(n35293) );
  NOR2HSV2 U40404 ( .A1(n35447), .A2(n57204), .ZN(n35291) );
  CLKNHSV2 U40405 ( .I(n35448), .ZN(n35290) );
  OAI22HSV4 U40406 ( .A1(n35288), .A2(n35287), .B1(n35286), .B2(n35449), .ZN(
        n35289) );
  AOI21HSV4 U40407 ( .A1(n35291), .A2(n35290), .B(n35289), .ZN(n35292) );
  XNOR2HSV4 U40408 ( .A1(n35293), .A2(n35292), .ZN(n35313) );
  INAND2HSV4 U40409 ( .A1(n35294), .B1(n35313), .ZN(n35308) );
  NOR2HSV4 U40410 ( .A1(n35296), .A2(n35295), .ZN(n35297) );
  NAND3HSV4 U40411 ( .A1(n35298), .A2(n35299), .A3(n35297), .ZN(n35301) );
  NAND2HSV2 U40412 ( .A1(n33167), .A2(\pe4/ti_7t [27]), .ZN(n35300) );
  INHSV4 U40413 ( .I(n44690), .ZN(n35304) );
  NAND2HSV4 U40414 ( .A1(n35304), .A2(n52755), .ZN(n46563) );
  XNOR2HSV4 U40415 ( .A1(n46563), .A2(n46564), .ZN(n35481) );
  INHSV3 U40416 ( .I(n35481), .ZN(n35480) );
  NAND2HSV2 U40417 ( .A1(n35307), .A2(n35306), .ZN(n35312) );
  INHSV2 U40418 ( .I(n35308), .ZN(n35309) );
  CLKNAND2HSV3 U40419 ( .A1(n35310), .A2(n35309), .ZN(n35458) );
  INHSV2 U40420 ( .I(n35313), .ZN(n45792) );
  CLKNHSV0 U40421 ( .I(\pe4/ti_7t [27]), .ZN(n35315) );
  AOI21HSV4 U40422 ( .A1(n35316), .A2(n35315), .B(n52696), .ZN(n35459) );
  CLKNAND2HSV1 U40423 ( .A1(n47842), .A2(n34020), .ZN(n35427) );
  NAND2HSV2 U40424 ( .A1(n35318), .A2(n50065), .ZN(n35426) );
  INAND2HSV2 U40425 ( .A1(n35319), .B1(n35577), .ZN(n35424) );
  NAND2HSV0 U40426 ( .A1(n35320), .A2(n57309), .ZN(n35422) );
  BUFHSV2 U40427 ( .I(n59526), .Z(n57984) );
  NAND2HSV2 U40428 ( .A1(n57984), .A2(n57567), .ZN(n35418) );
  NAND2HSV0 U40429 ( .A1(n44695), .A2(n35321), .ZN(n35414) );
  NAND2HSV0 U40430 ( .A1(n35489), .A2(n59353), .ZN(n35412) );
  NAND2HSV0 U40431 ( .A1(n57209), .A2(\pe4/got [16]), .ZN(n35409) );
  NAND2HSV0 U40432 ( .A1(n35322), .A2(n35490), .ZN(n35405) );
  CLKNAND2HSV0 U40433 ( .A1(n59667), .A2(n58153), .ZN(n35396) );
  NAND2HSV0 U40434 ( .A1(n47733), .A2(n57180), .ZN(n35392) );
  NAND2HSV0 U40435 ( .A1(n57251), .A2(n58216), .ZN(n35339) );
  BUFHSV2 U40436 ( .I(\pe4/bq[9] ), .Z(n57798) );
  NAND2HSV0 U40437 ( .A1(n57210), .A2(n57798), .ZN(n35325) );
  NAND2HSV0 U40438 ( .A1(n47709), .A2(n35323), .ZN(n35324) );
  XOR2HSV0 U40439 ( .A1(n35325), .A2(n35324), .Z(n35330) );
  NAND2HSV0 U40440 ( .A1(n35326), .A2(n58116), .ZN(n35328) );
  INHSV1 U40441 ( .I(n57775), .ZN(n58087) );
  NAND2HSV0 U40442 ( .A1(n58087), .A2(n33533), .ZN(n35327) );
  XOR2HSV0 U40443 ( .A1(n35328), .A2(n35327), .Z(n35329) );
  XOR2HSV0 U40444 ( .A1(n35330), .A2(n35329), .Z(n35337) );
  XOR2HSV0 U40445 ( .A1(n35331), .A2(n50355), .Z(n35335) );
  CLKNAND2HSV0 U40446 ( .A1(\pe4/aot [9]), .A2(n35194), .ZN(n35332) );
  XOR2HSV0 U40447 ( .A1(n35333), .A2(n35332), .Z(n35334) );
  XOR2HSV0 U40448 ( .A1(n35335), .A2(n35334), .Z(n35336) );
  XOR2HSV0 U40449 ( .A1(n35337), .A2(n35336), .Z(n35338) );
  XOR2HSV0 U40450 ( .A1(n35339), .A2(n35338), .Z(n35390) );
  NAND2HSV0 U40451 ( .A1(n35340), .A2(n57177), .ZN(n35389) );
  NAND2HSV0 U40452 ( .A1(n59683), .A2(n57460), .ZN(n35342) );
  NAND2HSV0 U40453 ( .A1(n59388), .A2(n34480), .ZN(n35341) );
  XOR2HSV0 U40454 ( .A1(n35342), .A2(n35341), .Z(n35346) );
  NAND2HSV0 U40455 ( .A1(n57138), .A2(n58130), .ZN(n35344) );
  NAND2HSV0 U40456 ( .A1(n59343), .A2(n57691), .ZN(n35343) );
  XOR2HSV0 U40457 ( .A1(n35344), .A2(n35343), .Z(n35345) );
  XOR2HSV0 U40458 ( .A1(n35346), .A2(n35345), .Z(n35355) );
  NAND2HSV0 U40459 ( .A1(n35347), .A2(\pe4/bq[22] ), .ZN(n35349) );
  NAND2HSV0 U40460 ( .A1(n57218), .A2(n57929), .ZN(n35348) );
  XOR2HSV0 U40461 ( .A1(n35349), .A2(n35348), .Z(n35353) );
  NAND2HSV0 U40462 ( .A1(n59951), .A2(\pe4/bq[16] ), .ZN(n35351) );
  NAND2HSV0 U40463 ( .A1(n50215), .A2(n57089), .ZN(n35350) );
  XOR2HSV0 U40464 ( .A1(n35351), .A2(n35350), .Z(n35352) );
  XOR2HSV0 U40465 ( .A1(n35353), .A2(n35352), .Z(n35354) );
  XOR2HSV0 U40466 ( .A1(n35355), .A2(n35354), .Z(n35367) );
  NAND2HSV0 U40467 ( .A1(n57463), .A2(n50007), .ZN(n35357) );
  NAND2HSV0 U40468 ( .A1(\pe4/aot [14]), .A2(n57476), .ZN(n35356) );
  XOR2HSV0 U40469 ( .A1(n35357), .A2(n35356), .Z(n35361) );
  NAND2HSV0 U40470 ( .A1(n57014), .A2(n57785), .ZN(n35359) );
  NAND2HSV0 U40471 ( .A1(\pe4/aot [7]), .A2(n57134), .ZN(n35358) );
  XOR2HSV0 U40472 ( .A1(n35359), .A2(n35358), .Z(n35360) );
  XOR2HSV0 U40473 ( .A1(n35361), .A2(n35360), .Z(n35365) );
  NAND2HSV0 U40474 ( .A1(n59486), .A2(\pe4/pvq [28]), .ZN(n35362) );
  XNOR2HSV1 U40475 ( .A1(n35362), .A2(\pe4/phq [28]), .ZN(n35363) );
  NAND2HSV0 U40476 ( .A1(n59838), .A2(\pe4/bq[12] ), .ZN(n57028) );
  XNOR2HSV1 U40477 ( .A1(n35363), .A2(n57028), .ZN(n35364) );
  XNOR2HSV1 U40478 ( .A1(n35365), .A2(n35364), .ZN(n35366) );
  XNOR2HSV1 U40479 ( .A1(n35367), .A2(n35366), .ZN(n35387) );
  NAND2HSV0 U40480 ( .A1(n47718), .A2(n34598), .ZN(n35369) );
  NAND2HSV0 U40481 ( .A1(n57234), .A2(\pe4/bq[21] ), .ZN(n35368) );
  XOR2HSV0 U40482 ( .A1(n35369), .A2(n35368), .Z(n35374) );
  NAND2HSV0 U40483 ( .A1(n57338), .A2(n34738), .ZN(n35372) );
  NAND2HSV0 U40484 ( .A1(n57677), .A2(n35370), .ZN(n35371) );
  XOR2HSV0 U40485 ( .A1(n35372), .A2(n35371), .Z(n35373) );
  XOR2HSV0 U40486 ( .A1(n35374), .A2(n35373), .Z(n35383) );
  NOR2HSV0 U40487 ( .A1(n49982), .A2(n47809), .ZN(n35376) );
  NAND2HSV0 U40488 ( .A1(n58306), .A2(n57098), .ZN(n35375) );
  XOR2HSV0 U40489 ( .A1(n35376), .A2(n35375), .Z(n35381) );
  NAND2HSV0 U40490 ( .A1(n33965), .A2(n34879), .ZN(n35379) );
  CLKNHSV0 U40491 ( .I(n50351), .ZN(n57784) );
  NAND2HSV0 U40492 ( .A1(n35377), .A2(n57784), .ZN(n35378) );
  XOR2HSV0 U40493 ( .A1(n35379), .A2(n35378), .Z(n35380) );
  XOR2HSV0 U40494 ( .A1(n35381), .A2(n35380), .Z(n35382) );
  XOR2HSV0 U40495 ( .A1(n35383), .A2(n35382), .Z(n35385) );
  NAND2HSV0 U40496 ( .A1(n35227), .A2(n58137), .ZN(n35384) );
  XNOR2HSV1 U40497 ( .A1(n35385), .A2(n35384), .ZN(n35386) );
  XOR2HSV0 U40498 ( .A1(n35387), .A2(n35386), .Z(n35388) );
  XOR3HSV2 U40499 ( .A1(n35390), .A2(n35389), .A3(n35388), .Z(n35391) );
  XOR2HSV0 U40500 ( .A1(n35392), .A2(n35391), .Z(n35394) );
  NAND2HSV0 U40501 ( .A1(n57526), .A2(n59663), .ZN(n35393) );
  XNOR2HSV1 U40502 ( .A1(n35394), .A2(n35393), .ZN(n35395) );
  XNOR2HSV1 U40503 ( .A1(n35396), .A2(n35395), .ZN(n35399) );
  NAND2HSV0 U40504 ( .A1(n35555), .A2(n35397), .ZN(n35398) );
  XNOR2HSV1 U40505 ( .A1(n35399), .A2(n35398), .ZN(n35403) );
  NAND2HSV0 U40506 ( .A1(n35401), .A2(n35400), .ZN(n35402) );
  XOR2HSV0 U40507 ( .A1(n35403), .A2(n35402), .Z(n35404) );
  XNOR2HSV1 U40508 ( .A1(n35405), .A2(n35404), .ZN(n35407) );
  NAND2HSV0 U40509 ( .A1(n57414), .A2(n59664), .ZN(n35406) );
  XNOR2HSV1 U40510 ( .A1(n35407), .A2(n35406), .ZN(n35408) );
  XNOR2HSV1 U40511 ( .A1(n35409), .A2(n35408), .ZN(n35411) );
  CLKNAND2HSV1 U40512 ( .A1(n57188), .A2(n34042), .ZN(n35410) );
  XOR3HSV2 U40513 ( .A1(n35412), .A2(n35411), .A3(n35410), .Z(n35413) );
  XNOR2HSV1 U40514 ( .A1(n35414), .A2(n35413), .ZN(n35416) );
  NAND2HSV0 U40515 ( .A1(n57985), .A2(n59386), .ZN(n35415) );
  XNOR2HSV1 U40516 ( .A1(n35416), .A2(n35415), .ZN(n35417) );
  XNOR2HSV1 U40517 ( .A1(n35418), .A2(n35417), .ZN(n35420) );
  CLKNAND2HSV0 U40518 ( .A1(n49951), .A2(n59601), .ZN(n35419) );
  XNOR2HSV1 U40519 ( .A1(n35420), .A2(n35419), .ZN(n35421) );
  XNOR2HSV1 U40520 ( .A1(n35422), .A2(n35421), .ZN(n35423) );
  XNOR2HSV1 U40521 ( .A1(n35424), .A2(n35423), .ZN(n35425) );
  NAND2HSV0 U40522 ( .A1(n35428), .A2(n59350), .ZN(n35429) );
  XNOR2HSV1 U40523 ( .A1(n35430), .A2(n35429), .ZN(n35433) );
  CLKNAND2HSV2 U40524 ( .A1(n59574), .A2(n57195), .ZN(n35432) );
  INHSV2 U40525 ( .I(n35434), .ZN(n35438) );
  NAND2HSV2 U40526 ( .A1(n35435), .A2(n59956), .ZN(n35436) );
  AOI21HSV2 U40527 ( .A1(n35437), .A2(n35438), .B(n35436), .ZN(n35442) );
  INHSV2 U40528 ( .I(n35438), .ZN(n35439) );
  NAND2HSV2 U40529 ( .A1(n35440), .A2(n35439), .ZN(n35441) );
  NAND2HSV2 U40530 ( .A1(n35442), .A2(n35441), .ZN(n35443) );
  XNOR2HSV4 U40531 ( .A1(n35444), .A2(n35443), .ZN(n35453) );
  INHSV2 U40532 ( .I(n33098), .ZN(n35445) );
  NOR2HSV1 U40533 ( .A1(n35449), .A2(n34416), .ZN(n35450) );
  XOR2HSV4 U40534 ( .A1(n35453), .A2(n35452), .Z(n47928) );
  OAI21HSV4 U40535 ( .A1(n35465), .A2(n35464), .B(n35463), .ZN(n59666) );
  NAND3HSV2 U40536 ( .A1(n59666), .A2(n59345), .A3(n35462), .ZN(n35456) );
  AOI21HSV2 U40537 ( .A1(n47928), .A2(n34718), .B(n34423), .ZN(n35455) );
  INHSV3 U40538 ( .I(n35458), .ZN(n35478) );
  NAND2HSV2 U40539 ( .A1(n35482), .A2(\pe4/ti_7t [28]), .ZN(n35472) );
  AND2HSV2 U40540 ( .A1(n35459), .A2(n35472), .Z(n35460) );
  CLKNAND2HSV2 U40541 ( .A1(n35461), .A2(n35460), .ZN(n35477) );
  INHSV2 U40542 ( .I(n59666), .ZN(n47853) );
  NOR2HSV2 U40543 ( .A1(n35465), .A2(n35464), .ZN(n35468) );
  INHSV4 U40544 ( .I(n47928), .ZN(n35471) );
  NAND2HSV0 U40545 ( .A1(n35472), .A2(n59345), .ZN(n35466) );
  NOR2HSV4 U40546 ( .A1(n35471), .A2(n35466), .ZN(n35467) );
  INOR2HSV1 U40547 ( .A1(n35472), .B1(n59345), .ZN(n35470) );
  CLKNAND2HSV2 U40548 ( .A1(n35474), .A2(n35473), .ZN(n35475) );
  AOI21HSV4 U40549 ( .A1(n29685), .A2(n47853), .B(n35475), .ZN(n35476) );
  OAI21HSV2 U40550 ( .A1(n47930), .A2(n35486), .B(n35485), .ZN(n35479) );
  NAND2HSV2 U40551 ( .A1(n35482), .A2(\pe4/ti_7t [29]), .ZN(n46566) );
  CLKNAND2HSV1 U40552 ( .A1(n46566), .A2(n35483), .ZN(n47774) );
  NAND2HSV2 U40553 ( .A1(n47774), .A2(n47772), .ZN(n35484) );
  NAND2HSV2 U40554 ( .A1(n35304), .A2(n35487), .ZN(n35602) );
  CLKNAND2HSV1 U40555 ( .A1(n50065), .A2(n57309), .ZN(n35582) );
  BUFHSV2 U40556 ( .I(n35489), .Z(n57324) );
  NAND2HSV2 U40557 ( .A1(n57324), .A2(n59664), .ZN(n35568) );
  NAND2HSV2 U40558 ( .A1(n57678), .A2(n35490), .ZN(n35565) );
  CLKNAND2HSV1 U40559 ( .A1(n59667), .A2(n57180), .ZN(n35554) );
  NAND2HSV0 U40560 ( .A1(n47733), .A2(n58102), .ZN(n35550) );
  NAND2HSV0 U40561 ( .A1(n57251), .A2(n57951), .ZN(n35500) );
  NAND2HSV0 U40562 ( .A1(n35491), .A2(n57851), .ZN(n47663) );
  XOR2HSV0 U40563 ( .A1(n35492), .A2(n47663), .Z(n35498) );
  INHSV2 U40564 ( .I(n35493), .ZN(n59486) );
  CLKNAND2HSV1 U40565 ( .A1(n57140), .A2(n49943), .ZN(n57235) );
  CLKNAND2HSV1 U40566 ( .A1(n47692), .A2(\pe4/bq[3] ), .ZN(n57105) );
  XOR3HSV2 U40567 ( .A1(n35498), .A2(n35497), .A3(n35496), .Z(n35499) );
  XOR2HSV0 U40568 ( .A1(n35500), .A2(n35499), .Z(n35548) );
  NOR2HSV0 U40569 ( .A1(n35501), .A2(n50214), .ZN(n35547) );
  NAND2HSV0 U40570 ( .A1(n59683), .A2(\pe4/bq[24] ), .ZN(n35503) );
  NAND2HSV0 U40571 ( .A1(n59343), .A2(\pe4/bq[23] ), .ZN(n35502) );
  XOR2HSV0 U40572 ( .A1(n35503), .A2(n35502), .Z(n35507) );
  INHSV2 U40573 ( .I(\pe4/aot [3]), .ZN(n58194) );
  NAND2HSV0 U40574 ( .A1(\pe4/aot [3]), .A2(n57098), .ZN(n35505) );
  CLKNHSV0 U40575 ( .I(\pe4/got [3]), .ZN(n47725) );
  NAND2HSV0 U40576 ( .A1(\pe4/got [3]), .A2(n47679), .ZN(n35504) );
  XOR2HSV0 U40577 ( .A1(n35505), .A2(n35504), .Z(n35506) );
  XOR2HSV0 U40578 ( .A1(n35507), .A2(n35506), .Z(n35516) );
  NAND2HSV0 U40579 ( .A1(n35508), .A2(n58130), .ZN(n35510) );
  NAND2HSV0 U40580 ( .A1(n47718), .A2(n57691), .ZN(n35509) );
  XOR2HSV0 U40581 ( .A1(n35510), .A2(n35509), .Z(n35514) );
  NAND2HSV0 U40582 ( .A1(n59831), .A2(n34021), .ZN(n35512) );
  CLKNAND2HSV1 U40583 ( .A1(\pe4/aot [14]), .A2(n34636), .ZN(n35511) );
  XOR2HSV0 U40584 ( .A1(n35512), .A2(n35511), .Z(n35513) );
  XOR2HSV0 U40585 ( .A1(n35514), .A2(n35513), .Z(n35515) );
  XOR2HSV0 U40586 ( .A1(n35516), .A2(n35515), .Z(n35532) );
  CLKNAND2HSV0 U40587 ( .A1(n58198), .A2(n35194), .ZN(n35518) );
  NAND2HSV0 U40588 ( .A1(n33867), .A2(n57926), .ZN(n35517) );
  XOR2HSV0 U40589 ( .A1(n35518), .A2(n35517), .Z(n35522) );
  NAND2HSV0 U40590 ( .A1(n57014), .A2(n57089), .ZN(n35520) );
  NAND2HSV0 U40591 ( .A1(n47709), .A2(n58155), .ZN(n35519) );
  XOR2HSV0 U40592 ( .A1(n35520), .A2(n35519), .Z(n35521) );
  XOR2HSV0 U40593 ( .A1(n35522), .A2(n35521), .Z(n35530) );
  NAND2HSV0 U40594 ( .A1(n57338), .A2(n57377), .ZN(n35524) );
  NAND2HSV0 U40595 ( .A1(n33947), .A2(n57135), .ZN(n35523) );
  XOR2HSV0 U40596 ( .A1(n35524), .A2(n35523), .Z(n35528) );
  NOR2HSV0 U40597 ( .A1(n50008), .A2(n57387), .ZN(n35526) );
  NAND2HSV0 U40598 ( .A1(\pe4/aot [20]), .A2(n58084), .ZN(n35525) );
  XOR2HSV0 U40599 ( .A1(n35526), .A2(n35525), .Z(n35527) );
  XNOR2HSV1 U40600 ( .A1(n35528), .A2(n35527), .ZN(n35529) );
  XNOR2HSV1 U40601 ( .A1(n35530), .A2(n35529), .ZN(n35531) );
  XNOR2HSV1 U40602 ( .A1(n35532), .A2(n35531), .ZN(n35545) );
  NAND2HSV0 U40603 ( .A1(n35533), .A2(n58197), .ZN(n35535) );
  NAND2HSV0 U40604 ( .A1(n57727), .A2(\pe4/bq[11] ), .ZN(n35534) );
  XOR2HSV0 U40605 ( .A1(n35535), .A2(n35534), .Z(n35539) );
  NAND2HSV0 U40606 ( .A1(n59668), .A2(n33427), .ZN(n35537) );
  NAND2HSV0 U40607 ( .A1(\pe4/aot [4]), .A2(n34738), .ZN(n35536) );
  XOR2HSV0 U40608 ( .A1(n35537), .A2(n35536), .Z(n35538) );
  XOR2HSV0 U40609 ( .A1(n35539), .A2(n35538), .Z(n35541) );
  CLKNHSV0 U40610 ( .I(n44338), .ZN(n57585) );
  XNOR2HSV1 U40611 ( .A1(n35541), .A2(n35540), .ZN(n35543) );
  NAND2HSV0 U40612 ( .A1(n34127), .A2(n58206), .ZN(n35542) );
  XNOR2HSV1 U40613 ( .A1(n35543), .A2(n35542), .ZN(n35544) );
  XNOR2HSV1 U40614 ( .A1(n35545), .A2(n35544), .ZN(n35546) );
  XOR3HSV2 U40615 ( .A1(n35548), .A2(n35547), .A3(n35546), .Z(n35549) );
  XNOR2HSV1 U40616 ( .A1(n35550), .A2(n35549), .ZN(n35552) );
  NAND2HSV0 U40617 ( .A1(n59662), .A2(n57177), .ZN(n35551) );
  XNOR2HSV1 U40618 ( .A1(n35552), .A2(n35551), .ZN(n35553) );
  XNOR2HSV1 U40619 ( .A1(n35554), .A2(n35553), .ZN(n35557) );
  BUFHSV2 U40620 ( .I(n35555), .Z(n57405) );
  NAND2HSV2 U40621 ( .A1(n57405), .A2(n59663), .ZN(n35556) );
  XNOR2HSV1 U40622 ( .A1(n35557), .A2(n35556), .ZN(n35559) );
  NAND2HSV0 U40623 ( .A1(n57679), .A2(n58153), .ZN(n35558) );
  XOR2HSV0 U40624 ( .A1(n35559), .A2(n35558), .Z(n35563) );
  CLKNAND2HSV0 U40625 ( .A1(n34352), .A2(n50189), .ZN(n35562) );
  CLKNAND2HSV1 U40626 ( .A1(n57183), .A2(n47657), .ZN(n35561) );
  XOR3HSV2 U40627 ( .A1(n35563), .A2(n35562), .A3(n35561), .Z(n35564) );
  XNOR2HSV1 U40628 ( .A1(n35565), .A2(n35564), .ZN(n35567) );
  NAND2HSV2 U40629 ( .A1(n59845), .A2(n47656), .ZN(n35566) );
  XOR3HSV2 U40630 ( .A1(n35568), .A2(n35567), .A3(n35566), .Z(n35573) );
  NAND2HSV2 U40631 ( .A1(n49966), .A2(n59353), .ZN(n35572) );
  NAND2HSV2 U40632 ( .A1(n57547), .A2(\pe4/got [18]), .ZN(n35571) );
  XOR3HSV2 U40633 ( .A1(n35573), .A2(n35572), .A3(n35571), .Z(n35576) );
  NAND2HSV2 U40634 ( .A1(n59526), .A2(n50404), .ZN(n35575) );
  NAND2HSV2 U40635 ( .A1(n57817), .A2(n57564), .ZN(n35574) );
  XOR3HSV2 U40636 ( .A1(n35576), .A2(n35575), .A3(n35574), .Z(n35580) );
  CLKNAND2HSV1 U40637 ( .A1(n35577), .A2(n59601), .ZN(n35579) );
  NAND2HSV2 U40638 ( .A1(n50288), .A2(n57567), .ZN(n35578) );
  XOR3HSV2 U40639 ( .A1(n35580), .A2(n35579), .A3(n35578), .Z(n35581) );
  XOR2HSV0 U40640 ( .A1(n35582), .A2(n35581), .Z(n35586) );
  INHSV4 U40641 ( .I(n35583), .ZN(n50400) );
  CLKNAND2HSV2 U40642 ( .A1(n58183), .A2(n59600), .ZN(n35585) );
  NAND2HSV2 U40643 ( .A1(n57560), .A2(n59603), .ZN(n35584) );
  XOR3HSV2 U40644 ( .A1(n35586), .A2(n35585), .A3(n35584), .Z(n35589) );
  CLKAND2HSV2 U40645 ( .A1(n58103), .A2(n34864), .Z(n35588) );
  XNOR2HSV4 U40646 ( .A1(n35589), .A2(n35588), .ZN(n35590) );
  INHSV2 U40647 ( .I(n50301), .ZN(n57310) );
  NAND2HSV2 U40648 ( .A1(n57310), .A2(n59350), .ZN(n35591) );
  CLKNAND2HSV2 U40649 ( .A1(n35590), .A2(n35591), .ZN(n35595) );
  INHSV3 U40650 ( .I(n35590), .ZN(n35593) );
  INHSV2 U40651 ( .I(n35591), .ZN(n35592) );
  CLKNAND2HSV3 U40652 ( .A1(n35593), .A2(n35592), .ZN(n35594) );
  CLKNAND2HSV3 U40653 ( .A1(n35595), .A2(n35594), .ZN(n35597) );
  CLKNAND2HSV1 U40654 ( .A1(n49921), .A2(n33461), .ZN(n35596) );
  XNOR2HSV4 U40655 ( .A1(n35597), .A2(n35596), .ZN(n35600) );
  CLKNAND2HSV1 U40656 ( .A1(n59666), .A2(n35598), .ZN(n35599) );
  XNOR2HSV4 U40657 ( .A1(n35600), .A2(n35599), .ZN(n35601) );
  XNOR2HSV4 U40658 ( .A1(n35602), .A2(n35601), .ZN(n35603) );
  CLKNAND2HSV1 U40659 ( .A1(n36102), .A2(n31861), .ZN(n35696) );
  BUFHSV2 U40660 ( .I(n49318), .Z(n36103) );
  NAND2HSV2 U40661 ( .A1(n36103), .A2(\pe6/got [24]), .ZN(n35694) );
  BUFHSV2 U40662 ( .I(n59914), .Z(n49667) );
  NAND2HSV2 U40663 ( .A1(n46632), .A2(n59328), .ZN(n35688) );
  BUFHSV2 U40664 ( .I(n44391), .Z(n36105) );
  CLKNAND2HSV1 U40665 ( .A1(n36105), .A2(n46818), .ZN(n35686) );
  BUFHSV2 U40666 ( .I(n59034), .Z(n44392) );
  NAND2HSV2 U40667 ( .A1(n44392), .A2(n35922), .ZN(n35684) );
  NAND2HSV0 U40668 ( .A1(n35722), .A2(n36104), .ZN(n35682) );
  CLKNAND2HSV0 U40669 ( .A1(n58815), .A2(n35723), .ZN(n35680) );
  BUFHSV2 U40670 ( .I(n26109), .Z(n49319) );
  CLKNAND2HSV1 U40671 ( .A1(n49319), .A2(n36106), .ZN(n35678) );
  BUFHSV2 U40672 ( .I(n59678), .Z(n36107) );
  CLKNAND2HSV1 U40673 ( .A1(n36107), .A2(\pe6/got [14]), .ZN(n35674) );
  NAND2HSV0 U40674 ( .A1(n59183), .A2(n58711), .ZN(n35672) );
  NAND2HSV2 U40675 ( .A1(n35724), .A2(\pe6/got [10]), .ZN(n35606) );
  BUFHSV2 U40676 ( .I(n59037), .Z(n58525) );
  NAND2HSV0 U40677 ( .A1(n59038), .A2(n58525), .ZN(n35605) );
  XOR2HSV0 U40678 ( .A1(n35606), .A2(n35605), .Z(n35665) );
  NAND2HSV0 U40679 ( .A1(n44453), .A2(n33024), .ZN(n59196) );
  NOR2HSV0 U40680 ( .A1(n44397), .A2(n58537), .ZN(n58871) );
  INHSV1 U40681 ( .I(n58537), .ZN(n59099) );
  CLKNHSV0 U40682 ( .I(n35607), .ZN(n49836) );
  AOI22HSV0 U40683 ( .A1(n59071), .A2(n59099), .B1(n59051), .B2(n49836), .ZN(
        n35608) );
  AOI21HSV0 U40684 ( .A1(n35609), .A2(n58871), .B(n35608), .ZN(n35611) );
  NOR2HSV0 U40685 ( .A1(n35837), .A2(n46637), .ZN(n35927) );
  NAND2HSV0 U40686 ( .A1(n36168), .A2(\pe6/aot [23]), .ZN(n49328) );
  XOR2HSV0 U40687 ( .A1(n35927), .A2(n49328), .Z(n35610) );
  XOR3HSV1 U40688 ( .A1(n59196), .A2(n35611), .A3(n35610), .Z(n35628) );
  NAND2HSV0 U40689 ( .A1(n35612), .A2(n59182), .ZN(n35627) );
  NOR2HSV0 U40690 ( .A1(n46688), .A2(n32373), .ZN(n35614) );
  NAND2HSV0 U40691 ( .A1(n44336), .A2(n46677), .ZN(n35613) );
  XOR2HSV0 U40692 ( .A1(n35614), .A2(n35613), .Z(n35618) );
  NAND2HSV0 U40693 ( .A1(n35760), .A2(\pe6/aot [11]), .ZN(n35616) );
  NAND2HSV0 U40694 ( .A1(n36143), .A2(n59272), .ZN(n35615) );
  XOR2HSV0 U40695 ( .A1(n35616), .A2(n35615), .Z(n35617) );
  XOR2HSV0 U40696 ( .A1(n35618), .A2(n35617), .Z(n35625) );
  NOR2HSV0 U40697 ( .A1(n31791), .A2(n58983), .ZN(n35620) );
  INHSV2 U40698 ( .I(\pe6/aot [7]), .ZN(n58392) );
  CLKNHSV2 U40699 ( .I(n58392), .ZN(n46792) );
  CLKNAND2HSV1 U40700 ( .A1(n46627), .A2(n46792), .ZN(n35619) );
  XOR2HSV0 U40701 ( .A1(n35620), .A2(n35619), .Z(n35623) );
  NAND2HSV0 U40702 ( .A1(n46176), .A2(n36109), .ZN(n35621) );
  XOR2HSV0 U40703 ( .A1(n35621), .A2(\pe6/phq [26]), .Z(n35622) );
  XOR2HSV0 U40704 ( .A1(n35623), .A2(n35622), .Z(n35624) );
  XOR2HSV0 U40705 ( .A1(n35625), .A2(n35624), .Z(n35626) );
  XOR3HSV2 U40706 ( .A1(n35628), .A2(n35627), .A3(n35626), .Z(n35663) );
  CLKNAND2HSV0 U40707 ( .A1(n59100), .A2(\pe6/aot [17]), .ZN(n35630) );
  INHSV2 U40708 ( .I(n44436), .ZN(n58628) );
  NAND2HSV0 U40709 ( .A1(n58628), .A2(n35925), .ZN(n35629) );
  XOR2HSV0 U40710 ( .A1(n35630), .A2(n35629), .Z(n35636) );
  CLKNAND2HSV1 U40711 ( .A1(n46658), .A2(n35632), .ZN(n35634) );
  NAND2HSV0 U40712 ( .A1(n59206), .A2(n49208), .ZN(n35633) );
  XOR2HSV0 U40713 ( .A1(n35634), .A2(n35633), .Z(n35635) );
  XOR2HSV0 U40714 ( .A1(n35636), .A2(n35635), .Z(n35644) );
  CLKNHSV0 U40715 ( .I(n50837), .ZN(n58749) );
  CLKNAND2HSV1 U40716 ( .A1(n58682), .A2(n58749), .ZN(n35638) );
  CLKNAND2HSV0 U40717 ( .A1(n59054), .A2(n35732), .ZN(n35637) );
  XOR2HSV0 U40718 ( .A1(n35638), .A2(n35637), .Z(n35642) );
  CLKNHSV0 U40719 ( .I(n59205), .ZN(n49862) );
  NAND2HSV0 U40720 ( .A1(n49862), .A2(n35726), .ZN(n35640) );
  NAND2HSV0 U40721 ( .A1(n46210), .A2(n58991), .ZN(n35639) );
  XOR2HSV0 U40722 ( .A1(n35640), .A2(n35639), .Z(n35641) );
  XOR2HSV0 U40723 ( .A1(n35642), .A2(n35641), .Z(n35643) );
  XOR2HSV0 U40724 ( .A1(n35644), .A2(n35643), .Z(n35661) );
  CLKNHSV0 U40725 ( .I(n46663), .ZN(n35956) );
  NAND2HSV2 U40726 ( .A1(n58668), .A2(n35956), .ZN(n35646) );
  CLKNAND2HSV0 U40727 ( .A1(n36150), .A2(\pe6/aot [21]), .ZN(n35645) );
  XOR2HSV0 U40728 ( .A1(n35646), .A2(n35645), .Z(n35651) );
  CLKNHSV0 U40729 ( .I(n35647), .ZN(n58965) );
  CLKNAND2HSV0 U40730 ( .A1(n58965), .A2(n32972), .ZN(n35649) );
  CLKNHSV0 U40731 ( .I(n31253), .ZN(n46230) );
  CLKNAND2HSV1 U40732 ( .A1(n59075), .A2(n46230), .ZN(n35648) );
  XOR2HSV0 U40733 ( .A1(n35649), .A2(n35648), .Z(n35650) );
  XOR2HSV0 U40734 ( .A1(n35651), .A2(n35650), .Z(n35659) );
  NAND2HSV0 U40735 ( .A1(n59246), .A2(n36114), .ZN(n35926) );
  NAND2HSV0 U40736 ( .A1(n59201), .A2(\pe6/pvq [26]), .ZN(n35652) );
  XOR2HSV0 U40737 ( .A1(n35926), .A2(n35652), .Z(n35657) );
  CLKNAND2HSV0 U40738 ( .A1(n35768), .A2(n58488), .ZN(n35655) );
  NAND2HSV0 U40739 ( .A1(n48051), .A2(n32981), .ZN(n35654) );
  XOR2HSV0 U40740 ( .A1(n35655), .A2(n35654), .Z(n35656) );
  XOR2HSV0 U40741 ( .A1(n35657), .A2(n35656), .Z(n35658) );
  XOR2HSV0 U40742 ( .A1(n35659), .A2(n35658), .Z(n35660) );
  XOR2HSV0 U40743 ( .A1(n35661), .A2(n35660), .Z(n35662) );
  XNOR2HSV1 U40744 ( .A1(n35663), .A2(n35662), .ZN(n35664) );
  XNOR2HSV1 U40745 ( .A1(n35665), .A2(n35664), .ZN(n35667) );
  CLKNHSV0 U40746 ( .I(n53110), .ZN(n44477) );
  CLKNAND2HSV1 U40747 ( .A1(n32900), .A2(n44477), .ZN(n35666) );
  XOR2HSV0 U40748 ( .A1(n35667), .A2(n35666), .Z(n35670) );
  NAND2HSV0 U40749 ( .A1(n36183), .A2(n58719), .ZN(n35669) );
  XNOR2HSV1 U40750 ( .A1(n35670), .A2(n35669), .ZN(n35671) );
  XNOR2HSV1 U40751 ( .A1(n35672), .A2(n35671), .ZN(n35673) );
  XNOR2HSV1 U40752 ( .A1(n35674), .A2(n35673), .ZN(n35676) );
  NAND2HSV0 U40753 ( .A1(n36185), .A2(\pe6/got [15]), .ZN(n35675) );
  XNOR2HSV1 U40754 ( .A1(n35676), .A2(n35675), .ZN(n35677) );
  XOR2HSV0 U40755 ( .A1(n35678), .A2(n35677), .Z(n35679) );
  XNOR2HSV1 U40756 ( .A1(n35680), .A2(n35679), .ZN(n35681) );
  XOR2HSV0 U40757 ( .A1(n35682), .A2(n35681), .Z(n35683) );
  XOR2HSV0 U40758 ( .A1(n35684), .A2(n35683), .Z(n35685) );
  XNOR2HSV1 U40759 ( .A1(n35686), .A2(n35685), .ZN(n35687) );
  XOR2HSV0 U40760 ( .A1(n35688), .A2(n35687), .Z(n35690) );
  NAND2HSV0 U40761 ( .A1(n58901), .A2(n59175), .ZN(n35689) );
  XOR2HSV0 U40762 ( .A1(n35690), .A2(n35689), .Z(n35692) );
  INHSV2 U40763 ( .I(n50805), .ZN(n59676) );
  CLKNAND2HSV1 U40764 ( .A1(n59676), .A2(n59174), .ZN(n35691) );
  XOR2HSV0 U40765 ( .A1(n35692), .A2(n35691), .Z(n35693) );
  XOR2HSV0 U40766 ( .A1(n35694), .A2(n35693), .Z(n35695) );
  XNOR2HSV1 U40767 ( .A1(n35696), .A2(n35695), .ZN(n35698) );
  CLKBUFHSV4 U40768 ( .I(n46170), .Z(n44390) );
  CLKNAND2HSV1 U40769 ( .A1(n44390), .A2(n32354), .ZN(n35697) );
  XNOR2HSV1 U40770 ( .A1(n35698), .A2(n35697), .ZN(n35700) );
  BUFHSV2 U40771 ( .I(n35788), .Z(n36196) );
  CLKNAND2HSV1 U40772 ( .A1(n36196), .A2(n49665), .ZN(n35699) );
  CLKNAND2HSV0 U40773 ( .A1(n46825), .A2(n46289), .ZN(n35701) );
  XNOR2HSV1 U40774 ( .A1(n35702), .A2(n35701), .ZN(n35707) );
  CLKNAND2HSV1 U40775 ( .A1(n25860), .A2(n35705), .ZN(n35706) );
  NAND3HSV4 U40776 ( .A1(n35904), .A2(n35709), .A3(n35903), .ZN(n36203) );
  XNOR2HSV4 U40777 ( .A1(n35714), .A2(n35713), .ZN(n35918) );
  INAND2HSV2 U40778 ( .A1(n32457), .B1(n35918), .ZN(n35711) );
  NAND2HSV2 U40779 ( .A1(n36206), .A2(n36207), .ZN(n35712) );
  OAI21HSV2 U40780 ( .A1(n36034), .A2(n46765), .B(n44519), .ZN(n35715) );
  AOI21HSV4 U40781 ( .A1(n35716), .A2(n35712), .B(n35715), .ZN(n44358) );
  INHSV4 U40782 ( .I(n35717), .ZN(n35718) );
  CLKNAND2HSV4 U40783 ( .A1(n35719), .A2(n35718), .ZN(n35720) );
  NAND2HSV2 U40784 ( .A1(n49319), .A2(n35723), .ZN(n35774) );
  NOR2HSV0 U40785 ( .A1(n46688), .A2(n49699), .ZN(n35728) );
  NAND2HSV0 U40786 ( .A1(n59100), .A2(n35726), .ZN(n35727) );
  XOR2HSV0 U40787 ( .A1(n35728), .A2(n35727), .Z(n35731) );
  NAND2HSV0 U40788 ( .A1(n46176), .A2(\pe6/got [8]), .ZN(n35729) );
  XOR2HSV0 U40789 ( .A1(n35729), .A2(\pe6/phq [25]), .Z(n35730) );
  CLKNAND2HSV1 U40790 ( .A1(n58962), .A2(n35732), .ZN(n49322) );
  OAI22HSV0 U40791 ( .A1(n32714), .A2(n49680), .B1(n59194), .B2(n46789), .ZN(
        n35733) );
  OAI21HSV0 U40792 ( .A1(n35734), .A2(n49322), .B(n35733), .ZN(n35738) );
  INHSV2 U40793 ( .I(\pe6/bq[9] ), .ZN(n50847) );
  OAI22HSV0 U40794 ( .A1(n31253), .A2(n48042), .B1(n50847), .B2(n32086), .ZN(
        n35735) );
  OAI21HSV1 U40795 ( .A1(n35926), .A2(n35736), .B(n35735), .ZN(n35737) );
  NOR2HSV0 U40796 ( .A1(n35837), .A2(n35607), .ZN(n58859) );
  NAND2HSV0 U40797 ( .A1(n59201), .A2(\pe6/pvq [25]), .ZN(n35742) );
  NAND2HSV0 U40798 ( .A1(n35740), .A2(\pe6/aot [10]), .ZN(n35741) );
  NAND2HSV0 U40799 ( .A1(n35743), .A2(n58857), .ZN(n35745) );
  NAND2HSV0 U40800 ( .A1(n59267), .A2(\pe6/aot [13]), .ZN(n35744) );
  XOR2HSV0 U40801 ( .A1(n35745), .A2(n35744), .Z(n35749) );
  NAND2HSV0 U40802 ( .A1(n58668), .A2(n59272), .ZN(n35747) );
  NAND2HSV0 U40803 ( .A1(n32568), .A2(\pe6/aot [19]), .ZN(n35746) );
  XOR2HSV0 U40804 ( .A1(n35747), .A2(n35746), .Z(n35748) );
  NAND2HSV0 U40805 ( .A1(n35750), .A2(n46677), .ZN(n35753) );
  NAND2HSV0 U40806 ( .A1(n35751), .A2(n59245), .ZN(n35752) );
  XOR2HSV0 U40807 ( .A1(n35753), .A2(n35752), .Z(n35757) );
  CLKNAND2HSV1 U40808 ( .A1(n36150), .A2(n33004), .ZN(n35755) );
  NAND2HSV0 U40809 ( .A1(n59206), .A2(n33024), .ZN(n35754) );
  XOR2HSV0 U40810 ( .A1(n35755), .A2(n35754), .Z(n35756) );
  NAND2HSV0 U40811 ( .A1(n36168), .A2(n59239), .ZN(n35759) );
  CLKNAND2HSV0 U40812 ( .A1(n32252), .A2(n49208), .ZN(n35758) );
  XOR2HSV0 U40813 ( .A1(n35759), .A2(n35758), .Z(n35765) );
  NAND2HSV0 U40814 ( .A1(n35760), .A2(n32972), .ZN(n35763) );
  NAND2HSV0 U40815 ( .A1(n35761), .A2(\pe6/aot [21]), .ZN(n35762) );
  XOR2HSV0 U40816 ( .A1(n35763), .A2(n35762), .Z(n35764) );
  CLKNAND2HSV0 U40817 ( .A1(n59054), .A2(\pe6/aot [17]), .ZN(n35767) );
  NAND2HSV0 U40818 ( .A1(n59240), .A2(n58991), .ZN(n35766) );
  XOR2HSV0 U40819 ( .A1(n35767), .A2(n35766), .Z(n35772) );
  CLKNAND2HSV1 U40820 ( .A1(n46658), .A2(n59099), .ZN(n35770) );
  NAND2HSV0 U40821 ( .A1(n35768), .A2(\pe6/aot [11]), .ZN(n35769) );
  XOR2HSV0 U40822 ( .A1(n35770), .A2(n35769), .Z(n35771) );
  INHSV2 U40823 ( .I(n35779), .ZN(n35783) );
  INHSV2 U40824 ( .I(n35777), .ZN(n46760) );
  CLKNAND2HSV0 U40825 ( .A1(n35783), .A2(n46760), .ZN(n35781) );
  NOR2HSV0 U40826 ( .A1(n35778), .A2(n35777), .ZN(n35780) );
  NOR2HSV1 U40827 ( .A1(n35783), .A2(n35782), .ZN(n35785) );
  NAND2HSV2 U40828 ( .A1(n49726), .A2(n46289), .ZN(n35791) );
  CLKNAND2HSV1 U40829 ( .A1(n44390), .A2(n35789), .ZN(n35790) );
  XOR2HSV0 U40830 ( .A1(n35791), .A2(n35790), .Z(n35792) );
  XOR2HSV2 U40831 ( .A1(n35793), .A2(n35792), .Z(n35794) );
  NAND2HSV4 U40832 ( .A1(n36203), .A2(n46567), .ZN(n35800) );
  XNOR2HSV4 U40833 ( .A1(n35801), .A2(n35800), .ZN(n36057) );
  NOR2HSV0 U40834 ( .A1(n35797), .A2(\pe6/ti_7t [25]), .ZN(n36214) );
  NOR2HSV2 U40835 ( .A1(n36214), .A2(n46549), .ZN(n35799) );
  OAI21HSV4 U40836 ( .A1(n35912), .A2(n36057), .B(n35799), .ZN(n36038) );
  XNOR2HSV4 U40837 ( .A1(n35801), .A2(n35800), .ZN(n35915) );
  CLKNHSV0 U40838 ( .I(n36053), .ZN(n35802) );
  INHSV4 U40839 ( .I(n35803), .ZN(n36039) );
  NOR2HSV8 U40840 ( .A1(n36038), .A2(n36039), .ZN(n44359) );
  NAND4HSV2 U40841 ( .A1(n44358), .A2(n29649), .A3(n59168), .A4(n44359), .ZN(
        n35811) );
  INHSV2 U40842 ( .I(n35918), .ZN(n35805) );
  NAND2HSV4 U40843 ( .A1(n36206), .A2(n36207), .ZN(n46824) );
  NOR2HSV2 U40844 ( .A1(n35805), .A2(n46824), .ZN(n35804) );
  NOR2HSV4 U40845 ( .A1(n44359), .A2(n35804), .ZN(n44355) );
  CLKNHSV3 U40846 ( .I(n35912), .ZN(n35910) );
  INHSV2 U40847 ( .I(n32530), .ZN(n36095) );
  NAND3HSV4 U40848 ( .A1(n35805), .A2(n35910), .A3(n36095), .ZN(n44352) );
  AOI21HSV4 U40849 ( .A1(n36034), .A2(n44372), .B(n35806), .ZN(n36090) );
  INHSV2 U40850 ( .I(n36090), .ZN(n44353) );
  NOR2HSV2 U40851 ( .A1(n44353), .A2(n35710), .ZN(n35807) );
  CLKAND2HSV2 U40852 ( .A1(n32329), .A2(\pe6/ti_7t [26]), .Z(n44357) );
  CLKNAND2HSV0 U40853 ( .A1(n44357), .A2(n35808), .ZN(n35809) );
  NAND3HSV3 U40854 ( .A1(n35811), .A2(n35810), .A3(n35809), .ZN(n36225) );
  CLKNAND2HSV0 U40855 ( .A1(n26152), .A2(n59025), .ZN(n35902) );
  CLKNAND2HSV1 U40856 ( .A1(n46769), .A2(n46283), .ZN(n35900) );
  BUFHSV2 U40857 ( .I(n46592), .Z(n58663) );
  BUFHSV2 U40858 ( .I(n49667), .Z(n58722) );
  CLKNHSV0 U40859 ( .I(n49666), .ZN(n46171) );
  CLKNAND2HSV0 U40860 ( .A1(n49743), .A2(n32596), .ZN(n35896) );
  BUFHSV2 U40861 ( .I(n32165), .Z(n49829) );
  NAND2HSV0 U40862 ( .A1(n49829), .A2(n35991), .ZN(n35894) );
  NAND2HSV0 U40863 ( .A1(n49319), .A2(n58711), .ZN(n35892) );
  CLKNAND2HSV1 U40864 ( .A1(n59678), .A2(n44477), .ZN(n35888) );
  NAND2HSV0 U40865 ( .A1(n59183), .A2(n58812), .ZN(n35886) );
  NAND2HSV0 U40866 ( .A1(n35724), .A2(n58814), .ZN(n35815) );
  BUFHSV2 U40867 ( .I(\pe6/got [6]), .Z(n58399) );
  NAND2HSV0 U40868 ( .A1(n59038), .A2(n58399), .ZN(n35814) );
  XOR2HSV0 U40869 ( .A1(n35815), .A2(n35814), .Z(n35880) );
  NAND2HSV0 U40870 ( .A1(n59246), .A2(n59065), .ZN(n35819) );
  NAND2HSV0 U40871 ( .A1(n58460), .A2(n59234), .ZN(n35818) );
  XOR2HSV0 U40872 ( .A1(n35819), .A2(n35818), .Z(n35823) );
  BUFHSV2 U40873 ( .I(n58537), .Z(n59193) );
  INHSV2 U40874 ( .I(n59193), .ZN(n46197) );
  NAND2HSV0 U40875 ( .A1(n58965), .A2(n46197), .ZN(n35821) );
  NAND2HSV0 U40876 ( .A1(n59247), .A2(n46792), .ZN(n35820) );
  XOR2HSV0 U40877 ( .A1(n35821), .A2(n35820), .Z(n35822) );
  XOR2HSV0 U40878 ( .A1(n35823), .A2(n35822), .Z(n35847) );
  BUFHSV2 U40879 ( .I(\pe6/got [5]), .Z(n58400) );
  NAND2HSV0 U40880 ( .A1(n44426), .A2(n58400), .ZN(n35846) );
  BUFHSV2 U40881 ( .I(\pe6/aot [6]), .Z(n59266) );
  NAND2HSV0 U40882 ( .A1(n46672), .A2(n59266), .ZN(n35825) );
  NAND2HSV0 U40883 ( .A1(n49862), .A2(\pe6/aot [15]), .ZN(n35824) );
  XOR2HSV0 U40884 ( .A1(n35825), .A2(n35824), .Z(n35829) );
  NAND2HSV0 U40885 ( .A1(n36150), .A2(n58760), .ZN(n35827) );
  NAND2HSV0 U40886 ( .A1(n36168), .A2(n44439), .ZN(n35826) );
  XOR2HSV0 U40887 ( .A1(n35827), .A2(n35826), .Z(n35828) );
  XOR2HSV0 U40888 ( .A1(n35829), .A2(n35828), .Z(n35845) );
  CLKNAND2HSV0 U40889 ( .A1(n59224), .A2(\pe6/aot [17]), .ZN(n35831) );
  NAND2HSV0 U40890 ( .A1(n46624), .A2(\pe6/aot [11]), .ZN(n35830) );
  XOR2HSV0 U40891 ( .A1(n35831), .A2(n35830), .Z(n35835) );
  NAND2HSV0 U40892 ( .A1(n58668), .A2(n33004), .ZN(n35833) );
  NAND2HSV0 U40893 ( .A1(n46210), .A2(n35956), .ZN(n35832) );
  XOR2HSV0 U40894 ( .A1(n35833), .A2(n35832), .Z(n35834) );
  XOR2HSV0 U40895 ( .A1(n35835), .A2(n35834), .Z(n35843) );
  NAND2HSV0 U40896 ( .A1(n46176), .A2(n46173), .ZN(n35836) );
  XOR2HSV0 U40897 ( .A1(n35836), .A2(\pe6/phq [29]), .Z(n35841) );
  CLKNAND2HSV0 U40898 ( .A1(n33005), .A2(n59250), .ZN(n58766) );
  CLKNAND2HSV0 U40899 ( .A1(n33005), .A2(n35732), .ZN(n44399) );
  OAI21HSV0 U40900 ( .A1(n58359), .A2(n44411), .B(n44399), .ZN(n35838) );
  OAI21HSV0 U40901 ( .A1(n35839), .A2(n58766), .B(n35838), .ZN(n35840) );
  XOR2HSV0 U40902 ( .A1(n35841), .A2(n35840), .Z(n35842) );
  XNOR2HSV1 U40903 ( .A1(n35843), .A2(n35842), .ZN(n35844) );
  XOR4HSV1 U40904 ( .A1(n35847), .A2(n35846), .A3(n35845), .A4(n35844), .Z(
        n35878) );
  NAND2HSV0 U40905 ( .A1(n58628), .A2(n32981), .ZN(n35849) );
  NAND2HSV0 U40906 ( .A1(n46627), .A2(\pe6/aot [4]), .ZN(n35848) );
  XOR2HSV0 U40907 ( .A1(n35849), .A2(n35848), .Z(n35853) );
  NAND2HSV0 U40908 ( .A1(n32252), .A2(n58488), .ZN(n35851) );
  INHSV2 U40909 ( .I(n46147), .ZN(n58618) );
  NAND2HSV0 U40910 ( .A1(n58618), .A2(n35925), .ZN(n35850) );
  XOR2HSV0 U40911 ( .A1(n35851), .A2(n35850), .Z(n35852) );
  XOR2HSV0 U40912 ( .A1(n35853), .A2(n35852), .Z(n35861) );
  NAND2HSV0 U40913 ( .A1(n44453), .A2(n53115), .ZN(n35855) );
  NAND2HSV0 U40914 ( .A1(n48051), .A2(n58749), .ZN(n35854) );
  XOR2HSV0 U40915 ( .A1(n35855), .A2(n35854), .Z(n35859) );
  INHSV2 U40916 ( .I(n46146), .ZN(n48037) );
  NAND2HSV0 U40917 ( .A1(n48037), .A2(n36114), .ZN(n35857) );
  NAND2HSV0 U40918 ( .A1(n59054), .A2(\pe6/aot [13]), .ZN(n35856) );
  XOR2HSV0 U40919 ( .A1(n35857), .A2(n35856), .Z(n35858) );
  XOR2HSV0 U40920 ( .A1(n35859), .A2(n35858), .Z(n35860) );
  XOR2HSV0 U40921 ( .A1(n35861), .A2(n35860), .Z(n35876) );
  CLKNAND2HSV0 U40922 ( .A1(\pe6/bq[10] ), .A2(n59272), .ZN(n35863) );
  NAND2HSV0 U40923 ( .A1(\pe6/bq[4] ), .A2(n46230), .ZN(n35862) );
  XOR2HSV0 U40924 ( .A1(n35863), .A2(n35862), .Z(n35868) );
  NAND2HSV0 U40925 ( .A1(n36143), .A2(n36153), .ZN(n35866) );
  NAND2HSV0 U40926 ( .A1(n35751), .A2(\pe6/aot [21]), .ZN(n35865) );
  XOR2HSV0 U40927 ( .A1(n35866), .A2(n35865), .Z(n35867) );
  XOR2HSV0 U40928 ( .A1(n35868), .A2(n35867), .Z(n35874) );
  NOR2HSV0 U40929 ( .A1(n46688), .A2(n46637), .ZN(n59191) );
  CLKNAND2HSV0 U40930 ( .A1(n35760), .A2(n58857), .ZN(n36126) );
  XOR2HSV0 U40931 ( .A1(n59191), .A2(n36126), .Z(n35872) );
  CLKNAND2HSV1 U40932 ( .A1(n48046), .A2(\pe6/pvq [29]), .ZN(n35870) );
  NAND2HSV0 U40933 ( .A1(n44435), .A2(n58943), .ZN(n35869) );
  XOR2HSV0 U40934 ( .A1(n35870), .A2(n35869), .Z(n35871) );
  XOR2HSV0 U40935 ( .A1(n35872), .A2(n35871), .Z(n35873) );
  XOR2HSV0 U40936 ( .A1(n35874), .A2(n35873), .Z(n35875) );
  XOR2HSV0 U40937 ( .A1(n35876), .A2(n35875), .Z(n35877) );
  XNOR2HSV1 U40938 ( .A1(n35878), .A2(n35877), .ZN(n35879) );
  XNOR2HSV1 U40939 ( .A1(n35880), .A2(n35879), .ZN(n35882) );
  NAND2HSV0 U40940 ( .A1(n32900), .A2(n58526), .ZN(n35881) );
  XNOR2HSV1 U40941 ( .A1(n35882), .A2(n35881), .ZN(n35884) );
  NAND2HSV0 U40942 ( .A1(n25218), .A2(n58525), .ZN(n35883) );
  XNOR2HSV1 U40943 ( .A1(n35884), .A2(n35883), .ZN(n35885) );
  XNOR2HSV1 U40944 ( .A1(n35886), .A2(n35885), .ZN(n35887) );
  XNOR2HSV1 U40945 ( .A1(n35888), .A2(n35887), .ZN(n35890) );
  NAND2HSV0 U40946 ( .A1(n36185), .A2(n58719), .ZN(n35889) );
  XNOR2HSV1 U40947 ( .A1(n35890), .A2(n35889), .ZN(n35891) );
  XOR2HSV0 U40948 ( .A1(n35892), .A2(n35891), .Z(n35893) );
  XOR2HSV0 U40949 ( .A1(n35894), .A2(n35893), .Z(n35895) );
  XOR2HSV0 U40950 ( .A1(n35896), .A2(n35895), .Z(n35897) );
  XNOR2HSV1 U40951 ( .A1(n35900), .A2(n35899), .ZN(n35901) );
  XNOR2HSV1 U40952 ( .A1(n35902), .A2(n35901), .ZN(n35906) );
  NAND3HSV2 U40953 ( .A1(n35709), .A2(n35904), .A3(n35903), .ZN(n44508) );
  BUFHSV2 U40954 ( .I(n44508), .Z(n59677) );
  NAND2HSV2 U40955 ( .A1(n59677), .A2(n49665), .ZN(n35905) );
  CLKNHSV0 U40956 ( .I(n35915), .ZN(n35909) );
  CLKNAND2HSV2 U40957 ( .A1(n35909), .A2(n32234), .ZN(n35911) );
  NOR2HSV0 U40958 ( .A1(n36214), .A2(n35777), .ZN(n35916) );
  XNOR2HSV4 U40959 ( .A1(n36225), .A2(n36224), .ZN(n36071) );
  CLKNHSV0 U40960 ( .I(n35917), .ZN(n46154) );
  BUFHSV2 U40961 ( .I(n46154), .Z(n46163) );
  CLKNAND2HSV2 U40962 ( .A1(n36053), .A2(n44344), .ZN(n36035) );
  NAND2HSV0 U40963 ( .A1(n35919), .A2(n49665), .ZN(n35920) );
  NOR2HSV1 U40964 ( .A1(n35921), .A2(n35920), .ZN(n36019) );
  CLKNAND2HSV1 U40965 ( .A1(n44390), .A2(n31861), .ZN(n36015) );
  CLKNAND2HSV0 U40966 ( .A1(n36102), .A2(\pe6/got [24]), .ZN(n36013) );
  INHSV2 U40967 ( .I(n49315), .ZN(n58808) );
  CLKNAND2HSV1 U40968 ( .A1(n36103), .A2(n58808), .ZN(n36011) );
  CLKNAND2HSV1 U40969 ( .A1(n46632), .A2(n59176), .ZN(n36005) );
  CLKNAND2HSV0 U40970 ( .A1(n36105), .A2(n35922), .ZN(n36003) );
  CLKNAND2HSV1 U40971 ( .A1(n44392), .A2(n36104), .ZN(n36001) );
  CLKNAND2HSV1 U40972 ( .A1(n49743), .A2(n49098), .ZN(n35999) );
  NAND2HSV0 U40973 ( .A1(n58815), .A2(n36106), .ZN(n35997) );
  CLKNAND2HSV0 U40974 ( .A1(n49319), .A2(\pe6/got [15]), .ZN(n35995) );
  CLKNAND2HSV0 U40975 ( .A1(n36107), .A2(\pe6/got [13]), .ZN(n35990) );
  NAND2HSV0 U40976 ( .A1(n32167), .A2(n59180), .ZN(n35988) );
  NAND2HSV0 U40977 ( .A1(n35724), .A2(n58525), .ZN(n35924) );
  CLKNAND2HSV0 U40978 ( .A1(n59038), .A2(n58526), .ZN(n35923) );
  XOR2HSV0 U40979 ( .A1(n35924), .A2(n35923), .Z(n35982) );
  NAND2HSV0 U40980 ( .A1(n59075), .A2(n35925), .ZN(n36127) );
  NAND2HSV2 U40981 ( .A1(n59224), .A2(n58760), .ZN(n36160) );
  CLKNAND2HSV1 U40982 ( .A1(n35768), .A2(n59099), .ZN(n36125) );
  XOR2HSV0 U40983 ( .A1(n35929), .A2(n36125), .Z(n35930) );
  XNOR2HSV1 U40984 ( .A1(n35931), .A2(n35930), .ZN(n35947) );
  NAND2HSV0 U40985 ( .A1(n44426), .A2(n36109), .ZN(n35946) );
  NOR2HSV2 U40986 ( .A1(n59094), .A2(n32877), .ZN(n35933) );
  CLKNAND2HSV0 U40987 ( .A1(n44336), .A2(n59065), .ZN(n35932) );
  XOR2HSV0 U40988 ( .A1(n35933), .A2(n35932), .Z(n35937) );
  NAND2HSV0 U40989 ( .A1(n46627), .A2(n59266), .ZN(n35935) );
  NAND2HSV0 U40990 ( .A1(n44453), .A2(n49208), .ZN(n35934) );
  XOR2HSV0 U40991 ( .A1(n35935), .A2(n35934), .Z(n35936) );
  XOR2HSV0 U40992 ( .A1(n35937), .A2(n35936), .Z(n35944) );
  NOR2HSV0 U40993 ( .A1(n46192), .A2(n49188), .ZN(n35939) );
  INHSV2 U40994 ( .I(n46147), .ZN(n48038) );
  NAND2HSV0 U40995 ( .A1(n48038), .A2(n46230), .ZN(n35938) );
  XOR2HSV0 U40996 ( .A1(n35939), .A2(n35938), .Z(n35942) );
  NAND2HSV0 U40997 ( .A1(n46176), .A2(n58399), .ZN(n35940) );
  XOR2HSV0 U40998 ( .A1(n35940), .A2(\pe6/phq [27]), .Z(n35941) );
  XOR2HSV0 U40999 ( .A1(n35942), .A2(n35941), .Z(n35943) );
  XOR2HSV0 U41000 ( .A1(n35944), .A2(n35943), .Z(n35945) );
  XOR3HSV2 U41001 ( .A1(n35947), .A2(n35946), .A3(n35945), .Z(n35980) );
  CLKNAND2HSV0 U41002 ( .A1(n59054), .A2(\pe6/aot [15]), .ZN(n35949) );
  NAND2HSV0 U41003 ( .A1(n32982), .A2(\pe6/aot [21]), .ZN(n35948) );
  XOR2HSV0 U41004 ( .A1(n35949), .A2(n35948), .Z(n35953) );
  NAND2HSV0 U41005 ( .A1(n35760), .A2(n58488), .ZN(n35951) );
  NAND2HSV0 U41006 ( .A1(n58682), .A2(n36153), .ZN(n35950) );
  XOR2HSV0 U41007 ( .A1(n35951), .A2(n35950), .Z(n35952) );
  XOR2HSV0 U41008 ( .A1(n35953), .A2(n35952), .Z(n35962) );
  CLKNAND2HSV0 U41009 ( .A1(n46658), .A2(n46792), .ZN(n35955) );
  NAND2HSV0 U41010 ( .A1(n58628), .A2(n46677), .ZN(n35954) );
  XOR2HSV0 U41011 ( .A1(n35955), .A2(n35954), .Z(n35960) );
  NAND2HSV2 U41012 ( .A1(n59206), .A2(\pe6/aot [13]), .ZN(n35958) );
  NAND2HSV0 U41013 ( .A1(n36143), .A2(n35956), .ZN(n35957) );
  XOR2HSV0 U41014 ( .A1(n35958), .A2(n35957), .Z(n35959) );
  XOR2HSV0 U41015 ( .A1(n35960), .A2(n35959), .Z(n35961) );
  XOR2HSV0 U41016 ( .A1(n35962), .A2(n35961), .Z(n35978) );
  NAND2HSV0 U41017 ( .A1(n58965), .A2(\pe6/aot [11]), .ZN(n35964) );
  NAND2HSV0 U41018 ( .A1(n59071), .A2(n58857), .ZN(n35963) );
  XOR2HSV0 U41019 ( .A1(n35964), .A2(n35963), .Z(n35968) );
  CLKNAND2HSV1 U41020 ( .A1(n44435), .A2(n59044), .ZN(n35966) );
  CLKNAND2HSV0 U41021 ( .A1(n49862), .A2(\pe6/aot [17]), .ZN(n35965) );
  XOR2HSV0 U41022 ( .A1(n35966), .A2(n35965), .Z(n35967) );
  XOR2HSV0 U41023 ( .A1(n35968), .A2(n35967), .Z(n35976) );
  NOR2HSV0 U41024 ( .A1(n46850), .A2(n32589), .ZN(n35970) );
  NAND2HSV2 U41025 ( .A1(n53214), .A2(\pe6/pvq [27]), .ZN(n35969) );
  XOR2HSV0 U41026 ( .A1(n35970), .A2(n35969), .Z(n35974) );
  CLKNAND2HSV1 U41027 ( .A1(n58668), .A2(n58749), .ZN(n35972) );
  NAND2HSV0 U41028 ( .A1(n36168), .A2(n33004), .ZN(n35971) );
  XOR2HSV0 U41029 ( .A1(n35972), .A2(n35971), .Z(n35973) );
  XOR2HSV0 U41030 ( .A1(n35974), .A2(n35973), .Z(n35975) );
  XOR2HSV0 U41031 ( .A1(n35976), .A2(n35975), .Z(n35977) );
  XOR2HSV0 U41032 ( .A1(n35978), .A2(n35977), .Z(n35979) );
  XNOR2HSV1 U41033 ( .A1(n35980), .A2(n35979), .ZN(n35981) );
  XNOR2HSV1 U41034 ( .A1(n35982), .A2(n35981), .ZN(n35984) );
  CLKNAND2HSV1 U41035 ( .A1(n32900), .A2(n58812), .ZN(n35983) );
  XNOR2HSV1 U41036 ( .A1(n35984), .A2(n35983), .ZN(n35986) );
  CLKNAND2HSV0 U41037 ( .A1(n36183), .A2(n44477), .ZN(n35985) );
  XNOR2HSV1 U41038 ( .A1(n35986), .A2(n35985), .ZN(n35987) );
  XNOR2HSV1 U41039 ( .A1(n35988), .A2(n35987), .ZN(n35989) );
  XNOR2HSV1 U41040 ( .A1(n35990), .A2(n35989), .ZN(n35993) );
  NAND2HSV0 U41041 ( .A1(n36185), .A2(n35991), .ZN(n35992) );
  XNOR2HSV1 U41042 ( .A1(n35993), .A2(n35992), .ZN(n35994) );
  XOR2HSV0 U41043 ( .A1(n35995), .A2(n35994), .Z(n35996) );
  XOR2HSV0 U41044 ( .A1(n35997), .A2(n35996), .Z(n35998) );
  XOR2HSV0 U41045 ( .A1(n35999), .A2(n35998), .Z(n36000) );
  XOR2HSV0 U41046 ( .A1(n36001), .A2(n36000), .Z(n36002) );
  XNOR2HSV1 U41047 ( .A1(n36003), .A2(n36002), .ZN(n36004) );
  XOR2HSV0 U41048 ( .A1(n36005), .A2(n36004), .Z(n36007) );
  CLKNAND2HSV1 U41049 ( .A1(n59317), .A2(n59328), .ZN(n36006) );
  XOR2HSV0 U41050 ( .A1(n36007), .A2(n36006), .Z(n36009) );
  CLKNAND2HSV1 U41051 ( .A1(n59676), .A2(n58714), .ZN(n36008) );
  XOR2HSV0 U41052 ( .A1(n36009), .A2(n36008), .Z(n36010) );
  XOR2HSV0 U41053 ( .A1(n36011), .A2(n36010), .Z(n36012) );
  XNOR2HSV1 U41054 ( .A1(n36013), .A2(n36012), .ZN(n36014) );
  XNOR2HSV1 U41055 ( .A1(n36015), .A2(n36014), .ZN(n36017) );
  CLKNAND2HSV1 U41056 ( .A1(n36196), .A2(n32242), .ZN(n36016) );
  XNOR2HSV1 U41057 ( .A1(n36017), .A2(n36016), .ZN(n36018) );
  XOR2HSV0 U41058 ( .A1(n36019), .A2(n36018), .Z(n36020) );
  XNOR2HSV4 U41059 ( .A1(n36022), .A2(n29690), .ZN(n36028) );
  NAND2HSV0 U41060 ( .A1(n36024), .A2(n36023), .ZN(n36048) );
  CLKNHSV2 U41061 ( .I(n36048), .ZN(n36025) );
  NOR2HSV2 U41062 ( .A1(n36025), .A2(n32651), .ZN(n36026) );
  OAI21HSV2 U41063 ( .A1(n36053), .A2(n36030), .B(n36026), .ZN(n36027) );
  IOA21HSV2 U41064 ( .A1(n36029), .A2(n44342), .B(n26462), .ZN(n36064) );
  CLKNHSV0 U41065 ( .I(n36034), .ZN(n36032) );
  CLKNAND2HSV0 U41066 ( .A1(n36030), .A2(n46574), .ZN(n36033) );
  CLKNAND2HSV1 U41067 ( .A1(n36032), .A2(n36031), .ZN(n36037) );
  NAND3HSV2 U41068 ( .A1(n36035), .A2(n36034), .A3(n36033), .ZN(n36036) );
  INHSV2 U41069 ( .I(n36038), .ZN(n36041) );
  CLKNHSV2 U41070 ( .I(n36039), .ZN(n36040) );
  NAND2HSV2 U41071 ( .A1(n36041), .A2(n36040), .ZN(n36042) );
  NAND2HSV2 U41072 ( .A1(n36044), .A2(n44359), .ZN(n36045) );
  NOR2HSV0 U41073 ( .A1(n46575), .A2(n46549), .ZN(n36047) );
  INHSV2 U41074 ( .I(n36057), .ZN(n47942) );
  INOR2HSV0 U41075 ( .A1(n36048), .B1(n51438), .ZN(n36054) );
  OR2HSV1 U41076 ( .A1(n36054), .A2(n44380), .Z(n36049) );
  OAI21HSV0 U41077 ( .A1(n36053), .A2(n36050), .B(n36049), .ZN(n36051) );
  CLKNAND2HSV1 U41078 ( .A1(n47942), .A2(n36051), .ZN(n36060) );
  CLKNHSV0 U41079 ( .I(\pe6/ti_7t [25]), .ZN(n36052) );
  OR2HSV1 U41080 ( .A1(n46591), .A2(n36052), .Z(n36059) );
  BUFHSV2 U41081 ( .I(n36053), .Z(n46585) );
  INHSV2 U41082 ( .I(n36054), .ZN(n47941) );
  NOR2HSV0 U41083 ( .A1(n47941), .A2(n36055), .ZN(n36056) );
  INHSV2 U41084 ( .I(n49317), .ZN(n44389) );
  NOR2HSV2 U41085 ( .A1(n44389), .A2(n48018), .ZN(n36062) );
  INHSV4 U41086 ( .I(n36087), .ZN(n36069) );
  INHSV4 U41087 ( .I(n36067), .ZN(n36088) );
  INHSV4 U41088 ( .I(n36088), .ZN(n36068) );
  NOR2HSV8 U41089 ( .A1(n36069), .A2(n36068), .ZN(n44692) );
  OAI22HSV2 U41090 ( .A1(n36070), .A2(n44692), .B1(n46765), .B2(n36071), .ZN(
        n36077) );
  INHSV2 U41091 ( .I(n36071), .ZN(n36072) );
  CLKNHSV0 U41092 ( .I(\pe6/ti_7t [28]), .ZN(n36073) );
  AOI21HSV2 U41093 ( .A1(n36073), .A2(n31350), .B(n48010), .ZN(n46568) );
  AND2HSV2 U41094 ( .A1(n46568), .A2(n32685), .Z(n36074) );
  CLKNAND2HSV2 U41095 ( .A1(n36075), .A2(n36074), .ZN(n36076) );
  NOR2HSV2 U41096 ( .A1(n36077), .A2(n36076), .ZN(n36222) );
  INHSV2 U41097 ( .I(n36080), .ZN(n36078) );
  NOR2HSV2 U41098 ( .A1(n36080), .A2(n36029), .ZN(n36082) );
  OAI21HSV1 U41099 ( .A1(\pe6/ti_7t [27]), .A2(n35797), .B(n36081), .ZN(n44339) );
  NAND2HSV0 U41100 ( .A1(n36083), .A2(n46587), .ZN(n36084) );
  NOR2HSV2 U41101 ( .A1(n46575), .A2(n36084), .ZN(n36085) );
  NAND2HSV4 U41102 ( .A1(n47940), .A2(n36085), .ZN(n44341) );
  CLKNAND2HSV1 U41103 ( .A1(n44352), .A2(n29710), .ZN(n36091) );
  INHSV2 U41104 ( .I(n36091), .ZN(n36092) );
  NAND2HSV0 U41105 ( .A1(n44357), .A2(n46765), .ZN(n36093) );
  CLKNAND2HSV1 U41106 ( .A1(n44358), .A2(n36095), .ZN(n36096) );
  NOR2HSV2 U41107 ( .A1(n36097), .A2(n36096), .ZN(n36098) );
  NOR2HSV4 U41108 ( .A1(n36099), .A2(n36098), .ZN(n36221) );
  INAND2HSV4 U41109 ( .A1(n31971), .B1(n26152), .ZN(n36202) );
  CLKNAND2HSV1 U41110 ( .A1(n46769), .A2(n36101), .ZN(n36200) );
  CLKNAND2HSV0 U41111 ( .A1(n44390), .A2(\pe6/got [24]), .ZN(n36195) );
  CLKNAND2HSV0 U41112 ( .A1(n36102), .A2(n59174), .ZN(n36193) );
  CLKNAND2HSV0 U41113 ( .A1(n36103), .A2(n58714), .ZN(n36191) );
  NAND2HSV0 U41114 ( .A1(n36108), .A2(n58526), .ZN(n36111) );
  NAND2HSV0 U41115 ( .A1(n59038), .A2(n36109), .ZN(n36110) );
  XOR2HSV0 U41116 ( .A1(n36111), .A2(n36110), .Z(n36180) );
  NAND2HSV0 U41117 ( .A1(n44453), .A2(\pe6/aot [13]), .ZN(n36113) );
  NAND2HSV0 U41118 ( .A1(n32252), .A2(\pe6/aot [11]), .ZN(n36112) );
  XOR2HSV0 U41119 ( .A1(n36113), .A2(n36112), .Z(n36118) );
  NAND2HSV0 U41120 ( .A1(n58618), .A2(n36114), .ZN(n36116) );
  NAND2HSV0 U41121 ( .A1(n48037), .A2(n46230), .ZN(n36115) );
  XOR2HSV0 U41122 ( .A1(n36116), .A2(n36115), .Z(n36117) );
  XOR2HSV0 U41123 ( .A1(n36118), .A2(n36117), .Z(n36142) );
  NAND2HSV0 U41124 ( .A1(n46176), .A2(n58400), .ZN(n36119) );
  XOR2HSV0 U41125 ( .A1(n36119), .A2(\pe6/phq [28]), .Z(n36122) );
  NAND2HSV0 U41126 ( .A1(n48051), .A2(n49208), .ZN(n58863) );
  XNOR2HSV1 U41127 ( .A1(n36122), .A2(n36121), .ZN(n36131) );
  CLKNHSV0 U41128 ( .I(n36127), .ZN(n36128) );
  XNOR2HSV1 U41129 ( .A1(n36129), .A2(n36128), .ZN(n36130) );
  XNOR2HSV1 U41130 ( .A1(n36131), .A2(n36130), .ZN(n36141) );
  NOR2HSV0 U41131 ( .A1(n36132), .A2(n49188), .ZN(n36134) );
  NAND2HSV0 U41132 ( .A1(n46627), .A2(n58378), .ZN(n36133) );
  XOR2HSV0 U41133 ( .A1(n36134), .A2(n36133), .Z(n36138) );
  NAND2HSV0 U41134 ( .A1(n46658), .A2(\pe6/aot [6]), .ZN(n36136) );
  NAND2HSV0 U41135 ( .A1(n58628), .A2(n59065), .ZN(n36135) );
  XOR2HSV0 U41136 ( .A1(n36136), .A2(n36135), .Z(n36137) );
  XOR2HSV0 U41137 ( .A1(n36138), .A2(n36137), .Z(n36140) );
  NAND2HSV0 U41138 ( .A1(n44426), .A2(n58399), .ZN(n36139) );
  XOR4HSV1 U41139 ( .A1(n36142), .A2(n36141), .A3(n36140), .A4(n36139), .Z(
        n36178) );
  NAND2HSV0 U41140 ( .A1(n36143), .A2(n58749), .ZN(n36145) );
  NAND2HSV0 U41141 ( .A1(n44435), .A2(\pe6/aot [15]), .ZN(n36144) );
  XOR2HSV0 U41142 ( .A1(n36145), .A2(n36144), .Z(n36149) );
  NAND2HSV0 U41143 ( .A1(n58682), .A2(n33004), .ZN(n36147) );
  NAND2HSV0 U41144 ( .A1(n59098), .A2(\pe6/aot [17]), .ZN(n36146) );
  XOR2HSV0 U41145 ( .A1(n36147), .A2(n36146), .Z(n36148) );
  XOR2HSV0 U41146 ( .A1(n36149), .A2(n36148), .Z(n36159) );
  NAND2HSV0 U41147 ( .A1(n36150), .A2(\pe6/aot [19]), .ZN(n36152) );
  NAND2HSV0 U41148 ( .A1(n58965), .A2(n58488), .ZN(n36151) );
  XOR2HSV0 U41149 ( .A1(n36152), .A2(n36151), .Z(n36157) );
  NAND2HSV0 U41150 ( .A1(n32982), .A2(n44439), .ZN(n36155) );
  NAND2HSV0 U41151 ( .A1(n58668), .A2(n36153), .ZN(n36154) );
  XOR2HSV0 U41152 ( .A1(n36155), .A2(n36154), .Z(n36156) );
  XOR2HSV0 U41153 ( .A1(n36157), .A2(n36156), .Z(n36158) );
  XOR2HSV0 U41154 ( .A1(n36159), .A2(n36158), .Z(n36176) );
  NAND2HSV0 U41155 ( .A1(n49862), .A2(n59044), .ZN(n49324) );
  XOR2HSV0 U41156 ( .A1(n36160), .A2(n49324), .Z(n36165) );
  NAND2HSV0 U41157 ( .A1(n36161), .A2(\pe6/pvq [28]), .ZN(n36162) );
  XOR2HSV0 U41158 ( .A1(n36163), .A2(n36162), .Z(n36164) );
  XOR2HSV0 U41159 ( .A1(n36165), .A2(n36164), .Z(n36174) );
  NAND2HSV0 U41160 ( .A1(n46672), .A2(n46792), .ZN(n36167) );
  NAND2HSV0 U41161 ( .A1(n59246), .A2(n59234), .ZN(n36166) );
  XOR2HSV0 U41162 ( .A1(n36167), .A2(n36166), .Z(n36172) );
  NAND2HSV0 U41163 ( .A1(n36168), .A2(\pe6/aot [21]), .ZN(n36170) );
  NAND2HSV0 U41164 ( .A1(n58962), .A2(n32981), .ZN(n36169) );
  XOR2HSV0 U41165 ( .A1(n36170), .A2(n36169), .Z(n36171) );
  XOR2HSV0 U41166 ( .A1(n36172), .A2(n36171), .Z(n36173) );
  XOR2HSV0 U41167 ( .A1(n36174), .A2(n36173), .Z(n36175) );
  XOR2HSV0 U41168 ( .A1(n36176), .A2(n36175), .Z(n36177) );
  XNOR2HSV1 U41169 ( .A1(n36178), .A2(n36177), .ZN(n36179) );
  XNOR2HSV1 U41170 ( .A1(n36180), .A2(n36179), .ZN(n36182) );
  NAND2HSV0 U41171 ( .A1(n32900), .A2(n58525), .ZN(n36181) );
  XOR2HSV0 U41172 ( .A1(n36182), .A2(n36181), .Z(n36184) );
  CLKNAND2HSV0 U41173 ( .A1(n59317), .A2(n59176), .ZN(n36186) );
  XOR2HSV0 U41174 ( .A1(n36187), .A2(n36186), .Z(n36189) );
  CLKNAND2HSV0 U41175 ( .A1(n59676), .A2(\pe6/got [21]), .ZN(n36188) );
  XOR2HSV0 U41176 ( .A1(n36189), .A2(n36188), .Z(n36190) );
  XNOR2HSV1 U41177 ( .A1(n36191), .A2(n36190), .ZN(n36192) );
  XNOR2HSV1 U41178 ( .A1(n36193), .A2(n36192), .ZN(n36194) );
  XNOR2HSV1 U41179 ( .A1(n36195), .A2(n36194), .ZN(n36198) );
  CLKNAND2HSV0 U41180 ( .A1(n36196), .A2(\pe6/got [25]), .ZN(n36197) );
  XNOR2HSV1 U41181 ( .A1(n36198), .A2(n36197), .ZN(n36199) );
  XOR2HSV2 U41182 ( .A1(n36200), .A2(n36199), .Z(n36201) );
  XNOR2HSV4 U41183 ( .A1(n36202), .A2(n36201), .ZN(n36204) );
  NOR2HSV1 U41184 ( .A1(n44362), .A2(n46824), .ZN(n36213) );
  XOR3HSV2 U41185 ( .A1(n46760), .A2(n36205), .A3(n36204), .Z(n36211) );
  CLKNHSV2 U41186 ( .I(n36206), .ZN(n36209) );
  CLKNHSV0 U41187 ( .I(n36207), .ZN(n36208) );
  NOR2HSV4 U41188 ( .A1(n36209), .A2(n36208), .ZN(n36210) );
  NOR2HSV4 U41189 ( .A1(n36211), .A2(n36210), .ZN(n36212) );
  NOR2HSV2 U41190 ( .A1(n36213), .A2(n36212), .ZN(n36219) );
  NOR2HSV0 U41191 ( .A1(n36214), .A2(n32651), .ZN(n36215) );
  CLKAND2HSV2 U41192 ( .A1(n36216), .A2(n36215), .Z(n36217) );
  CLKNAND2HSV3 U41193 ( .A1(n36218), .A2(n36217), .ZN(n44365) );
  XNOR2HSV4 U41194 ( .A1(n36221), .A2(n36220), .ZN(n47933) );
  CLKNAND2HSV3 U41195 ( .A1(n36223), .A2(n29727), .ZN(n46144) );
  INHSV4 U41196 ( .I(n46144), .ZN(n36236) );
  XNOR2HSV4 U41197 ( .A1(n36225), .A2(n36224), .ZN(n46569) );
  INHSV2 U41198 ( .I(n46569), .ZN(n36228) );
  NAND2HSV2 U41199 ( .A1(n36228), .A2(n46574), .ZN(n36227) );
  INHSV1 U41200 ( .I(n44692), .ZN(n36226) );
  CLKNAND2HSV2 U41201 ( .A1(n36227), .A2(n36226), .ZN(n36233) );
  CLKNAND2HSV1 U41202 ( .A1(n36228), .A2(n44692), .ZN(n36232) );
  NAND2HSV0 U41203 ( .A1(n46569), .A2(n36229), .ZN(n36230) );
  CLKNAND2HSV1 U41204 ( .A1(n36230), .A2(n44519), .ZN(n36231) );
  AOI21HSV4 U41205 ( .A1(n36233), .A2(n36232), .B(n36231), .ZN(n36234) );
  CLKNAND2HSV4 U41206 ( .A1(n36236), .A2(n46151), .ZN(n59570) );
  INHSV4 U41207 ( .I(\pe2/aot [30]), .ZN(n38404) );
  INHSV4 U41208 ( .I(n38404), .ZN(n36604) );
  CLKNHSV2 U41209 ( .I(\pe2/bq[31] ), .ZN(n36237) );
  INHSV4 U41210 ( .I(n36237), .ZN(n36385) );
  NAND2HSV2 U41211 ( .A1(n36604), .A2(n36385), .ZN(n36239) );
  CLKBUFHSV4 U41212 ( .I(n36458), .Z(n36553) );
  INHSV4 U41213 ( .I(n36350), .ZN(n45008) );
  NAND2HSV2 U41214 ( .A1(n36377), .A2(n45008), .ZN(n36238) );
  CLKXOR2HSV4 U41215 ( .A1(n36239), .A2(n36238), .Z(n36244) );
  INHSV2 U41216 ( .I(n38787), .ZN(n52941) );
  CLKNHSV4 U41217 ( .I(\pe2/bq[32] ), .ZN(n38418) );
  NAND2HSV2 U41218 ( .A1(n52941), .A2(n36590), .ZN(n36242) );
  INHSV4 U41219 ( .I(n36240), .ZN(n36433) );
  NOR2HSV2 U41220 ( .A1(n36240), .A2(n36389), .ZN(n36241) );
  XOR2HSV2 U41221 ( .A1(n36242), .A2(n36241), .Z(n36243) );
  XNOR2HSV4 U41222 ( .A1(n36244), .A2(n36243), .ZN(n36248) );
  NAND2HSV2 U41223 ( .A1(n37952), .A2(\pe2/pvq [4]), .ZN(n36245) );
  XNOR2HSV1 U41224 ( .A1(n36245), .A2(\pe2/phq [4]), .ZN(n36247) );
  INHSV2 U41225 ( .I(\pe2/aot [31]), .ZN(n36274) );
  BUFHSV2 U41226 ( .I(n36274), .Z(n44889) );
  INHSV4 U41227 ( .I(\pe2/bq[30] ), .ZN(n36294) );
  BUFHSV4 U41228 ( .I(n36294), .Z(n36388) );
  BUFHSV8 U41229 ( .I(n36388), .Z(n38823) );
  NOR2HSV2 U41230 ( .A1(n44889), .A2(n38823), .ZN(n36246) );
  XNOR2HSV4 U41231 ( .A1(n36248), .A2(n29687), .ZN(n36264) );
  BUFHSV8 U41232 ( .I(n36350), .Z(n36443) );
  INHSV2 U41233 ( .I(\pe2/phq [1]), .ZN(n36249) );
  INHSV6 U41234 ( .I(\pe2/got [32]), .ZN(n36665) );
  INHSV4 U41235 ( .I(n36260), .ZN(n36257) );
  CLKNAND2HSV1 U41236 ( .A1(\pe2/bq[32] ), .A2(\pe2/aot [32]), .ZN(n36255) );
  INHSV4 U41237 ( .I(\pe2/ctrq ), .ZN(n44884) );
  NOR2HSV2 U41238 ( .A1(n36240), .A2(n44884), .ZN(n36254) );
  CLKNHSV2 U41239 ( .I(\pe2/bq[32] ), .ZN(n36251) );
  NOR2HSV4 U41240 ( .A1(n36252), .A2(n36251), .ZN(n36253) );
  AOI22HSV4 U41241 ( .A1(n36255), .A2(n36252), .B1(n36254), .B2(n36253), .ZN(
        n36259) );
  CLKNAND2HSV2 U41242 ( .A1(n36255), .A2(n44884), .ZN(n36258) );
  CLKNAND2HSV2 U41243 ( .A1(n36259), .A2(n36258), .ZN(n36256) );
  NAND2HSV4 U41244 ( .A1(n36257), .A2(n36256), .ZN(n36362) );
  CLKBUFHSV4 U41245 ( .I(ctro2), .Z(n36574) );
  CLKAND2HSV2 U41246 ( .A1(n36574), .A2(\pe2/ti_7t [1]), .Z(n36365) );
  INHSV2 U41247 ( .I(n36365), .ZN(n36261) );
  NAND3HSV4 U41248 ( .A1(n36362), .A2(n36363), .A3(n36261), .ZN(n36263) );
  BUFHSV2 U41249 ( .I(n38899), .Z(n37931) );
  NAND2HSV2 U41250 ( .A1(n36261), .A2(n38099), .ZN(n36262) );
  CLKNAND2HSV4 U41251 ( .A1(n36263), .A2(n36262), .ZN(n36299) );
  INHSV2 U41252 ( .I(n38733), .ZN(n38742) );
  INHSV2 U41253 ( .I(n38742), .ZN(n38738) );
  NOR2HSV4 U41254 ( .A1(n36376), .A2(n38738), .ZN(n36265) );
  NAND2HSV2 U41255 ( .A1(n36264), .A2(n36265), .ZN(n36268) );
  INHSV3 U41256 ( .I(n36264), .ZN(n36267) );
  INHSV2 U41257 ( .I(n36265), .ZN(n36266) );
  INHSV4 U41258 ( .I(n36341), .ZN(n36310) );
  BUFHSV2 U41259 ( .I(n36350), .Z(n38126) );
  NOR2HSV4 U41260 ( .A1(n36319), .A2(n38126), .ZN(n36273) );
  NAND2HSV4 U41261 ( .A1(\pe2/aot [32]), .A2(\pe2/bq[31] ), .ZN(n36271) );
  INHSV4 U41262 ( .I(\pe2/phq [2]), .ZN(n36270) );
  XNOR2HSV4 U41263 ( .A1(n36271), .A2(n36270), .ZN(n36272) );
  XNOR2HSV4 U41264 ( .A1(n36273), .A2(n36272), .ZN(n36305) );
  NAND2HSV2 U41265 ( .A1(n36380), .A2(\pe2/pvq [2]), .ZN(n36276) );
  INHSV3 U41266 ( .I(n36274), .ZN(n52449) );
  XOR2HSV2 U41267 ( .A1(n36276), .A2(n36275), .Z(n36304) );
  XNOR2HSV4 U41268 ( .A1(n36305), .A2(n36304), .ZN(n36281) );
  CLKNHSV6 U41269 ( .I(n36281), .ZN(n36408) );
  BUFHSV2 U41270 ( .I(n36665), .Z(n37871) );
  BUFHSV2 U41271 ( .I(n38899), .Z(n38195) );
  INHSV2 U41272 ( .I(n38335), .ZN(n45409) );
  NAND3HSV2 U41273 ( .A1(n36310), .A2(n36408), .A3(n45409), .ZN(n36280) );
  NOR2HSV2 U41274 ( .A1(n36408), .A2(n36277), .ZN(n36402) );
  BUFHSV2 U41275 ( .I(n38899), .Z(n38272) );
  INHSV2 U41276 ( .I(n38272), .ZN(n36473) );
  NOR2HSV2 U41277 ( .A1(n36473), .A2(\pe2/ti_7t [2]), .ZN(n36403) );
  OR2HSV1 U41278 ( .A1(n36403), .A2(n45267), .Z(n36278) );
  NOR2HSV2 U41279 ( .A1(n36402), .A2(n36278), .ZN(n36279) );
  CLKNHSV2 U41280 ( .I(n36287), .ZN(n36284) );
  INHSV2 U41281 ( .I(n36376), .ZN(n52981) );
  INAND2HSV2 U41282 ( .A1(n38886), .B1(n36281), .ZN(n36282) );
  NOR2HSV4 U41283 ( .A1(n52981), .A2(n36282), .ZN(n36406) );
  NAND3HSV4 U41284 ( .A1(n36284), .A2(n36285), .A3(n36283), .ZN(n36289) );
  INHSV4 U41285 ( .I(n36285), .ZN(n36286) );
  OAI21HSV4 U41286 ( .A1(n36287), .A2(n25871), .B(n36286), .ZN(n36288) );
  NAND2HSV4 U41287 ( .A1(n36289), .A2(n36288), .ZN(n36430) );
  NAND2HSV2 U41288 ( .A1(\pe2/bq[31] ), .A2(\pe2/aot [31]), .ZN(n36291) );
  CLKAND2HSV4 U41289 ( .A1(\pe2/bq[32] ), .A2(\pe2/aot [30]), .Z(n36290) );
  BUFHSV4 U41290 ( .I(\pe2/ctrq ), .Z(n46623) );
  NAND2HSV2 U41291 ( .A1(n46623), .A2(\pe2/pvq [3]), .ZN(n36292) );
  INHSV1 U41292 ( .I(\pe2/phq [3]), .ZN(n36293) );
  BUFHSV8 U41293 ( .I(n36294), .Z(n36296) );
  OAI21HSV4 U41294 ( .A1(n36296), .A2(n36240), .B(\pe2/phq [3]), .ZN(n36295)
         );
  XNOR2HSV4 U41295 ( .A1(n36300), .A2(n36301), .ZN(n36317) );
  INHSV4 U41296 ( .I(n36317), .ZN(n36321) );
  INHSV2 U41297 ( .I(\pe2/got [31]), .ZN(n38523) );
  CLKNHSV0 U41298 ( .I(n38523), .ZN(n53094) );
  CLKNAND2HSV2 U41299 ( .A1(n36321), .A2(n53094), .ZN(n36298) );
  INHSV2 U41300 ( .I(n36298), .ZN(n36303) );
  BUFHSV2 U41301 ( .I(n36574), .Z(n38099) );
  AOI21HSV4 U41302 ( .A1(n36303), .A2(n52981), .B(n36302), .ZN(n36328) );
  XNOR2HSV4 U41303 ( .A1(n36305), .A2(n36304), .ZN(n36368) );
  INHSV4 U41304 ( .I(n36368), .ZN(n36306) );
  NOR2HSV4 U41305 ( .A1(n36306), .A2(n38886), .ZN(n36308) );
  BUFHSV2 U41306 ( .I(n37871), .Z(n45130) );
  OR2HSV1 U41307 ( .A1(n36403), .A2(n45130), .Z(n36307) );
  AOI21HSV4 U41308 ( .A1(n36308), .A2(n36341), .B(n36307), .ZN(n36314) );
  CLKNAND2HSV4 U41309 ( .A1(n36408), .A2(n45265), .ZN(n36309) );
  NAND2HSV4 U41310 ( .A1(n36314), .A2(n36313), .ZN(n36312) );
  INHSV6 U41311 ( .I(n36312), .ZN(n53375) );
  CLKNAND2HSV2 U41312 ( .A1(n36328), .A2(n53375), .ZN(n36325) );
  NAND2HSV4 U41313 ( .A1(n36314), .A2(n36313), .ZN(n36330) );
  INHSV2 U41314 ( .I(n38523), .ZN(n38603) );
  CLKNAND2HSV1 U41315 ( .A1(n38264), .A2(n38108), .ZN(n36316) );
  NOR2HSV2 U41316 ( .A1(n36331), .A2(n36316), .ZN(n36322) );
  INHSV2 U41317 ( .I(n36317), .ZN(n53374) );
  BUFHSV2 U41318 ( .I(n36376), .Z(n36318) );
  NAND2HSV4 U41319 ( .A1(n53374), .A2(n36318), .ZN(n36332) );
  NOR2HSV4 U41320 ( .A1(n36587), .A2(n36320), .ZN(n53373) );
  INAND2HSV4 U41321 ( .A1(n36321), .B1(n53373), .ZN(n36329) );
  NAND4HSV4 U41322 ( .A1(n36330), .A2(n36322), .A3(n36332), .A4(n36329), .ZN(
        n36324) );
  BUFHSV2 U41323 ( .I(n36560), .Z(n38344) );
  NAND2HSV2 U41324 ( .A1(n38344), .A2(\pe2/ti_7t [3]), .ZN(n36326) );
  OR2HSV1 U41325 ( .A1(n36326), .A2(n38013), .Z(n36323) );
  XNOR2HSV4 U41326 ( .A1(n36430), .A2(n36429), .ZN(n59509) );
  INHSV1 U41327 ( .I(n37931), .ZN(n38627) );
  NAND2HSV2 U41328 ( .A1(n38454), .A2(\pe2/ti_7t [4]), .ZN(n36501) );
  INHSV2 U41329 ( .I(\pe2/got [27]), .ZN(n36493) );
  CLKBUFHSV4 U41330 ( .I(n36493), .Z(n38472) );
  BUFHSV2 U41331 ( .I(n38472), .Z(n38902) );
  CLKNAND2HSV0 U41332 ( .A1(n44906), .A2(\pe2/got [27]), .ZN(n36375) );
  INHSV2 U41333 ( .I(n36326), .ZN(n36327) );
  AOI21HSV4 U41334 ( .A1(n36328), .A2(n53375), .B(n36327), .ZN(n36413) );
  CLKAND2HSV4 U41335 ( .A1(n36330), .A2(n36329), .Z(n36335) );
  CLKAND2HSV4 U41336 ( .A1(n36333), .A2(n36332), .Z(n36334) );
  INHSV2 U41337 ( .I(n38042), .ZN(n49492) );
  NAND2HSV2 U41338 ( .A1(n36619), .A2(n49492), .ZN(n36361) );
  CLKNHSV0 U41339 ( .I(n38404), .ZN(n38055) );
  CLKNAND2HSV1 U41340 ( .A1(n38055), .A2(n44987), .ZN(n36340) );
  BUFHSV2 U41341 ( .I(n37952), .Z(n48078) );
  INHSV4 U41342 ( .I(n38787), .ZN(n37792) );
  CLKNAND2HSV0 U41343 ( .A1(n37792), .A2(n38064), .ZN(n36337) );
  INHSV2 U41344 ( .I(n44049), .ZN(n59970) );
  NAND2HSV0 U41345 ( .A1(n59970), .A2(n36608), .ZN(n36336) );
  XOR2HSV0 U41346 ( .A1(n36337), .A2(n36336), .Z(n36338) );
  XOR3HSV2 U41347 ( .A1(n36340), .A2(n36339), .A3(n36338), .Z(n36359) );
  INHSV2 U41348 ( .I(n36341), .ZN(n43950) );
  NAND2HSV2 U41349 ( .A1(n43950), .A2(n59584), .ZN(n36358) );
  INHSV2 U41350 ( .I(\pe2/aot [25]), .ZN(n38664) );
  CLKNAND2HSV0 U41351 ( .A1(n38048), .A2(n38043), .ZN(n36343) );
  CLKNAND2HSV0 U41352 ( .A1(n59972), .A2(n36607), .ZN(n36342) );
  XOR2HSV0 U41353 ( .A1(n36343), .A2(n36342), .Z(n36347) );
  CLKNAND2HSV0 U41354 ( .A1(n50930), .A2(n36590), .ZN(n36345) );
  INHSV2 U41355 ( .I(n36240), .ZN(n59582) );
  CLKNAND2HSV0 U41356 ( .A1(n59582), .A2(\pe2/bq[23] ), .ZN(n36344) );
  XOR2HSV0 U41357 ( .A1(n36345), .A2(n36344), .Z(n36346) );
  XOR2HSV0 U41358 ( .A1(n36347), .A2(n36346), .Z(n36356) );
  CLKNAND2HSV0 U41359 ( .A1(n52310), .A2(n36588), .ZN(n36349) );
  INHSV2 U41360 ( .I(n44212), .ZN(n36589) );
  CLKNAND2HSV0 U41361 ( .A1(n36589), .A2(n38394), .ZN(n36348) );
  XOR2HSV0 U41362 ( .A1(n36349), .A2(n36348), .Z(n36354) );
  INHSV2 U41363 ( .I(\pe2/aot [31]), .ZN(n37941) );
  CLKNHSV0 U41364 ( .I(n37941), .ZN(n38061) );
  CLKNAND2HSV1 U41365 ( .A1(n38061), .A2(n38053), .ZN(n36352) );
  INHSV2 U41366 ( .I(n38275), .ZN(n38080) );
  BUFHSV2 U41367 ( .I(n36350), .Z(n38213) );
  CLKNAND2HSV0 U41368 ( .A1(n38080), .A2(n38401), .ZN(n36351) );
  XOR2HSV0 U41369 ( .A1(n36352), .A2(n36351), .Z(n36353) );
  XOR2HSV0 U41370 ( .A1(n36354), .A2(n36353), .Z(n36355) );
  XOR2HSV0 U41371 ( .A1(n36356), .A2(n36355), .Z(n36357) );
  XOR3HSV2 U41372 ( .A1(n36359), .A2(n36358), .A3(n36357), .Z(n36360) );
  XNOR2HSV1 U41373 ( .A1(n36361), .A2(n36360), .ZN(n36373) );
  CLKAND2HSV0 U41374 ( .A1(n38264), .A2(n45265), .Z(n36364) );
  NAND2HSV2 U41375 ( .A1(n60102), .A2(n36364), .ZN(n36367) );
  NAND2HSV0 U41376 ( .A1(n36365), .A2(n36250), .ZN(n36366) );
  NAND2HSV2 U41377 ( .A1(n36367), .A2(n36366), .ZN(n36369) );
  XNOR2HSV4 U41378 ( .A1(n36369), .A2(n36368), .ZN(n60003) );
  NAND2HSV2 U41379 ( .A1(n60003), .A2(n36654), .ZN(n36371) );
  CLKNAND2HSV0 U41380 ( .A1(n38886), .A2(\pe2/ti_7t [2]), .ZN(n36370) );
  CLKNAND2HSV1 U41381 ( .A1(n36614), .A2(n38324), .ZN(n36372) );
  XNOR2HSV1 U41382 ( .A1(n36373), .A2(n36372), .ZN(n36374) );
  XNOR2HSV1 U41383 ( .A1(n36375), .A2(n36374), .ZN(n36428) );
  INHSV2 U41384 ( .I(n36376), .ZN(n36396) );
  INHSV4 U41385 ( .I(n36396), .ZN(n38907) );
  INHSV2 U41386 ( .I(n36377), .ZN(n36397) );
  NOR2HSV2 U41387 ( .A1(n45411), .A2(n38213), .ZN(n36379) );
  CLKNAND2HSV0 U41388 ( .A1(n59759), .A2(n36590), .ZN(n36378) );
  XOR2HSV2 U41389 ( .A1(n36379), .A2(n36378), .Z(n36384) );
  CLKNAND2HSV1 U41390 ( .A1(n36380), .A2(\pe2/pvq [5]), .ZN(n36382) );
  INHSV2 U41391 ( .I(\pe2/phq [5]), .ZN(n36381) );
  XOR2HSV0 U41392 ( .A1(n36382), .A2(n36381), .Z(n36383) );
  XNOR2HSV4 U41393 ( .A1(n36384), .A2(n36383), .ZN(n36394) );
  NAND2HSV2 U41394 ( .A1(n37792), .A2(n36385), .ZN(n36387) );
  NAND2HSV2 U41395 ( .A1(n36433), .A2(n36588), .ZN(n36386) );
  XOR2HSV0 U41396 ( .A1(n36387), .A2(n36386), .Z(n36392) );
  CLKNHSV2 U41397 ( .I(n38404), .ZN(n59969) );
  INHSV4 U41398 ( .I(n36388), .ZN(n36475) );
  NAND2HSV4 U41399 ( .A1(n59969), .A2(n36475), .ZN(n38671) );
  INHSV2 U41400 ( .I(n37941), .ZN(n44976) );
  INHSV4 U41401 ( .I(n36389), .ZN(n44759) );
  NAND2HSV2 U41402 ( .A1(n44976), .A2(n44759), .ZN(n36390) );
  CLKXOR2HSV2 U41403 ( .A1(n38671), .A2(n36390), .Z(n36391) );
  XOR2HSV2 U41404 ( .A1(n36392), .A2(n36391), .Z(n36393) );
  XNOR2HSV4 U41405 ( .A1(n36394), .A2(n36393), .ZN(n36399) );
  INHSV4 U41406 ( .I(n36399), .ZN(n36395) );
  OAI21HSV4 U41407 ( .A1(n38907), .A2(n36397), .B(n36395), .ZN(n36401) );
  INHSV4 U41408 ( .I(n36396), .ZN(n37876) );
  INHSV2 U41409 ( .I(n36402), .ZN(n36405) );
  INHSV2 U41410 ( .I(\pe2/got [30]), .ZN(n45091) );
  NOR2HSV0 U41411 ( .A1(n36403), .A2(n45091), .ZN(n36404) );
  BUFHSV8 U41412 ( .I(n36587), .Z(n44053) );
  CLKNAND2HSV2 U41413 ( .A1(n36409), .A2(n29703), .ZN(n36410) );
  XNOR2HSV4 U41414 ( .A1(n36421), .A2(n36422), .ZN(n52718) );
  CLKNAND2HSV4 U41415 ( .A1(n36413), .A2(n36412), .ZN(n36415) );
  INHSV2 U41416 ( .I(n38523), .ZN(n43919) );
  INHSV2 U41417 ( .I(n45267), .ZN(n36414) );
  INHSV2 U41418 ( .I(n38335), .ZN(n37846) );
  INHSV2 U41419 ( .I(n36416), .ZN(n36417) );
  INHSV2 U41420 ( .I(n36560), .ZN(n38183) );
  CLKAND2HSV2 U41421 ( .A1(n38184), .A2(\pe2/ti_7t [5]), .Z(n36419) );
  AOI21HSV4 U41422 ( .A1(n36420), .A2(n59509), .B(n36419), .ZN(n36470) );
  BUFHSV2 U41423 ( .I(n36665), .Z(n53098) );
  INHSV2 U41424 ( .I(n53098), .ZN(n52745) );
  NAND2HSV2 U41425 ( .A1(n59509), .A2(n52745), .ZN(n36426) );
  INHSV4 U41426 ( .I(n36421), .ZN(n36423) );
  XOR2HSV4 U41427 ( .A1(n36424), .A2(n52719), .Z(n36425) );
  NAND3HSV4 U41428 ( .A1(n36426), .A2(n36425), .A3(n38627), .ZN(n36471) );
  BUFHSV4 U41429 ( .I(n44780), .Z(n38841) );
  INHSV2 U41430 ( .I(n45411), .ZN(n52415) );
  BUFHSV2 U41431 ( .I(n38630), .Z(n38184) );
  INHSV2 U41432 ( .I(n38184), .ZN(n44041) );
  CLKNAND2HSV0 U41433 ( .A1(n36513), .A2(n44041), .ZN(n36511) );
  XNOR2HSV4 U41434 ( .A1(n36430), .A2(n36429), .ZN(n36504) );
  BUFHSV2 U41435 ( .I(n45267), .Z(n44831) );
  BUFHSV2 U41436 ( .I(n38195), .Z(n45129) );
  NOR2HSV2 U41437 ( .A1(n44831), .A2(n45129), .ZN(n45100) );
  INHSV2 U41438 ( .I(n45100), .ZN(n44314) );
  INHSV2 U41439 ( .I(n44314), .ZN(n36432) );
  NOR2HSV2 U41440 ( .A1(n36501), .A2(n45267), .ZN(n36431) );
  AOI21HSV4 U41441 ( .A1(n36504), .A2(n36432), .B(n36431), .ZN(n36466) );
  INHSV2 U41442 ( .I(n36466), .ZN(n36465) );
  INHSV2 U41443 ( .I(n38733), .ZN(n36661) );
  INHSV2 U41444 ( .I(n45411), .ZN(n36623) );
  INHSV2 U41445 ( .I(n36623), .ZN(n38993) );
  NOR2HSV4 U41446 ( .A1(n37876), .A2(n38993), .ZN(n36451) );
  INHSV2 U41447 ( .I(n37941), .ZN(n59968) );
  NAND2HSV2 U41448 ( .A1(n59968), .A2(n38565), .ZN(n36435) );
  XOR3HSV2 U41449 ( .A1(\pe2/phq [6]), .A2(n36436), .A3(n36435), .Z(n36440) );
  CLKNAND2HSV2 U41450 ( .A1(n38549), .A2(n49530), .ZN(n36438) );
  NAND2HSV2 U41451 ( .A1(n36380), .A2(\pe2/pvq [6]), .ZN(n36437) );
  XNOR2HSV4 U41452 ( .A1(n36438), .A2(n36437), .ZN(n36439) );
  XNOR2HSV4 U41453 ( .A1(n36440), .A2(n36439), .ZN(n36449) );
  NOR2HSV4 U41454 ( .A1(n37940), .A2(n37953), .ZN(n36441) );
  XOR2HSV2 U41455 ( .A1(n36442), .A2(n36441), .Z(n36447) );
  INAND2HSV2 U41456 ( .A1(n38404), .B1(n44759), .ZN(n36445) );
  XNOR2HSV4 U41457 ( .A1(n36445), .A2(n36444), .ZN(n36446) );
  XNOR2HSV4 U41458 ( .A1(n36447), .A2(n36446), .ZN(n36448) );
  XNOR2HSV4 U41459 ( .A1(n36449), .A2(n36448), .ZN(n36452) );
  CLKNHSV2 U41460 ( .I(n36452), .ZN(n36450) );
  INHSV2 U41461 ( .I(n36451), .ZN(n36453) );
  NAND2HSV2 U41462 ( .A1(n36453), .A2(n36452), .ZN(n36454) );
  NAND2HSV4 U41463 ( .A1(n36455), .A2(n36454), .ZN(n36461) );
  INHSV2 U41464 ( .I(\pe2/ti_7t [2]), .ZN(n36456) );
  NOR2HSV2 U41465 ( .A1(n44041), .A2(n36456), .ZN(n36457) );
  AOI21HSV4 U41466 ( .A1(n60003), .A2(n44041), .B(n36457), .ZN(n36496) );
  BUFHSV2 U41467 ( .I(n36458), .Z(n44184) );
  INHSV2 U41468 ( .I(n44145), .ZN(n38644) );
  NOR2HSV4 U41469 ( .A1(n36496), .A2(n38644), .ZN(n36460) );
  NOR2HSV4 U41470 ( .A1(n36461), .A2(n36460), .ZN(n36459) );
  AOI21HSV4 U41471 ( .A1(n36461), .A2(n36460), .B(n36459), .ZN(n36462) );
  XNOR2HSV4 U41472 ( .A1(n36463), .A2(n36462), .ZN(n36467) );
  INHSV3 U41473 ( .I(n36467), .ZN(n36464) );
  CLKNAND2HSV3 U41474 ( .A1(n36465), .A2(n36464), .ZN(n36469) );
  INHSV2 U41475 ( .I(n36560), .ZN(n38383) );
  NAND3HSV2 U41476 ( .A1(n36631), .A2(n44780), .A3(n38383), .ZN(n36528) );
  INHSV2 U41477 ( .I(n36528), .ZN(n36642) );
  CLKNAND2HSV3 U41478 ( .A1(n36472), .A2(n36630), .ZN(n36645) );
  NOR2HSV2 U41479 ( .A1(n36473), .A2(\pe2/ti_7t [6]), .ZN(n36632) );
  NOR2HSV2 U41480 ( .A1(n36632), .A2(n36519), .ZN(n36640) );
  CLKNAND2HSV0 U41481 ( .A1(n36645), .A2(n36640), .ZN(n36474) );
  NOR2HSV2 U41482 ( .A1(n36474), .A2(n36642), .ZN(n36507) );
  NAND2HSV4 U41483 ( .A1(n36557), .A2(n38026), .ZN(n36638) );
  NAND2HSV2 U41484 ( .A1(n36604), .A2(\pe2/bq[28] ), .ZN(n36477) );
  NAND2HSV2 U41485 ( .A1(n36589), .A2(n36475), .ZN(n36476) );
  CLKNAND2HSV2 U41486 ( .A1(n37952), .A2(\pe2/pvq [7]), .ZN(n36478) );
  XNOR2HSV4 U41487 ( .A1(n36478), .A2(\pe2/phq [7]), .ZN(n36479) );
  CLKNHSV2 U41488 ( .I(n38126), .ZN(n36602) );
  CLKNAND2HSV0 U41489 ( .A1(n36602), .A2(n49492), .ZN(n36481) );
  XNOR2HSV4 U41490 ( .A1(n36482), .A2(n36481), .ZN(n36483) );
  XNOR2HSV4 U41491 ( .A1(n36484), .A2(n36483), .ZN(n36492) );
  NAND2HSV2 U41492 ( .A1(n36603), .A2(n38047), .ZN(n36486) );
  INHSV2 U41493 ( .I(n38787), .ZN(n52485) );
  CLKNAND2HSV1 U41494 ( .A1(n52485), .A2(n36608), .ZN(n36485) );
  XOR2HSV0 U41495 ( .A1(n36486), .A2(n36485), .Z(n36490) );
  NAND2HSV2 U41496 ( .A1(n59582), .A2(\pe2/bq[26] ), .ZN(n36488) );
  CLKNAND2HSV1 U41497 ( .A1(\pe2/aot [26]), .A2(n36590), .ZN(n36487) );
  XOR2HSV0 U41498 ( .A1(n36488), .A2(n36487), .Z(n36489) );
  XNOR2HSV1 U41499 ( .A1(n36490), .A2(n36489), .ZN(n36491) );
  XNOR2HSV4 U41500 ( .A1(n36492), .A2(n36491), .ZN(n36495) );
  BUFHSV2 U41501 ( .I(n36493), .Z(n44969) );
  XNOR2HSV4 U41502 ( .A1(n36495), .A2(n36494), .ZN(n36498) );
  NOR2HSV2 U41503 ( .A1(n36496), .A2(n38163), .ZN(n36497) );
  CLKXOR2HSV4 U41504 ( .A1(n36498), .A2(n36497), .Z(n36500) );
  NAND2HSV2 U41505 ( .A1(n36619), .A2(n36377), .ZN(n36499) );
  XNOR2HSV4 U41506 ( .A1(n36500), .A2(n36499), .ZN(n36506) );
  BUFHSV2 U41507 ( .I(n38733), .Z(n45281) );
  NOR2HSV1 U41508 ( .A1(n45281), .A2(n36560), .ZN(n36503) );
  NOR2HSV1 U41509 ( .A1(n36501), .A2(n38514), .ZN(n36502) );
  AOI21HSV4 U41510 ( .A1(n36504), .A2(n36503), .B(n36502), .ZN(n36505) );
  XNOR2HSV4 U41511 ( .A1(n36506), .A2(n36505), .ZN(n36639) );
  XNOR2HSV4 U41512 ( .A1(n36507), .A2(n36647), .ZN(n60005) );
  INHSV2 U41513 ( .I(\pe2/ti_7t [7]), .ZN(n36508) );
  BUFHSV2 U41514 ( .I(n38272), .Z(n38529) );
  NAND2HSV2 U41515 ( .A1(n36508), .A2(n38529), .ZN(n37827) );
  CLKNAND2HSV1 U41516 ( .A1(n37827), .A2(n36661), .ZN(n36512) );
  OR2HSV1 U41517 ( .A1(n36512), .A2(n44041), .Z(n36515) );
  MUX2NHSV1 U41518 ( .I0(n36515), .I1(n36514), .S(n36513), .ZN(n36516) );
  NOR2HSV4 U41519 ( .A1(n36517), .A2(n36516), .ZN(n36522) );
  CLKNAND2HSV2 U41520 ( .A1(n44780), .A2(n52745), .ZN(n36629) );
  NOR2HSV2 U41521 ( .A1(n36630), .A2(n38529), .ZN(n36518) );
  NOR2HSV1 U41522 ( .A1(n45129), .A2(n36519), .ZN(n36521) );
  CLKNHSV0 U41523 ( .I(n48896), .ZN(n38119) );
  XNOR2HSV4 U41524 ( .A1(n36522), .A2(n29673), .ZN(n36581) );
  CLKNAND2HSV1 U41525 ( .A1(n37827), .A2(n47997), .ZN(n36561) );
  INHSV2 U41526 ( .I(n36640), .ZN(n36526) );
  NOR2HSV1 U41527 ( .A1(n36526), .A2(n45129), .ZN(n36527) );
  NAND3HSV2 U41528 ( .A1(n36528), .A2(n36645), .A3(n36527), .ZN(n36529) );
  NOR2HSV4 U41529 ( .A1(n36529), .A2(n36647), .ZN(n36635) );
  NOR2HSV4 U41530 ( .A1(n36573), .A2(n36635), .ZN(n36578) );
  INHSV3 U41531 ( .I(n36614), .ZN(n44971) );
  NOR2HSV2 U41532 ( .A1(n44971), .A2(n44969), .ZN(n36550) );
  NAND2HSV2 U41533 ( .A1(n59970), .A2(n36607), .ZN(n36532) );
  NAND2HSV2 U41534 ( .A1(n36604), .A2(n38394), .ZN(n36531) );
  XOR2HSV0 U41535 ( .A1(n36532), .A2(n36531), .Z(n36536) );
  NAND2HSV2 U41536 ( .A1(n52310), .A2(n39020), .ZN(n36534) );
  CLKNAND2HSV1 U41537 ( .A1(n52485), .A2(n36588), .ZN(n36533) );
  XOR2HSV0 U41538 ( .A1(n36534), .A2(n36533), .Z(n36535) );
  XOR2HSV0 U41539 ( .A1(n36536), .A2(n36535), .Z(n36548) );
  INHSV2 U41540 ( .I(n49492), .ZN(n52164) );
  NOR2HSV4 U41541 ( .A1(n37876), .A2(n52164), .ZN(n36537) );
  NAND2HSV2 U41542 ( .A1(n59582), .A2(\pe2/bq[25] ), .ZN(n36539) );
  CLKNAND2HSV1 U41543 ( .A1(n36589), .A2(n36608), .ZN(n36538) );
  XOR2HSV0 U41544 ( .A1(n36539), .A2(n36538), .Z(n36543) );
  INHSV4 U41545 ( .I(\pe2/aot [25]), .ZN(n48934) );
  NAND2HSV2 U41546 ( .A1(n52998), .A2(n36590), .ZN(n36541) );
  CLKNAND2HSV0 U41547 ( .A1(\pe2/got [25]), .A2(n36602), .ZN(n36540) );
  XOR2HSV0 U41548 ( .A1(n36541), .A2(n36540), .Z(n36542) );
  BUFHSV2 U41549 ( .I(n37952), .Z(n45811) );
  XNOR2HSV1 U41550 ( .A1(n36545), .A2(n36544), .ZN(n36546) );
  XOR3HSV2 U41551 ( .A1(n36548), .A2(n36547), .A3(n36546), .Z(n36549) );
  XNOR2HSV1 U41552 ( .A1(n36550), .A2(n36549), .ZN(n36552) );
  BUFHSV4 U41553 ( .I(n36619), .Z(n38081) );
  NAND2HSV2 U41554 ( .A1(n38081), .A2(n36623), .ZN(n36551) );
  XNOR2HSV4 U41555 ( .A1(n36552), .A2(n36551), .ZN(n36555) );
  INHSV2 U41556 ( .I(n36555), .ZN(n36556) );
  INHSV2 U41557 ( .I(n36553), .ZN(n52916) );
  NAND2HSV2 U41558 ( .A1(n44906), .A2(n52916), .ZN(n36554) );
  MUX2NHSV2 U41559 ( .I0(n36556), .I1(n36555), .S(n36554), .ZN(n36559) );
  XNOR2HSV4 U41560 ( .A1(n36559), .A2(n36558), .ZN(n36577) );
  NOR2HSV1 U41561 ( .A1(n44827), .A2(n45129), .ZN(n36565) );
  CLKNAND2HSV3 U41562 ( .A1(n36578), .A2(n29678), .ZN(n36656) );
  AND2HSV2 U41563 ( .A1(n36560), .A2(\pe2/ti_7t [8]), .Z(n36568) );
  OR2HSV1 U41564 ( .A1(n36561), .A2(n36568), .Z(n36564) );
  INOR2HSV0 U41565 ( .A1(n36564), .B1(n37846), .ZN(n36566) );
  INHSV2 U41566 ( .I(n36568), .ZN(n36569) );
  NAND2HSV2 U41567 ( .A1(n36570), .A2(n36569), .ZN(n36571) );
  INHSV1 U41568 ( .I(n38523), .ZN(n38340) );
  XNOR2HSV4 U41569 ( .A1(n36573), .A2(n36577), .ZN(n36584) );
  INHSV4 U41570 ( .I(n37791), .ZN(n45290) );
  NOR2HSV2 U41571 ( .A1(n45290), .A2(n38454), .ZN(n36583) );
  CLKNAND2HSV1 U41572 ( .A1(n36583), .A2(n59979), .ZN(n36576) );
  XNOR2HSV4 U41573 ( .A1(n36578), .A2(n26874), .ZN(n53381) );
  CLKNHSV2 U41574 ( .I(n37791), .ZN(n52053) );
  CLKAND2HSV2 U41575 ( .A1(n52053), .A2(n45100), .Z(n37786) );
  XNOR2HSV4 U41576 ( .A1(n36581), .A2(n36580), .ZN(n38023) );
  CLKNHSV4 U41577 ( .I(n36582), .ZN(n36585) );
  NAND2HSV4 U41578 ( .A1(n36586), .A2(n37918), .ZN(n37975) );
  INHSV2 U41579 ( .I(n36587), .ZN(n38291) );
  NAND2HSV2 U41580 ( .A1(n38291), .A2(n44711), .ZN(n36601) );
  CLKNAND2HSV0 U41581 ( .A1(n36589), .A2(n36588), .ZN(n36592) );
  INHSV2 U41582 ( .I(n38655), .ZN(n50956) );
  CLKNAND2HSV1 U41583 ( .A1(n50956), .A2(n36590), .ZN(n36591) );
  XOR2HSV0 U41584 ( .A1(n36592), .A2(n36591), .Z(n36595) );
  NAND2HSV2 U41585 ( .A1(n53014), .A2(\pe2/pvq [9]), .ZN(n36593) );
  XNOR2HSV1 U41586 ( .A1(n36593), .A2(\pe2/phq [9]), .ZN(n36594) );
  XNOR2HSV1 U41587 ( .A1(n36595), .A2(n36594), .ZN(n36599) );
  NOR2HSV2 U41588 ( .A1(n44049), .A2(n44699), .ZN(n36597) );
  INHSV2 U41589 ( .I(n38687), .ZN(n45015) );
  CLKNAND2HSV1 U41590 ( .A1(n59582), .A2(n45015), .ZN(n36596) );
  XOR2HSV0 U41591 ( .A1(n36597), .A2(n36596), .Z(n36598) );
  XNOR2HSV1 U41592 ( .A1(n36599), .A2(n36598), .ZN(n36600) );
  XNOR2HSV1 U41593 ( .A1(n36601), .A2(n36600), .ZN(n36622) );
  CLKNAND2HSV1 U41594 ( .A1(\pe2/got [24]), .A2(n36602), .ZN(n36613) );
  CLKNAND2HSV1 U41595 ( .A1(n36603), .A2(n44987), .ZN(n36606) );
  NAND2HSV2 U41596 ( .A1(n36604), .A2(n38064), .ZN(n36605) );
  XNOR2HSV1 U41597 ( .A1(n36606), .A2(n36605), .ZN(n36612) );
  CLKNAND2HSV1 U41598 ( .A1(n37792), .A2(n38047), .ZN(n38499) );
  CLKNAND2HSV1 U41599 ( .A1(n59971), .A2(n36607), .ZN(n36610) );
  CLKNAND2HSV0 U41600 ( .A1(n49530), .A2(n36608), .ZN(n36609) );
  XOR2HSV0 U41601 ( .A1(n36610), .A2(n36609), .Z(n36611) );
  XOR4HSV1 U41602 ( .A1(n36613), .A2(n36612), .A3(n38499), .A4(n36611), .Z(
        n36615) );
  OAI21HSV2 U41603 ( .A1(n44971), .A2(n52285), .B(n36615), .ZN(n36618) );
  NOR2HSV0 U41604 ( .A1(n36615), .A2(n38042), .ZN(n36616) );
  NAND2HSV2 U41605 ( .A1(n59349), .A2(n36616), .ZN(n36617) );
  NAND2HSV2 U41606 ( .A1(n36618), .A2(n36617), .ZN(n36621) );
  BUFHSV2 U41607 ( .I(n36619), .Z(n44187) );
  INHSV1 U41608 ( .I(n38472), .ZN(n59981) );
  NAND2HSV2 U41609 ( .A1(n44187), .A2(n59981), .ZN(n36620) );
  XOR3HSV2 U41610 ( .A1(n36622), .A2(n36621), .A3(n36620), .Z(n36625) );
  CLKNAND2HSV1 U41611 ( .A1(n44906), .A2(n36623), .ZN(n36624) );
  CLKNHSV2 U41612 ( .I(n36626), .ZN(n36627) );
  XNOR2HSV4 U41613 ( .A1(n36628), .A2(n36627), .ZN(n36664) );
  BUFHSV2 U41614 ( .I(n38629), .Z(n59586) );
  NOR2HSV2 U41615 ( .A1(n36632), .A2(n38514), .ZN(n36633) );
  XNOR2HSV4 U41616 ( .A1(n36664), .A2(n36634), .ZN(n36652) );
  CLKNHSV0 U41617 ( .I(n37827), .ZN(n36636) );
  NOR2HSV0 U41618 ( .A1(n36636), .A2(n45267), .ZN(n36637) );
  OAI31HSV0 U41619 ( .A1(n36638), .A2(n36639), .A3(n38629), .B(n36637), .ZN(
        n36644) );
  NAND2HSV0 U41620 ( .A1(n36640), .A2(n45100), .ZN(n36641) );
  CLKNHSV0 U41621 ( .I(n36645), .ZN(n36646) );
  CLKNAND2HSV0 U41622 ( .A1(n36646), .A2(n36647), .ZN(n36648) );
  NAND2HSV2 U41623 ( .A1(n36649), .A2(n36648), .ZN(n37835) );
  INHSV2 U41624 ( .I(n37835), .ZN(n36651) );
  NAND2HSV2 U41625 ( .A1(n36653), .A2(n36652), .ZN(n37845) );
  NAND2HSV4 U41626 ( .A1(n37847), .A2(n37845), .ZN(n47998) );
  NOR2HSV2 U41627 ( .A1(n47998), .A2(n37923), .ZN(n36668) );
  INHSV2 U41628 ( .I(n36657), .ZN(n36658) );
  NAND3HSV3 U41629 ( .A1(n36659), .A2(n29694), .A3(n36658), .ZN(n37832) );
  INHSV2 U41630 ( .I(n37832), .ZN(n37919) );
  CLKNAND2HSV2 U41631 ( .A1(n36660), .A2(n37919), .ZN(n36667) );
  NAND2HSV2 U41632 ( .A1(n52934), .A2(n36661), .ZN(n36663) );
  BUFHSV2 U41633 ( .I(n36665), .Z(n38013) );
  AOI22HSV4 U41634 ( .A1(n37927), .A2(n36668), .B1(n36667), .B2(n36666), .ZN(
        n36669) );
  CLKBUFHSV4 U41635 ( .I(n36682), .Z(n37168) );
  BUFHSV2 U41636 ( .I(n37168), .Z(n36692) );
  INHSV2 U41637 ( .I(\pe3/ti_7t [1]), .ZN(n36670) );
  CLKBUFHSV4 U41638 ( .I(n36682), .Z(n36724) );
  CLKAND2HSV4 U41639 ( .A1(n36671), .A2(n36724), .Z(n36672) );
  INHSV4 U41640 ( .I(n36672), .ZN(n45621) );
  INHSV2 U41641 ( .I(n36672), .ZN(n42609) );
  INHSV2 U41642 ( .I(\pe3/ctrq ), .ZN(n36791) );
  INHSV2 U41643 ( .I(n36791), .ZN(n48075) );
  NAND2HSV2 U41644 ( .A1(n48075), .A2(\pe3/pvq [3]), .ZN(n36681) );
  INHSV2 U41645 ( .I(\pe3/phq [3]), .ZN(n36673) );
  XNOR2HSV4 U41646 ( .A1(n36674), .A2(n36673), .ZN(n36680) );
  INHSV4 U41647 ( .I(\pe3/bq[32] ), .ZN(n43623) );
  NOR2HSV2 U41648 ( .A1(n43757), .A2(n43623), .ZN(n36679) );
  INHSV4 U41649 ( .I(\pe3/got [30]), .ZN(n36751) );
  OAI21HSV4 U41650 ( .A1(n36677), .A2(n42821), .B(n36676), .ZN(n36678) );
  CLKBUFHSV4 U41651 ( .I(n36682), .Z(n43870) );
  INHSV2 U41652 ( .I(n43870), .ZN(n43591) );
  NOR2HSV2 U41653 ( .A1(n43591), .A2(n36719), .ZN(n36902) );
  AOI22HSV2 U41654 ( .A1(n36696), .A2(\pe3/got [31]), .B1(n49001), .B2(n36902), 
        .ZN(n36684) );
  INHSV3 U41655 ( .I(n36683), .ZN(n36686) );
  INHSV2 U41656 ( .I(n36684), .ZN(n36685) );
  CLKNAND2HSV3 U41657 ( .A1(n36686), .A2(n36685), .ZN(n36687) );
  INHSV3 U41658 ( .I(n43467), .ZN(n36877) );
  AOI21HSV4 U41659 ( .A1(n48893), .A2(n36877), .B(n36689), .ZN(n36690) );
  INHSV2 U41660 ( .I(\pe3/ti_7t [3]), .ZN(n36691) );
  NOR2HSV2 U41661 ( .A1(n36692), .A2(n36691), .ZN(n36782) );
  INHSV2 U41662 ( .I(n36782), .ZN(n36709) );
  INHSV4 U41663 ( .I(n36693), .ZN(n37020) );
  INHSV2 U41664 ( .I(n37265), .ZN(n45612) );
  INHSV2 U41665 ( .I(n36989), .ZN(n36710) );
  INHSV2 U41666 ( .I(n43623), .ZN(n36795) );
  INHSV4 U41667 ( .I(n42643), .ZN(n59609) );
  INHSV4 U41668 ( .I(n59606), .ZN(n59614) );
  INHSV4 U41669 ( .I(n36694), .ZN(n37298) );
  INHSV2 U41670 ( .I(n36791), .ZN(n46139) );
  INHSV2 U41671 ( .I(n36999), .ZN(n59608) );
  INHSV2 U41672 ( .I(\pe3/bq[30] ), .ZN(n37185) );
  NAND2HSV2 U41673 ( .A1(n59608), .A2(n36789), .ZN(n42651) );
  CLKNAND2HSV2 U41674 ( .A1(n49001), .A2(n43021), .ZN(n36698) );
  INHSV2 U41675 ( .I(n36696), .ZN(n36697) );
  NAND2HSV4 U41676 ( .A1(n36698), .A2(n36697), .ZN(n43185) );
  INHSV2 U41677 ( .I(n36751), .ZN(n43464) );
  NAND2HSV2 U41678 ( .A1(n43185), .A2(n43464), .ZN(n36699) );
  XNOR2HSV4 U41679 ( .A1(n36700), .A2(n36699), .ZN(n36749) );
  INHSV2 U41680 ( .I(n45625), .ZN(n45932) );
  INHSV1 U41681 ( .I(\pe3/ti_7t [2]), .ZN(n36701) );
  CLKBUFHSV4 U41682 ( .I(n36682), .Z(n36972) );
  INHSV2 U41683 ( .I(n36972), .ZN(n43242) );
  INHSV4 U41684 ( .I(\pe3/got [31]), .ZN(n37348) );
  AOI21HSV2 U41685 ( .A1(n36701), .A2(n43242), .B(n37348), .ZN(n36702) );
  OAI21HSV2 U41686 ( .A1(n48893), .A2(n45932), .B(n36702), .ZN(n36703) );
  XNOR2HSV4 U41687 ( .A1(n36749), .A2(n36703), .ZN(n36705) );
  INHSV2 U41688 ( .I(n36877), .ZN(n36704) );
  NOR2HSV4 U41689 ( .A1(n36705), .A2(n36704), .ZN(n36706) );
  NAND2HSV4 U41690 ( .A1(n36708), .A2(n36707), .ZN(n36775) );
  CLKNHSV2 U41691 ( .I(n36724), .ZN(n37454) );
  NOR2HSV2 U41692 ( .A1(\pe3/got [32]), .A2(n43743), .ZN(n36901) );
  INHSV2 U41693 ( .I(n45622), .ZN(n37447) );
  NAND2HSV2 U41694 ( .A1(n43743), .A2(\pe3/ti_7t [5]), .ZN(n36864) );
  INHSV2 U41695 ( .I(n36864), .ZN(n36839) );
  NOR2HSV0 U41696 ( .A1(n37447), .A2(n36839), .ZN(n36737) );
  INHSV2 U41697 ( .I(n45555), .ZN(n59809) );
  INHSV3 U41698 ( .I(n36711), .ZN(n46141) );
  INHSV2 U41699 ( .I(\pe3/got [29]), .ZN(n37784) );
  INHSV2 U41700 ( .I(n37784), .ZN(n36788) );
  NAND2HSV2 U41701 ( .A1(n43185), .A2(n36788), .ZN(n36713) );
  NAND2HSV2 U41702 ( .A1(n36712), .A2(n36713), .ZN(n36716) );
  INHSV2 U41703 ( .I(n36713), .ZN(n36714) );
  NAND2HSV4 U41704 ( .A1(n36716), .A2(n36715), .ZN(n36727) );
  NOR2HSV2 U41705 ( .A1(n36727), .A2(n43880), .ZN(n36717) );
  INHSV2 U41706 ( .I(n36727), .ZN(n36730) );
  BUFHSV2 U41707 ( .I(n36719), .Z(n36721) );
  INHSV2 U41708 ( .I(n36721), .ZN(n36729) );
  NAND2HSV2 U41709 ( .A1(\pe3/ti_7t [2]), .A2(n36689), .ZN(n36725) );
  INHSV2 U41710 ( .I(n43464), .ZN(n43744) );
  NAND2HSV4 U41711 ( .A1(n37017), .A2(n42697), .ZN(n36733) );
  OAI22HSV4 U41712 ( .A1(n36732), .A2(n36731), .B1(n36730), .B2(n36729), .ZN(
        n36734) );
  NOR2HSV4 U41713 ( .A1(n36734), .A2(n36733), .ZN(n36736) );
  INHSV2 U41714 ( .I(n37348), .ZN(n36924) );
  CLKNAND2HSV1 U41715 ( .A1(n36738), .A2(n36924), .ZN(n36741) );
  INHSV2 U41716 ( .I(n37238), .ZN(n36898) );
  CLKAND2HSV1 U41717 ( .A1(n36729), .A2(n36844), .Z(n36739) );
  CLKNAND2HSV0 U41718 ( .A1(n36775), .A2(n36739), .ZN(n36740) );
  CLKNAND2HSV1 U41719 ( .A1(n36741), .A2(n36740), .ZN(n36742) );
  NAND2HSV4 U41720 ( .A1(n36746), .A2(n46107), .ZN(n36750) );
  CLKAND2HSV2 U41721 ( .A1(n36925), .A2(n43898), .Z(n36754) );
  CLKAND2HSV2 U41722 ( .A1(n43604), .A2(n44669), .Z(n36747) );
  BUFHSV2 U41723 ( .I(n36751), .Z(n46084) );
  INHSV2 U41724 ( .I(n43752), .ZN(n46082) );
  NAND2HSV2 U41725 ( .A1(n47428), .A2(\pe3/ti_7t [4]), .ZN(n36926) );
  OAI22HSV4 U41726 ( .A1(n36780), .A2(n36752), .B1(n46084), .B2(n36926), .ZN(
        n36753) );
  AOI21HSV4 U41727 ( .A1(n36779), .A2(n36754), .B(n36753), .ZN(n36771) );
  BUFHSV4 U41728 ( .I(n43185), .Z(n37012) );
  BUFHSV2 U41729 ( .I(n42683), .Z(n43235) );
  NAND2HSV2 U41730 ( .A1(n37012), .A2(n36958), .ZN(n36767) );
  INHSV3 U41731 ( .I(n25889), .ZN(n46133) );
  CLKNHSV1 U41732 ( .I(n36989), .ZN(n46463) );
  INHSV2 U41733 ( .I(n36694), .ZN(n48527) );
  NAND2HSV2 U41734 ( .A1(n46463), .A2(n48527), .ZN(n36947) );
  INHSV2 U41735 ( .I(n42843), .ZN(n36755) );
  CLKNAND2HSV1 U41736 ( .A1(n36755), .A2(\pe3/bq[31] ), .ZN(n36756) );
  XOR2HSV0 U41737 ( .A1(n36947), .A2(n36756), .Z(n36757) );
  INHSV2 U41738 ( .I(n45525), .ZN(n43780) );
  CLKNAND2HSV0 U41739 ( .A1(n59608), .A2(n43780), .ZN(n36759) );
  INHSV2 U41740 ( .I(n45555), .ZN(n55750) );
  INHSV2 U41741 ( .I(n37185), .ZN(n37112) );
  CLKNAND2HSV1 U41742 ( .A1(n55750), .A2(n37112), .ZN(n36758) );
  XOR2HSV0 U41743 ( .A1(n36759), .A2(n36758), .Z(n36763) );
  NAND2HSV2 U41744 ( .A1(n55988), .A2(n37180), .ZN(n36761) );
  CLKNAND2HSV1 U41745 ( .A1(n59614), .A2(\pe3/bq[26] ), .ZN(n36760) );
  XOR2HSV0 U41746 ( .A1(n36761), .A2(n36760), .Z(n36762) );
  XOR2HSV0 U41747 ( .A1(n36763), .A2(n36762), .Z(n36764) );
  INHSV2 U41748 ( .I(n45941), .ZN(n46309) );
  XOR3HSV2 U41749 ( .A1(n36767), .A2(n36766), .A3(n36765), .Z(n36768) );
  XNOR2HSV4 U41750 ( .A1(n36769), .A2(n36768), .ZN(n36770) );
  XNOR2HSV4 U41751 ( .A1(n36771), .A2(n36770), .ZN(n36772) );
  XNOR2HSV4 U41752 ( .A1(n36773), .A2(n36772), .ZN(n36884) );
  NOR2HSV4 U41753 ( .A1(n36774), .A2(n36861), .ZN(n36858) );
  BUFHSV2 U41754 ( .I(n37168), .Z(n42806) );
  INHSV2 U41755 ( .I(n36775), .ZN(n36841) );
  NAND2HSV2 U41756 ( .A1(n36776), .A2(n36777), .ZN(n36805) );
  NOR2HSV3 U41757 ( .A1(n36858), .A2(n36778), .ZN(n36963) );
  NOR2HSV2 U41758 ( .A1(n36926), .A2(n43880), .ZN(n36781) );
  INHSV2 U41759 ( .I(n46084), .ZN(n42697) );
  INHSV2 U41760 ( .I(n36784), .ZN(n36785) );
  INHSV2 U41761 ( .I(n46084), .ZN(n37081) );
  CLKNAND2HSV1 U41762 ( .A1(n37274), .A2(n36788), .ZN(n36802) );
  INHSV2 U41763 ( .I(n45555), .ZN(n37109) );
  INHSV2 U41764 ( .I(n45649), .ZN(n37280) );
  INHSV2 U41765 ( .I(n42843), .ZN(n55987) );
  INHSV2 U41766 ( .I(n36799), .ZN(n37041) );
  CLKNAND2HSV1 U41767 ( .A1(n43185), .A2(n55940), .ZN(n36800) );
  XNOR2HSV4 U41768 ( .A1(n36802), .A2(n36801), .ZN(n36803) );
  XNOR2HSV4 U41769 ( .A1(n36857), .A2(n36856), .ZN(n36804) );
  MUX2NHSV4 U41770 ( .I0(n36805), .I1(n36963), .S(n36804), .ZN(n36883) );
  OAI21HSV2 U41771 ( .A1(n42806), .A2(\pe3/ti_7t [6]), .B(n59962), .ZN(n36806)
         );
  NOR2HSV4 U41772 ( .A1(n36883), .A2(n36806), .ZN(n36807) );
  XNOR2HSV4 U41773 ( .A1(n36884), .A2(n36807), .ZN(n36916) );
  NAND2HSV2 U41774 ( .A1(n37017), .A2(n36958), .ZN(n36808) );
  INHSV2 U41775 ( .I(n36808), .ZN(n36832) );
  INHSV1 U41776 ( .I(n42843), .ZN(n36809) );
  NAND2HSV2 U41777 ( .A1(n36809), .A2(n37112), .ZN(n36811) );
  CLKNAND2HSV0 U41778 ( .A1(n59614), .A2(n42527), .ZN(n36810) );
  XOR2HSV0 U41779 ( .A1(n36811), .A2(n36810), .Z(n36815) );
  INHSV2 U41780 ( .I(n45555), .ZN(n37374) );
  NAND2HSV2 U41781 ( .A1(n37374), .A2(n48527), .ZN(n36813) );
  CLKNAND2HSV1 U41782 ( .A1(\pe3/aot [25]), .A2(n37180), .ZN(n36812) );
  XOR2HSV0 U41783 ( .A1(n36813), .A2(n36812), .Z(n36814) );
  XOR2HSV0 U41784 ( .A1(n36815), .A2(n36814), .Z(n36830) );
  INHSV2 U41785 ( .I(n45525), .ZN(n37050) );
  CLKNAND2HSV1 U41786 ( .A1(n48496), .A2(n37050), .ZN(n36818) );
  INHSV1 U41787 ( .I(n45948), .ZN(n43855) );
  CLKNAND2HSV0 U41788 ( .A1(n43855), .A2(n36816), .ZN(n36817) );
  CLKNAND2HSV0 U41789 ( .A1(n59608), .A2(\pe3/bq[26] ), .ZN(n36820) );
  CLKNAND2HSV1 U41790 ( .A1(\pe3/aot [26]), .A2(n37186), .ZN(n36819) );
  XOR2HSV0 U41791 ( .A1(n36820), .A2(n36819), .Z(n36821) );
  XOR2HSV0 U41792 ( .A1(n36822), .A2(n36821), .Z(n36827) );
  NAND2HSV2 U41793 ( .A1(n46133), .A2(\pe3/pvq [8]), .ZN(n36823) );
  XNOR2HSV1 U41794 ( .A1(n36823), .A2(\pe3/phq [8]), .ZN(n36825) );
  CLKNAND2HSV1 U41795 ( .A1(n37373), .A2(n42634), .ZN(n36824) );
  XNOR2HSV1 U41796 ( .A1(n36825), .A2(n36824), .ZN(n36826) );
  XNOR2HSV1 U41797 ( .A1(n36827), .A2(n36826), .ZN(n36828) );
  XOR3HSV2 U41798 ( .A1(n36830), .A2(n36829), .A3(n36828), .Z(n36831) );
  XNOR2HSV1 U41799 ( .A1(n36832), .A2(n36831), .ZN(n36834) );
  INHSV2 U41800 ( .I(n37273), .ZN(n55940) );
  NAND2HSV2 U41801 ( .A1(n37312), .A2(n55940), .ZN(n36833) );
  XNOR2HSV4 U41802 ( .A1(n36834), .A2(n36833), .ZN(n36849) );
  CLKNAND2HSV1 U41803 ( .A1(n36925), .A2(n59963), .ZN(n36835) );
  INHSV2 U41804 ( .I(\pe3/got [29]), .ZN(n43866) );
  OAI22HSV2 U41805 ( .A1(n36835), .A2(n36930), .B1(n43866), .B2(n36926), .ZN(
        n36838) );
  NOR2HSV2 U41806 ( .A1(n36925), .A2(n43866), .ZN(n36836) );
  CLKAND2HSV2 U41807 ( .A1(n36928), .A2(n36836), .Z(n36837) );
  NOR2HSV4 U41808 ( .A1(n36838), .A2(n36837), .ZN(n36848) );
  XNOR2HSV4 U41809 ( .A1(n36849), .A2(n36848), .ZN(n36889) );
  BUFHSV2 U41810 ( .I(n46090), .Z(n37241) );
  OAI22HSV4 U41811 ( .A1(n36964), .A2(n37241), .B1(n36842), .B2(n36863), .ZN(
        n36875) );
  INHSV3 U41812 ( .I(n36875), .ZN(n36874) );
  NOR2HSV2 U41813 ( .A1(n37241), .A2(n36861), .ZN(n36843) );
  INHSV2 U41814 ( .I(n36845), .ZN(n36846) );
  CLKNAND2HSV3 U41815 ( .A1(n36874), .A2(n36847), .ZN(n36891) );
  NAND2HSV2 U41816 ( .A1(n36851), .A2(n36891), .ZN(n36907) );
  NOR2HSV2 U41817 ( .A1(n36876), .A2(n36875), .ZN(n36852) );
  XNOR2HSV4 U41818 ( .A1(n36849), .A2(n36848), .ZN(n36885) );
  NAND2HSV2 U41819 ( .A1(n36852), .A2(n36885), .ZN(n36900) );
  NAND2HSV2 U41820 ( .A1(n36907), .A2(n36900), .ZN(n36895) );
  INHSV2 U41821 ( .I(n36895), .ZN(n36850) );
  CLKNHSV1 U41822 ( .I(n36885), .ZN(n36851) );
  NAND2HSV2 U41823 ( .A1(n36891), .A2(n36851), .ZN(n36854) );
  CLKNAND2HSV1 U41824 ( .A1(n36885), .A2(n36852), .ZN(n36853) );
  NAND2HSV2 U41825 ( .A1(n36854), .A2(n36853), .ZN(n52739) );
  INHSV2 U41826 ( .I(n43483), .ZN(n37264) );
  CLKAND2HSV2 U41827 ( .A1(n52739), .A2(n37264), .Z(n36855) );
  NAND2HSV2 U41828 ( .A1(n36855), .A2(n36916), .ZN(n36881) );
  XNOR2HSV4 U41829 ( .A1(n36857), .A2(n36856), .ZN(n36871) );
  INHSV2 U41830 ( .I(n36871), .ZN(n36869) );
  BUFHSV2 U41831 ( .I(n45931), .Z(n45628) );
  INHSV2 U41832 ( .I(n45628), .ZN(n36859) );
  CLKNAND2HSV2 U41833 ( .A1(n36858), .A2(n36859), .ZN(n36870) );
  AND2HSV2 U41834 ( .A1(n42806), .A2(n36859), .Z(n36860) );
  NAND2HSV2 U41835 ( .A1(n36861), .A2(n36860), .ZN(n36862) );
  INHSV2 U41836 ( .I(n36862), .ZN(n36867) );
  INHSV2 U41837 ( .I(n36863), .ZN(n36866) );
  NOR2HSV2 U41838 ( .A1(n36864), .A2(n45628), .ZN(n36865) );
  AOI21HSV4 U41839 ( .A1(n36867), .A2(n36866), .B(n36865), .ZN(n36872) );
  NAND2HSV2 U41840 ( .A1(n36870), .A2(n36872), .ZN(n36868) );
  CLKNHSV0 U41841 ( .I(n36902), .ZN(n43359) );
  INHSV2 U41842 ( .I(n43359), .ZN(n43608) );
  NOR2HSV2 U41843 ( .A1(n36876), .A2(n36875), .ZN(n36890) );
  NOR2HSV1 U41844 ( .A1(n36890), .A2(n36877), .ZN(n36878) );
  CLKNAND2HSV1 U41845 ( .A1(n36878), .A2(n36889), .ZN(n36879) );
  CLKNHSV2 U41846 ( .I(n36909), .ZN(n36888) );
  INAND2HSV0 U41847 ( .A1(n36889), .B1(n36891), .ZN(n36887) );
  AOI21HSV0 U41848 ( .A1(n36890), .A2(n36885), .B(n43467), .ZN(n36886) );
  MUX2NHSV2 U41849 ( .I0(n36891), .I1(n36890), .S(n36889), .ZN(n36899) );
  INHSV2 U41850 ( .I(n36893), .ZN(n36894) );
  NAND2HSV2 U41851 ( .A1(n36909), .A2(n36895), .ZN(n36896) );
  INHSV2 U41852 ( .I(n36898), .ZN(n43905) );
  INHSV2 U41853 ( .I(n37447), .ZN(n37089) );
  INHSV2 U41854 ( .I(n36900), .ZN(n36905) );
  INHSV2 U41855 ( .I(n36902), .ZN(n45624) );
  INHSV2 U41856 ( .I(n45624), .ZN(n43355) );
  NOR2HSV0 U41857 ( .A1(n42806), .A2(\pe3/ti_7t [8]), .ZN(n36903) );
  OR2HSV1 U41858 ( .A1(n43355), .A2(n36903), .Z(n36904) );
  CLKAND2HSV2 U41859 ( .A1(n52739), .A2(n43126), .Z(n36910) );
  CLKNAND2HSV1 U41860 ( .A1(n36910), .A2(n36909), .ZN(n36911) );
  NAND3HSV4 U41861 ( .A1(n36915), .A2(n36914), .A3(n36913), .ZN(n36923) );
  INHSV4 U41862 ( .I(n36923), .ZN(n37085) );
  INHSV4 U41863 ( .I(n37085), .ZN(n37106) );
  INHSV2 U41864 ( .I(n37784), .ZN(n37340) );
  CLKNAND2HSV3 U41865 ( .A1(n37106), .A2(n37340), .ZN(n36984) );
  CLKNHSV0 U41866 ( .I(\pe3/got [30]), .ZN(n43752) );
  CLKNAND2HSV2 U41867 ( .A1(n36916), .A2(n36979), .ZN(n36919) );
  INHSV2 U41868 ( .I(\pe3/ti_7t [7]), .ZN(n36917) );
  OR2HSV1 U41869 ( .A1(n42806), .A2(n36917), .Z(n36918) );
  INHSV2 U41870 ( .I(n37170), .ZN(n36921) );
  NAND2HSV2 U41871 ( .A1(n37161), .A2(n59962), .ZN(n36920) );
  NOR2HSV4 U41872 ( .A1(n36921), .A2(n36920), .ZN(n36922) );
  NAND2HSV2 U41873 ( .A1(n37170), .A2(n36924), .ZN(n48619) );
  INHSV2 U41874 ( .I(n36925), .ZN(n36931) );
  CLKNHSV1 U41875 ( .I(n36926), .ZN(n36927) );
  AOI21HSV2 U41876 ( .A1(n36928), .A2(n36931), .B(n36927), .ZN(n36929) );
  OAI21HSV2 U41877 ( .A1(n36931), .A2(n36930), .B(n36929), .ZN(n42874) );
  INHSV2 U41878 ( .I(n42874), .ZN(n37043) );
  INHSV2 U41879 ( .I(n37043), .ZN(n37316) );
  INAND2HSV2 U41880 ( .A1(n37273), .B1(n37316), .ZN(n36962) );
  CLKNAND2HSV1 U41881 ( .A1(n48496), .A2(\pe3/bq[26] ), .ZN(n36933) );
  BUFHSV2 U41882 ( .I(\pe3/aot [26]), .Z(n59610) );
  CLKNAND2HSV0 U41883 ( .A1(n59610), .A2(n37112), .ZN(n36932) );
  XOR2HSV0 U41884 ( .A1(n36933), .A2(n36932), .Z(n36937) );
  NAND2HSV0 U41885 ( .A1(n59608), .A2(n42527), .ZN(n36935) );
  CLKNAND2HSV0 U41886 ( .A1(n43034), .A2(n46614), .ZN(n36934) );
  XOR2HSV0 U41887 ( .A1(n36935), .A2(n36934), .Z(n36936) );
  XOR2HSV0 U41888 ( .A1(n36937), .A2(n36936), .Z(n36954) );
  INHSV2 U41889 ( .I(n45948), .ZN(n45634) );
  NAND2HSV2 U41890 ( .A1(n37012), .A2(n45634), .ZN(n36953) );
  CLKNAND2HSV1 U41891 ( .A1(n37109), .A2(n43539), .ZN(n36939) );
  INHSV2 U41892 ( .I(n55714), .ZN(n37279) );
  CLKNAND2HSV1 U41893 ( .A1(n37279), .A2(n37186), .ZN(n36938) );
  XOR2HSV0 U41894 ( .A1(n36939), .A2(n36938), .Z(n36944) );
  CLKNAND2HSV0 U41895 ( .A1(n59614), .A2(n42530), .ZN(n36942) );
  CLKBUFHSV4 U41896 ( .I(n36940), .Z(n46126) );
  CLKNAND2HSV1 U41897 ( .A1(n43452), .A2(n37051), .ZN(n36941) );
  XOR2HSV0 U41898 ( .A1(n36942), .A2(n36941), .Z(n36943) );
  XOR2HSV0 U41899 ( .A1(n36944), .A2(n36943), .Z(n36951) );
  INHSV2 U41900 ( .I(n46141), .ZN(n37378) );
  INHSV2 U41901 ( .I(n37378), .ZN(n46616) );
  NAND2HSV2 U41902 ( .A1(n46616), .A2(\pe3/pvq [9]), .ZN(n36945) );
  XOR2HSV0 U41903 ( .A1(n36945), .A2(\pe3/phq [9]), .Z(n36949) );
  NAND2HSV2 U41904 ( .A1(n37050), .A2(n59622), .ZN(n37122) );
  OAI22HSV1 U41905 ( .A1(n36694), .A2(n42843), .B1(n36989), .B2(n45525), .ZN(
        n36946) );
  OAI21HSV1 U41906 ( .A1(n37122), .A2(n36947), .B(n36946), .ZN(n36948) );
  XOR2HSV0 U41907 ( .A1(n36949), .A2(n36948), .Z(n36950) );
  XNOR2HSV1 U41908 ( .A1(n36951), .A2(n36950), .ZN(n36952) );
  XOR3HSV2 U41909 ( .A1(n36954), .A2(n36953), .A3(n36952), .Z(n36957) );
  CLKNAND2HSV0 U41910 ( .A1(n37017), .A2(n36955), .ZN(n36956) );
  XNOR2HSV1 U41911 ( .A1(n36957), .A2(n36956), .ZN(n36960) );
  CLKNAND2HSV1 U41912 ( .A1(n37312), .A2(n36958), .ZN(n36959) );
  XNOR2HSV1 U41913 ( .A1(n36960), .A2(n36959), .ZN(n36961) );
  XNOR2HSV1 U41914 ( .A1(n36962), .A2(n36961), .ZN(n36966) );
  NAND2HSV2 U41915 ( .A1(n36964), .A2(n36963), .ZN(n59613) );
  CLKBUFHSV4 U41916 ( .I(n59613), .Z(n55951) );
  NAND2HSV2 U41917 ( .A1(n55951), .A2(n36788), .ZN(n36965) );
  XNOR2HSV1 U41918 ( .A1(n36966), .A2(n36965), .ZN(n36971) );
  BUFHSV2 U41919 ( .I(n37168), .Z(n43604) );
  NAND2HSV2 U41920 ( .A1(n36967), .A2(\pe3/ti_7t [6]), .ZN(n36968) );
  NAND2HSV4 U41921 ( .A1(n36969), .A2(n36968), .ZN(n52738) );
  NAND2HSV2 U41922 ( .A1(n52738), .A2(n37081), .ZN(n36970) );
  XNOR2HSV4 U41923 ( .A1(n36971), .A2(n36970), .ZN(n48620) );
  INHSV2 U41924 ( .I(\pe3/ti_7t [9]), .ZN(n36973) );
  NOR2HSV2 U41925 ( .A1(n45615), .A2(n36973), .ZN(n37099) );
  INHSV2 U41926 ( .I(n46084), .ZN(n37272) );
  NAND2HSV0 U41927 ( .A1(n37099), .A2(n37272), .ZN(n36983) );
  CLKNHSV1 U41928 ( .I(n36983), .ZN(n36974) );
  INAND2HSV2 U41929 ( .A1(n42697), .B1(n36986), .ZN(n36976) );
  NAND2HSV2 U41930 ( .A1(n36977), .A2(n36976), .ZN(n37033) );
  NOR2HSV2 U41931 ( .A1(n48620), .A2(n36980), .ZN(n36981) );
  CLKNAND2HSV3 U41932 ( .A1(n37104), .A2(n37103), .ZN(n37236) );
  NAND3HSV2 U41933 ( .A1(n37236), .A2(n36986), .A3(n37101), .ZN(n37035) );
  CLKBUFHSV4 U41934 ( .I(n52738), .Z(n49405) );
  CLKNAND2HSV1 U41935 ( .A1(n45949), .A2(n37107), .ZN(n37028) );
  CLKBUFHSV4 U41936 ( .I(n59613), .Z(n37176) );
  BUFHSV2 U41937 ( .I(n42938), .Z(n37457) );
  NAND2HSV2 U41938 ( .A1(n37457), .A2(n59616), .ZN(n37026) );
  BUFHSV2 U41939 ( .I(n45948), .Z(n37785) );
  INHSV2 U41940 ( .I(n37785), .ZN(n37175) );
  CLKNAND2HSV0 U41941 ( .A1(n37316), .A2(n37175), .ZN(n37024) );
  NAND2HSV0 U41942 ( .A1(n59612), .A2(n37112), .ZN(n36988) );
  CLKNAND2HSV1 U41943 ( .A1(n36809), .A2(\pe3/bq[26] ), .ZN(n36987) );
  XOR2HSV0 U41944 ( .A1(n36988), .A2(n36987), .Z(n36993) );
  NAND2HSV0 U41945 ( .A1(n37279), .A2(n37280), .ZN(n36991) );
  INHSV2 U41946 ( .I(n36989), .ZN(n37373) );
  CLKNAND2HSV0 U41947 ( .A1(n37373), .A2(n42530), .ZN(n36990) );
  XOR2HSV0 U41948 ( .A1(n36991), .A2(n36990), .Z(n36992) );
  XOR2HSV0 U41949 ( .A1(n36993), .A2(n36992), .Z(n37016) );
  NAND2HSV0 U41950 ( .A1(n37374), .A2(n42527), .ZN(n36995) );
  NAND2HSV0 U41951 ( .A1(n43034), .A2(n37298), .ZN(n36994) );
  XOR2HSV0 U41952 ( .A1(n36995), .A2(n36994), .Z(n36998) );
  CLKNHSV0 U41953 ( .I(n37378), .ZN(n46130) );
  NAND2HSV2 U41954 ( .A1(n46130), .A2(\pe3/pvq [12]), .ZN(n36996) );
  XNOR2HSV1 U41955 ( .A1(n36996), .A2(\pe3/phq [12]), .ZN(n36997) );
  XNOR2HSV1 U41956 ( .A1(n36998), .A2(n36997), .ZN(n37004) );
  INHSV2 U41957 ( .I(n37196), .ZN(n45807) );
  NAND2HSV2 U41958 ( .A1(n56182), .A2(n45807), .ZN(n43071) );
  BUFHSV2 U41959 ( .I(n43623), .Z(n42833) );
  BUFHSV2 U41960 ( .I(n36999), .Z(n43392) );
  OAI22HSV1 U41961 ( .A1(n42833), .A2(n42539), .B1(n43392), .B2(n37196), .ZN(
        n37000) );
  OAI21HSV0 U41962 ( .A1(n43071), .A2(n37001), .B(n37000), .ZN(n37002) );
  NOR2HSV2 U41963 ( .A1(n42821), .A2(n43039), .ZN(n43420) );
  XNOR2HSV1 U41964 ( .A1(n37002), .A2(n43420), .ZN(n37003) );
  XNOR2HSV1 U41965 ( .A1(n37004), .A2(n37003), .ZN(n37015) );
  CLKNHSV0 U41966 ( .I(n45525), .ZN(n37276) );
  CLKNAND2HSV0 U41967 ( .A1(n59610), .A2(n37276), .ZN(n37006) );
  CLKNAND2HSV1 U41968 ( .A1(n37362), .A2(n56213), .ZN(n37005) );
  XOR2HSV0 U41969 ( .A1(n37006), .A2(n37005), .Z(n37011) );
  NAND2HSV0 U41970 ( .A1(n59618), .A2(n37186), .ZN(n37009) );
  INHSV2 U41971 ( .I(n37275), .ZN(n42520) );
  CLKNAND2HSV1 U41972 ( .A1(n42520), .A2(n37007), .ZN(n37008) );
  XOR2HSV0 U41973 ( .A1(n37009), .A2(n37008), .Z(n37010) );
  XOR2HSV0 U41974 ( .A1(n37011), .A2(n37010), .Z(n37014) );
  BUFHSV2 U41975 ( .I(n37012), .Z(n37131) );
  CLKNAND2HSV1 U41976 ( .A1(n37131), .A2(n48485), .ZN(n37013) );
  XOR4HSV1 U41977 ( .A1(n37016), .A2(n37015), .A3(n37014), .A4(n37013), .Z(
        n37019) );
  CLKNAND2HSV0 U41978 ( .A1(n37177), .A2(n42673), .ZN(n37018) );
  XNOR2HSV1 U41979 ( .A1(n37019), .A2(n37018), .ZN(n37022) );
  CLKNAND2HSV1 U41980 ( .A1(n59617), .A2(n37312), .ZN(n37021) );
  XNOR2HSV1 U41981 ( .A1(n37022), .A2(n37021), .ZN(n37023) );
  XOR2HSV0 U41982 ( .A1(n37024), .A2(n37023), .Z(n37025) );
  XOR2HSV0 U41983 ( .A1(n37026), .A2(n37025), .Z(n37027) );
  XOR2HSV0 U41984 ( .A1(n37028), .A2(n37027), .Z(n37030) );
  INHSV2 U41985 ( .I(n37273), .ZN(n37169) );
  CLKNAND2HSV1 U41986 ( .A1(n59364), .A2(n37169), .ZN(n37029) );
  XOR2HSV0 U41987 ( .A1(n37030), .A2(n37029), .Z(n37036) );
  INHSV1 U41988 ( .I(n37036), .ZN(n37031) );
  INHSV1 U41989 ( .I(n37033), .ZN(n37037) );
  NAND4HSV2 U41990 ( .A1(n37037), .A2(n37036), .A3(n37035), .A4(n37034), .ZN(
        n37038) );
  CLKNAND2HSV0 U41991 ( .A1(n55951), .A2(n37041), .ZN(n37077) );
  CLKNHSV1 U41992 ( .I(n37176), .ZN(n37042) );
  NOR2HSV2 U41993 ( .A1(n37042), .A2(n45941), .ZN(n37076) );
  INHSV2 U41994 ( .I(n37043), .ZN(n37353) );
  INAND2HSV2 U41995 ( .A1(n43235), .B1(n37353), .ZN(n37074) );
  NAND2HSV0 U41996 ( .A1(n59609), .A2(n42527), .ZN(n37049) );
  INHSV2 U41997 ( .I(n37378), .ZN(n46132) );
  NAND2HSV2 U41998 ( .A1(n46132), .A2(\pe3/pvq [10]), .ZN(n37044) );
  XNOR2HSV1 U41999 ( .A1(n37044), .A2(\pe3/phq [10]), .ZN(n37048) );
  NAND2HSV0 U42000 ( .A1(n36809), .A2(n43539), .ZN(n37046) );
  NAND2HSV0 U42001 ( .A1(n46463), .A2(\pe3/bq[26] ), .ZN(n37045) );
  XOR2HSV0 U42002 ( .A1(n37046), .A2(n37045), .Z(n37047) );
  XOR3HSV2 U42003 ( .A1(n37049), .A2(n37048), .A3(n37047), .Z(n37068) );
  CLKNAND2HSV1 U42004 ( .A1(n37131), .A2(n55701), .ZN(n37067) );
  NAND2HSV0 U42005 ( .A1(n37109), .A2(n37050), .ZN(n37053) );
  INHSV2 U42006 ( .I(n42827), .ZN(n48483) );
  CLKNAND2HSV1 U42007 ( .A1(n48483), .A2(n37051), .ZN(n37052) );
  XOR2HSV0 U42008 ( .A1(n37053), .A2(n37052), .Z(n37057) );
  NAND2HSV0 U42009 ( .A1(\pe3/aot [23]), .A2(n37180), .ZN(n37055) );
  INHSV2 U42010 ( .I(n55714), .ZN(n59368) );
  NAND2HSV0 U42011 ( .A1(n59368), .A2(n37112), .ZN(n37054) );
  XOR2HSV0 U42012 ( .A1(n37055), .A2(n37054), .Z(n37056) );
  XOR2HSV0 U42013 ( .A1(n37057), .A2(n37056), .Z(n37065) );
  NAND2HSV0 U42014 ( .A1(n59610), .A2(n37298), .ZN(n37059) );
  NAND2HSV0 U42015 ( .A1(n45695), .A2(n37186), .ZN(n37058) );
  XOR2HSV0 U42016 ( .A1(n37059), .A2(n37058), .Z(n37063) );
  NAND2HSV0 U42017 ( .A1(n59608), .A2(n42530), .ZN(n37061) );
  INHSV2 U42018 ( .I(n42821), .ZN(n45572) );
  CLKNAND2HSV0 U42019 ( .A1(n45572), .A2(\pe3/bq[23] ), .ZN(n37060) );
  XOR2HSV0 U42020 ( .A1(n37061), .A2(n37060), .Z(n37062) );
  XOR2HSV0 U42021 ( .A1(n37063), .A2(n37062), .Z(n37064) );
  XOR2HSV0 U42022 ( .A1(n37065), .A2(n37064), .Z(n37066) );
  XOR3HSV2 U42023 ( .A1(n37068), .A2(n37067), .A3(n37066), .Z(n37070) );
  CLKNAND2HSV0 U42024 ( .A1(n37177), .A2(n37175), .ZN(n37069) );
  XNOR2HSV1 U42025 ( .A1(n37070), .A2(n37069), .ZN(n37072) );
  NAND2HSV0 U42026 ( .A1(n37312), .A2(n59616), .ZN(n37071) );
  XNOR2HSV1 U42027 ( .A1(n37072), .A2(n37071), .ZN(n37073) );
  XNOR2HSV1 U42028 ( .A1(n37074), .A2(n37073), .ZN(n37075) );
  MUX2NHSV1 U42029 ( .I0(n37077), .I1(n37076), .S(n37075), .ZN(n37078) );
  XNOR2HSV4 U42030 ( .A1(n37079), .A2(n37078), .ZN(n37082) );
  AOI21HSV4 U42031 ( .A1(n59364), .A2(n37081), .B(n37082), .ZN(n37080) );
  CLKNAND2HSV2 U42032 ( .A1(n37084), .A2(n37083), .ZN(n37087) );
  XNOR2HSV4 U42033 ( .A1(n37087), .A2(n37086), .ZN(n37335) );
  INHSV2 U42034 ( .I(\pe3/ti_7t [10]), .ZN(n37091) );
  NOR2HSV2 U42035 ( .A1(n45615), .A2(n37091), .ZN(n37239) );
  CLKAND2HSV2 U42036 ( .A1(n37239), .A2(n37161), .Z(n37092) );
  CLKNHSV0 U42037 ( .I(n37092), .ZN(n37095) );
  NOR2HSV0 U42038 ( .A1(n42609), .A2(n43880), .ZN(n37093) );
  NOR2HSV2 U42039 ( .A1(n37093), .A2(n37092), .ZN(n37094) );
  AOI31HSV2 U42040 ( .A1(n37236), .A2(n37237), .A3(n37095), .B(n37094), .ZN(
        n37096) );
  NAND2HSV2 U42041 ( .A1(n29707), .A2(n37096), .ZN(n37097) );
  INHSV2 U42042 ( .I(n37099), .ZN(n37100) );
  AOI21HSV4 U42043 ( .A1(n37104), .A2(n37103), .B(n37102), .ZN(n37149) );
  XNOR2HSV4 U42044 ( .A1(n37335), .A2(n37149), .ZN(n37105) );
  CLKAND2HSV2 U42045 ( .A1(n52738), .A2(n37169), .Z(n37145) );
  NAND2HSV2 U42046 ( .A1(n37176), .A2(n37107), .ZN(n37143) );
  INHSV2 U42047 ( .I(n59616), .ZN(n37108) );
  INAND2HSV2 U42048 ( .A1(n37108), .B1(n37353), .ZN(n37141) );
  CLKNAND2HSV0 U42049 ( .A1(n48500), .A2(n42527), .ZN(n37111) );
  CLKNAND2HSV0 U42050 ( .A1(n37109), .A2(\pe3/bq[26] ), .ZN(n37110) );
  XOR2HSV0 U42051 ( .A1(n37111), .A2(n37110), .Z(n37116) );
  INHSV2 U42052 ( .I(n43392), .ZN(n37354) );
  NAND2HSV2 U42053 ( .A1(n37354), .A2(n56213), .ZN(n37114) );
  CLKNAND2HSV0 U42054 ( .A1(\pe3/aot [24]), .A2(n37112), .ZN(n37113) );
  XOR2HSV0 U42055 ( .A1(n37114), .A2(n37113), .Z(n37115) );
  XOR2HSV0 U42056 ( .A1(n37116), .A2(n37115), .Z(n37135) );
  NAND2HSV0 U42057 ( .A1(n42530), .A2(n48496), .ZN(n37118) );
  CLKNAND2HSV1 U42058 ( .A1(n55821), .A2(n37007), .ZN(n37117) );
  XOR2HSV0 U42059 ( .A1(n37118), .A2(n37117), .Z(n37121) );
  INHSV2 U42060 ( .I(n37378), .ZN(n45808) );
  NAND2HSV2 U42061 ( .A1(n45808), .A2(\pe3/pvq [11]), .ZN(n37119) );
  XNOR2HSV1 U42062 ( .A1(n37119), .A2(\pe3/phq [11]), .ZN(n37120) );
  XNOR2HSV1 U42063 ( .A1(n37121), .A2(n37120), .ZN(n37124) );
  CLKNAND2HSV1 U42064 ( .A1(n59618), .A2(n37180), .ZN(n37493) );
  XOR2HSV0 U42065 ( .A1(n37122), .A2(n37493), .Z(n37123) );
  XNOR2HSV1 U42066 ( .A1(n37124), .A2(n37123), .ZN(n37134) );
  NOR2HSV1 U42067 ( .A1(n59606), .A2(n37196), .ZN(n37126) );
  NAND2HSV0 U42068 ( .A1(n59368), .A2(n37298), .ZN(n37125) );
  XOR2HSV0 U42069 ( .A1(n37126), .A2(n37125), .Z(n37130) );
  CLKNAND2HSV1 U42070 ( .A1(n59610), .A2(n43539), .ZN(n37128) );
  CLKNAND2HSV1 U42071 ( .A1(n59612), .A2(n37186), .ZN(n37127) );
  XOR2HSV0 U42072 ( .A1(n37128), .A2(n37127), .Z(n37129) );
  XOR2HSV0 U42073 ( .A1(n37130), .A2(n37129), .Z(n37133) );
  NAND2HSV2 U42074 ( .A1(n37131), .A2(n42673), .ZN(n37132) );
  XOR4HSV1 U42075 ( .A1(n37135), .A2(n37134), .A3(n37133), .A4(n37132), .Z(
        n37137) );
  NAND2HSV2 U42076 ( .A1(n37177), .A2(n59617), .ZN(n37136) );
  XNOR2HSV1 U42077 ( .A1(n37137), .A2(n37136), .ZN(n37139) );
  INHSV2 U42078 ( .I(n43231), .ZN(n42508) );
  XNOR2HSV1 U42079 ( .A1(n37139), .A2(n37138), .ZN(n37140) );
  XOR2HSV0 U42080 ( .A1(n37141), .A2(n37140), .Z(n37142) );
  XOR2HSV0 U42081 ( .A1(n37143), .A2(n37142), .Z(n37144) );
  INHSV4 U42082 ( .I(n37148), .ZN(n53369) );
  INHSV4 U42083 ( .I(n37149), .ZN(n37174) );
  INHSV4 U42084 ( .I(n37174), .ZN(n37222) );
  NOR2HSV4 U42085 ( .A1(n53369), .A2(n37151), .ZN(n37246) );
  NOR2HSV4 U42086 ( .A1(n37148), .A2(n37268), .ZN(n37152) );
  AOI21HSV4 U42087 ( .A1(n37148), .A2(n43469), .B(n43132), .ZN(n37245) );
  INHSV2 U42088 ( .I(n37153), .ZN(n37154) );
  CLKNAND2HSV1 U42089 ( .A1(n37162), .A2(n37161), .ZN(n37159) );
  INHSV2 U42090 ( .I(n37174), .ZN(n37158) );
  INHSV4 U42091 ( .I(n37158), .ZN(n59519) );
  NAND2HSV4 U42092 ( .A1(n37159), .A2(n59519), .ZN(n37160) );
  OAI21HSV4 U42093 ( .A1(n37151), .A2(n53369), .B(n37160), .ZN(n37249) );
  INHSV2 U42094 ( .I(n37248), .ZN(n37163) );
  NAND3HSV4 U42095 ( .A1(n37251), .A2(n37249), .A3(n37163), .ZN(n37267) );
  NAND2HSV2 U42096 ( .A1(n25882), .A2(n37267), .ZN(n42512) );
  XNOR2HSV4 U42097 ( .A1(n37166), .A2(n37165), .ZN(n37414) );
  BUFHSV2 U42098 ( .I(n37168), .Z(n42698) );
  NOR2HSV2 U42099 ( .A1(n42698), .A2(\pe3/ti_7t [12]), .ZN(n42684) );
  NOR2HSV2 U42100 ( .A1(n42684), .A2(n45607), .ZN(n52750) );
  AOI31HSV2 U42101 ( .A1(n37262), .A2(n37261), .A3(n52750), .B(n46559), .ZN(
        n37259) );
  CLKNAND2HSV0 U42102 ( .A1(n37106), .A2(n37169), .ZN(n37172) );
  CLKNAND2HSV0 U42103 ( .A1(n42767), .A2(n37516), .ZN(n37171) );
  BUFHSV2 U42104 ( .I(n43866), .Z(n43613) );
  CLKNAND2HSV1 U42105 ( .A1(n37223), .A2(n43866), .ZN(n37226) );
  BUFHSV2 U42106 ( .I(n55825), .Z(n45949) );
  NAND2HSV2 U42107 ( .A1(n45949), .A2(n36955), .ZN(n37220) );
  CLKNAND2HSV0 U42108 ( .A1(n37176), .A2(n37175), .ZN(n37218) );
  NAND2HSV0 U42109 ( .A1(n37177), .A2(n42770), .ZN(n37214) );
  NAND2HSV0 U42110 ( .A1(n37279), .A2(n37276), .ZN(n37179) );
  NAND2HSV0 U42111 ( .A1(n45695), .A2(n37280), .ZN(n37178) );
  XOR2HSV0 U42112 ( .A1(n37179), .A2(n37178), .Z(n37184) );
  NAND2HSV0 U42113 ( .A1(n56204), .A2(n37180), .ZN(n37182) );
  INHSV2 U42114 ( .I(n45635), .ZN(n55823) );
  CLKNAND2HSV0 U42115 ( .A1(n55823), .A2(n37007), .ZN(n37181) );
  XOR2HSV0 U42116 ( .A1(n37182), .A2(n37181), .Z(n37183) );
  XOR2HSV0 U42117 ( .A1(n37184), .A2(n37183), .Z(n37193) );
  BUFHSV2 U42118 ( .I(n37185), .Z(n42649) );
  INHSV2 U42119 ( .I(n42649), .ZN(n45663) );
  NAND2HSV2 U42120 ( .A1(n59618), .A2(n45663), .ZN(n37188) );
  NAND2HSV0 U42121 ( .A1(n42940), .A2(n37186), .ZN(n37187) );
  XOR2HSV0 U42122 ( .A1(n37188), .A2(n37187), .Z(n37191) );
  CLKNHSV0 U42123 ( .I(n37378), .ZN(n45809) );
  NAND2HSV2 U42124 ( .A1(n45809), .A2(\pe3/pvq [13]), .ZN(n37189) );
  XOR2HSV0 U42125 ( .A1(n37189), .A2(\pe3/phq [13]), .Z(n37190) );
  XOR2HSV0 U42126 ( .A1(n37191), .A2(n37190), .Z(n37192) );
  XOR2HSV0 U42127 ( .A1(n37193), .A2(n37192), .Z(n37195) );
  BUFHSV2 U42128 ( .I(n59648), .Z(n42725) );
  INHSV2 U42129 ( .I(n37275), .ZN(n42999) );
  CLKNAND2HSV1 U42130 ( .A1(n42725), .A2(n42999), .ZN(n37194) );
  XNOR2HSV1 U42131 ( .A1(n37195), .A2(n37194), .ZN(n37211) );
  INHSV1 U42132 ( .I(n37196), .ZN(n56222) );
  CLKNAND2HSV1 U42133 ( .A1(n37362), .A2(n56222), .ZN(n37198) );
  CLKNAND2HSV0 U42134 ( .A1(n37354), .A2(n56218), .ZN(n37197) );
  XOR2HSV0 U42135 ( .A1(n37198), .A2(n37197), .Z(n37202) );
  NAND2HSV0 U42136 ( .A1(n59612), .A2(n37298), .ZN(n37200) );
  CLKNAND2HSV0 U42137 ( .A1(n37373), .A2(n56213), .ZN(n37199) );
  XOR2HSV0 U42138 ( .A1(n37200), .A2(n37199), .Z(n37201) );
  XOR2HSV0 U42139 ( .A1(n37202), .A2(n37201), .Z(n37209) );
  CLKNAND2HSV0 U42140 ( .A1(n36809), .A2(\pe3/bq[25] ), .ZN(n37204) );
  NAND2HSV0 U42141 ( .A1(n37374), .A2(n42530), .ZN(n37203) );
  XOR2HSV0 U42142 ( .A1(n37204), .A2(n37203), .Z(n37207) );
  NAND2HSV2 U42143 ( .A1(n45572), .A2(n42971), .ZN(n42745) );
  NAND2HSV0 U42144 ( .A1(n59610), .A2(\pe3/bq[26] ), .ZN(n37205) );
  XOR2HSV0 U42145 ( .A1(n42745), .A2(n37205), .Z(n37206) );
  XOR2HSV0 U42146 ( .A1(n37207), .A2(n37206), .Z(n37208) );
  XOR2HSV0 U42147 ( .A1(n37209), .A2(n37208), .Z(n37210) );
  XNOR2HSV1 U42148 ( .A1(n37211), .A2(n37210), .ZN(n37213) );
  CLKNAND2HSV0 U42149 ( .A1(n37312), .A2(n42673), .ZN(n37212) );
  XOR3HSV2 U42150 ( .A1(n37214), .A2(n37213), .A3(n37212), .Z(n37216) );
  NAND2HSV0 U42151 ( .A1(n37353), .A2(n59617), .ZN(n37215) );
  XOR2HSV0 U42152 ( .A1(n37216), .A2(n37215), .Z(n37217) );
  XOR2HSV0 U42153 ( .A1(n37218), .A2(n37217), .Z(n37219) );
  XOR2HSV0 U42154 ( .A1(n37220), .A2(n37219), .Z(n37228) );
  CLKNAND2HSV0 U42155 ( .A1(n37226), .A2(n37228), .ZN(n37221) );
  INOR2HSV1 U42156 ( .A1(n37227), .B1(n37221), .ZN(n37225) );
  INHSV4 U42157 ( .I(n37222), .ZN(n47991) );
  INHSV2 U42158 ( .I(n47991), .ZN(n37231) );
  CLKNAND2HSV1 U42159 ( .A1(n37231), .A2(n37223), .ZN(n37224) );
  CLKNAND2HSV1 U42160 ( .A1(n37225), .A2(n37224), .ZN(n37235) );
  CLKNAND2HSV1 U42161 ( .A1(n37227), .A2(n37226), .ZN(n37233) );
  CLKNHSV0 U42162 ( .I(n37228), .ZN(n37232) );
  NOR2HSV1 U42163 ( .A1(n37229), .A2(n37228), .ZN(n37230) );
  AOI22HSV2 U42164 ( .A1(n37233), .A2(n37232), .B1(n37231), .B2(n37230), .ZN(
        n37234) );
  INHSV2 U42165 ( .I(n37239), .ZN(n37331) );
  CLKNAND2HSV2 U42166 ( .A1(n37338), .A2(n37331), .ZN(n37512) );
  CLKNAND2HSV2 U42167 ( .A1(n37240), .A2(n36844), .ZN(n37242) );
  AOI31HSV2 U42168 ( .A1(n37332), .A2(n37242), .A3(n37331), .B(n37241), .ZN(
        n37243) );
  INHSV2 U42169 ( .I(n37251), .ZN(n53372) );
  NOR2HSV0 U42170 ( .A1(n37248), .A2(n37268), .ZN(n37250) );
  NAND3HSV2 U42171 ( .A1(n37251), .A2(n37250), .A3(n37249), .ZN(n37254) );
  INHSV2 U42172 ( .I(\pe3/ti_7t [11]), .ZN(n37252) );
  NOR2HSV2 U42173 ( .A1(n42698), .A2(n37252), .ZN(n42513) );
  CLKNAND2HSV1 U42174 ( .A1(n42513), .A2(n42815), .ZN(n37253) );
  CLKNAND2HSV2 U42175 ( .A1(n37254), .A2(n37253), .ZN(n37255) );
  AOI21HSV4 U42176 ( .A1(n37256), .A2(n53372), .B(n37255), .ZN(n37257) );
  CLKNAND2HSV1 U42177 ( .A1(n47428), .A2(\pe3/ti_7t [13]), .ZN(n37260) );
  CLKNAND2HSV1 U42178 ( .A1(n37262), .A2(n37261), .ZN(n52751) );
  BUFHSV2 U42179 ( .I(n42698), .Z(n43360) );
  NAND2HSV2 U42180 ( .A1(n52750), .A2(n43360), .ZN(n37263) );
  NOR2HSV4 U42181 ( .A1(n52751), .A2(n37263), .ZN(n37347) );
  CLKNAND2HSV2 U42182 ( .A1(n52752), .A2(n37347), .ZN(n37430) );
  CLKNAND2HSV4 U42183 ( .A1(n42584), .A2(n37264), .ZN(n42692) );
  CLKNHSV0 U42184 ( .I(n42692), .ZN(n37345) );
  CLKAND2HSV2 U42185 ( .A1(n37414), .A2(n43360), .Z(n37266) );
  INHSV2 U42186 ( .I(n42513), .ZN(n42509) );
  INHSV2 U42187 ( .I(n36859), .ZN(n43891) );
  NAND3HSV2 U42188 ( .A1(n25882), .A2(n37267), .A3(n42509), .ZN(n37520) );
  NAND3HSV3 U42189 ( .A1(n37520), .A2(n29704), .A3(n43905), .ZN(n37415) );
  INHSV2 U42190 ( .I(n42684), .ZN(n42507) );
  CLKAND2HSV2 U42191 ( .A1(n42507), .A2(n37161), .Z(n37269) );
  NOR2HSV8 U42192 ( .A1(n37271), .A2(n37270), .ZN(n37428) );
  INHSV2 U42193 ( .I(n37273), .ZN(n42936) );
  NAND2HSV2 U42194 ( .A1(n47991), .A2(n42936), .ZN(n37330) );
  BUFHSV3 U42195 ( .I(n55825), .Z(n59626) );
  NAND2HSV2 U42196 ( .A1(n59626), .A2(n42508), .ZN(n37322) );
  NAND2HSV2 U42197 ( .A1(n37457), .A2(n59617), .ZN(n37320) );
  INHSV2 U42198 ( .I(n37275), .ZN(n43262) );
  CLKNAND2HSV1 U42199 ( .A1(n37177), .A2(n43262), .ZN(n37315) );
  NAND2HSV0 U42200 ( .A1(n43034), .A2(n37276), .ZN(n37278) );
  NAND2HSV0 U42201 ( .A1(n37373), .A2(n56222), .ZN(n37277) );
  XOR2HSV0 U42202 ( .A1(n37278), .A2(n37277), .Z(n37284) );
  NAND2HSV0 U42203 ( .A1(n37279), .A2(\pe3/bq[26] ), .ZN(n37282) );
  NAND2HSV0 U42204 ( .A1(n59612), .A2(n37280), .ZN(n37281) );
  XOR2HSV0 U42205 ( .A1(n37282), .A2(n37281), .Z(n37283) );
  XOR2HSV0 U42206 ( .A1(n37284), .A2(n37283), .Z(n37292) );
  INHSV2 U42207 ( .I(\pe3/bq[19] ), .ZN(n46131) );
  CLKNAND2HSV0 U42208 ( .A1(n45572), .A2(\pe3/bq[19] ), .ZN(n37286) );
  NAND2HSV0 U42209 ( .A1(n59610), .A2(\pe3/bq[25] ), .ZN(n37285) );
  XOR2HSV0 U42210 ( .A1(n37286), .A2(n37285), .Z(n37290) );
  NAND2HSV0 U42211 ( .A1(n36809), .A2(\pe3/bq[24] ), .ZN(n37288) );
  NAND2HSV0 U42212 ( .A1(n37354), .A2(\pe3/bq[20] ), .ZN(n37287) );
  XOR2HSV0 U42213 ( .A1(n37288), .A2(n37287), .Z(n37289) );
  XOR2HSV0 U42214 ( .A1(n37290), .A2(n37289), .Z(n37291) );
  XOR2HSV0 U42215 ( .A1(n37292), .A2(n37291), .Z(n37294) );
  CLKNAND2HSV0 U42216 ( .A1(n42725), .A2(n42996), .ZN(n37293) );
  XNOR2HSV1 U42217 ( .A1(n37294), .A2(n37293), .ZN(n37311) );
  INHSV2 U42218 ( .I(n43039), .ZN(n37472) );
  CLKNAND2HSV0 U42219 ( .A1(n37362), .A2(n37472), .ZN(n37296) );
  INHSV2 U42220 ( .I(n42649), .ZN(n43389) );
  NAND2HSV2 U42221 ( .A1(n42940), .A2(n43389), .ZN(n37295) );
  XOR2HSV0 U42222 ( .A1(n37296), .A2(n37295), .Z(n37309) );
  CLKNAND2HSV1 U42223 ( .A1(n46132), .A2(\pe3/pvq [14]), .ZN(n37297) );
  XNOR2HSV1 U42224 ( .A1(n37297), .A2(\pe3/phq [14]), .ZN(n37300) );
  NAND2HSV0 U42225 ( .A1(n59618), .A2(n37298), .ZN(n37299) );
  XNOR2HSV1 U42226 ( .A1(n37300), .A2(n37299), .ZN(n37308) );
  NAND2HSV0 U42227 ( .A1(n37374), .A2(n56213), .ZN(n37302) );
  BUFHSV2 U42228 ( .I(\pe3/bq[31] ), .Z(n48538) );
  NAND2HSV2 U42229 ( .A1(n56204), .A2(n48538), .ZN(n37301) );
  XOR2HSV0 U42230 ( .A1(n37302), .A2(n37301), .Z(n37306) );
  INHSV2 U42231 ( .I(n42833), .ZN(n42540) );
  NAND2HSV2 U42232 ( .A1(n56464), .A2(n42540), .ZN(n37304) );
  CLKNHSV0 U42233 ( .I(n46126), .ZN(n45955) );
  CLKNAND2HSV0 U42234 ( .A1(\pe3/got [19]), .A2(n45955), .ZN(n37303) );
  XOR2HSV0 U42235 ( .A1(n37304), .A2(n37303), .Z(n37305) );
  XOR2HSV0 U42236 ( .A1(n37306), .A2(n37305), .Z(n37307) );
  XOR3HSV2 U42237 ( .A1(n37309), .A2(n37308), .A3(n37307), .Z(n37310) );
  XNOR2HSV1 U42238 ( .A1(n37311), .A2(n37310), .ZN(n37314) );
  NAND2HSV0 U42239 ( .A1(n37312), .A2(n42770), .ZN(n37313) );
  XOR3HSV2 U42240 ( .A1(n37315), .A2(n37314), .A3(n37313), .Z(n37318) );
  NAND2HSV0 U42241 ( .A1(n37316), .A2(n42673), .ZN(n37317) );
  XOR2HSV0 U42242 ( .A1(n37318), .A2(n37317), .Z(n37319) );
  XOR2HSV0 U42243 ( .A1(n37320), .A2(n37319), .Z(n37321) );
  XOR2HSV0 U42244 ( .A1(n37322), .A2(n37321), .Z(n37324) );
  BUFHSV2 U42245 ( .I(n46031), .Z(n42767) );
  CLKNAND2HSV1 U42246 ( .A1(n42767), .A2(n36955), .ZN(n37323) );
  CLKNHSV2 U42247 ( .I(n37106), .ZN(n37326) );
  INHSV2 U42248 ( .I(n37326), .ZN(n59581) );
  INAND2HSV2 U42249 ( .A1(n37326), .B1(n37516), .ZN(n37327) );
  XNOR2HSV1 U42250 ( .A1(n37328), .A2(n37327), .ZN(n37329) );
  XOR2HSV2 U42251 ( .A1(n37330), .A2(n37329), .Z(n37341) );
  CLKNHSV0 U42252 ( .I(n37334), .ZN(n37336) );
  NAND2HSV2 U42253 ( .A1(n37336), .A2(n47992), .ZN(n37337) );
  XNOR2HSV4 U42254 ( .A1(n37343), .A2(n37342), .ZN(n37427) );
  XNOR2HSV4 U42255 ( .A1(n37428), .A2(n37427), .ZN(n37423) );
  CLKNHSV2 U42256 ( .I(n37423), .ZN(n37344) );
  INHSV4 U42257 ( .I(n37344), .ZN(n42690) );
  CLKNAND2HSV3 U42258 ( .A1(n52752), .A2(n37347), .ZN(n37420) );
  INHSV2 U42259 ( .I(n37348), .ZN(n43468) );
  CLKNAND2HSV4 U42260 ( .A1(n37349), .A2(n37430), .ZN(n42706) );
  AND2HSV2 U42261 ( .A1(n42507), .A2(n37272), .Z(n37416) );
  CLKNAND2HSV1 U42262 ( .A1(n37415), .A2(n37416), .ZN(n37350) );
  INHSV2 U42263 ( .I(n37350), .ZN(n37352) );
  NAND2HSV2 U42264 ( .A1(n37352), .A2(n37351), .ZN(n37413) );
  NAND2HSV2 U42265 ( .A1(n47991), .A2(n37516), .ZN(n37407) );
  CLKNAND2HSV1 U42266 ( .A1(n37457), .A2(n42673), .ZN(n37399) );
  BUFHSV2 U42267 ( .I(n37353), .Z(n59621) );
  NAND2HSV2 U42268 ( .A1(n59621), .A2(n55821), .ZN(n37397) );
  BUFHSV2 U42269 ( .I(n37177), .Z(n42710) );
  CLKNAND2HSV1 U42270 ( .A1(n42710), .A2(n55823), .ZN(n37395) );
  CLKNHSV0 U42271 ( .I(n42843), .ZN(n59622) );
  NAND2HSV0 U42272 ( .A1(n59622), .A2(n56213), .ZN(n37356) );
  NAND2HSV0 U42273 ( .A1(n37354), .A2(\pe3/bq[19] ), .ZN(n37355) );
  XOR2HSV0 U42274 ( .A1(n37356), .A2(n37355), .Z(n37361) );
  NAND2HSV0 U42275 ( .A1(n59610), .A2(\pe3/bq[24] ), .ZN(n37359) );
  CLKNAND2HSV0 U42276 ( .A1(\pe3/aot [20]), .A2(n43389), .ZN(n37358) );
  XOR2HSV0 U42277 ( .A1(n37359), .A2(n37358), .Z(n37360) );
  XOR2HSV0 U42278 ( .A1(n37361), .A2(n37360), .Z(n37370) );
  NAND2HSV0 U42279 ( .A1(n45695), .A2(\pe3/bq[26] ), .ZN(n37364) );
  NAND2HSV0 U42280 ( .A1(n37362), .A2(\pe3/bq[20] ), .ZN(n37363) );
  XOR2HSV0 U42281 ( .A1(n37364), .A2(n37363), .Z(n37368) );
  NAND2HSV0 U42282 ( .A1(n59368), .A2(\pe3/bq[25] ), .ZN(n37366) );
  CLKNAND2HSV1 U42283 ( .A1(n56349), .A2(n42540), .ZN(n37365) );
  XOR2HSV0 U42284 ( .A1(n37366), .A2(n37365), .Z(n37367) );
  XOR2HSV0 U42285 ( .A1(n37368), .A2(n37367), .Z(n37369) );
  XOR2HSV0 U42286 ( .A1(n37370), .A2(n37369), .Z(n37372) );
  CLKNAND2HSV0 U42287 ( .A1(n42725), .A2(n42937), .ZN(n37371) );
  XNOR2HSV1 U42288 ( .A1(n37372), .A2(n37371), .ZN(n37392) );
  CLKNAND2HSV1 U42289 ( .A1(n37373), .A2(n37472), .ZN(n42549) );
  NAND2HSV0 U42290 ( .A1(n37374), .A2(n56222), .ZN(n37375) );
  XOR2HSV0 U42291 ( .A1(n42549), .A2(n37375), .Z(n37390) );
  NAND2HSV0 U42292 ( .A1(n59618), .A2(n42634), .ZN(n37377) );
  CLKNAND2HSV0 U42293 ( .A1(\pe3/aot [19]), .A2(n48538), .ZN(n37376) );
  XOR2HSV0 U42294 ( .A1(n37377), .A2(n37376), .Z(n37381) );
  CLKNHSV0 U42295 ( .I(n37378), .ZN(n46129) );
  NAND2HSV2 U42296 ( .A1(n46129), .A2(\pe3/pvq [15]), .ZN(n37379) );
  XNOR2HSV1 U42297 ( .A1(n37379), .A2(\pe3/phq [15]), .ZN(n37380) );
  XNOR2HSV1 U42298 ( .A1(n37381), .A2(n37380), .ZN(n37389) );
  NAND2HSV0 U42299 ( .A1(n42940), .A2(n48527), .ZN(n37383) );
  NAND2HSV0 U42300 ( .A1(n43374), .A2(n37007), .ZN(n37382) );
  XOR2HSV0 U42301 ( .A1(n37383), .A2(n37382), .Z(n37387) );
  CLKNHSV0 U42302 ( .I(n45525), .ZN(n42653) );
  NAND2HSV0 U42303 ( .A1(n59612), .A2(n42653), .ZN(n37385) );
  NAND2HSV0 U42304 ( .A1(n45572), .A2(\pe3/bq[18] ), .ZN(n37384) );
  XOR2HSV0 U42305 ( .A1(n37385), .A2(n37384), .Z(n37386) );
  XOR2HSV0 U42306 ( .A1(n37387), .A2(n37386), .Z(n37388) );
  XOR3HSV2 U42307 ( .A1(n37390), .A2(n37389), .A3(n37388), .Z(n37391) );
  XNOR2HSV1 U42308 ( .A1(n37392), .A2(n37391), .ZN(n37394) );
  BUFHSV2 U42309 ( .I(n37312), .Z(n59671) );
  BUFHSV2 U42310 ( .I(n59671), .Z(n43516) );
  CLKNAND2HSV1 U42311 ( .A1(n43516), .A2(n42520), .ZN(n37393) );
  XOR3HSV2 U42312 ( .A1(n37395), .A2(n37394), .A3(n37393), .Z(n37396) );
  XNOR2HSV1 U42313 ( .A1(n37397), .A2(n37396), .ZN(n37398) );
  XNOR2HSV1 U42314 ( .A1(n37399), .A2(n37398), .ZN(n37401) );
  CLKAND2HSV1 U42315 ( .A1(n55825), .A2(\pe3/got [24]), .Z(n37400) );
  XNOR2HSV1 U42316 ( .A1(n37401), .A2(n37400), .ZN(n37403) );
  CLKNAND2HSV1 U42317 ( .A1(n42767), .A2(n42508), .ZN(n37402) );
  INAND2HSV2 U42318 ( .A1(n37326), .B1(n46311), .ZN(n37404) );
  XNOR2HSV1 U42319 ( .A1(n37407), .A2(n37406), .ZN(n37410) );
  CLKNAND2HSV1 U42320 ( .A1(n37408), .A2(n42936), .ZN(n37409) );
  XOR2HSV0 U42321 ( .A1(n37410), .A2(n37409), .Z(n37411) );
  NAND2HSV2 U42322 ( .A1(n42682), .A2(n37414), .ZN(n37455) );
  NAND3HSV2 U42323 ( .A1(n37455), .A2(n37416), .A3(n37415), .ZN(n37417) );
  OAI21HSV2 U42324 ( .A1(n37433), .A2(n43468), .B(n36972), .ZN(n37418) );
  CLKNHSV1 U42325 ( .I(n42700), .ZN(n42496) );
  NOR2HSV0 U42326 ( .A1(n42599), .A2(n42496), .ZN(n37442) );
  INHSV2 U42327 ( .I(n37422), .ZN(n37429) );
  CLKNHSV0 U42328 ( .I(\pe3/ti_7t [14]), .ZN(n37424) );
  NAND2HSV0 U42329 ( .A1(n37424), .A2(n45618), .ZN(n42702) );
  AND2HSV2 U42330 ( .A1(n42702), .A2(n36671), .Z(n37425) );
  CLKNAND2HSV4 U42331 ( .A1(n37426), .A2(n37425), .ZN(n42594) );
  INHSV4 U42332 ( .I(n42594), .ZN(n37432) );
  XNOR2HSV4 U42333 ( .A1(n37428), .A2(n37427), .ZN(n37443) );
  INHSV4 U42334 ( .I(n37443), .ZN(n42592) );
  CLKNAND2HSV1 U42335 ( .A1(n37430), .A2(n37429), .ZN(n42591) );
  INHSV2 U42336 ( .I(n42600), .ZN(n53378) );
  INHSV2 U42337 ( .I(n53378), .ZN(n37441) );
  CLKNHSV0 U42338 ( .I(n45931), .ZN(n52726) );
  OAI21HSV0 U42339 ( .A1(n42600), .A2(n42496), .B(n52726), .ZN(n37440) );
  INHSV2 U42340 ( .I(n37433), .ZN(n37434) );
  NOR2HSV1 U42341 ( .A1(n42492), .A2(n43483), .ZN(n37438) );
  INHSV2 U42342 ( .I(n42595), .ZN(n37436) );
  CLKNHSV0 U42343 ( .I(n42493), .ZN(n37437) );
  CLKNAND2HSV2 U42344 ( .A1(n37438), .A2(n37437), .ZN(n37439) );
  AOI22HSV4 U42345 ( .A1(n37442), .A2(n37441), .B1(n37440), .B2(n37439), .ZN(
        n37527) );
  NOR2HSV4 U42346 ( .A1(n37443), .A2(n42609), .ZN(n37444) );
  CLKNAND2HSV3 U42347 ( .A1(n37444), .A2(n42706), .ZN(n42500) );
  CLKNHSV1 U42348 ( .I(n42702), .ZN(n42501) );
  NOR2HSV1 U42349 ( .A1(n42501), .A2(n59615), .ZN(n37445) );
  CLKNAND2HSV2 U42350 ( .A1(n42500), .A2(n37445), .ZN(n37446) );
  NAND2HSV2 U42351 ( .A1(n42693), .A2(n46519), .ZN(n37448) );
  CLKNAND2HSV1 U42352 ( .A1(n29704), .A2(n42698), .ZN(n37451) );
  BUFHSV2 U42353 ( .I(n37784), .Z(n43873) );
  NOR2HSV2 U42354 ( .A1(n42684), .A2(n43873), .ZN(n37452) );
  NOR2HSV2 U42355 ( .A1(n37455), .A2(n37454), .ZN(n42506) );
  NOR2HSV2 U42356 ( .A1(n37456), .A2(n42506), .ZN(n37524) );
  CLKNAND2HSV1 U42357 ( .A1(n37151), .A2(n59616), .ZN(n37519) );
  NAND2HSV0 U42358 ( .A1(n49405), .A2(n42673), .ZN(n37466) );
  CLKNAND2HSV0 U42359 ( .A1(n37457), .A2(n42770), .ZN(n37464) );
  CLKNAND2HSV1 U42360 ( .A1(n59621), .A2(n42520), .ZN(n37462) );
  NAND2HSV2 U42361 ( .A1(n42710), .A2(n56489), .ZN(n37458) );
  XNOR2HSV1 U42362 ( .A1(n37458), .A2(\pe3/phq [16]), .ZN(n37460) );
  CLKNAND2HSV1 U42363 ( .A1(n43516), .A2(n55823), .ZN(n37459) );
  XOR2HSV0 U42364 ( .A1(n37460), .A2(n37459), .Z(n37461) );
  XOR2HSV0 U42365 ( .A1(n37462), .A2(n37461), .Z(n37463) );
  XOR2HSV0 U42366 ( .A1(n37464), .A2(n37463), .Z(n37465) );
  XNOR2HSV1 U42367 ( .A1(n37466), .A2(n37465), .ZN(n37469) );
  CLKNHSV0 U42368 ( .I(n37469), .ZN(n37467) );
  NOR2HSV1 U42369 ( .A1(n37467), .A2(n37785), .ZN(n37471) );
  NOR2HSV0 U42370 ( .A1(n37326), .A2(n37785), .ZN(n37468) );
  NOR2HSV1 U42371 ( .A1(n37469), .A2(n37468), .ZN(n37470) );
  AOI21HSV2 U42372 ( .A1(n37471), .A2(n59581), .B(n37470), .ZN(n37510) );
  CLKNAND2HSV1 U42373 ( .A1(n42767), .A2(n43452), .ZN(n37508) );
  CLKNHSV0 U42374 ( .I(n45555), .ZN(n45554) );
  NAND2HSV2 U42375 ( .A1(n45554), .A2(n37472), .ZN(n37474) );
  CLKNHSV0 U42376 ( .I(n42821), .ZN(n43528) );
  INHSV2 U42377 ( .I(n55755), .ZN(n42642) );
  CLKNAND2HSV1 U42378 ( .A1(n43528), .A2(n42642), .ZN(n37473) );
  XOR2HSV0 U42379 ( .A1(n37474), .A2(n37473), .Z(n37478) );
  NAND2HSV2 U42380 ( .A1(\pe3/aot [24]), .A2(n42527), .ZN(n37476) );
  CLKNAND2HSV0 U42381 ( .A1(n42743), .A2(n56213), .ZN(n37475) );
  XOR2HSV0 U42382 ( .A1(n37476), .A2(n37475), .Z(n37477) );
  XOR2HSV0 U42383 ( .A1(n37478), .A2(n37477), .Z(n37486) );
  NAND2HSV2 U42384 ( .A1(n43547), .A2(\pe3/bq[18] ), .ZN(n37480) );
  NAND2HSV0 U42385 ( .A1(n59368), .A2(\pe3/bq[24] ), .ZN(n37479) );
  XOR2HSV0 U42386 ( .A1(n37480), .A2(n37479), .Z(n37484) );
  CLKNAND2HSV1 U42387 ( .A1(n42818), .A2(\pe3/bq[26] ), .ZN(n37482) );
  NAND2HSV2 U42388 ( .A1(n42950), .A2(n48538), .ZN(n37481) );
  XOR2HSV0 U42389 ( .A1(n37482), .A2(n37481), .Z(n37483) );
  XOR2HSV0 U42390 ( .A1(n37484), .A2(n37483), .Z(n37485) );
  XOR2HSV0 U42391 ( .A1(n37486), .A2(n37485), .Z(n37488) );
  CLKNAND2HSV1 U42392 ( .A1(n42725), .A2(\pe3/got [18]), .ZN(n37487) );
  XNOR2HSV1 U42393 ( .A1(n37488), .A2(n37487), .ZN(n37506) );
  CLKNHSV0 U42394 ( .I(n43757), .ZN(n43650) );
  NAND2HSV2 U42395 ( .A1(n43650), .A2(\pe3/bq[19] ), .ZN(n42738) );
  INHSV2 U42396 ( .I(n42835), .ZN(n42728) );
  INHSV2 U42397 ( .I(n42649), .ZN(n48522) );
  NAND2HSV2 U42398 ( .A1(n42728), .A2(n48522), .ZN(n37489) );
  XOR2HSV0 U42399 ( .A1(n42738), .A2(n37489), .Z(n37504) );
  NAND2HSV0 U42400 ( .A1(n56204), .A2(n48527), .ZN(n37491) );
  BUFHSV2 U42401 ( .I(n46141), .Z(n43059) );
  INHSV2 U42402 ( .I(n46613), .ZN(n46124) );
  NAND2HSV2 U42403 ( .A1(n46124), .A2(\pe3/pvq [16]), .ZN(n37490) );
  XOR2HSV0 U42404 ( .A1(n37491), .A2(n37490), .Z(n37495) );
  NAND2HSV2 U42405 ( .A1(n46363), .A2(n42653), .ZN(n42842) );
  OAI22HSV0 U42406 ( .A1(n42833), .A2(n43527), .B1(n45567), .B2(n45525), .ZN(
        n37492) );
  OAI21HSV0 U42407 ( .A1(n37493), .A2(n42842), .B(n37492), .ZN(n37494) );
  XNOR2HSV1 U42408 ( .A1(n37495), .A2(n37494), .ZN(n37503) );
  NOR2HSV0 U42409 ( .A1(n42539), .A2(n45649), .ZN(n37497) );
  CLKNAND2HSV1 U42410 ( .A1(n56064), .A2(n45955), .ZN(n37496) );
  XOR2HSV0 U42411 ( .A1(n37497), .A2(n37496), .Z(n37501) );
  INHSV2 U42412 ( .I(n37196), .ZN(n43146) );
  NAND2HSV2 U42413 ( .A1(n59622), .A2(n43146), .ZN(n37499) );
  INHSV2 U42414 ( .I(n36989), .ZN(n45648) );
  CLKNAND2HSV1 U42415 ( .A1(n45648), .A2(n42971), .ZN(n37498) );
  XOR2HSV0 U42416 ( .A1(n37499), .A2(n37498), .Z(n37500) );
  XOR2HSV0 U42417 ( .A1(n37501), .A2(n37500), .Z(n37502) );
  XOR3HSV2 U42418 ( .A1(n37504), .A2(n37503), .A3(n37502), .Z(n37505) );
  XNOR2HSV1 U42419 ( .A1(n37506), .A2(n37505), .ZN(n37507) );
  XNOR2HSV1 U42420 ( .A1(n37508), .A2(n37507), .ZN(n37509) );
  XOR2HSV0 U42421 ( .A1(n37510), .A2(n37509), .Z(n37511) );
  CLKNHSV2 U42422 ( .I(n37511), .ZN(n37518) );
  INHSV2 U42423 ( .I(n37512), .ZN(n37515) );
  CLKNAND2HSV1 U42424 ( .A1(n37513), .A2(n47992), .ZN(n37514) );
  NAND2HSV4 U42425 ( .A1(n37515), .A2(n37514), .ZN(n43622) );
  CLKNAND2HSV2 U42426 ( .A1(n43622), .A2(n37516), .ZN(n37517) );
  XOR3HSV2 U42427 ( .A1(n37519), .A2(n37518), .A3(n37517), .Z(n37522) );
  XNOR2HSV4 U42428 ( .A1(n37522), .A2(n37521), .ZN(n37523) );
  XNOR2HSV4 U42429 ( .A1(n37524), .A2(n37523), .ZN(n37526) );
  NOR2HSV1 U42430 ( .A1(n37529), .A2(n39379), .ZN(n37764) );
  CLKNHSV2 U42431 ( .I(n37530), .ZN(n37542) );
  NOR2HSV2 U42432 ( .A1(n37532), .A2(n37534), .ZN(n37539) );
  CLKNHSV2 U42433 ( .I(n37533), .ZN(n37538) );
  INHSV2 U42434 ( .I(n37534), .ZN(n37535) );
  NAND3HSV4 U42435 ( .A1(n37545), .A2(n37542), .A3(n37765), .ZN(n39413) );
  CLKNHSV0 U42436 ( .I(\pe5/ti_7t [21]), .ZN(n37543) );
  CLKNAND2HSV0 U42437 ( .A1(n37543), .A2(n39239), .ZN(n37771) );
  NAND2HSV0 U42438 ( .A1(n37771), .A2(n37544), .ZN(n39354) );
  NOR2HSV2 U42439 ( .A1(n39354), .A2(n37638), .ZN(n39390) );
  CLKNAND2HSV2 U42440 ( .A1(n39413), .A2(n39390), .ZN(n37649) );
  NOR2HSV3 U42441 ( .A1(n37545), .A2(n37766), .ZN(n37546) );
  CLKNAND2HSV3 U42442 ( .A1(n37546), .A2(n37769), .ZN(n37547) );
  NOR2HSV2 U42443 ( .A1(n37754), .A2(n37551), .ZN(n37552) );
  NAND2HSV2 U42444 ( .A1(n37552), .A2(n37756), .ZN(n37553) );
  NAND2HSV2 U42445 ( .A1(n39251), .A2(n37554), .ZN(n39218) );
  INHSV2 U42446 ( .I(n39118), .ZN(n59525) );
  NAND2HSV2 U42447 ( .A1(n59525), .A2(n48742), .ZN(n37634) );
  BUFHSV2 U42448 ( .I(n39120), .Z(n45820) );
  NAND2HSV2 U42449 ( .A1(n45820), .A2(n31148), .ZN(n37629) );
  NAND2HSV0 U42450 ( .A1(n37657), .A2(\pe5/got [22]), .ZN(n37627) );
  CLKNAND2HSV1 U42451 ( .A1(n30781), .A2(n37656), .ZN(n37625) );
  CLKNAND2HSV1 U42452 ( .A1(n40172), .A2(n45816), .ZN(n37623) );
  NAND2HSV0 U42453 ( .A1(n39258), .A2(n37556), .ZN(n37621) );
  CLKNAND2HSV0 U42454 ( .A1(n37558), .A2(n37557), .ZN(n37616) );
  NAND2HSV2 U42455 ( .A1(n31151), .A2(n39516), .ZN(n37614) );
  NAND2HSV2 U42456 ( .A1(n39466), .A2(n39259), .ZN(n37577) );
  XOR2HSV0 U42457 ( .A1(n37560), .A2(n37559), .Z(n37573) );
  OAI22HSV0 U42458 ( .A1(n44704), .A2(n46134), .B1(n45451), .B2(n45460), .ZN(
        n37561) );
  OAI21HSV1 U42459 ( .A1(n37562), .A2(n39263), .B(n37561), .ZN(n37563) );
  NOR2HSV0 U42460 ( .A1(n48204), .A2(n39166), .ZN(n48812) );
  XNOR2HSV1 U42461 ( .A1(n37563), .A2(n48812), .ZN(n37572) );
  NAND2HSV0 U42462 ( .A1(n39446), .A2(n30692), .ZN(n37566) );
  NAND2HSV0 U42463 ( .A1(n30788), .A2(n47305), .ZN(n37565) );
  XOR2HSV0 U42464 ( .A1(n37566), .A2(n37565), .Z(n37570) );
  CLKNHSV0 U42465 ( .I(n45844), .ZN(n39480) );
  CLKNAND2HSV0 U42466 ( .A1(n37700), .A2(n39480), .ZN(n37568) );
  NAND2HSV0 U42467 ( .A1(n59640), .A2(n48787), .ZN(n37567) );
  XOR2HSV0 U42468 ( .A1(n37568), .A2(n37567), .Z(n37569) );
  XOR2HSV0 U42469 ( .A1(n37570), .A2(n37569), .Z(n37571) );
  XOR3HSV2 U42470 ( .A1(n37573), .A2(n37572), .A3(n37571), .Z(n37575) );
  NAND2HSV0 U42471 ( .A1(n39278), .A2(n48167), .ZN(n37574) );
  XNOR2HSV1 U42472 ( .A1(n37575), .A2(n37574), .ZN(n37576) );
  XNOR2HSV1 U42473 ( .A1(n37577), .A2(n37576), .ZN(n37612) );
  NAND2HSV0 U42474 ( .A1(n59366), .A2(n39592), .ZN(n37579) );
  NAND2HSV0 U42475 ( .A1(n48658), .A2(n39436), .ZN(n37578) );
  XOR2HSV0 U42476 ( .A1(n37579), .A2(n37578), .Z(n37583) );
  NAND2HSV0 U42477 ( .A1(n51022), .A2(n40207), .ZN(n37581) );
  CLKNAND2HSV0 U42478 ( .A1(\pe5/aot [23]), .A2(n37685), .ZN(n37580) );
  XOR2HSV0 U42479 ( .A1(n37581), .A2(n37580), .Z(n37582) );
  XOR2HSV0 U42480 ( .A1(n37583), .A2(n37582), .Z(n37592) );
  CLKNAND2HSV1 U42481 ( .A1(n39266), .A2(n53314), .ZN(n37586) );
  NAND2HSV0 U42482 ( .A1(\pe5/got [11]), .A2(n37584), .ZN(n37585) );
  XOR2HSV0 U42483 ( .A1(n37586), .A2(n37585), .Z(n37590) );
  CLKNAND2HSV0 U42484 ( .A1(n39269), .A2(n39921), .ZN(n37588) );
  NAND2HSV0 U42485 ( .A1(n39490), .A2(n39130), .ZN(n37587) );
  XOR2HSV0 U42486 ( .A1(n37588), .A2(n37587), .Z(n37589) );
  XOR2HSV0 U42487 ( .A1(n37590), .A2(n37589), .Z(n37591) );
  XOR2HSV0 U42488 ( .A1(n37592), .A2(n37591), .Z(n37607) );
  NOR2HSV0 U42489 ( .A1(n48175), .A2(n39796), .ZN(n37594) );
  NAND2HSV0 U42490 ( .A1(\pe5/aot [13]), .A2(n39495), .ZN(n37593) );
  XOR2HSV0 U42491 ( .A1(n37594), .A2(n37593), .Z(n37599) );
  NAND2HSV0 U42492 ( .A1(n59943), .A2(n45470), .ZN(n37597) );
  CLKNAND2HSV1 U42493 ( .A1(n59938), .A2(n40221), .ZN(n37596) );
  XOR2HSV0 U42494 ( .A1(n37597), .A2(n37596), .Z(n37598) );
  XOR2HSV0 U42495 ( .A1(n37599), .A2(n37598), .Z(n37605) );
  NAND2HSV0 U42496 ( .A1(n37707), .A2(\pe5/pvq [22]), .ZN(n37600) );
  XOR2HSV0 U42497 ( .A1(n37600), .A2(\pe5/phq [22]), .Z(n37603) );
  CLKNAND2HSV1 U42498 ( .A1(n39629), .A2(n52619), .ZN(n37662) );
  OAI22HSV0 U42499 ( .A1(n39779), .A2(n50428), .B1(n39123), .B2(n48050), .ZN(
        n37601) );
  OAI21HSV1 U42500 ( .A1(n37662), .A2(n40045), .B(n37601), .ZN(n37602) );
  XOR2HSV0 U42501 ( .A1(n37603), .A2(n37602), .Z(n37604) );
  XNOR2HSV1 U42502 ( .A1(n37605), .A2(n37604), .ZN(n37606) );
  XNOR2HSV1 U42503 ( .A1(n37607), .A2(n37606), .ZN(n37610) );
  BUFHSV2 U42504 ( .I(n37608), .Z(n48014) );
  CLKNHSV0 U42505 ( .I(n45817), .ZN(n39435) );
  CLKNAND2HSV1 U42506 ( .A1(n48014), .A2(n39435), .ZN(n37609) );
  XNOR2HSV1 U42507 ( .A1(n37610), .A2(n37609), .ZN(n37611) );
  XNOR2HSV1 U42508 ( .A1(n37612), .A2(n37611), .ZN(n37613) );
  XNOR2HSV1 U42509 ( .A1(n37614), .A2(n37613), .ZN(n37615) );
  XNOR2HSV1 U42510 ( .A1(n37616), .A2(n37615), .ZN(n37619) );
  CLKNAND2HSV1 U42511 ( .A1(n37723), .A2(n37725), .ZN(n37618) );
  NAND2HSV0 U42512 ( .A1(n47058), .A2(n37658), .ZN(n37617) );
  XOR3HSV2 U42513 ( .A1(n37619), .A2(n37618), .A3(n37617), .Z(n37620) );
  XNOR2HSV1 U42514 ( .A1(n37621), .A2(n37620), .ZN(n37622) );
  XNOR2HSV1 U42515 ( .A1(n37623), .A2(n37622), .ZN(n37624) );
  XOR2HSV0 U42516 ( .A1(n37625), .A2(n37624), .Z(n37626) );
  XNOR2HSV1 U42517 ( .A1(n37627), .A2(n37626), .ZN(n37628) );
  XOR2HSV0 U42518 ( .A1(n37629), .A2(n37628), .Z(n37633) );
  BUFHSV2 U42519 ( .I(n45819), .Z(n39257) );
  NAND2HSV2 U42520 ( .A1(n39257), .A2(n37631), .ZN(n37632) );
  CLKNHSV0 U42521 ( .I(n30596), .ZN(n37635) );
  XNOR2HSV4 U42522 ( .A1(n37637), .A2(n37636), .ZN(n37641) );
  NOR2HSV2 U42523 ( .A1(n40130), .A2(n37638), .ZN(n40133) );
  AOI22HSV2 U42524 ( .A1(n30142), .A2(n37639), .B1(n60054), .B2(n40133), .ZN(
        n37640) );
  XNOR2HSV4 U42525 ( .A1(n37641), .A2(n37640), .ZN(n37644) );
  XNOR2HSV4 U42526 ( .A1(n37644), .A2(n37643), .ZN(n39228) );
  XNOR2HSV4 U42527 ( .A1(n39228), .A2(n39218), .ZN(n37646) );
  NOR2HSV2 U42528 ( .A1(n37645), .A2(\pe5/ti_7t [22]), .ZN(n39418) );
  NOR2HSV2 U42529 ( .A1(n39418), .A2(n39733), .ZN(n37647) );
  CLKNAND2HSV2 U42530 ( .A1(n37646), .A2(n37647), .ZN(n37650) );
  CLKNAND2HSV1 U42531 ( .A1(n37647), .A2(n39730), .ZN(n37648) );
  NAND2HSV3 U42532 ( .A1(n37650), .A2(n29693), .ZN(n39680) );
  NOR2HSV4 U42533 ( .A1(n39389), .A2(n39671), .ZN(n37651) );
  INHSV4 U42534 ( .I(n37651), .ZN(n39681) );
  INHSV2 U42535 ( .I(n37652), .ZN(n39431) );
  INHSV2 U42536 ( .I(n39431), .ZN(n39256) );
  NAND2HSV2 U42537 ( .A1(n39256), .A2(n30596), .ZN(n37748) );
  CLKNAND2HSV1 U42538 ( .A1(n59525), .A2(n48739), .ZN(n37744) );
  BUFHSV2 U42539 ( .I(n37653), .Z(n39840) );
  CLKNHSV0 U42540 ( .I(n37654), .ZN(n37655) );
  NOR2HSV2 U42541 ( .A1(n39840), .A2(n37655), .ZN(n37742) );
  CLKNAND2HSV1 U42542 ( .A1(n39257), .A2(n31148), .ZN(n37740) );
  CLKNAND2HSV1 U42543 ( .A1(n45820), .A2(n39532), .ZN(n37738) );
  NAND2HSV0 U42544 ( .A1(n37657), .A2(n37656), .ZN(n37736) );
  CLKNAND2HSV1 U42545 ( .A1(n40171), .A2(n45816), .ZN(n37734) );
  CLKNAND2HSV0 U42546 ( .A1(n40172), .A2(n39432), .ZN(n37732) );
  NAND2HSV0 U42547 ( .A1(n39258), .A2(n37658), .ZN(n37730) );
  CLKNAND2HSV1 U42548 ( .A1(n48168), .A2(n39516), .ZN(n37722) );
  CLKNAND2HSV1 U42549 ( .A1(n59639), .A2(n39259), .ZN(n37720) );
  CLKNAND2HSV0 U42550 ( .A1(n39466), .A2(n39435), .ZN(n37682) );
  INHSV2 U42551 ( .I(n50507), .ZN(n59896) );
  NAND2HSV0 U42552 ( .A1(n59896), .A2(n39495), .ZN(n48657) );
  CLKNHSV0 U42553 ( .I(n48822), .ZN(n39443) );
  NAND2HSV0 U42554 ( .A1(n37660), .A2(n39443), .ZN(n37661) );
  XOR2HSV0 U42555 ( .A1(n48657), .A2(n37661), .Z(n37678) );
  CLKNAND2HSV1 U42556 ( .A1(\pe5/aot [11]), .A2(n52619), .ZN(n46932) );
  OAI21HSV0 U42557 ( .A1(n30223), .A2(n48204), .B(n37662), .ZN(n37663) );
  OAI21HSV0 U42558 ( .A1(n37664), .A2(n46932), .B(n37663), .ZN(n37669) );
  CLKNAND2HSV0 U42559 ( .A1(\pe5/aot [13]), .A2(\pe5/bq[15] ), .ZN(n47225) );
  NOR2HSV0 U42560 ( .A1(n37665), .A2(n47225), .ZN(n37667) );
  INHSV2 U42561 ( .I(n51057), .ZN(n50500) );
  AOI22HSV0 U42562 ( .A1(n39801), .A2(n50500), .B1(n39130), .B2(\pe5/aot [13]), 
        .ZN(n37666) );
  NOR2HSV2 U42563 ( .A1(n37667), .A2(n37666), .ZN(n37668) );
  XNOR2HSV1 U42564 ( .A1(n37669), .A2(n37668), .ZN(n37677) );
  INHSV2 U42565 ( .I(n46961), .ZN(n52571) );
  NAND2HSV0 U42566 ( .A1(n52571), .A2(n37584), .ZN(n37671) );
  NAND2HSV0 U42567 ( .A1(n59366), .A2(n48170), .ZN(n37670) );
  XOR2HSV0 U42568 ( .A1(n37671), .A2(n37670), .Z(n37675) );
  NAND2HSV0 U42569 ( .A1(\pe5/aot [16]), .A2(n52594), .ZN(n37673) );
  NAND2HSV0 U42570 ( .A1(n51022), .A2(n52585), .ZN(n37672) );
  XOR2HSV0 U42571 ( .A1(n37673), .A2(n37672), .Z(n37674) );
  XOR2HSV0 U42572 ( .A1(n37675), .A2(n37674), .Z(n37676) );
  XOR3HSV2 U42573 ( .A1(n37678), .A2(n37677), .A3(n37676), .Z(n37680) );
  NAND2HSV0 U42574 ( .A1(n39278), .A2(n59643), .ZN(n37679) );
  XNOR2HSV1 U42575 ( .A1(n37680), .A2(n37679), .ZN(n37681) );
  XNOR2HSV1 U42576 ( .A1(n37682), .A2(n37681), .ZN(n37718) );
  CLKNAND2HSV0 U42577 ( .A1(n59642), .A2(n31192), .ZN(n37684) );
  NAND2HSV0 U42578 ( .A1(n39490), .A2(n45470), .ZN(n37683) );
  XOR2HSV0 U42579 ( .A1(n37684), .A2(n37683), .Z(n37689) );
  CLKNAND2HSV0 U42580 ( .A1(n39473), .A2(\pe5/bq[16] ), .ZN(n37687) );
  NAND2HSV0 U42581 ( .A1(n39444), .A2(n37685), .ZN(n37686) );
  XOR2HSV0 U42582 ( .A1(n37687), .A2(n37686), .Z(n37688) );
  XOR2HSV0 U42583 ( .A1(n37689), .A2(n37688), .Z(n37697) );
  NAND2HSV0 U42584 ( .A1(n39269), .A2(n52595), .ZN(n37691) );
  NAND2HSV0 U42585 ( .A1(\pe5/aot [23]), .A2(n39454), .ZN(n37690) );
  XOR2HSV0 U42586 ( .A1(n37691), .A2(n37690), .Z(n37695) );
  NAND2HSV0 U42587 ( .A1(n30788), .A2(n39480), .ZN(n37693) );
  NAND2HSV0 U42588 ( .A1(n39446), .A2(n31160), .ZN(n37692) );
  XOR2HSV0 U42589 ( .A1(n37693), .A2(n37692), .Z(n37694) );
  XOR2HSV0 U42590 ( .A1(n37695), .A2(n37694), .Z(n37696) );
  XOR2HSV0 U42591 ( .A1(n37697), .A2(n37696), .Z(n37714) );
  NAND2HSV0 U42592 ( .A1(n39266), .A2(n39472), .ZN(n37699) );
  NAND2HSV0 U42593 ( .A1(n50653), .A2(n48787), .ZN(n37698) );
  XOR2HSV0 U42594 ( .A1(n37699), .A2(n37698), .Z(n37704) );
  NAND2HSV0 U42595 ( .A1(\pe5/aot [18]), .A2(n30692), .ZN(n37702) );
  CLKNAND2HSV1 U42596 ( .A1(n48242), .A2(n39445), .ZN(n37701) );
  XOR2HSV0 U42597 ( .A1(n37702), .A2(n37701), .Z(n37703) );
  XOR2HSV0 U42598 ( .A1(n37704), .A2(n37703), .Z(n37712) );
  CLKNAND2HSV0 U42599 ( .A1(n59938), .A2(n39471), .ZN(n37706) );
  CLKNHSV0 U42600 ( .I(n39779), .ZN(n39455) );
  CLKNAND2HSV0 U42601 ( .A1(n39455), .A2(n39592), .ZN(n37705) );
  XOR2HSV0 U42602 ( .A1(n37706), .A2(n37705), .Z(n37710) );
  NAND2HSV0 U42603 ( .A1(n37707), .A2(\pe5/pvq [23]), .ZN(n37708) );
  XOR2HSV0 U42604 ( .A1(n37708), .A2(\pe5/phq [23]), .Z(n37709) );
  XOR2HSV0 U42605 ( .A1(n37710), .A2(n37709), .Z(n37711) );
  XOR2HSV0 U42606 ( .A1(n37712), .A2(n37711), .Z(n37713) );
  XOR2HSV0 U42607 ( .A1(n37714), .A2(n37713), .Z(n37716) );
  NAND2HSV0 U42608 ( .A1(n48014), .A2(n48167), .ZN(n37715) );
  XNOR2HSV1 U42609 ( .A1(n37716), .A2(n37715), .ZN(n37717) );
  XNOR2HSV1 U42610 ( .A1(n37718), .A2(n37717), .ZN(n37719) );
  XNOR2HSV1 U42611 ( .A1(n37720), .A2(n37719), .ZN(n37721) );
  XNOR2HSV1 U42612 ( .A1(n37722), .A2(n37721), .ZN(n37728) );
  CLKNAND2HSV0 U42613 ( .A1(n37723), .A2(n39434), .ZN(n37727) );
  BUFHSV2 U42614 ( .I(n37724), .Z(n48848) );
  CLKNAND2HSV0 U42615 ( .A1(n48848), .A2(n37725), .ZN(n37726) );
  XOR3HSV2 U42616 ( .A1(n37728), .A2(n37727), .A3(n37726), .Z(n37729) );
  XNOR2HSV1 U42617 ( .A1(n37730), .A2(n37729), .ZN(n37731) );
  XNOR2HSV1 U42618 ( .A1(n37732), .A2(n37731), .ZN(n37733) );
  XOR2HSV0 U42619 ( .A1(n37734), .A2(n37733), .Z(n37735) );
  XNOR2HSV1 U42620 ( .A1(n37736), .A2(n37735), .ZN(n37737) );
  XOR2HSV0 U42621 ( .A1(n37738), .A2(n37737), .Z(n37739) );
  XNOR2HSV1 U42622 ( .A1(n37740), .A2(n37739), .ZN(n37741) );
  XNOR2HSV1 U42623 ( .A1(n37742), .A2(n37741), .ZN(n37743) );
  XNOR2HSV1 U42624 ( .A1(n37744), .A2(n37743), .ZN(n37746) );
  CLKNAND2HSV0 U42625 ( .A1(n39537), .A2(n48742), .ZN(n37745) );
  NAND2HSV2 U42626 ( .A1(n39542), .A2(n30513), .ZN(n37749) );
  XNOR2HSV4 U42627 ( .A1(n37750), .A2(n37749), .ZN(n37752) );
  NAND2HSV0 U42628 ( .A1(n39116), .A2(n30046), .ZN(n37751) );
  XNOR2HSV4 U42629 ( .A1(n37752), .A2(n37751), .ZN(n39388) );
  NOR2HSV4 U42630 ( .A1(n37754), .A2(n37753), .ZN(n39255) );
  NAND3HSV2 U42631 ( .A1(n39255), .A2(n30881), .A3(n39117), .ZN(n37758) );
  CLKNAND2HSV1 U42632 ( .A1(n39251), .A2(n40008), .ZN(n37755) );
  XNOR2HSV4 U42633 ( .A1(n39388), .A2(n39387), .ZN(n39399) );
  XNOR2HSV4 U42634 ( .A1(n37761), .A2(n37760), .ZN(n37768) );
  CLKNHSV0 U42635 ( .I(n37762), .ZN(n37763) );
  NOR2HSV4 U42636 ( .A1(n37768), .A2(n37763), .ZN(n37774) );
  NOR2HSV4 U42637 ( .A1(n39399), .A2(n29664), .ZN(n37772) );
  CLKNAND2HSV3 U42638 ( .A1(n37768), .A2(n37767), .ZN(n37770) );
  CLKNAND2HSV2 U42639 ( .A1(n37772), .A2(n39401), .ZN(n37777) );
  NAND2HSV2 U42640 ( .A1(n37775), .A2(n39399), .ZN(n37776) );
  CLKNAND2HSV3 U42641 ( .A1(n37777), .A2(n37776), .ZN(n37780) );
  OAI21HSV4 U42642 ( .A1(n39675), .A2(n39676), .B(n37778), .ZN(n37783) );
  NAND3HSV4 U42643 ( .A1(n37781), .A2(n37780), .A3(n37779), .ZN(n37782) );
  CLKNAND2HSV8 U42644 ( .A1(n37783), .A2(n37782), .ZN(n59573) );
  INHSV1 U42645 ( .I(n37273), .ZN(n59964) );
  INHSV2 U42646 ( .I(n37785), .ZN(n59384) );
  INHSV2 U42647 ( .I(n56906), .ZN(n59356) );
  INHSV2 U42648 ( .I(\pe1/got [16]), .ZN(n53793) );
  CLKNHSV4 U42649 ( .I(n53381), .ZN(n37788) );
  CLKNHSV1 U42650 ( .I(n37786), .ZN(n37787) );
  NOR2HSV4 U42651 ( .A1(n37788), .A2(n37787), .ZN(n37790) );
  INHSV2 U42652 ( .I(n38738), .ZN(n53092) );
  NAND2HSV2 U42653 ( .A1(n48896), .A2(n52415), .ZN(n37831) );
  BUFHSV2 U42654 ( .I(n44906), .Z(n38276) );
  INHSV2 U42655 ( .I(n38042), .ZN(n38389) );
  NAND2HSV2 U42656 ( .A1(n38276), .A2(n38389), .ZN(n37824) );
  CLKNAND2HSV1 U42657 ( .A1(n59349), .A2(n52416), .ZN(n37820) );
  CLKNAND2HSV0 U42658 ( .A1(n37792), .A2(\pe2/bq[25] ), .ZN(n37794) );
  CLKNAND2HSV0 U42659 ( .A1(n59970), .A2(n52987), .ZN(n37793) );
  XOR2HSV0 U42660 ( .A1(n37794), .A2(n37793), .Z(n37798) );
  NAND2HSV2 U42661 ( .A1(n59759), .A2(n38064), .ZN(n37796) );
  CLKNAND2HSV1 U42662 ( .A1(\pe2/aot [23]), .A2(n38046), .ZN(n37795) );
  XOR2HSV0 U42663 ( .A1(n37796), .A2(n37795), .Z(n37797) );
  XOR2HSV0 U42664 ( .A1(n37798), .A2(n37797), .Z(n37807) );
  INHSV2 U42665 ( .I(n38655), .ZN(n38122) );
  CLKNAND2HSV0 U42666 ( .A1(n38122), .A2(n38043), .ZN(n37800) );
  CLKNAND2HSV0 U42667 ( .A1(n52310), .A2(n38047), .ZN(n37799) );
  XOR2HSV0 U42668 ( .A1(n37800), .A2(n37799), .Z(n37805) );
  NAND2HSV2 U42669 ( .A1(n37801), .A2(n38549), .ZN(n37803) );
  INHSV2 U42670 ( .I(n45248), .ZN(n49591) );
  CLKNAND2HSV0 U42671 ( .A1(n49591), .A2(n38401), .ZN(n37802) );
  XOR2HSV0 U42672 ( .A1(n37803), .A2(n37802), .Z(n37804) );
  XOR2HSV0 U42673 ( .A1(n37805), .A2(n37804), .Z(n37806) );
  XOR2HSV0 U42674 ( .A1(n37807), .A2(n37806), .Z(n37816) );
  CLKNAND2HSV1 U42675 ( .A1(n38055), .A2(n38053), .ZN(n37809) );
  CLKNAND2HSV1 U42676 ( .A1(n38061), .A2(\pe2/bq[23] ), .ZN(n37808) );
  XOR2HSV0 U42677 ( .A1(n37809), .A2(n37808), .Z(n37812) );
  NAND2HSV2 U42678 ( .A1(n45811), .A2(\pe2/pvq [11]), .ZN(n37810) );
  XNOR2HSV1 U42679 ( .A1(n37810), .A2(\pe2/phq [11]), .ZN(n37811) );
  XNOR2HSV1 U42680 ( .A1(n37812), .A2(n37811), .ZN(n37814) );
  NOR2HSV2 U42681 ( .A1(n36240), .A2(n52430), .ZN(n44206) );
  NAND2HSV2 U42682 ( .A1(n38048), .A2(n36608), .ZN(n37896) );
  XOR2HSV0 U42683 ( .A1(n44206), .A2(n37896), .Z(n37813) );
  XNOR2HSV1 U42684 ( .A1(n37814), .A2(n37813), .ZN(n37815) );
  XNOR2HSV1 U42685 ( .A1(n37816), .A2(n37815), .ZN(n37818) );
  NAND2HSV2 U42686 ( .A1(n39061), .A2(n38080), .ZN(n37817) );
  XOR2HSV0 U42687 ( .A1(n37818), .A2(n37817), .Z(n37819) );
  XNOR2HSV1 U42688 ( .A1(n37820), .A2(n37819), .ZN(n37822) );
  CLKNAND2HSV0 U42689 ( .A1(n38081), .A2(n38324), .ZN(n37821) );
  XNOR2HSV1 U42690 ( .A1(n37822), .A2(n37821), .ZN(n37823) );
  XOR2HSV2 U42691 ( .A1(n37824), .A2(n37823), .Z(n37826) );
  NAND2HSV2 U42692 ( .A1(n38841), .A2(\pe2/got [27]), .ZN(n37825) );
  XNOR2HSV4 U42693 ( .A1(n37826), .A2(n37825), .ZN(n37830) );
  INHSV2 U42694 ( .I(n44184), .ZN(n59635) );
  CLKAND2HSV1 U42695 ( .A1(n37827), .A2(n59635), .Z(n37828) );
  OAI21HSV2 U42696 ( .A1(n60005), .A2(n38454), .B(n37828), .ZN(n37829) );
  NOR2HSV2 U42697 ( .A1(\pe2/got [32]), .A2(n38184), .ZN(n44316) );
  INHSV1 U42698 ( .I(n36277), .ZN(n37834) );
  CLKNHSV0 U42699 ( .I(n37836), .ZN(n37838) );
  NAND2HSV2 U42700 ( .A1(n37838), .A2(n37837), .ZN(n37840) );
  CLKNHSV0 U42701 ( .I(n37923), .ZN(n37839) );
  CLKAND2HSV2 U42702 ( .A1(n37840), .A2(n37839), .Z(n37842) );
  OR2HSV1 U42703 ( .A1(n37845), .A2(n36277), .Z(n37841) );
  CLKNAND2HSV2 U42704 ( .A1(n37842), .A2(n37841), .ZN(n37843) );
  NOR2HSV4 U42705 ( .A1(n37844), .A2(n37843), .ZN(n37854) );
  AND3HSV0 U42706 ( .A1(n37847), .A2(n37846), .A3(n37845), .Z(n37848) );
  CLKNAND2HSV4 U42707 ( .A1(n37854), .A2(n37855), .ZN(n37978) );
  INHSV3 U42708 ( .I(n37863), .ZN(n53384) );
  INHSV4 U42709 ( .I(n29632), .ZN(n37850) );
  CLKNHSV0 U42710 ( .I(n37864), .ZN(n53385) );
  INHSV4 U42711 ( .I(n37978), .ZN(n38972) );
  BUFHSV8 U42712 ( .I(n38972), .Z(n44264) );
  NAND2HSV4 U42713 ( .A1(n53385), .A2(n38972), .ZN(n37992) );
  NAND3HSV4 U42714 ( .A1(n37992), .A2(n37850), .A3(n37849), .ZN(n38022) );
  INHSV2 U42715 ( .I(n52746), .ZN(n37859) );
  CLKNAND2HSV3 U42716 ( .A1(n38022), .A2(n37859), .ZN(n37862) );
  NAND2HSV2 U42717 ( .A1(n37978), .A2(n45399), .ZN(n37851) );
  INHSV2 U42718 ( .I(n37854), .ZN(n37857) );
  CLKNAND2HSV2 U42719 ( .A1(n37855), .A2(n45399), .ZN(n37856) );
  NOR2HSV4 U42720 ( .A1(n37857), .A2(n37856), .ZN(n37858) );
  CLKNAND2HSV2 U42721 ( .A1(n38023), .A2(n37858), .ZN(n38025) );
  NOR2HSV2 U42722 ( .A1(n44315), .A2(\pe2/ti_7t [10]), .ZN(n37874) );
  NOR2HSV2 U42723 ( .A1(n37874), .A2(n37871), .ZN(n38034) );
  INHSV2 U42724 ( .I(n38034), .ZN(n37865) );
  INHSV2 U42725 ( .I(n37865), .ZN(n38004) );
  CLKAND2HSV2 U42726 ( .A1(n37859), .A2(n38004), .Z(n37860) );
  CLKNAND2HSV4 U42727 ( .A1(n37862), .A2(n37861), .ZN(n38106) );
  INHSV2 U42728 ( .I(n38007), .ZN(n37985) );
  INAND2HSV2 U42729 ( .A1(n37978), .B1(n37864), .ZN(n37983) );
  INHSV2 U42730 ( .I(n38529), .ZN(n38885) );
  NOR2HSV2 U42731 ( .A1(n38006), .A2(n37870), .ZN(n37868) );
  NOR2HSV3 U42732 ( .A1(n38005), .A2(n38007), .ZN(n37867) );
  NAND2HSV2 U42733 ( .A1(n38025), .A2(n38034), .ZN(n37869) );
  INHSV2 U42734 ( .I(n37869), .ZN(n37866) );
  NAND3HSV4 U42735 ( .A1(n37868), .A2(n37867), .A3(n37866), .ZN(n52747) );
  BUFHSV2 U42736 ( .I(n37871), .Z(n44307) );
  NAND3HSV4 U42737 ( .A1(n37873), .A2(n25870), .A3(n37872), .ZN(n52748) );
  NOR2HSV2 U42738 ( .A1(n37874), .A2(n39105), .ZN(n37875) );
  MUX2NHSV1 U42739 ( .I0(n60005), .I1(\pe2/ti_7t [7]), .S(n44821), .ZN(n37933)
         );
  INHSV2 U42740 ( .I(n37933), .ZN(n38041) );
  NAND2HSV2 U42741 ( .A1(n45150), .A2(n59981), .ZN(n37912) );
  CLKNAND2HSV1 U42742 ( .A1(n39061), .A2(n49591), .ZN(n37905) );
  CLKNAND2HSV1 U42743 ( .A1(\pe2/aot [22]), .A2(n38046), .ZN(n37878) );
  NAND2HSV0 U42744 ( .A1(n38061), .A2(n38054), .ZN(n37877) );
  XOR2HSV0 U42745 ( .A1(n37878), .A2(n37877), .Z(n37882) );
  NAND2HSV2 U42746 ( .A1(n59585), .A2(n38043), .ZN(n37880) );
  NAND2HSV0 U42747 ( .A1(n38055), .A2(\pe2/bq[23] ), .ZN(n37879) );
  XOR2HSV0 U42748 ( .A1(n37880), .A2(n37879), .Z(n37881) );
  XOR2HSV0 U42749 ( .A1(n37882), .A2(n37881), .Z(n37890) );
  CLKNHSV0 U42750 ( .I(n38787), .ZN(n38134) );
  CLKNAND2HSV1 U42751 ( .A1(n38134), .A2(n38053), .ZN(n37884) );
  NAND2HSV0 U42752 ( .A1(\pe2/aot [26]), .A2(n38047), .ZN(n37883) );
  XOR2HSV0 U42753 ( .A1(n37884), .A2(n37883), .Z(n37888) );
  CLKNAND2HSV1 U42754 ( .A1(n59759), .A2(n44987), .ZN(n37886) );
  CLKNHSV0 U42755 ( .I(n49518), .ZN(n52952) );
  NAND2HSV0 U42756 ( .A1(n52310), .A2(n52952), .ZN(n37885) );
  XOR2HSV0 U42757 ( .A1(n37886), .A2(n37885), .Z(n37887) );
  XOR2HSV0 U42758 ( .A1(n37888), .A2(n37887), .Z(n37889) );
  XOR2HSV0 U42759 ( .A1(n37890), .A2(n37889), .Z(n37902) );
  CLKNAND2HSV1 U42760 ( .A1(n52104), .A2(n43972), .ZN(n37892) );
  INHSV2 U42761 ( .I(\pe2/got [21]), .ZN(n38711) );
  CLKNAND2HSV0 U42762 ( .A1(\pe2/got [21]), .A2(n38401), .ZN(n37891) );
  XOR2HSV0 U42763 ( .A1(n37892), .A2(n37891), .Z(n37895) );
  CLKNAND2HSV1 U42764 ( .A1(n45811), .A2(\pe2/pvq [12]), .ZN(n37893) );
  XNOR2HSV1 U42765 ( .A1(n37893), .A2(\pe2/phq [12]), .ZN(n37894) );
  XNOR2HSV1 U42766 ( .A1(n37895), .A2(n37894), .ZN(n37900) );
  CLKNAND2HSV0 U42767 ( .A1(n38122), .A2(n36588), .ZN(n45192) );
  CLKNHSV0 U42768 ( .I(n36240), .ZN(n38558) );
  INHSV2 U42769 ( .I(\pe2/bq[21] ), .ZN(n47608) );
  CLKNAND2HSV1 U42770 ( .A1(n38558), .A2(\pe2/bq[21] ), .ZN(n37897) );
  XNOR2HSV1 U42771 ( .A1(n37898), .A2(n37897), .ZN(n37899) );
  XNOR2HSV1 U42772 ( .A1(n37900), .A2(n37899), .ZN(n37901) );
  XNOR2HSV1 U42773 ( .A1(n37902), .A2(n37901), .ZN(n37904) );
  INHSV2 U42774 ( .I(n38205), .ZN(n39008) );
  CLKNAND2HSV0 U42775 ( .A1(n38081), .A2(n39008), .ZN(n37903) );
  XOR3HSV2 U42776 ( .A1(n37905), .A2(n37904), .A3(n37903), .Z(n37907) );
  INHSV2 U42777 ( .I(n59349), .ZN(n52420) );
  NOR2HSV2 U42778 ( .A1(n52420), .A2(n38275), .ZN(n37906) );
  XNOR2HSV1 U42779 ( .A1(n37907), .A2(n37906), .ZN(n37910) );
  NAND2HSV2 U42780 ( .A1(n38276), .A2(n38324), .ZN(n37909) );
  BUFHSV2 U42781 ( .I(n38841), .Z(n38151) );
  INHSV2 U42782 ( .I(n38042), .ZN(n38512) );
  NAND2HSV2 U42783 ( .A1(n38151), .A2(n38512), .ZN(n37908) );
  XOR3HSV2 U42784 ( .A1(n37910), .A2(n37909), .A3(n37908), .Z(n37911) );
  XOR2HSV0 U42785 ( .A1(n37912), .A2(n37911), .Z(n37913) );
  XNOR2HSV1 U42786 ( .A1(n37914), .A2(n37913), .ZN(n37916) );
  NAND2HSV0 U42787 ( .A1(n36398), .A2(n37975), .ZN(n37915) );
  CLKNHSV0 U42788 ( .I(n47998), .ZN(n37917) );
  CLKNAND2HSV0 U42789 ( .A1(n37917), .A2(n38742), .ZN(n37926) );
  NAND2HSV0 U42790 ( .A1(n37919), .A2(n37918), .ZN(n37920) );
  NAND2HSV1 U42791 ( .A1(n37920), .A2(n36277), .ZN(n37922) );
  CLKAND2HSV2 U42792 ( .A1(n47998), .A2(n53092), .Z(n37921) );
  CLKNAND2HSV1 U42793 ( .A1(n37922), .A2(n37921), .ZN(n37925) );
  NAND2HSV0 U42794 ( .A1(n37923), .A2(n38742), .ZN(n37924) );
  CLKNAND2HSV1 U42795 ( .A1(\pe2/ti_7t [12]), .A2(n38099), .ZN(n37929) );
  INHSV2 U42796 ( .I(n37929), .ZN(n38114) );
  NAND3HSV2 U42797 ( .A1(n52748), .A2(n52747), .A3(n37929), .ZN(n37930) );
  CLKNAND2HSV0 U42798 ( .A1(\pe2/ti_7t [10]), .A2(n37931), .ZN(n38098) );
  INHSV2 U42799 ( .I(n38098), .ZN(n38101) );
  INHSV2 U42800 ( .I(n38101), .ZN(n37932) );
  CLKNAND2HSV3 U42801 ( .A1(n38016), .A2(n37932), .ZN(n38001) );
  CLKNAND2HSV2 U42802 ( .A1(n38001), .A2(n44145), .ZN(n37982) );
  CLKNAND2HSV1 U42803 ( .A1(n45149), .A2(n38389), .ZN(n37974) );
  CLKNAND2HSV0 U42804 ( .A1(n45150), .A2(n38324), .ZN(n37972) );
  CLKNAND2HSV0 U42805 ( .A1(n38276), .A2(n38080), .ZN(n37968) );
  CLKNAND2HSV1 U42806 ( .A1(n52294), .A2(n38303), .ZN(n37935) );
  NAND2HSV0 U42807 ( .A1(\pe2/aot [22]), .A2(n36608), .ZN(n37934) );
  XOR2HSV0 U42808 ( .A1(n37935), .A2(n37934), .Z(n37939) );
  CLKNHSV0 U42809 ( .I(n38687), .ZN(n38542) );
  NAND2HSV0 U42810 ( .A1(n49530), .A2(n38542), .ZN(n37937) );
  NAND2HSV0 U42811 ( .A1(n59982), .A2(n38401), .ZN(n37936) );
  XOR2HSV0 U42812 ( .A1(n37937), .A2(n37936), .Z(n37938) );
  XOR2HSV0 U42813 ( .A1(n37939), .A2(n37938), .Z(n37949) );
  NAND2HSV0 U42814 ( .A1(n44081), .A2(n52179), .ZN(n37943) );
  INHSV2 U42815 ( .I(n47599), .ZN(n51998) );
  CLKNAND2HSV1 U42816 ( .A1(n38061), .A2(n51998), .ZN(n37942) );
  XOR2HSV0 U42817 ( .A1(n37943), .A2(n37942), .Z(n37947) );
  NAND2HSV0 U42818 ( .A1(n59758), .A2(n38043), .ZN(n37945) );
  NAND2HSV0 U42819 ( .A1(n52974), .A2(n52950), .ZN(n37944) );
  XOR2HSV0 U42820 ( .A1(n37945), .A2(n37944), .Z(n37946) );
  XOR2HSV0 U42821 ( .A1(n37947), .A2(n37946), .Z(n37948) );
  XOR2HSV0 U42822 ( .A1(n37949), .A2(n37948), .Z(n37951) );
  INHSV2 U42823 ( .I(n44327), .ZN(n38390) );
  NAND2HSV0 U42824 ( .A1(n38291), .A2(n38390), .ZN(n37950) );
  XNOR2HSV1 U42825 ( .A1(n37951), .A2(n37950), .ZN(n37966) );
  NOR2HSV1 U42826 ( .A1(n52420), .A2(n38711), .ZN(n37965) );
  NAND2HSV0 U42827 ( .A1(n38048), .A2(\pe2/bq[26] ), .ZN(n38123) );
  CLKNAND2HSV0 U42828 ( .A1(n38134), .A2(\pe2/bq[22] ), .ZN(n52940) );
  XOR2HSV0 U42829 ( .A1(n38123), .A2(n52940), .Z(n37962) );
  BUFHSV4 U42830 ( .I(n37952), .Z(n53014) );
  INHSV2 U42831 ( .I(\pe2/bq[19] ), .ZN(n52429) );
  NOR2HSV1 U42832 ( .A1(n36240), .A2(n52429), .ZN(n52938) );
  INHSV2 U42833 ( .I(n50947), .ZN(n59587) );
  CLKNAND2HSV1 U42834 ( .A1(n59587), .A2(n36480), .ZN(n37955) );
  INHSV2 U42835 ( .I(n38404), .ZN(n44207) );
  CLKNAND2HSV1 U42836 ( .A1(n44207), .A2(\pe2/bq[21] ), .ZN(n37954) );
  XOR2HSV0 U42837 ( .A1(n37955), .A2(n37954), .Z(n37959) );
  NAND2HSV0 U42838 ( .A1(n38122), .A2(n38047), .ZN(n37957) );
  NAND2HSV0 U42839 ( .A1(n59585), .A2(\pe2/bq[28] ), .ZN(n37956) );
  XOR2HSV0 U42840 ( .A1(n37957), .A2(n37956), .Z(n37958) );
  XOR2HSV0 U42841 ( .A1(n37959), .A2(n37958), .Z(n37960) );
  XOR3HSV2 U42842 ( .A1(n37962), .A2(n37961), .A3(n37960), .Z(n37964) );
  CLKNHSV0 U42843 ( .I(n45248), .ZN(n45287) );
  CLKNAND2HSV0 U42844 ( .A1(n38081), .A2(n45287), .ZN(n37963) );
  XOR4HSV1 U42845 ( .A1(n37966), .A2(n37965), .A3(n37964), .A4(n37963), .Z(
        n37967) );
  XNOR2HSV1 U42846 ( .A1(n37968), .A2(n37967), .ZN(n37970) );
  CLKNAND2HSV0 U42847 ( .A1(n38151), .A2(n59584), .ZN(n37969) );
  XNOR2HSV1 U42848 ( .A1(n37970), .A2(n37969), .ZN(n37971) );
  XNOR2HSV1 U42849 ( .A1(n37972), .A2(n37971), .ZN(n37973) );
  XNOR2HSV1 U42850 ( .A1(n37974), .A2(n37973), .ZN(n37977) );
  BUFHSV2 U42851 ( .I(n37975), .Z(n38323) );
  NAND2HSV2 U42852 ( .A1(n38323), .A2(n59981), .ZN(n37976) );
  XOR2HSV2 U42853 ( .A1(n37977), .A2(n37976), .Z(n37980) );
  NAND2HSV2 U42854 ( .A1(n38024), .A2(n38327), .ZN(n37979) );
  CLKXOR2HSV4 U42855 ( .A1(n37980), .A2(n37979), .Z(n37981) );
  XNOR2HSV4 U42856 ( .A1(n37982), .A2(n37981), .ZN(n38000) );
  INHSV3 U42857 ( .I(n38000), .ZN(n37998) );
  NAND2HSV0 U42858 ( .A1(n37983), .A2(n53092), .ZN(n37984) );
  NOR2HSV2 U42859 ( .A1(n37984), .A2(n38005), .ZN(n37986) );
  AND3HSV4 U42860 ( .A1(n37987), .A2(n37986), .A3(n37985), .Z(n37996) );
  INHSV2 U42861 ( .I(n52746), .ZN(n38035) );
  AOI21HSV2 U42862 ( .A1(n29632), .A2(n38035), .B(n52411), .ZN(n37988) );
  IOA21HSV2 U42863 ( .A1(n25869), .A2(n38035), .B(n37988), .ZN(n37994) );
  NAND2HSV0 U42864 ( .A1(n38034), .A2(n38035), .ZN(n37990) );
  OAI22HSV2 U42865 ( .A1(n37992), .A2(n52746), .B1(n37991), .B2(n37990), .ZN(
        n37993) );
  NOR2HSV3 U42866 ( .A1(n37994), .A2(n37993), .ZN(n37995) );
  NOR2HSV4 U42867 ( .A1(n37996), .A2(n37995), .ZN(n37999) );
  INHSV2 U42868 ( .I(n37999), .ZN(n37997) );
  CLKNAND2HSV2 U42869 ( .A1(n38336), .A2(n38383), .ZN(n52772) );
  CLKNAND2HSV3 U42870 ( .A1(n38001), .A2(n38340), .ZN(n38003) );
  XNOR2HSV4 U42871 ( .A1(n38003), .A2(n38002), .ZN(n38109) );
  INHSV2 U42872 ( .I(n38005), .ZN(n38009) );
  NOR2HSV2 U42873 ( .A1(n53386), .A2(n38033), .ZN(n38010) );
  INHSV2 U42874 ( .I(n38010), .ZN(n38011) );
  CLKNAND2HSV3 U42875 ( .A1(n38106), .A2(n38011), .ZN(n38328) );
  OAI21HSV0 U42876 ( .A1(n38183), .A2(\pe2/ti_7t [12]), .B(n47997), .ZN(n47978) );
  NAND2HSV0 U42877 ( .A1(n47978), .A2(n38627), .ZN(n38178) );
  INHSV2 U42878 ( .I(\pe2/ti_7t [13]), .ZN(n38014) );
  NOR2HSV2 U42879 ( .A1(n38108), .A2(n38014), .ZN(n38180) );
  INHSV2 U42880 ( .I(n38180), .ZN(n38177) );
  CLKAND2HSV1 U42881 ( .A1(n38178), .A2(n38177), .Z(n38015) );
  MUX2NHSV2 U42882 ( .I0(n38018), .I1(n38017), .S(n38388), .ZN(n38020) );
  AO21HSV1 U42883 ( .A1(n38002), .A2(n39105), .B(n44821), .Z(n38019) );
  NOR2HSV2 U42884 ( .A1(n38020), .A2(n38019), .ZN(n38021) );
  CLKNAND2HSV2 U42885 ( .A1(n38021), .A2(n59583), .ZN(n38176) );
  INHSV2 U42886 ( .I(n38176), .ZN(n38191) );
  NOR2HSV4 U42887 ( .A1(n38022), .A2(n36575), .ZN(n38040) );
  NAND2HSV2 U42888 ( .A1(n37853), .A2(n38024), .ZN(n38030) );
  CLKNHSV0 U42889 ( .I(n38025), .ZN(n38028) );
  NAND2HSV0 U42890 ( .A1(n38034), .A2(n38026), .ZN(n38027) );
  NOR2HSV2 U42891 ( .A1(n38028), .A2(n38027), .ZN(n38029) );
  NAND2HSV2 U42892 ( .A1(n38030), .A2(n38029), .ZN(n38032) );
  OR2HSV1 U42893 ( .A1(n38035), .A2(n44156), .Z(n38031) );
  CLKNAND2HSV2 U42894 ( .A1(n38032), .A2(n38031), .ZN(n38039) );
  INHSV4 U42895 ( .I(n38033), .ZN(n38104) );
  NAND2HSV0 U42896 ( .A1(n38035), .A2(n38034), .ZN(n38037) );
  INAND2HSV4 U42897 ( .A1(n38037), .B1(n38036), .ZN(n38038) );
  CLKNAND2HSV0 U42898 ( .A1(n38041), .A2(\pe2/got [27]), .ZN(n38093) );
  NAND2HSV2 U42899 ( .A1(n52288), .A2(n38778), .ZN(n38091) );
  CLKNAND2HSV0 U42900 ( .A1(n37801), .A2(n38043), .ZN(n38045) );
  NAND2HSV0 U42901 ( .A1(n59585), .A2(n36608), .ZN(n38044) );
  XOR2HSV0 U42902 ( .A1(n38045), .A2(n38044), .Z(n38052) );
  NAND2HSV0 U42903 ( .A1(n59758), .A2(n38046), .ZN(n38050) );
  NAND2HSV0 U42904 ( .A1(n38048), .A2(n38047), .ZN(n38049) );
  XOR2HSV0 U42905 ( .A1(n38050), .A2(n38049), .Z(n38051) );
  XOR2HSV0 U42906 ( .A1(n38052), .A2(n38051), .Z(n38060) );
  CLKNAND2HSV0 U42907 ( .A1(n59759), .A2(n38053), .ZN(n38300) );
  NAND2HSV0 U42908 ( .A1(n52310), .A2(\pe2/bq[25] ), .ZN(n38297) );
  XOR2HSV0 U42909 ( .A1(n38300), .A2(n38297), .Z(n38058) );
  NAND2HSV0 U42910 ( .A1(n38055), .A2(n38054), .ZN(n38056) );
  XOR2HSV0 U42911 ( .A1(n45192), .A2(n38056), .Z(n38057) );
  XOR2HSV0 U42912 ( .A1(n38058), .A2(n38057), .Z(n38059) );
  XOR2HSV0 U42913 ( .A1(n38060), .A2(n38059), .Z(n38077) );
  CLKNAND2HSV0 U42914 ( .A1(\pe2/aot [20]), .A2(n38549), .ZN(n38063) );
  NAND2HSV0 U42915 ( .A1(n38061), .A2(\pe2/bq[21] ), .ZN(n38062) );
  XOR2HSV0 U42916 ( .A1(n38063), .A2(n38062), .Z(n38068) );
  CLKNAND2HSV0 U42917 ( .A1(n59970), .A2(n38064), .ZN(n38066) );
  NAND2HSV0 U42918 ( .A1(n38558), .A2(n51998), .ZN(n38065) );
  XOR2HSV0 U42919 ( .A1(n38066), .A2(n38065), .Z(n38067) );
  XOR2HSV0 U42920 ( .A1(n38068), .A2(n38067), .Z(n38075) );
  NOR2HSV0 U42921 ( .A1(n44327), .A2(n38213), .ZN(n38070) );
  NAND2HSV0 U42922 ( .A1(n38134), .A2(\pe2/bq[23] ), .ZN(n38069) );
  XOR2HSV0 U42923 ( .A1(n38070), .A2(n38069), .Z(n38073) );
  CLKNAND2HSV0 U42924 ( .A1(n45811), .A2(\pe2/pvq [13]), .ZN(n38071) );
  XOR2HSV0 U42925 ( .A1(n38071), .A2(\pe2/phq [13]), .Z(n38072) );
  XOR2HSV0 U42926 ( .A1(n38073), .A2(n38072), .Z(n38074) );
  XOR2HSV0 U42927 ( .A1(n38075), .A2(n38074), .Z(n38076) );
  XOR2HSV0 U42928 ( .A1(n38077), .A2(n38076), .Z(n38079) );
  NAND2HSV0 U42929 ( .A1(n38291), .A2(n52922), .ZN(n38078) );
  XNOR2HSV1 U42930 ( .A1(n38079), .A2(n38078), .ZN(n38083) );
  NAND2HSV0 U42931 ( .A1(n38081), .A2(n38080), .ZN(n38082) );
  XNOR2HSV1 U42932 ( .A1(n38083), .A2(n38082), .ZN(n38085) );
  CLKNAND2HSV0 U42933 ( .A1(n59349), .A2(n49591), .ZN(n38084) );
  XNOR2HSV1 U42934 ( .A1(n38085), .A2(n38084), .ZN(n38087) );
  CLKNAND2HSV0 U42935 ( .A1(n38276), .A2(n59584), .ZN(n38086) );
  XOR2HSV0 U42936 ( .A1(n38087), .A2(n38086), .Z(n38089) );
  CLKNAND2HSV1 U42937 ( .A1(n38151), .A2(n44711), .ZN(n38088) );
  XNOR2HSV1 U42938 ( .A1(n38089), .A2(n38088), .ZN(n38090) );
  XNOR2HSV1 U42939 ( .A1(n38091), .A2(n38090), .ZN(n38092) );
  XNOR2HSV1 U42940 ( .A1(n38093), .A2(n38092), .ZN(n38094) );
  CLKNAND2HSV3 U42941 ( .A1(n38024), .A2(n45388), .ZN(n38096) );
  AOI21HSV1 U42942 ( .A1(n38099), .A2(n38098), .B(n38738), .ZN(n38100) );
  OAI21HSV4 U42943 ( .A1(n60019), .A2(n38101), .B(n38100), .ZN(n38102) );
  XNOR2HSV4 U42944 ( .A1(n38175), .A2(n38174), .ZN(n38190) );
  INHSV2 U42945 ( .I(n38177), .ZN(n38189) );
  OAI22HSV4 U42946 ( .A1(n38192), .A2(n38191), .B1(n38190), .B2(n38189), .ZN(
        n38201) );
  INHSV2 U42947 ( .I(n53386), .ZN(n38105) );
  NAND2HSV2 U42948 ( .A1(n38107), .A2(n38106), .ZN(n38167) );
  NOR2HSV0 U42949 ( .A1(n38454), .A2(n47978), .ZN(n38199) );
  INHSV2 U42950 ( .I(n38199), .ZN(n38110) );
  NOR2HSV4 U42951 ( .A1(n38198), .A2(n38110), .ZN(n38111) );
  INAND3HSV4 U42952 ( .A1(n38190), .B1(n38111), .B2(n25851), .ZN(n38193) );
  NAND2HSV4 U42953 ( .A1(n38201), .A2(n38193), .ZN(n38387) );
  INHSV2 U42954 ( .I(n38269), .ZN(n38441) );
  INHSV2 U42955 ( .I(n38112), .ZN(n38113) );
  NAND2HSV2 U42956 ( .A1(n52748), .A2(n52747), .ZN(n38116) );
  INHSV2 U42957 ( .I(n39080), .ZN(n38173) );
  NAND2HSV0 U42958 ( .A1(n45150), .A2(n59584), .ZN(n38155) );
  CLKNAND2HSV0 U42959 ( .A1(n38276), .A2(n43925), .ZN(n38150) );
  NAND2HSV2 U42960 ( .A1(n36603), .A2(n43961), .ZN(n38228) );
  CLKNAND2HSV1 U42961 ( .A1(\pe2/aot [19]), .A2(n52444), .ZN(n38120) );
  XOR2HSV0 U42962 ( .A1(n38228), .A2(n38120), .Z(n38133) );
  NAND2HSV0 U42963 ( .A1(n48078), .A2(\pe2/pvq [15]), .ZN(n38121) );
  XOR2HSV0 U42964 ( .A1(n38121), .A2(\pe2/phq [15]), .Z(n38125) );
  NAND2HSV0 U42965 ( .A1(n38122), .A2(n52950), .ZN(n38295) );
  XNOR2HSV1 U42966 ( .A1(n38125), .A2(n38124), .ZN(n38132) );
  BUFHSV2 U42967 ( .I(n47648), .Z(n38973) );
  NAND2HSV2 U42968 ( .A1(n49530), .A2(n52300), .ZN(n38128) );
  NAND2HSV0 U42969 ( .A1(n38558), .A2(n52988), .ZN(n38127) );
  XOR2HSV0 U42970 ( .A1(n38128), .A2(n38127), .Z(n38129) );
  XOR2HSV0 U42971 ( .A1(n38130), .A2(n38129), .Z(n38131) );
  XOR3HSV2 U42972 ( .A1(n38133), .A2(n38132), .A3(n38131), .Z(n38148) );
  CLKNHSV0 U42973 ( .I(n59349), .ZN(n38489) );
  NOR2HSV2 U42974 ( .A1(n38489), .A2(n44327), .ZN(n38147) );
  INHSV2 U42975 ( .I(n52103), .ZN(n51639) );
  NAND2HSV0 U42976 ( .A1(\pe2/aot [22]), .A2(\pe2/bq[28] ), .ZN(n38136) );
  NAND2HSV0 U42977 ( .A1(n59585), .A2(n38394), .ZN(n38135) );
  XOR2HSV0 U42978 ( .A1(n38136), .A2(n38135), .Z(n38140) );
  CLKNAND2HSV0 U42979 ( .A1(n52995), .A2(\pe2/bq[22] ), .ZN(n38138) );
  INHSV2 U42980 ( .I(n47599), .ZN(n38419) );
  CLKNAND2HSV1 U42981 ( .A1(n44207), .A2(n38419), .ZN(n38137) );
  XOR2HSV0 U42982 ( .A1(n38138), .A2(n38137), .Z(n38139) );
  XOR2HSV0 U42983 ( .A1(n38140), .A2(n38139), .Z(n38141) );
  XOR2HSV0 U42984 ( .A1(n38142), .A2(n38141), .Z(n38144) );
  NAND2HSV0 U42985 ( .A1(n38291), .A2(n39075), .ZN(n38143) );
  XNOR2HSV1 U42986 ( .A1(n38144), .A2(n38143), .ZN(n38146) );
  CLKNAND2HSV0 U42987 ( .A1(n44187), .A2(n52167), .ZN(n38145) );
  XOR4HSV1 U42988 ( .A1(n38148), .A2(n38147), .A3(n38146), .A4(n38145), .Z(
        n38149) );
  XNOR2HSV1 U42989 ( .A1(n38150), .A2(n38149), .ZN(n38153) );
  NAND2HSV0 U42990 ( .A1(n38151), .A2(n45249), .ZN(n38152) );
  XNOR2HSV1 U42991 ( .A1(n38153), .A2(n38152), .ZN(n38154) );
  XNOR2HSV1 U42992 ( .A1(n38155), .A2(n38154), .ZN(n38158) );
  NAND2HSV2 U42993 ( .A1(n45149), .A2(n38324), .ZN(n38157) );
  XOR3HSV2 U42994 ( .A1(n38158), .A2(n38157), .A3(n38156), .Z(n38161) );
  CLKNHSV2 U42995 ( .I(n59981), .ZN(n38159) );
  NOR2HSV4 U42996 ( .A1(n44264), .A2(n38159), .ZN(n38160) );
  XNOR2HSV4 U42997 ( .A1(n38161), .A2(n38160), .ZN(n38164) );
  CLKNAND2HSV1 U42998 ( .A1(n38162), .A2(n50929), .ZN(n38166) );
  INHSV2 U42999 ( .I(n38206), .ZN(n38274) );
  OAI21HSV2 U43000 ( .A1(n38274), .A2(n44143), .B(n38164), .ZN(n38165) );
  CLKNAND2HSV2 U43001 ( .A1(n38167), .A2(n36398), .ZN(n38168) );
  INHSV2 U43002 ( .I(n38733), .ZN(n38382) );
  CLKNAND2HSV2 U43003 ( .A1(n38171), .A2(n38382), .ZN(n38172) );
  AND2HSV2 U43004 ( .A1(n38178), .A2(n38177), .Z(n38179) );
  XNOR2HSV4 U43005 ( .A1(n38182), .A2(n38181), .ZN(n38444) );
  CLKNHSV0 U43006 ( .I(\pe2/ti_7t [14]), .ZN(n38185) );
  CLKNAND2HSV0 U43007 ( .A1(n38185), .A2(n38184), .ZN(n38341) );
  NAND2HSV2 U43008 ( .A1(n38341), .A2(n47997), .ZN(n38196) );
  NOR2HSV2 U43009 ( .A1(n38196), .A2(n59586), .ZN(n38186) );
  OAI21HSV2 U43010 ( .A1(n38337), .A2(n38387), .B(n38186), .ZN(n38268) );
  INHSV2 U43011 ( .I(n38268), .ZN(n38442) );
  INHSV2 U43012 ( .I(n38442), .ZN(n38187) );
  INHSV2 U43013 ( .I(n38270), .ZN(n38448) );
  OAI21HSV4 U43014 ( .A1(n38188), .A2(n38187), .B(n38448), .ZN(n38456) );
  OAI22HSV2 U43015 ( .A1(n38192), .A2(n38191), .B1(n38190), .B2(n38189), .ZN(
        n38194) );
  INHSV2 U43016 ( .I(n38196), .ZN(n52771) );
  NAND3HSV2 U43017 ( .A1(n52772), .A2(n38471), .A3(n52771), .ZN(n38447) );
  INHSV4 U43018 ( .I(n38444), .ZN(n38443) );
  INHSV4 U43019 ( .I(n38443), .ZN(n52775) );
  NOR2HSV8 U43020 ( .A1(n38197), .A2(n52775), .ZN(n38455) );
  CLKNHSV0 U43021 ( .I(n38198), .ZN(n47980) );
  NAND2HSV2 U43022 ( .A1(n25851), .A2(n47980), .ZN(n38203) );
  NOR2HSV2 U43023 ( .A1(n47981), .A2(n38110), .ZN(n38200) );
  INHSV2 U43024 ( .I(n38200), .ZN(n38202) );
  OAI22HSV4 U43025 ( .A1(n38203), .A2(n38202), .B1(n38201), .B2(n38375), .ZN(
        n38204) );
  CLKXOR2HSV4 U43026 ( .A1(n38204), .A2(n38336), .Z(n60020) );
  NAND2HSV2 U43027 ( .A1(\pe2/ti_7t [14]), .A2(n38529), .ZN(n38470) );
  CLKNAND2HSV1 U43028 ( .A1(n26098), .A2(n38723), .ZN(n38261) );
  CLKNHSV0 U43029 ( .I(n38471), .ZN(n45148) );
  INHSV2 U43030 ( .I(n45148), .ZN(n39009) );
  NAND2HSV2 U43031 ( .A1(n39009), .A2(n38512), .ZN(n38259) );
  INHSV4 U43032 ( .I(n59583), .ZN(n38779) );
  NAND2HSV2 U43033 ( .A1(\pe2/got [24]), .A2(n51966), .ZN(n38257) );
  BUFHSV2 U43034 ( .I(n50929), .Z(n38780) );
  INHSV3 U43035 ( .I(n44327), .ZN(n39010) );
  CLKNHSV0 U43036 ( .I(n59349), .ZN(n53033) );
  NOR2HSV1 U43037 ( .A1(n53033), .A2(n47573), .ZN(n38253) );
  BUFHSV2 U43038 ( .I(n44187), .Z(n38539) );
  CLKNAND2HSV0 U43039 ( .A1(n38539), .A2(\pe2/got [16]), .ZN(n38252) );
  NAND2HSV0 U43040 ( .A1(n39052), .A2(n52950), .ZN(n38208) );
  INHSV2 U43041 ( .I(n38822), .ZN(n51921) );
  NAND2HSV0 U43042 ( .A1(n51921), .A2(n53015), .ZN(n38207) );
  XOR2HSV0 U43043 ( .A1(n38208), .A2(n38207), .Z(n38212) );
  NAND2HSV0 U43044 ( .A1(n59971), .A2(n44197), .ZN(n38210) );
  NAND2HSV0 U43045 ( .A1(n52995), .A2(n44074), .ZN(n38209) );
  XOR2HSV0 U43046 ( .A1(n38210), .A2(n38209), .Z(n38211) );
  XOR2HSV0 U43047 ( .A1(n38212), .A2(n38211), .Z(n38221) );
  CLKNHSV1 U43048 ( .I(n52103), .ZN(n38678) );
  CLKNAND2HSV0 U43049 ( .A1(n38678), .A2(n38394), .ZN(n38215) );
  INHSV2 U43050 ( .I(n51607), .ZN(n59375) );
  NAND2HSV0 U43051 ( .A1(n59375), .A2(n38401), .ZN(n38214) );
  XOR2HSV0 U43052 ( .A1(n38215), .A2(n38214), .Z(n38219) );
  NAND2HSV0 U43053 ( .A1(n45295), .A2(\pe2/bq[18] ), .ZN(n38217) );
  INHSV2 U43054 ( .I(\pe2/aot [16]), .ZN(n38482) );
  INHSV2 U43055 ( .I(n38482), .ZN(n45024) );
  NAND2HSV0 U43056 ( .A1(n45024), .A2(n44759), .ZN(n38216) );
  XOR2HSV0 U43057 ( .A1(n38217), .A2(n38216), .Z(n38218) );
  XOR2HSV0 U43058 ( .A1(n38219), .A2(n38218), .Z(n38220) );
  XOR2HSV0 U43059 ( .A1(n38221), .A2(n38220), .Z(n38233) );
  CLKNAND2HSV0 U43060 ( .A1(\pe2/aot [17]), .A2(n38565), .ZN(n38223) );
  NAND2HSV0 U43061 ( .A1(n59974), .A2(n38043), .ZN(n38222) );
  XOR2HSV0 U43062 ( .A1(n38223), .A2(n38222), .Z(n38226) );
  NAND2HSV0 U43063 ( .A1(n38576), .A2(\pe2/pvq [20]), .ZN(n38224) );
  XNOR2HSV1 U43064 ( .A1(n38224), .A2(\pe2/phq [20]), .ZN(n38225) );
  XNOR2HSV1 U43065 ( .A1(n38226), .A2(n38225), .ZN(n38231) );
  CLKNAND2HSV1 U43066 ( .A1(n52974), .A2(\pe2/bq[14] ), .ZN(n43932) );
  OAI22HSV0 U43067 ( .A1(n44889), .A2(n47580), .B1(n44049), .B2(n45199), .ZN(
        n38227) );
  OAI21HSV0 U43068 ( .A1(n43932), .A2(n38228), .B(n38227), .ZN(n38229) );
  NAND2HSV0 U43069 ( .A1(n38479), .A2(\pe2/bq[21] ), .ZN(n50955) );
  XNOR2HSV1 U43070 ( .A1(n38229), .A2(n50955), .ZN(n38230) );
  XNOR2HSV1 U43071 ( .A1(n38231), .A2(n38230), .ZN(n38232) );
  XNOR2HSV1 U43072 ( .A1(n38233), .A2(n38232), .ZN(n38250) );
  NAND2HSV0 U43073 ( .A1(n39029), .A2(n38542), .ZN(n38235) );
  INHSV2 U43074 ( .I(n49628), .ZN(n51839) );
  CLKNAND2HSV1 U43075 ( .A1(n44892), .A2(n51839), .ZN(n38234) );
  XOR2HSV0 U43076 ( .A1(n38235), .A2(n38234), .Z(n38239) );
  CLKNAND2HSV1 U43077 ( .A1(n51920), .A2(n36480), .ZN(n38237) );
  NAND2HSV0 U43078 ( .A1(\pe2/aot [23]), .A2(n52299), .ZN(n38236) );
  XOR2HSV0 U43079 ( .A1(n38237), .A2(n38236), .Z(n38238) );
  XOR2HSV0 U43080 ( .A1(n38239), .A2(n38238), .Z(n38246) );
  BUFHSV2 U43081 ( .I(n38787), .Z(n48935) );
  NOR2HSV2 U43082 ( .A1(n48935), .A2(n48063), .ZN(n44729) );
  NOR2HSV2 U43083 ( .A1(n38404), .A2(n48066), .ZN(n38495) );
  CLKNHSV0 U43084 ( .I(n38495), .ZN(n38240) );
  XOR2HSV0 U43085 ( .A1(n44729), .A2(n38240), .Z(n38244) );
  NAND2HSV0 U43086 ( .A1(\pe2/aot [22]), .A2(n52300), .ZN(n38242) );
  NAND2HSV0 U43087 ( .A1(\pe2/aot [19]), .A2(n52952), .ZN(n38241) );
  XOR2HSV0 U43088 ( .A1(n38242), .A2(n38241), .Z(n38243) );
  XOR2HSV0 U43089 ( .A1(n38244), .A2(n38243), .Z(n38245) );
  XOR2HSV0 U43090 ( .A1(n38246), .A2(n38245), .Z(n38248) );
  INHSV4 U43091 ( .I(n47498), .ZN(n59354) );
  NAND2HSV0 U43092 ( .A1(n39061), .A2(n59354), .ZN(n38247) );
  XNOR2HSV1 U43093 ( .A1(n38248), .A2(n38247), .ZN(n38249) );
  XOR2HSV0 U43094 ( .A1(n38250), .A2(n38249), .Z(n38251) );
  BUFHSV2 U43095 ( .I(n44906), .Z(n44715) );
  BUFHSV2 U43096 ( .I(n44715), .Z(n43928) );
  CLKNAND2HSV0 U43097 ( .A1(n43928), .A2(n38782), .ZN(n38254) );
  BUFHSV2 U43098 ( .I(n38841), .Z(n38702) );
  BUFHSV2 U43099 ( .I(n47648), .Z(n52169) );
  INHSV2 U43100 ( .I(n52169), .ZN(n38781) );
  BUFHSV2 U43101 ( .I(n38323), .Z(n52367) );
  INHSV1 U43102 ( .I(n38972), .ZN(n45218) );
  INHSV2 U43103 ( .I(n45248), .ZN(n38904) );
  INAND2HSV2 U43104 ( .A1(n39088), .B1(n25940), .ZN(n38255) );
  XOR3HSV2 U43105 ( .A1(n38257), .A2(n38256), .A3(n38255), .Z(n38258) );
  XNOR2HSV1 U43106 ( .A1(n38259), .A2(n38258), .ZN(n38260) );
  XNOR2HSV1 U43107 ( .A1(n38261), .A2(n38260), .ZN(n38263) );
  INHSV2 U43108 ( .I(n44710), .ZN(n38777) );
  XNOR2HSV4 U43109 ( .A1(n38263), .A2(n38262), .ZN(n38370) );
  NAND2HSV2 U43110 ( .A1(n38447), .A2(n38264), .ZN(n38266) );
  INHSV2 U43111 ( .I(n38445), .ZN(n38265) );
  NOR2HSV4 U43112 ( .A1(n38265), .A2(n38266), .ZN(n38267) );
  CLKNAND2HSV1 U43113 ( .A1(n38270), .A2(n47997), .ZN(n38271) );
  CLKNAND2HSV0 U43114 ( .A1(\pe2/ti_7t [16]), .A2(n38272), .ZN(n38347) );
  CLKNHSV1 U43115 ( .I(n38347), .ZN(n38273) );
  NOR2HSV4 U43116 ( .A1(n52777), .A2(n38273), .ZN(n38352) );
  NAND2HSV2 U43117 ( .A1(n39080), .A2(n59635), .ZN(n38332) );
  CLKNAND2HSV2 U43118 ( .A1(n38206), .A2(n38723), .ZN(n38326) );
  CLKNAND2HSV1 U43119 ( .A1(n45149), .A2(n39008), .ZN(n38322) );
  INHSV2 U43120 ( .I(n38275), .ZN(n43924) );
  NAND2HSV0 U43121 ( .A1(n52288), .A2(n43924), .ZN(n38320) );
  NAND2HSV0 U43122 ( .A1(n38276), .A2(n52167), .ZN(n38316) );
  NAND2HSV0 U43123 ( .A1(\pe2/aot [22]), .A2(n38394), .ZN(n38278) );
  NAND2HSV0 U43124 ( .A1(n59983), .A2(n38401), .ZN(n38277) );
  XOR2HSV0 U43125 ( .A1(n38278), .A2(n38277), .Z(n38282) );
  CLKNHSV0 U43126 ( .I(n38787), .ZN(n45005) );
  CLKNAND2HSV1 U43127 ( .A1(n45005), .A2(n38419), .ZN(n38280) );
  CLKNAND2HSV0 U43128 ( .A1(\pe2/aot [19]), .A2(n38393), .ZN(n38279) );
  XOR2HSV0 U43129 ( .A1(n38280), .A2(n38279), .Z(n38281) );
  XOR2HSV0 U43130 ( .A1(n38282), .A2(n38281), .Z(n38290) );
  CLKNAND2HSV1 U43131 ( .A1(n59968), .A2(\pe2/bq[18] ), .ZN(n38284) );
  CLKNAND2HSV1 U43132 ( .A1(n44207), .A2(n38792), .ZN(n38283) );
  XOR2HSV0 U43133 ( .A1(n38284), .A2(n38283), .Z(n38288) );
  NAND2HSV2 U43134 ( .A1(\pe2/aot [21]), .A2(\pe2/bq[28] ), .ZN(n38286) );
  NAND2HSV0 U43135 ( .A1(n59585), .A2(\pe2/bq[26] ), .ZN(n38285) );
  XOR2HSV0 U43136 ( .A1(n38286), .A2(n38285), .Z(n38287) );
  XOR2HSV0 U43137 ( .A1(n38288), .A2(n38287), .Z(n38289) );
  XOR2HSV0 U43138 ( .A1(n38290), .A2(n38289), .Z(n38293) );
  NAND2HSV0 U43139 ( .A1(n38291), .A2(n38781), .ZN(n38292) );
  XNOR2HSV1 U43140 ( .A1(n38293), .A2(n38292), .ZN(n38314) );
  NOR2HSV2 U43141 ( .A1(n38489), .A2(n47570), .ZN(n38313) );
  NAND2HSV2 U43142 ( .A1(n38576), .A2(\pe2/pvq [16]), .ZN(n38294) );
  XOR2HSV0 U43143 ( .A1(n38294), .A2(\pe2/phq [16]), .Z(n38299) );
  NAND2HSV0 U43144 ( .A1(n38479), .A2(\pe2/bq[22] ), .ZN(n38547) );
  OAI21HSV0 U43145 ( .A1(n52430), .A2(n44095), .B(n38295), .ZN(n38296) );
  OAI21HSV0 U43146 ( .A1(n38547), .A2(n38297), .B(n38296), .ZN(n38298) );
  XNOR2HSV1 U43147 ( .A1(n38299), .A2(n38298), .ZN(n38302) );
  CLKNAND2HSV1 U43148 ( .A1(n59971), .A2(\pe2/bq[21] ), .ZN(n38548) );
  NOR2HSV0 U43149 ( .A1(n36240), .A2(n44844), .ZN(n38494) );
  XNOR2HSV1 U43150 ( .A1(n38302), .A2(n38301), .ZN(n38310) );
  CLKNAND2HSV1 U43151 ( .A1(n52974), .A2(\pe2/bq[23] ), .ZN(n38305) );
  CLKNAND2HSV0 U43152 ( .A1(n51759), .A2(n38303), .ZN(n38304) );
  XOR2HSV0 U43153 ( .A1(n38305), .A2(n38304), .Z(n38308) );
  NAND2HSV0 U43154 ( .A1(n39052), .A2(n36608), .ZN(n52437) );
  CLKNAND2HSV0 U43155 ( .A1(n44062), .A2(n52444), .ZN(n38306) );
  XOR2HSV0 U43156 ( .A1(n52437), .A2(n38306), .Z(n38307) );
  XOR2HSV0 U43157 ( .A1(n38308), .A2(n38307), .Z(n38309) );
  XNOR2HSV1 U43158 ( .A1(n38310), .A2(n38309), .ZN(n38312) );
  NAND2HSV2 U43159 ( .A1(n38539), .A2(n38390), .ZN(n38311) );
  XOR4HSV1 U43160 ( .A1(n38314), .A2(n38313), .A3(n38312), .A4(n38311), .Z(
        n38315) );
  XNOR2HSV1 U43161 ( .A1(n38316), .A2(n38315), .ZN(n38318) );
  NAND2HSV0 U43162 ( .A1(n44254), .A2(n38904), .ZN(n38317) );
  XNOR2HSV1 U43163 ( .A1(n38318), .A2(n38317), .ZN(n38319) );
  XNOR2HSV1 U43164 ( .A1(n38320), .A2(n38319), .ZN(n38321) );
  XNOR2HSV1 U43165 ( .A1(n38322), .A2(n38321), .ZN(n38325) );
  BUFHSV2 U43166 ( .I(n38323), .Z(n38510) );
  NAND2HSV2 U43167 ( .A1(n38328), .A2(n38327), .ZN(n38329) );
  XNOR2HSV4 U43168 ( .A1(n38330), .A2(n38329), .ZN(n38331) );
  XOR2HSV2 U43169 ( .A1(n38332), .A2(n38331), .Z(n38333) );
  XNOR2HSV4 U43170 ( .A1(n38334), .A2(n38333), .ZN(n38362) );
  CLKAND2HSV2 U43171 ( .A1(n38362), .A2(n39007), .Z(n38343) );
  NAND3HSV2 U43172 ( .A1(n38387), .A2(n38336), .A3(n44312), .ZN(n38357) );
  INHSV2 U43173 ( .I(n38357), .ZN(n38339) );
  NAND2HSV2 U43174 ( .A1(n38341), .A2(n38340), .ZN(n38353) );
  INHSV2 U43175 ( .I(n38353), .ZN(n38345) );
  CLKNAND2HSV2 U43176 ( .A1(n38346), .A2(n38345), .ZN(n38342) );
  CLKNAND2HSV1 U43177 ( .A1(n38343), .A2(n38342), .ZN(n38351) );
  OAI21HSV2 U43178 ( .A1(n38348), .A2(n38362), .B(n38347), .ZN(n38349) );
  INHSV2 U43179 ( .I(n38349), .ZN(n38350) );
  NAND2HSV2 U43180 ( .A1(n38357), .A2(n38356), .ZN(n38360) );
  NOR2HSV2 U43181 ( .A1(n38338), .A2(n38360), .ZN(n38358) );
  NOR2HSV2 U43182 ( .A1(n38360), .A2(n38338), .ZN(n38361) );
  CLKNAND2HSV4 U43183 ( .A1(n52776), .A2(n38364), .ZN(n38365) );
  NOR2HSV4 U43184 ( .A1(n38377), .A2(n38365), .ZN(n38366) );
  NOR2HSV4 U43185 ( .A1(n38367), .A2(n38366), .ZN(n38536) );
  INHSV2 U43186 ( .I(n38536), .ZN(n38368) );
  NAND2HSV2 U43187 ( .A1(n38368), .A2(n36377), .ZN(n38369) );
  XNOR2HSV4 U43188 ( .A1(n38370), .A2(n38369), .ZN(n38467) );
  NAND3HSV4 U43189 ( .A1(n38374), .A2(n38373), .A3(n38372), .ZN(n38458) );
  CLKNHSV4 U43190 ( .I(n38458), .ZN(n46120) );
  NOR2HSV2 U43191 ( .A1(n46121), .A2(n38184), .ZN(n38376) );
  NOR2HSV4 U43192 ( .A1(n46120), .A2(n38376), .ZN(n38381) );
  INHSV2 U43193 ( .I(n38378), .ZN(n38379) );
  CLKNAND2HSV4 U43194 ( .A1(n38381), .A2(n38380), .ZN(n38601) );
  CLKNHSV0 U43195 ( .I(n38470), .ZN(n38386) );
  OAI21HSV0 U43196 ( .A1(n38383), .A2(n38386), .B(n38382), .ZN(n38384) );
  INHSV2 U43197 ( .I(n38384), .ZN(n38385) );
  OAI21HSV4 U43198 ( .A1(n60020), .A2(n38386), .B(n38385), .ZN(n38440) );
  CLKNAND2HSV0 U43199 ( .A1(n45149), .A2(n43924), .ZN(n38439) );
  INHSV2 U43200 ( .I(n45248), .ZN(n43925) );
  NAND2HSV0 U43201 ( .A1(n52288), .A2(n43925), .ZN(n38437) );
  CLKNAND2HSV1 U43202 ( .A1(n44715), .A2(n38390), .ZN(n38433) );
  NOR2HSV0 U43203 ( .A1(n44049), .A2(n52430), .ZN(n38392) );
  NAND2HSV0 U43204 ( .A1(n36603), .A2(n44074), .ZN(n38391) );
  XOR2HSV0 U43205 ( .A1(n38392), .A2(n38391), .Z(n38398) );
  CLKNAND2HSV0 U43206 ( .A1(n38678), .A2(n38393), .ZN(n38396) );
  NAND2HSV0 U43207 ( .A1(n52104), .A2(n38394), .ZN(n38395) );
  XNOR2HSV1 U43208 ( .A1(n38396), .A2(n38395), .ZN(n38397) );
  XNOR2HSV1 U43209 ( .A1(n38398), .A2(n38397), .ZN(n38400) );
  XNOR2HSV1 U43210 ( .A1(n38400), .A2(n38399), .ZN(n38409) );
  NAND2HSV0 U43211 ( .A1(\pe2/aot [19]), .A2(n36608), .ZN(n38403) );
  INHSV2 U43212 ( .I(n43999), .ZN(n51726) );
  NAND2HSV0 U43213 ( .A1(n51726), .A2(n38401), .ZN(n38402) );
  XOR2HSV0 U43214 ( .A1(n38403), .A2(n38402), .Z(n38407) );
  CLKNAND2HSV1 U43215 ( .A1(n59971), .A2(\pe2/bq[23] ), .ZN(n45184) );
  CLKNAND2HSV1 U43216 ( .A1(n52289), .A2(n52988), .ZN(n38405) );
  XOR2HSV0 U43217 ( .A1(n45184), .A2(n38405), .Z(n38406) );
  XOR2HSV0 U43218 ( .A1(n38407), .A2(n38406), .Z(n38408) );
  XNOR2HSV1 U43219 ( .A1(n38409), .A2(n38408), .ZN(n38431) );
  NOR2HSV1 U43220 ( .A1(n38489), .A2(n38973), .ZN(n38430) );
  NAND2HSV2 U43221 ( .A1(n59587), .A2(\pe2/bq[28] ), .ZN(n38411) );
  NAND2HSV0 U43222 ( .A1(\pe2/aot [22]), .A2(\pe2/bq[26] ), .ZN(n38410) );
  XOR2HSV0 U43223 ( .A1(n38411), .A2(n38410), .Z(n38415) );
  NAND2HSV0 U43224 ( .A1(n59585), .A2(n52950), .ZN(n38413) );
  CLKNAND2HSV1 U43225 ( .A1(n51759), .A2(n52444), .ZN(n38412) );
  XOR2HSV0 U43226 ( .A1(n38413), .A2(n38412), .Z(n38414) );
  XOR2HSV0 U43227 ( .A1(n38415), .A2(n38414), .Z(n38425) );
  CLKNAND2HSV1 U43228 ( .A1(\pe2/aot [27]), .A2(\pe2/bq[21] ), .ZN(n38417) );
  NAND2HSV0 U43229 ( .A1(n38479), .A2(n38542), .ZN(n38416) );
  XOR2HSV0 U43230 ( .A1(n38417), .A2(n38416), .Z(n38423) );
  INHSV2 U43231 ( .I(\pe2/aot [16]), .ZN(n52226) );
  NAND2HSV2 U43232 ( .A1(n51743), .A2(n38549), .ZN(n38421) );
  NAND2HSV0 U43233 ( .A1(n52995), .A2(n38419), .ZN(n38420) );
  XOR2HSV0 U43234 ( .A1(n38421), .A2(n38420), .Z(n38422) );
  XOR2HSV0 U43235 ( .A1(n38423), .A2(n38422), .Z(n38424) );
  XOR2HSV0 U43236 ( .A1(n38425), .A2(n38424), .Z(n38427) );
  NAND2HSV0 U43237 ( .A1(n43950), .A2(n59983), .ZN(n38426) );
  XNOR2HSV1 U43238 ( .A1(n38427), .A2(n38426), .ZN(n38429) );
  CLKNAND2HSV1 U43239 ( .A1(n38539), .A2(n52533), .ZN(n38428) );
  XOR4HSV1 U43240 ( .A1(n38431), .A2(n38430), .A3(n38429), .A4(n38428), .Z(
        n38432) );
  XNOR2HSV1 U43241 ( .A1(n38433), .A2(n38432), .ZN(n38435) );
  CLKNAND2HSV1 U43242 ( .A1(n38702), .A2(n52167), .ZN(n38434) );
  XNOR2HSV1 U43243 ( .A1(n38435), .A2(n38434), .ZN(n38436) );
  XNOR2HSV1 U43244 ( .A1(n38437), .A2(n38436), .ZN(n38438) );
  NAND2HSV2 U43245 ( .A1(n38447), .A2(n38603), .ZN(n38449) );
  OAI22HSV4 U43246 ( .A1(n38450), .A2(n38449), .B1(n36319), .B2(n38448), .ZN(
        n38451) );
  CLKNAND2HSV1 U43247 ( .A1(n38454), .A2(\pe2/ti_7t [17]), .ZN(n38611) );
  NOR2HSV4 U43248 ( .A1(n38456), .A2(n38455), .ZN(n38515) );
  CLKNHSV2 U43249 ( .I(n38518), .ZN(n38465) );
  INHSV2 U43250 ( .I(n38459), .ZN(n38461) );
  XNOR2HSV4 U43251 ( .A1(n38467), .A2(n38466), .ZN(n38887) );
  INHSV1 U43252 ( .I(n38889), .ZN(n38535) );
  CLKNAND2HSV2 U43253 ( .A1(n38607), .A2(n38264), .ZN(n38468) );
  NAND2HSV4 U43254 ( .A1(n38469), .A2(n38601), .ZN(n52809) );
  INHSV4 U43255 ( .I(n52809), .ZN(n38517) );
  NAND2HSV4 U43256 ( .A1(n38903), .A2(n45388), .ZN(n38614) );
  INHSV2 U43257 ( .I(n38471), .ZN(n52773) );
  INHSV2 U43258 ( .I(n52773), .ZN(n51802) );
  NAND2HSV2 U43259 ( .A1(n39011), .A2(n43925), .ZN(n38509) );
  NAND2HSV0 U43260 ( .A1(\pe2/aot [22]), .A2(n52950), .ZN(n38474) );
  CLKNAND2HSV0 U43261 ( .A1(n59971), .A2(n52299), .ZN(n38473) );
  XOR2HSV0 U43262 ( .A1(n38474), .A2(n38473), .Z(n38478) );
  CLKNAND2HSV1 U43263 ( .A1(n52070), .A2(n38549), .ZN(n38476) );
  CLKNAND2HSV1 U43264 ( .A1(\pe2/aot [17]), .A2(n38043), .ZN(n38475) );
  XOR2HSV0 U43265 ( .A1(n38476), .A2(n38475), .Z(n38477) );
  XOR2HSV0 U43266 ( .A1(n38478), .A2(n38477), .Z(n38488) );
  NAND2HSV0 U43267 ( .A1(n59970), .A2(\pe2/bq[21] ), .ZN(n38481) );
  NAND2HSV0 U43268 ( .A1(n38479), .A2(n52179), .ZN(n38480) );
  XOR2HSV0 U43269 ( .A1(n38481), .A2(n38480), .Z(n38486) );
  CLKNAND2HSV0 U43270 ( .A1(\pe2/aot [19]), .A2(n38565), .ZN(n38484) );
  INHSV2 U43271 ( .I(n38482), .ZN(n39014) );
  CLKNAND2HSV0 U43272 ( .A1(n39014), .A2(n52444), .ZN(n38483) );
  XOR2HSV0 U43273 ( .A1(n38484), .A2(n38483), .Z(n38485) );
  XOR2HSV0 U43274 ( .A1(n38486), .A2(n38485), .Z(n38487) );
  BUFHSV2 U43275 ( .I(n44002), .Z(n53064) );
  NAND2HSV2 U43276 ( .A1(n44976), .A2(n52984), .ZN(n38491) );
  NAND2HSV0 U43277 ( .A1(n38678), .A2(n44759), .ZN(n38490) );
  CLKNAND2HSV1 U43278 ( .A1(n38576), .A2(\pe2/pvq [18]), .ZN(n38492) );
  XOR2HSV0 U43279 ( .A1(n38492), .A2(\pe2/phq [18]), .Z(n38497) );
  CLKNHSV0 U43280 ( .I(n36240), .ZN(n44750) );
  INHSV2 U43281 ( .I(n48066), .ZN(n52215) );
  AOI22HSV0 U43282 ( .A1(n44750), .A2(n52215), .B1(n59969), .B2(n44074), .ZN(
        n38493) );
  AOI21HSV0 U43283 ( .A1(n38495), .A2(n38494), .B(n38493), .ZN(n38496) );
  NAND2HSV0 U43284 ( .A1(n59587), .A2(\pe2/bq[18] ), .ZN(n44238) );
  OAI22HSV0 U43285 ( .A1(n38787), .A2(n48064), .B1(n50947), .B2(n36530), .ZN(
        n38498) );
  OAI21HSV0 U43286 ( .A1(n44238), .A2(n38499), .B(n38498), .ZN(n38501) );
  NOR2HSV1 U43287 ( .A1(n37940), .A2(n45199), .ZN(n38500) );
  NOR2HSV0 U43288 ( .A1(n47573), .A2(n38213), .ZN(n38503) );
  NAND2HSV0 U43289 ( .A1(n59585), .A2(n38542), .ZN(n38502) );
  XOR2HSV0 U43290 ( .A1(n38503), .A2(n38502), .Z(n38507) );
  CLKNAND2HSV0 U43291 ( .A1(\pe2/aot [27]), .A2(n38920), .ZN(n38505) );
  NAND2HSV0 U43292 ( .A1(n52104), .A2(n52952), .ZN(n38504) );
  XOR2HSV0 U43293 ( .A1(n38505), .A2(n38504), .Z(n38506) );
  NAND2HSV2 U43294 ( .A1(n38510), .A2(n43924), .ZN(n38511) );
  XNOR2HSV4 U43295 ( .A1(n38614), .A2(n38513), .ZN(n38516) );
  NOR2HSV4 U43296 ( .A1(n38515), .A2(n38514), .ZN(n38615) );
  XNOR2HSV4 U43297 ( .A1(n38516), .A2(n38615), .ZN(n38613) );
  INHSV4 U43298 ( .I(n38613), .ZN(n38525) );
  NOR2HSV4 U43299 ( .A1(n38517), .A2(n38525), .ZN(n38521) );
  OR2HSV1 U43300 ( .A1(n38611), .A2(n44307), .Z(n38520) );
  INHSV4 U43301 ( .I(n38524), .ZN(n38526) );
  BUFHSV8 U43302 ( .I(n38526), .Z(n52808) );
  NAND2HSV2 U43303 ( .A1(n38526), .A2(n52809), .ZN(n38522) );
  INHSV2 U43304 ( .I(n38890), .ZN(n52559) );
  NOR2HSV4 U43305 ( .A1(n38536), .A2(n52559), .ZN(n38616) );
  NOR2HSV2 U43306 ( .A1(n38616), .A2(n37931), .ZN(n38732) );
  CLKNAND2HSV3 U43307 ( .A1(n38736), .A2(n38732), .ZN(n38531) );
  NAND2HSV2 U43308 ( .A1(n38524), .A2(n38613), .ZN(n38527) );
  CLKNHSV0 U43309 ( .I(n38616), .ZN(n38528) );
  NOR2HSV2 U43310 ( .A1(n38528), .A2(n59586), .ZN(n38737) );
  INHSV2 U43311 ( .I(\pe2/ti_7t [18]), .ZN(n38612) );
  NOR2HSV2 U43312 ( .A1(n44309), .A2(n38612), .ZN(n38741) );
  AOI21HSV4 U43313 ( .A1(n38739), .A2(n38737), .B(n38741), .ZN(n38530) );
  AOI21HSV0 U43314 ( .A1(n44043), .A2(n38340), .B(n38889), .ZN(n38532) );
  INHSV2 U43315 ( .I(n38532), .ZN(n38533) );
  OAI21HSV4 U43316 ( .A1(n38535), .A2(n38534), .B(n38533), .ZN(n38772) );
  AND2HSV4 U43317 ( .A1(n38645), .A2(n36661), .Z(n38600) );
  CLKNHSV2 U43318 ( .I(n38538), .ZN(n38597) );
  CLKNAND2HSV2 U43319 ( .A1(n26098), .A2(\pe2/got [28]), .ZN(n38596) );
  NOR2HSV2 U43320 ( .A1(n45148), .A2(n38902), .ZN(n38594) );
  CLKNAND2HSV0 U43321 ( .A1(n44711), .A2(n51966), .ZN(n38592) );
  CLKBUFHSV4 U43322 ( .I(n43999), .Z(n52526) );
  NOR2HSV0 U43323 ( .A1(n53033), .A2(n52526), .ZN(n38588) );
  CLKNAND2HSV0 U43324 ( .A1(n38539), .A2(n38782), .ZN(n38587) );
  NAND2HSV0 U43325 ( .A1(n52995), .A2(\pe2/bq[18] ), .ZN(n38541) );
  INHSV2 U43326 ( .I(n48066), .ZN(n52337) );
  CLKNAND2HSV0 U43327 ( .A1(n38061), .A2(n52337), .ZN(n38540) );
  XOR2HSV0 U43328 ( .A1(n38541), .A2(n38540), .Z(n38546) );
  NAND2HSV0 U43329 ( .A1(\pe2/aot [22]), .A2(n38542), .ZN(n38544) );
  CLKNAND2HSV0 U43330 ( .A1(n45024), .A2(n39020), .ZN(n38543) );
  XOR2HSV0 U43331 ( .A1(n38544), .A2(n38543), .Z(n38545) );
  XOR2HSV0 U43332 ( .A1(n38546), .A2(n38545), .Z(n38555) );
  XOR2HSV0 U43333 ( .A1(n38548), .A2(n38547), .Z(n38553) );
  NOR2HSV0 U43334 ( .A1(n44095), .A2(n52429), .ZN(n38551) );
  NAND2HSV0 U43335 ( .A1(n51920), .A2(n38549), .ZN(n38550) );
  XOR2HSV0 U43336 ( .A1(n38551), .A2(n38550), .Z(n38552) );
  XOR2HSV0 U43337 ( .A1(n38553), .A2(n38552), .Z(n38554) );
  XOR2HSV0 U43338 ( .A1(n38555), .A2(n38554), .Z(n38557) );
  INHSV2 U43339 ( .I(n47573), .ZN(n43926) );
  NAND2HSV0 U43340 ( .A1(n43950), .A2(n43926), .ZN(n38556) );
  XNOR2HSV1 U43341 ( .A1(n38557), .A2(n38556), .ZN(n38585) );
  NAND2HSV0 U43342 ( .A1(n45005), .A2(n44074), .ZN(n38560) );
  NAND2HSV0 U43343 ( .A1(n38558), .A2(\pe2/bq[14] ), .ZN(n38559) );
  XOR2HSV0 U43344 ( .A1(n38560), .A2(n38559), .Z(n38564) );
  NAND2HSV0 U43345 ( .A1(\pe2/aot [26]), .A2(n44197), .ZN(n38562) );
  NAND2HSV0 U43346 ( .A1(n59585), .A2(\pe2/bq[23] ), .ZN(n38561) );
  XOR2HSV0 U43347 ( .A1(n38562), .A2(n38561), .Z(n38563) );
  XOR2HSV0 U43348 ( .A1(n38564), .A2(n38563), .Z(n38573) );
  CLKNAND2HSV0 U43349 ( .A1(n38678), .A2(n38565), .ZN(n38567) );
  NAND2HSV0 U43350 ( .A1(\pe2/aot [19]), .A2(n38394), .ZN(n38566) );
  XOR2HSV0 U43351 ( .A1(n38567), .A2(n38566), .Z(n38571) );
  CLKNAND2HSV0 U43352 ( .A1(n44207), .A2(n38803), .ZN(n38569) );
  NAND2HSV0 U43353 ( .A1(n59354), .A2(n38401), .ZN(n38568) );
  XOR2HSV0 U43354 ( .A1(n38569), .A2(n38568), .Z(n38570) );
  XOR2HSV0 U43355 ( .A1(n38571), .A2(n38570), .Z(n38572) );
  XOR2HSV0 U43356 ( .A1(n38573), .A2(n38572), .Z(n38583) );
  NAND2HSV0 U43357 ( .A1(n59587), .A2(n52952), .ZN(n38575) );
  NAND2HSV0 U43358 ( .A1(\pe2/aot [17]), .A2(n44759), .ZN(n38574) );
  XOR2HSV0 U43359 ( .A1(n38575), .A2(n38574), .Z(n38579) );
  NAND2HSV0 U43360 ( .A1(n38576), .A2(\pe2/pvq [19]), .ZN(n38577) );
  XNOR2HSV1 U43361 ( .A1(n38577), .A2(\pe2/phq [19]), .ZN(n38578) );
  XNOR2HSV1 U43362 ( .A1(n38579), .A2(n38578), .ZN(n38581) );
  NAND2HSV0 U43363 ( .A1(\pe2/aot [21]), .A2(n44987), .ZN(n45189) );
  CLKNAND2HSV0 U43364 ( .A1(n59974), .A2(n52444), .ZN(n38810) );
  XOR2HSV0 U43365 ( .A1(n45189), .A2(n38810), .Z(n38580) );
  XNOR2HSV1 U43366 ( .A1(n38581), .A2(n38580), .ZN(n38582) );
  XNOR2HSV1 U43367 ( .A1(n38583), .A2(n38582), .ZN(n38584) );
  XOR2HSV0 U43368 ( .A1(n38585), .A2(n38584), .Z(n38586) );
  XOR3HSV2 U43369 ( .A1(n38588), .A2(n38587), .A3(n38586), .Z(n38589) );
  INAND2HSV2 U43370 ( .A1(n52164), .B1(n25940), .ZN(n38590) );
  XOR3HSV2 U43371 ( .A1(n38592), .A2(n38591), .A3(n38590), .Z(n38593) );
  XNOR2HSV4 U43372 ( .A1(n38594), .A2(n38593), .ZN(n38595) );
  XNOR2HSV4 U43373 ( .A1(n38600), .A2(n38599), .ZN(n38634) );
  NAND2HSV0 U43374 ( .A1(n38604), .A2(n38603), .ZN(n38605) );
  OR2HSV1 U43375 ( .A1(n38611), .A2(n39105), .Z(n38608) );
  NAND3HSV4 U43376 ( .A1(n38610), .A2(n38609), .A3(n38608), .ZN(n38633) );
  XNOR2HSV4 U43377 ( .A1(n38634), .A2(n38633), .ZN(n38624) );
  AOI21HSV2 U43378 ( .A1(n38612), .A2(n38099), .B(n38013), .ZN(n52811) );
  NAND2HSV2 U43379 ( .A1(n38625), .A2(n52811), .ZN(n38747) );
  NAND3HSV2 U43380 ( .A1(n38618), .A2(n38617), .A3(n52811), .ZN(n38750) );
  OAI21HSV2 U43381 ( .A1(n38626), .A2(n38750), .B(n44309), .ZN(n38619) );
  NOR2HSV4 U43382 ( .A1(n38620), .A2(n38619), .ZN(n38635) );
  INHSV2 U43383 ( .I(\pe2/ti_7t [19]), .ZN(n38621) );
  NOR2HSV2 U43384 ( .A1(n45265), .A2(n38621), .ZN(n38752) );
  INHSV2 U43385 ( .I(n38752), .ZN(n38622) );
  NOR2HSV2 U43386 ( .A1(n38623), .A2(n38629), .ZN(n38749) );
  NOR2HSV3 U43387 ( .A1(n38624), .A2(n38759), .ZN(n38628) );
  CLKNAND2HSV2 U43388 ( .A1(n38626), .A2(n44309), .ZN(n52813) );
  NAND2HSV1 U43389 ( .A1(n52811), .A2(n38627), .ZN(n38757) );
  NAND2HSV4 U43390 ( .A1(n38628), .A2(n38876), .ZN(n38872) );
  CLKNAND2HSV4 U43391 ( .A1(n38871), .A2(n38872), .ZN(n44807) );
  NOR2HSV4 U43392 ( .A1(n44807), .A2(n38629), .ZN(n38773) );
  CLKNAND2HSV1 U43393 ( .A1(n38772), .A2(n38773), .ZN(n38643) );
  NOR2HSV2 U43394 ( .A1(n38887), .A2(n44827), .ZN(n38767) );
  CLKNHSV0 U43395 ( .I(n52824), .ZN(n38631) );
  INHSV2 U43396 ( .I(n38630), .ZN(n39007) );
  NAND2HSV0 U43397 ( .A1(n38631), .A2(n39007), .ZN(n38636) );
  CLKNHSV2 U43398 ( .I(n38636), .ZN(n38632) );
  OR2HSV1 U43399 ( .A1(n38767), .A2(n38632), .Z(n38640) );
  CLKNHSV0 U43400 ( .I(n38872), .ZN(n38639) );
  CLKNAND2HSV0 U43401 ( .A1(n38635), .A2(n52815), .ZN(n38637) );
  CLKNAND2HSV1 U43402 ( .A1(n38637), .A2(n38636), .ZN(n38638) );
  OAI22HSV2 U43403 ( .A1(n38641), .A2(n38640), .B1(n38639), .B2(n38638), .ZN(
        n38642) );
  NAND2HSV2 U43404 ( .A1(n38643), .A2(n38642), .ZN(n38766) );
  NOR2HSV2 U43405 ( .A1(n44331), .A2(n38644), .ZN(n38728) );
  INHSV1 U43406 ( .I(n38645), .ZN(n38646) );
  NAND2HSV2 U43407 ( .A1(n59505), .A2(n38777), .ZN(n38727) );
  CLKNAND2HSV1 U43408 ( .A1(n39009), .A2(n38324), .ZN(n38720) );
  CLKNHSV2 U43409 ( .I(n38779), .ZN(n52419) );
  CLKNAND2HSV1 U43410 ( .A1(\pe2/got [23]), .A2(n52419), .ZN(n38718) );
  CLKNAND2HSV0 U43411 ( .A1(n38780), .A2(n38904), .ZN(n38715) );
  NAND2HSV0 U43412 ( .A1(n39011), .A2(n52533), .ZN(n38708) );
  NAND2HSV0 U43413 ( .A1(n48896), .A2(n38781), .ZN(n38706) );
  NOR2HSV0 U43414 ( .A1(n53033), .A2(n47498), .ZN(n38699) );
  BUFHSV2 U43415 ( .I(n44187), .Z(n44046) );
  CLKNAND2HSV0 U43416 ( .A1(n44046), .A2(n43926), .ZN(n38698) );
  NAND2HSV0 U43417 ( .A1(n51759), .A2(n38394), .ZN(n38648) );
  NAND2HSV0 U43418 ( .A1(\pe2/got [12]), .A2(n38401), .ZN(n38647) );
  XOR2HSV0 U43419 ( .A1(n38648), .A2(n38647), .Z(n38652) );
  NAND2HSV0 U43420 ( .A1(n59974), .A2(n44759), .ZN(n38650) );
  NAND2HSV0 U43421 ( .A1(\pe2/aot [22]), .A2(\pe2/bq[22] ), .ZN(n38649) );
  XOR2HSV0 U43422 ( .A1(n38650), .A2(n38649), .Z(n38651) );
  XOR2HSV0 U43423 ( .A1(n38652), .A2(n38651), .Z(n38661) );
  CLKNAND2HSV0 U43424 ( .A1(n45024), .A2(n38565), .ZN(n38654) );
  NAND2HSV0 U43425 ( .A1(\pe2/aot [19]), .A2(n52950), .ZN(n38653) );
  XOR2HSV0 U43426 ( .A1(n38654), .A2(n38653), .Z(n38659) );
  INHSV2 U43427 ( .I(n47599), .ZN(n38920) );
  CLKNAND2HSV0 U43428 ( .A1(n50956), .A2(n38920), .ZN(n38657) );
  NAND2HSV0 U43429 ( .A1(\pe2/aot [12]), .A2(n53015), .ZN(n38656) );
  XOR2HSV0 U43430 ( .A1(n38657), .A2(n38656), .Z(n38658) );
  XOR2HSV0 U43431 ( .A1(n38659), .A2(n38658), .Z(n38660) );
  XOR2HSV0 U43432 ( .A1(n38661), .A2(n38660), .Z(n38677) );
  NAND2HSV0 U43433 ( .A1(n44081), .A2(n38803), .ZN(n38663) );
  INHSV2 U43434 ( .I(n38822), .ZN(n45034) );
  CLKNAND2HSV0 U43435 ( .A1(n45034), .A2(n36480), .ZN(n38662) );
  XOR2HSV0 U43436 ( .A1(n38663), .A2(n38662), .Z(n38668) );
  NAND2HSV0 U43437 ( .A1(n38048), .A2(n38792), .ZN(n38666) );
  CLKNAND2HSV0 U43438 ( .A1(n39029), .A2(n52179), .ZN(n38665) );
  XOR2HSV0 U43439 ( .A1(n38666), .A2(n38665), .Z(n38667) );
  XOR2HSV0 U43440 ( .A1(n38668), .A2(n38667), .Z(n38675) );
  NAND2HSV0 U43441 ( .A1(n46623), .A2(\pe2/pvq [21]), .ZN(n38669) );
  XOR2HSV0 U43442 ( .A1(n38669), .A2(\pe2/phq [21]), .Z(n38673) );
  CLKNAND2HSV0 U43443 ( .A1(n59636), .A2(\pe2/bq[14] ), .ZN(n49541) );
  OAI22HSV1 U43444 ( .A1(n38404), .A2(n47580), .B1(n45165), .B2(n44699), .ZN(
        n38670) );
  OAI21HSV2 U43445 ( .A1(n38671), .A2(n49541), .B(n38670), .ZN(n38672) );
  XOR2HSV0 U43446 ( .A1(n38673), .A2(n38672), .Z(n38674) );
  XNOR2HSV1 U43447 ( .A1(n38675), .A2(n38674), .ZN(n38676) );
  XNOR2HSV1 U43448 ( .A1(n38677), .A2(n38676), .ZN(n38696) );
  CLKNAND2HSV0 U43449 ( .A1(n44892), .A2(n53006), .ZN(n38680) );
  NAND2HSV0 U43450 ( .A1(n38678), .A2(n52952), .ZN(n38679) );
  XOR2HSV0 U43451 ( .A1(n38680), .A2(n38679), .Z(n38684) );
  NAND2HSV0 U43452 ( .A1(n45005), .A2(n52337), .ZN(n38682) );
  INHSV2 U43453 ( .I(n49628), .ZN(n52472) );
  NAND2HSV0 U43454 ( .A1(n36603), .A2(n52472), .ZN(n38681) );
  XOR2HSV0 U43455 ( .A1(n38682), .A2(n38681), .Z(n38683) );
  XOR2HSV0 U43456 ( .A1(n38684), .A2(n38683), .Z(n38692) );
  NOR2HSV0 U43457 ( .A1(n44095), .A2(n44844), .ZN(n38686) );
  NAND2HSV0 U43458 ( .A1(n52974), .A2(\pe2/bq[18] ), .ZN(n38685) );
  XOR2HSV0 U43459 ( .A1(n38686), .A2(n38685), .Z(n38690) );
  NAND2HSV0 U43460 ( .A1(n59585), .A2(\pe2/bq[21] ), .ZN(n38820) );
  NAND2HSV0 U43461 ( .A1(n39052), .A2(\pe2/bq[24] ), .ZN(n38688) );
  XOR2HSV0 U43462 ( .A1(n38820), .A2(n38688), .Z(n38689) );
  XOR2HSV0 U43463 ( .A1(n38690), .A2(n38689), .Z(n38691) );
  XOR2HSV0 U43464 ( .A1(n38692), .A2(n38691), .Z(n38694) );
  CLKNHSV0 U43465 ( .I(n51607), .ZN(n39089) );
  NAND2HSV0 U43466 ( .A1(n39061), .A2(n39089), .ZN(n38693) );
  XNOR2HSV1 U43467 ( .A1(n38694), .A2(n38693), .ZN(n38695) );
  XOR2HSV0 U43468 ( .A1(n38696), .A2(n38695), .Z(n38697) );
  XOR3HSV2 U43469 ( .A1(n38699), .A2(n38698), .A3(n38697), .Z(n38701) );
  NAND2HSV0 U43470 ( .A1(n43928), .A2(\pe2/got [16]), .ZN(n38700) );
  XOR2HSV0 U43471 ( .A1(n38701), .A2(n38700), .Z(n38704) );
  NAND2HSV0 U43472 ( .A1(n38702), .A2(n59983), .ZN(n38703) );
  XNOR2HSV1 U43473 ( .A1(n38704), .A2(n38703), .ZN(n38705) );
  XNOR2HSV1 U43474 ( .A1(n38706), .A2(n38705), .ZN(n38707) );
  XNOR2HSV1 U43475 ( .A1(n38708), .A2(n38707), .ZN(n38710) );
  CLKNAND2HSV0 U43476 ( .A1(n38510), .A2(n39010), .ZN(n38709) );
  XOR2HSV0 U43477 ( .A1(n38710), .A2(n38709), .Z(n38713) );
  NAND2HSV0 U43478 ( .A1(n45218), .A2(n52167), .ZN(n38712) );
  XNOR2HSV1 U43479 ( .A1(n38713), .A2(n38712), .ZN(n38714) );
  XNOR2HSV1 U43480 ( .A1(n38715), .A2(n38714), .ZN(n38717) );
  NAND2HSV2 U43481 ( .A1(n25940), .A2(\pe2/got [24]), .ZN(n38716) );
  XOR3HSV2 U43482 ( .A1(n38718), .A2(n38717), .A3(n38716), .Z(n38719) );
  XOR2HSV0 U43483 ( .A1(n38720), .A2(n38719), .Z(n38721) );
  XNOR2HSV1 U43484 ( .A1(n38722), .A2(n38721), .ZN(n38725) );
  XNOR2HSV1 U43485 ( .A1(n38725), .A2(n38724), .ZN(n38726) );
  XNOR2HSV1 U43486 ( .A1(n38727), .A2(n38726), .ZN(n38729) );
  CLKNHSV0 U43487 ( .I(n38732), .ZN(n38734) );
  NOR2HSV2 U43488 ( .A1(n38734), .A2(n38733), .ZN(n38735) );
  CLKNAND2HSV2 U43489 ( .A1(n38736), .A2(n38735), .ZN(n38744) );
  AOI22HSV2 U43490 ( .A1(n38742), .A2(n38741), .B1(n38740), .B2(n38739), .ZN(
        n38743) );
  CLKNAND2HSV3 U43491 ( .A1(n38743), .A2(n38744), .ZN(n38745) );
  XNOR2HSV4 U43492 ( .A1(n38746), .A2(n38745), .ZN(n38765) );
  CLKNHSV0 U43493 ( .I(n38747), .ZN(n38748) );
  INAND2HSV2 U43494 ( .A1(n38749), .B1(n38748), .ZN(n38755) );
  CLKNHSV0 U43495 ( .I(n38750), .ZN(n38751) );
  AOI21HSV1 U43496 ( .A1(n52813), .A2(n38751), .B(n44314), .ZN(n38754) );
  AND2HSV2 U43497 ( .A1(n38752), .A2(n38890), .Z(n38753) );
  AOI31HSV2 U43498 ( .A1(n52815), .A2(n38755), .A3(n38754), .B(n38753), .ZN(
        n38763) );
  OR2HSV1 U43499 ( .A1(n38757), .A2(n39105), .Z(n38758) );
  NOR2HSV2 U43500 ( .A1(n38759), .A2(n38758), .ZN(n38760) );
  NAND2HSV2 U43501 ( .A1(n38762), .A2(n38763), .ZN(n38764) );
  XNOR2HSV4 U43502 ( .A1(n38765), .A2(n38764), .ZN(n38775) );
  INHSV4 U43503 ( .I(n38775), .ZN(n52822) );
  NAND2HSV4 U43504 ( .A1(n38766), .A2(n52822), .ZN(n44032) );
  NOR2HSV2 U43505 ( .A1(n38768), .A2(n38767), .ZN(n38770) );
  NAND2HSV2 U43506 ( .A1(n52824), .A2(n44309), .ZN(n38771) );
  NOR2HSV4 U43507 ( .A1(n52823), .A2(n38771), .ZN(n38774) );
  CLKNAND2HSV2 U43508 ( .A1(n38773), .A2(n38772), .ZN(n52825) );
  NAND3HSV4 U43509 ( .A1(n38775), .A2(n38774), .A3(n52825), .ZN(n44031) );
  NAND2HSV2 U43510 ( .A1(n44821), .A2(\pe2/ti_7t [21]), .ZN(n39006) );
  NAND3HSV3 U43511 ( .A1(n44032), .A2(n44031), .A3(n39006), .ZN(n44022) );
  NAND2HSV2 U43512 ( .A1(n44022), .A2(n47997), .ZN(n38884) );
  INHSV2 U43513 ( .I(n44043), .ZN(n45235) );
  CLKNHSV2 U43514 ( .I(n45235), .ZN(n38776) );
  CLKNHSV2 U43515 ( .I(n38776), .ZN(n38870) );
  INHSV2 U43516 ( .I(n44331), .ZN(n52173) );
  CLKNAND2HSV4 U43517 ( .A1(n51801), .A2(n38777), .ZN(n38866) );
  BUFHSV2 U43518 ( .I(n38903), .Z(n51965) );
  NAND2HSV2 U43519 ( .A1(n51965), .A2(n38324), .ZN(n38860) );
  CLKNAND2HSV1 U43520 ( .A1(n44713), .A2(n52416), .ZN(n38858) );
  CLKNHSV2 U43521 ( .I(n38779), .ZN(n52929) );
  NAND2HSV2 U43522 ( .A1(n38904), .A2(n52929), .ZN(n38856) );
  CLKNAND2HSV0 U43523 ( .A1(n38780), .A2(n52167), .ZN(n38853) );
  CLKNAND2HSV0 U43524 ( .A1(n39011), .A2(n38781), .ZN(n38847) );
  NAND2HSV2 U43525 ( .A1(n52053), .A2(n38782), .ZN(n38845) );
  CLKNAND2HSV0 U43526 ( .A1(n43928), .A2(n43926), .ZN(n38840) );
  INHSV2 U43527 ( .I(n47498), .ZN(n43927) );
  CLKNAND2HSV0 U43528 ( .A1(n44046), .A2(n43927), .ZN(n38784) );
  NOR2HSV0 U43529 ( .A1(n53033), .A2(n51607), .ZN(n38783) );
  XNOR2HSV1 U43530 ( .A1(n38784), .A2(n38783), .ZN(n38838) );
  CLKNHSV0 U43531 ( .I(n52103), .ZN(n44062) );
  CLKNAND2HSV0 U43532 ( .A1(n44062), .A2(n52950), .ZN(n38786) );
  NAND2HSV0 U43533 ( .A1(n39052), .A2(n52179), .ZN(n38785) );
  XOR2HSV0 U43534 ( .A1(n38786), .A2(n38785), .Z(n38791) );
  CLKNAND2HSV0 U43535 ( .A1(n39014), .A2(n39032), .ZN(n38789) );
  CLKNAND2HSV0 U43536 ( .A1(n59588), .A2(\pe2/bq[14] ), .ZN(n38788) );
  XOR2HSV0 U43537 ( .A1(n38789), .A2(n38788), .Z(n38790) );
  XOR2HSV0 U43538 ( .A1(n38791), .A2(n38790), .Z(n38800) );
  NAND2HSV0 U43539 ( .A1(n50956), .A2(n38792), .ZN(n38794) );
  NAND2HSV0 U43540 ( .A1(n44745), .A2(n44759), .ZN(n38793) );
  XOR2HSV0 U43541 ( .A1(n38794), .A2(n38793), .Z(n38798) );
  CLKNAND2HSV0 U43542 ( .A1(n44892), .A2(\pe2/bq[11] ), .ZN(n38796) );
  NAND2HSV0 U43543 ( .A1(n59968), .A2(n53006), .ZN(n38795) );
  XOR2HSV0 U43544 ( .A1(n38796), .A2(n38795), .Z(n38797) );
  XOR2HSV0 U43545 ( .A1(n38798), .A2(n38797), .Z(n38799) );
  XOR2HSV0 U43546 ( .A1(n38800), .A2(n38799), .Z(n38816) );
  NAND2HSV0 U43547 ( .A1(n39029), .A2(\pe2/bq[22] ), .ZN(n38802) );
  CLKNHSV0 U43548 ( .I(n49656), .ZN(n52374) );
  NAND2HSV0 U43549 ( .A1(n52374), .A2(n36602), .ZN(n38801) );
  XOR2HSV0 U43550 ( .A1(n38802), .A2(n38801), .Z(n38807) );
  CLKNAND2HSV1 U43551 ( .A1(n45295), .A2(n38803), .ZN(n38805) );
  CLKNAND2HSV0 U43552 ( .A1(n38048), .A2(n52988), .ZN(n38804) );
  XOR2HSV0 U43553 ( .A1(n38805), .A2(n38804), .Z(n38806) );
  XOR2HSV0 U43554 ( .A1(n38807), .A2(n38806), .Z(n38814) );
  NAND2HSV0 U43555 ( .A1(n46623), .A2(\pe2/pvq [22]), .ZN(n38808) );
  XOR2HSV0 U43556 ( .A1(n38808), .A2(\pe2/phq [22]), .Z(n38812) );
  CLKNAND2HSV1 U43557 ( .A1(n53005), .A2(n38565), .ZN(n43931) );
  OAI22HSV0 U43558 ( .A1(n36237), .A2(n51736), .B1(n47503), .B2(n36434), .ZN(
        n38809) );
  OAI21HSV1 U43559 ( .A1(n38810), .A2(n43931), .B(n38809), .ZN(n38811) );
  XOR2HSV0 U43560 ( .A1(n38812), .A2(n38811), .Z(n38813) );
  XNOR2HSV1 U43561 ( .A1(n38814), .A2(n38813), .ZN(n38815) );
  XNOR2HSV1 U43562 ( .A1(n38816), .A2(n38815), .ZN(n38836) );
  NAND2HSV0 U43563 ( .A1(\pe2/aot [19]), .A2(\pe2/bq[24] ), .ZN(n38818) );
  NAND2HSV0 U43564 ( .A1(\pe2/aot [11]), .A2(n38303), .ZN(n38817) );
  XOR2HSV0 U43565 ( .A1(n38818), .A2(n38817), .Z(n38832) );
  NAND2HSV0 U43566 ( .A1(\pe2/aot [22]), .A2(n38920), .ZN(n39058) );
  OAI22HSV0 U43567 ( .A1(n47574), .A2(n47599), .B1(n44871), .B2(n47608), .ZN(
        n38819) );
  OAI21HSV2 U43568 ( .A1(n38820), .A2(n39058), .B(n38819), .ZN(n38821) );
  NOR2HSV2 U43569 ( .A1(n44049), .A2(n44844), .ZN(n48943) );
  XNOR2HSV1 U43570 ( .A1(n38821), .A2(n48943), .ZN(n38831) );
  CLKNHSV0 U43571 ( .I(n48066), .ZN(n43956) );
  NAND2HSV0 U43572 ( .A1(n44081), .A2(n43956), .ZN(n38825) );
  INHSV2 U43573 ( .I(n38822), .ZN(n59975) );
  CLKNAND2HSV0 U43574 ( .A1(n59975), .A2(n39020), .ZN(n38824) );
  XOR2HSV0 U43575 ( .A1(n38825), .A2(n38824), .Z(n38829) );
  NAND2HSV0 U43576 ( .A1(n51759), .A2(n52952), .ZN(n38827) );
  NAND2HSV0 U43577 ( .A1(n44207), .A2(n51839), .ZN(n38826) );
  XOR2HSV0 U43578 ( .A1(n38827), .A2(n38826), .Z(n38828) );
  XOR2HSV0 U43579 ( .A1(n38829), .A2(n38828), .Z(n38830) );
  XOR3HSV2 U43580 ( .A1(n38832), .A2(n38831), .A3(n38830), .Z(n38834) );
  CLKNAND2HSV0 U43581 ( .A1(n39061), .A2(n52172), .ZN(n38833) );
  XNOR2HSV1 U43582 ( .A1(n38834), .A2(n38833), .ZN(n38835) );
  XOR2HSV0 U43583 ( .A1(n38836), .A2(n38835), .Z(n38837) );
  XNOR2HSV1 U43584 ( .A1(n38838), .A2(n38837), .ZN(n38839) );
  XNOR2HSV1 U43585 ( .A1(n38840), .A2(n38839), .ZN(n38843) );
  BUFHSV2 U43586 ( .I(n38841), .Z(n44254) );
  CLKNAND2HSV0 U43587 ( .A1(n44254), .A2(n51726), .ZN(n38842) );
  XNOR2HSV1 U43588 ( .A1(n38843), .A2(n38842), .ZN(n38844) );
  XNOR2HSV1 U43589 ( .A1(n38845), .A2(n38844), .ZN(n38846) );
  XNOR2HSV1 U43590 ( .A1(n38847), .A2(n38846), .ZN(n38849) );
  CLKBUFHSV4 U43591 ( .I(n52367), .Z(n45055) );
  NAND2HSV2 U43592 ( .A1(n45055), .A2(n39075), .ZN(n38848) );
  XOR2HSV0 U43593 ( .A1(n38849), .A2(n38848), .Z(n38851) );
  CLKNAND2HSV0 U43594 ( .A1(n45218), .A2(n39010), .ZN(n38850) );
  XNOR2HSV1 U43595 ( .A1(n38851), .A2(n38850), .ZN(n38852) );
  XNOR2HSV1 U43596 ( .A1(n38853), .A2(n38852), .ZN(n38855) );
  NAND2HSV2 U43597 ( .A1(n25939), .A2(\pe2/got [23]), .ZN(n38854) );
  XOR3HSV2 U43598 ( .A1(n38856), .A2(n38855), .A3(n38854), .Z(n38857) );
  XNOR2HSV1 U43599 ( .A1(n38858), .A2(n38857), .ZN(n38859) );
  XNOR2HSV1 U43600 ( .A1(n38860), .A2(n38859), .ZN(n38863) );
  INHSV4 U43601 ( .I(n38861), .ZN(n52251) );
  NAND2HSV2 U43602 ( .A1(n52251), .A2(n44944), .ZN(n38862) );
  XOR3HSV2 U43603 ( .A1(n38864), .A2(n38863), .A3(n38862), .Z(n38865) );
  XNOR2HSV4 U43604 ( .A1(n38866), .A2(n38865), .ZN(n38867) );
  CLKNAND2HSV4 U43605 ( .A1(n38867), .A2(n45388), .ZN(n38869) );
  XNOR2HSV2 U43606 ( .A1(n44043), .A2(n38887), .ZN(n38877) );
  XNOR2HSV4 U43607 ( .A1(n38877), .A2(n38894), .ZN(n38880) );
  NAND2HSV2 U43608 ( .A1(n38878), .A2(n38890), .ZN(n38879) );
  INHSV2 U43609 ( .I(n38882), .ZN(n38883) );
  XNOR2HSV4 U43610 ( .A1(n38884), .A2(n44034), .ZN(n60095) );
  INHSV2 U43611 ( .I(\pe2/ti_7t [22]), .ZN(n44027) );
  CLKNHSV1 U43612 ( .I(n38894), .ZN(n38892) );
  NOR2HSV1 U43613 ( .A1(n38887), .A2(n52559), .ZN(n38888) );
  NAND2HSV0 U43614 ( .A1(n38888), .A2(n44043), .ZN(n38893) );
  INHSV2 U43615 ( .I(n38895), .ZN(n38891) );
  NAND3HSV2 U43616 ( .A1(n38892), .A2(n38893), .A3(n38891), .ZN(n38898) );
  CLKNHSV0 U43617 ( .I(n38893), .ZN(n38896) );
  OAI21HSV2 U43618 ( .A1(n38896), .A2(n38895), .B(n38894), .ZN(n38897) );
  CLKNAND2HSV3 U43619 ( .A1(n38898), .A2(n38897), .ZN(n60021) );
  NAND2HSV0 U43620 ( .A1(\pe2/ti_7t [20]), .A2(n38899), .ZN(n43923) );
  CLKNHSV1 U43621 ( .I(n43923), .ZN(n39102) );
  OAI21HSV0 U43622 ( .A1(n38627), .A2(n39102), .B(n52916), .ZN(n38900) );
  INHSV2 U43623 ( .I(n38900), .ZN(n38901) );
  OAI21HSV1 U43624 ( .A1(n60021), .A2(n39102), .B(n38901), .ZN(n38999) );
  NAND2HSV2 U43625 ( .A1(n52924), .A2(n44944), .ZN(n38991) );
  CLKNAND2HSV0 U43626 ( .A1(n38778), .A2(n25824), .ZN(n38989) );
  CLKNAND2HSV1 U43627 ( .A1(n59773), .A2(n52416), .ZN(n38987) );
  BUFHSV2 U43628 ( .I(n26098), .Z(n45288) );
  CLKNAND2HSV1 U43629 ( .A1(n45288), .A2(\pe2/got [23]), .ZN(n38984) );
  CLKNAND2HSV0 U43630 ( .A1(n39009), .A2(n38904), .ZN(n38982) );
  NAND2HSV0 U43631 ( .A1(n39010), .A2(n51966), .ZN(n38980) );
  CLKNAND2HSV1 U43632 ( .A1(n38780), .A2(n39075), .ZN(n38977) );
  CLKNAND2HSV1 U43633 ( .A1(n44185), .A2(n51726), .ZN(n38969) );
  CLKNAND2HSV0 U43634 ( .A1(n52288), .A2(n43926), .ZN(n38967) );
  NAND2HSV0 U43635 ( .A1(n43928), .A2(n39089), .ZN(n38963) );
  NAND2HSV0 U43636 ( .A1(n44046), .A2(n52172), .ZN(n38906) );
  NOR2HSV0 U43637 ( .A1(n52420), .A2(n49656), .ZN(n38905) );
  XNOR2HSV1 U43638 ( .A1(n38906), .A2(n38905), .ZN(n38961) );
  INHSV2 U43639 ( .I(\pe2/got [10]), .ZN(n44045) );
  NOR2HSV1 U43640 ( .A1(n38907), .A2(n44045), .ZN(n38959) );
  NOR2HSV0 U43641 ( .A1(n44049), .A2(n48066), .ZN(n38909) );
  INHSV2 U43642 ( .I(\pe2/got [9]), .ZN(n44835) );
  NAND2HSV0 U43643 ( .A1(\pe2/got [9]), .A2(n45303), .ZN(n38908) );
  XOR2HSV0 U43644 ( .A1(n38909), .A2(n38908), .Z(n38913) );
  NAND2HSV0 U43645 ( .A1(\pe2/aot [20]), .A2(\pe2/bq[21] ), .ZN(n38911) );
  NAND2HSV0 U43646 ( .A1(n59972), .A2(n44074), .ZN(n38910) );
  XOR2HSV0 U43647 ( .A1(n38911), .A2(n38910), .Z(n38912) );
  XOR2HSV0 U43648 ( .A1(n38913), .A2(n38912), .Z(n38917) );
  NAND2HSV0 U43649 ( .A1(n48078), .A2(\pe2/pvq [24]), .ZN(n38914) );
  XNOR2HSV1 U43650 ( .A1(n38914), .A2(\pe2/phq [24]), .ZN(n38915) );
  INHSV2 U43651 ( .I(n49515), .ZN(n44090) );
  NAND2HSV0 U43652 ( .A1(n59968), .A2(n44090), .ZN(n52447) );
  XNOR2HSV1 U43653 ( .A1(n38915), .A2(n52447), .ZN(n38916) );
  XNOR2HSV1 U43654 ( .A1(n38917), .A2(n38916), .ZN(n38925) );
  NOR2HSV0 U43655 ( .A1(n44095), .A2(n47580), .ZN(n38919) );
  INHSV2 U43656 ( .I(n47511), .ZN(n52481) );
  CLKNAND2HSV0 U43657 ( .A1(n44892), .A2(n52481), .ZN(n38918) );
  XOR2HSV0 U43658 ( .A1(n38919), .A2(n38918), .Z(n38923) );
  CLKNAND2HSV0 U43659 ( .A1(n39029), .A2(n38920), .ZN(n45334) );
  NAND2HSV0 U43660 ( .A1(n38048), .A2(n52984), .ZN(n38921) );
  XOR2HSV0 U43661 ( .A1(n45334), .A2(n38921), .Z(n38922) );
  XOR2HSV0 U43662 ( .A1(n38923), .A2(n38922), .Z(n38924) );
  XNOR2HSV1 U43663 ( .A1(n38925), .A2(n38924), .ZN(n38958) );
  NAND2HSV0 U43664 ( .A1(n59588), .A2(n52438), .ZN(n38927) );
  CLKNHSV0 U43665 ( .I(n38418), .ZN(n43972) );
  NAND2HSV0 U43666 ( .A1(n53019), .A2(n43972), .ZN(n38926) );
  XOR2HSV0 U43667 ( .A1(n38927), .A2(n38926), .Z(n38931) );
  NAND2HSV0 U43668 ( .A1(n44062), .A2(n52179), .ZN(n38929) );
  INHSV2 U43669 ( .I(\pe2/aot [10]), .ZN(n43933) );
  INHSV2 U43670 ( .I(n43933), .ZN(n53009) );
  NAND2HSV0 U43671 ( .A1(n53009), .A2(n38046), .ZN(n38928) );
  XOR2HSV0 U43672 ( .A1(n38929), .A2(n38928), .Z(n38930) );
  XOR2HSV0 U43673 ( .A1(n38931), .A2(n38930), .Z(n38939) );
  NAND2HSV0 U43674 ( .A1(\pe2/aot [19]), .A2(\pe2/bq[22] ), .ZN(n38933) );
  NAND2HSV0 U43675 ( .A1(n53005), .A2(n36608), .ZN(n38932) );
  XOR2HSV0 U43676 ( .A1(n38933), .A2(n38932), .Z(n38937) );
  NAND2HSV0 U43677 ( .A1(n44745), .A2(n39032), .ZN(n38935) );
  NAND2HSV0 U43678 ( .A1(n50930), .A2(n52988), .ZN(n38934) );
  XOR2HSV0 U43679 ( .A1(n38935), .A2(n38934), .Z(n38936) );
  XOR2HSV0 U43680 ( .A1(n38937), .A2(n38936), .Z(n38938) );
  XOR2HSV0 U43681 ( .A1(n38939), .A2(n38938), .Z(n38956) );
  CLKNAND2HSV1 U43682 ( .A1(n52289), .A2(\pe2/bq[11] ), .ZN(n38941) );
  CLKNHSV0 U43683 ( .I(n44212), .ZN(n44081) );
  NAND2HSV0 U43684 ( .A1(n44081), .A2(n51839), .ZN(n38940) );
  XOR2HSV0 U43685 ( .A1(n38941), .A2(n38940), .Z(n38945) );
  NAND2HSV0 U43686 ( .A1(n39019), .A2(n39020), .ZN(n38943) );
  NAND2HSV0 U43687 ( .A1(\pe2/aot [22]), .A2(n43961), .ZN(n38942) );
  XOR2HSV0 U43688 ( .A1(n38943), .A2(n38942), .Z(n38944) );
  XOR2HSV0 U43689 ( .A1(n38945), .A2(n38944), .Z(n38954) );
  NAND2HSV0 U43690 ( .A1(\pe2/aot [17]), .A2(\pe2/bq[24] ), .ZN(n38948) );
  NAND2HSV0 U43691 ( .A1(n39014), .A2(n52950), .ZN(n38947) );
  XOR2HSV0 U43692 ( .A1(n38948), .A2(n38947), .Z(n38952) );
  NAND2HSV0 U43693 ( .A1(n59974), .A2(n38064), .ZN(n38950) );
  CLKNAND2HSV0 U43694 ( .A1(n45034), .A2(n52987), .ZN(n38949) );
  XOR2HSV0 U43695 ( .A1(n38950), .A2(n38949), .Z(n38951) );
  XOR2HSV0 U43696 ( .A1(n38952), .A2(n38951), .Z(n38953) );
  XOR2HSV0 U43697 ( .A1(n38954), .A2(n38953), .Z(n38955) );
  XOR2HSV0 U43698 ( .A1(n38956), .A2(n38955), .Z(n38957) );
  XOR3HSV2 U43699 ( .A1(n38959), .A2(n38958), .A3(n38957), .Z(n38960) );
  XNOR2HSV1 U43700 ( .A1(n38961), .A2(n38960), .ZN(n38962) );
  XNOR2HSV1 U43701 ( .A1(n38963), .A2(n38962), .ZN(n38965) );
  INHSV2 U43702 ( .I(n47498), .ZN(n48084) );
  NAND2HSV0 U43703 ( .A1(n44254), .A2(n48084), .ZN(n38964) );
  XNOR2HSV1 U43704 ( .A1(n38965), .A2(n38964), .ZN(n38966) );
  XNOR2HSV1 U43705 ( .A1(n38967), .A2(n38966), .ZN(n38968) );
  XNOR2HSV1 U43706 ( .A1(n38969), .A2(n38968), .ZN(n38971) );
  CLKNAND2HSV0 U43707 ( .A1(n45055), .A2(n59983), .ZN(n38970) );
  XOR2HSV0 U43708 ( .A1(n38971), .A2(n38970), .Z(n38975) );
  CLKNHSV0 U43709 ( .I(n44264), .ZN(n44120) );
  INHSV2 U43710 ( .I(n38973), .ZN(n52925) );
  CLKNAND2HSV0 U43711 ( .A1(n44120), .A2(n52925), .ZN(n38974) );
  XNOR2HSV1 U43712 ( .A1(n38975), .A2(n38974), .ZN(n38976) );
  XNOR2HSV1 U43713 ( .A1(n38977), .A2(n38976), .ZN(n38979) );
  BUFHSV4 U43714 ( .I(n29749), .Z(n51610) );
  NAND2HSV2 U43715 ( .A1(n51610), .A2(\pe2/got [21]), .ZN(n38978) );
  XOR3HSV2 U43716 ( .A1(n38980), .A2(n38979), .A3(n38978), .Z(n38981) );
  XNOR2HSV1 U43717 ( .A1(n38982), .A2(n38981), .ZN(n38983) );
  XNOR2HSV1 U43718 ( .A1(n38984), .A2(n38983), .ZN(n38986) );
  NOR2HSV2 U43719 ( .A1(n45071), .A2(n39088), .ZN(n38985) );
  XOR3HSV2 U43720 ( .A1(n38987), .A2(n38986), .A3(n38985), .Z(n38988) );
  XNOR2HSV1 U43721 ( .A1(n38989), .A2(n38988), .ZN(n38990) );
  XNOR2HSV1 U43722 ( .A1(n38991), .A2(n38990), .ZN(n38992) );
  OAI21HSV2 U43723 ( .A1(n44283), .A2(n38993), .B(n38992), .ZN(n38997) );
  CLKNHSV0 U43724 ( .I(n38992), .ZN(n38995) );
  NOR2HSV2 U43725 ( .A1(n44283), .A2(n38993), .ZN(n38994) );
  CLKNAND2HSV1 U43726 ( .A1(n38995), .A2(n38994), .ZN(n38996) );
  NAND2HSV2 U43727 ( .A1(n38997), .A2(n38996), .ZN(n38998) );
  XNOR2HSV2 U43728 ( .A1(n38999), .A2(n38998), .ZN(n39001) );
  NAND2HSV0 U43729 ( .A1(n44022), .A2(n59980), .ZN(n39000) );
  XNOR2HSV4 U43730 ( .A1(n39001), .A2(n39000), .ZN(n39002) );
  NAND3HSV4 U43731 ( .A1(n44032), .A2(n44031), .A3(n39006), .ZN(n60002) );
  NAND2HSV2 U43732 ( .A1(n45288), .A2(n39008), .ZN(n39087) );
  CLKNAND2HSV0 U43733 ( .A1(n39009), .A2(n45249), .ZN(n39085) );
  CLKNAND2HSV0 U43734 ( .A1(\pe2/got [21]), .A2(n51966), .ZN(n39083) );
  NAND2HSV2 U43735 ( .A1(n52176), .A2(n39010), .ZN(n39079) );
  NAND2HSV0 U43736 ( .A1(n39011), .A2(n59983), .ZN(n39072) );
  CLKNAND2HSV1 U43737 ( .A1(n45150), .A2(n51726), .ZN(n39070) );
  CLKNAND2HSV1 U43738 ( .A1(n44254), .A2(n43926), .ZN(n39068) );
  CLKNAND2HSV1 U43739 ( .A1(\pe2/aot [14]), .A2(n36588), .ZN(n39013) );
  CLKNAND2HSV1 U43740 ( .A1(n59975), .A2(n36608), .ZN(n39012) );
  XOR2HSV0 U43741 ( .A1(n39013), .A2(n39012), .Z(n39018) );
  NAND2HSV0 U43742 ( .A1(n39014), .A2(n38064), .ZN(n39016) );
  CLKNAND2HSV0 U43743 ( .A1(n51759), .A2(n52950), .ZN(n39015) );
  XOR2HSV0 U43744 ( .A1(n39016), .A2(n39015), .Z(n39017) );
  XOR2HSV0 U43745 ( .A1(n39018), .A2(n39017), .Z(n39028) );
  CLKNAND2HSV1 U43746 ( .A1(n39019), .A2(n36480), .ZN(n39022) );
  CLKNAND2HSV1 U43747 ( .A1(n53005), .A2(n39020), .ZN(n39021) );
  XOR2HSV0 U43748 ( .A1(n39022), .A2(n39021), .Z(n39026) );
  NAND2HSV2 U43749 ( .A1(n52974), .A2(n51732), .ZN(n39024) );
  CLKNAND2HSV1 U43750 ( .A1(n44062), .A2(\pe2/bq[24] ), .ZN(n39023) );
  XOR2HSV0 U43751 ( .A1(n39024), .A2(n39023), .Z(n39025) );
  XOR2HSV0 U43752 ( .A1(n39026), .A2(n39025), .Z(n39027) );
  XOR2HSV0 U43753 ( .A1(n39028), .A2(n39027), .Z(n39046) );
  CLKNAND2HSV1 U43754 ( .A1(n39029), .A2(\pe2/bq[21] ), .ZN(n39031) );
  INHSV2 U43755 ( .I(\pe2/aot [10]), .ZN(n52431) );
  CLKNAND2HSV1 U43756 ( .A1(n51460), .A2(n43972), .ZN(n39030) );
  XOR2HSV0 U43757 ( .A1(n39031), .A2(n39030), .Z(n39036) );
  CLKNAND2HSV1 U43758 ( .A1(n45295), .A2(n43956), .ZN(n39034) );
  CLKNAND2HSV0 U43759 ( .A1(n59974), .A2(n39032), .ZN(n39033) );
  XOR2HSV0 U43760 ( .A1(n39034), .A2(n39033), .Z(n39035) );
  XOR2HSV0 U43761 ( .A1(n39036), .A2(n39035), .Z(n39044) );
  NAND2HSV0 U43762 ( .A1(\pe2/aot [19]), .A2(n52179), .ZN(n39038) );
  NAND2HSV0 U43763 ( .A1(n44207), .A2(n52438), .ZN(n39037) );
  XOR2HSV0 U43764 ( .A1(n39038), .A2(n39037), .Z(n39042) );
  CLKNAND2HSV0 U43765 ( .A1(n59971), .A2(n44074), .ZN(n39040) );
  CLKNAND2HSV1 U43766 ( .A1(n59972), .A2(n52988), .ZN(n39039) );
  XOR2HSV0 U43767 ( .A1(n39040), .A2(n39039), .Z(n39041) );
  XOR2HSV0 U43768 ( .A1(n39042), .A2(n39041), .Z(n39043) );
  XOR2HSV0 U43769 ( .A1(n39044), .A2(n39043), .Z(n39045) );
  XOR2HSV0 U43770 ( .A1(n39046), .A2(n39045), .Z(n39066) );
  CLKNAND2HSV1 U43771 ( .A1(n59588), .A2(n51839), .ZN(n39048) );
  CLKNAND2HSV0 U43772 ( .A1(\pe2/got [10]), .A2(n36602), .ZN(n39047) );
  XOR2HSV0 U43773 ( .A1(n39048), .A2(n39047), .Z(n39051) );
  CLKNAND2HSV1 U43774 ( .A1(n44892), .A2(n44090), .ZN(n45294) );
  NAND2HSV0 U43775 ( .A1(\pe2/aot [23]), .A2(n43961), .ZN(n39049) );
  XOR2HSV0 U43776 ( .A1(n45294), .A2(n39049), .Z(n39050) );
  XOR2HSV0 U43777 ( .A1(n39051), .A2(n39050), .Z(n39064) );
  NAND2HSV0 U43778 ( .A1(n59968), .A2(n52073), .ZN(n39054) );
  NAND2HSV0 U43779 ( .A1(n39052), .A2(\pe2/bq[22] ), .ZN(n39053) );
  XOR2HSV0 U43780 ( .A1(n39054), .A2(n39053), .Z(n39057) );
  NAND2HSV0 U43781 ( .A1(n48078), .A2(\pe2/pvq [23]), .ZN(n39055) );
  XNOR2HSV1 U43782 ( .A1(n39055), .A2(\pe2/phq [23]), .ZN(n39056) );
  XNOR2HSV1 U43783 ( .A1(n39057), .A2(n39056), .ZN(n39060) );
  NAND2HSV2 U43784 ( .A1(n44081), .A2(\pe2/bq[14] ), .ZN(n44996) );
  XOR2HSV0 U43785 ( .A1(n39058), .A2(n44996), .Z(n39059) );
  XNOR2HSV1 U43786 ( .A1(n39060), .A2(n39059), .ZN(n39063) );
  CLKNHSV0 U43787 ( .I(n49656), .ZN(n44044) );
  CLKNAND2HSV1 U43788 ( .A1(n39061), .A2(n44044), .ZN(n39062) );
  XOR3HSV2 U43789 ( .A1(n39064), .A2(n39063), .A3(n39062), .Z(n39065) );
  XOR2HSV0 U43790 ( .A1(n39066), .A2(n39065), .Z(n39067) );
  XNOR2HSV1 U43791 ( .A1(n39068), .A2(n39067), .ZN(n39069) );
  XNOR2HSV1 U43792 ( .A1(n39070), .A2(n39069), .ZN(n39071) );
  XNOR2HSV1 U43793 ( .A1(n39072), .A2(n39071), .ZN(n39074) );
  CLKNAND2HSV1 U43794 ( .A1(n45055), .A2(n52925), .ZN(n39073) );
  XOR2HSV0 U43795 ( .A1(n39074), .A2(n39073), .Z(n39077) );
  CLKNAND2HSV1 U43796 ( .A1(n44120), .A2(n39075), .ZN(n39076) );
  XNOR2HSV1 U43797 ( .A1(n39077), .A2(n39076), .ZN(n39078) );
  XNOR2HSV1 U43798 ( .A1(n39079), .A2(n39078), .ZN(n39082) );
  CLKNAND2HSV1 U43799 ( .A1(n39080), .A2(n49591), .ZN(n39081) );
  XOR3HSV2 U43800 ( .A1(n39083), .A2(n39082), .A3(n39081), .Z(n39084) );
  XNOR2HSV1 U43801 ( .A1(n39085), .A2(n39084), .ZN(n39086) );
  XNOR2HSV1 U43802 ( .A1(n39087), .A2(n39086), .ZN(n39097) );
  NAND2HSV2 U43803 ( .A1(n43928), .A2(n43927), .ZN(n39093) );
  NAND2HSV2 U43804 ( .A1(n44046), .A2(n39089), .ZN(n39091) );
  NOR2HSV0 U43805 ( .A1(n52420), .A2(n47555), .ZN(n39090) );
  XOR2HSV0 U43806 ( .A1(n39091), .A2(n39090), .Z(n39092) );
  XOR2HSV0 U43807 ( .A1(n39093), .A2(n39092), .Z(n39094) );
  INHSV2 U43808 ( .I(n44331), .ZN(n51801) );
  NAND2HSV2 U43809 ( .A1(n44944), .A2(n52173), .ZN(n39095) );
  XOR3HSV2 U43810 ( .A1(n39097), .A2(n39096), .A3(n39095), .Z(n39098) );
  XNOR2HSV2 U43811 ( .A1(n39099), .A2(n39098), .ZN(n39101) );
  NAND2HSV2 U43812 ( .A1(n44807), .A2(n44145), .ZN(n39100) );
  XNOR2HSV4 U43813 ( .A1(n39101), .A2(n39100), .ZN(n39104) );
  OAI21HSV4 U43814 ( .A1(n60021), .A2(n39102), .B(n29723), .ZN(n39103) );
  XNOR2HSV4 U43815 ( .A1(n39104), .A2(n39103), .ZN(n39107) );
  XNOR2HSV4 U43816 ( .A1(n39107), .A2(n39106), .ZN(n39110) );
  XOR2HSV4 U43817 ( .A1(n39107), .A2(n39106), .Z(n39112) );
  CLKNAND2HSV4 U43818 ( .A1(n60095), .A2(n44312), .ZN(n44150) );
  AOI31HSV2 U43819 ( .A1(n26883), .A2(n44150), .A3(n44315), .B(n44316), .ZN(
        n39108) );
  CLKNAND2HSV2 U43820 ( .A1(n39109), .A2(n39108), .ZN(n44157) );
  INAND2HSV4 U43821 ( .A1(n52827), .B1(n44157), .ZN(n44176) );
  NOR2HSV4 U43822 ( .A1(n39110), .A2(n43916), .ZN(n44295) );
  INHSV2 U43823 ( .I(n43920), .ZN(n44149) );
  INHSV2 U43824 ( .I(n44149), .ZN(n39111) );
  NOR2HSV8 U43825 ( .A1(n44295), .A2(n39111), .ZN(n44183) );
  INHSV2 U43826 ( .I(n44150), .ZN(n39114) );
  CLKNAND2HSV4 U43827 ( .A1(n39114), .A2(n26883), .ZN(n44300) );
  CLKNAND2HSV0 U43828 ( .A1(n44821), .A2(\pe2/ti_7t [24]), .ZN(n44296) );
  INHSV2 U43829 ( .I(n44296), .ZN(n44298) );
  INHSV2 U43830 ( .I(n44298), .ZN(n44174) );
  INHSV3 U43831 ( .I(n44817), .ZN(n44943) );
  BUFHSV4 U43832 ( .I(n44943), .Z(n51894) );
  CLKNAND2HSV2 U43833 ( .A1(n60025), .A2(n39548), .ZN(n39115) );
  INAND2HSV4 U43834 ( .A1(n29722), .B1(n39115), .ZN(n40278) );
  INHSV2 U43835 ( .I(n30297), .ZN(n39879) );
  NAND2HSV2 U43836 ( .A1(n40278), .A2(n39879), .ZN(n39214) );
  NAND2HSV2 U43837 ( .A1(n40007), .A2(\pe5/ti_7t [20]), .ZN(n39428) );
  BUFHSV2 U43838 ( .I(n45900), .Z(n40020) );
  INHSV2 U43839 ( .I(n40020), .ZN(n48743) );
  CLKNAND2HSV1 U43840 ( .A1(n39256), .A2(n48743), .ZN(n39211) );
  CLKNHSV2 U43841 ( .I(n39118), .ZN(n45417) );
  BUFHSV2 U43842 ( .I(n45417), .Z(n40021) );
  NAND2HSV2 U43843 ( .A1(n40021), .A2(n39532), .ZN(n39207) );
  CLKBUFHSV2 U43844 ( .I(n45819), .Z(n51160) );
  CLKNAND2HSV0 U43845 ( .A1(n51160), .A2(n45816), .ZN(n39203) );
  CLKNAND2HSV1 U43846 ( .A1(n45820), .A2(n51103), .ZN(n39201) );
  CLKNAND2HSV1 U43847 ( .A1(n48748), .A2(n39433), .ZN(n39199) );
  INHSV2 U43848 ( .I(n50422), .ZN(n46974) );
  CLKNAND2HSV0 U43849 ( .A1(n30781), .A2(n46974), .ZN(n39197) );
  NAND2HSV0 U43850 ( .A1(n48624), .A2(n39881), .ZN(n39195) );
  NAND2HSV0 U43851 ( .A1(n59381), .A2(n39516), .ZN(n39193) );
  CLKNAND2HSV1 U43852 ( .A1(n48168), .A2(n48167), .ZN(n39188) );
  NAND2HSV0 U43853 ( .A1(n59639), .A2(n51305), .ZN(n39186) );
  NAND2HSV2 U43854 ( .A1(n39496), .A2(n50533), .ZN(n40227) );
  BUFHSV2 U43855 ( .I(n39122), .Z(n59427) );
  INHSV2 U43856 ( .I(\pe5/bq[7] ), .ZN(n47207) );
  CLKNAND2HSV1 U43857 ( .A1(n59427), .A2(\pe5/bq[7] ), .ZN(n40238) );
  CLKNAND2HSV0 U43858 ( .A1(n59366), .A2(\pe5/bq[7] ), .ZN(n39800) );
  OAI21HSV0 U43859 ( .A1(n47162), .A2(n39123), .B(n39800), .ZN(n39124) );
  OAI21HSV2 U43860 ( .A1(n40227), .A2(n40238), .B(n39124), .ZN(n39125) );
  NAND2HSV0 U43861 ( .A1(n39490), .A2(n46622), .ZN(n48680) );
  XNOR2HSV1 U43862 ( .A1(n39125), .A2(n48680), .ZN(n39129) );
  NAND2HSV2 U43863 ( .A1(n30788), .A2(n39454), .ZN(n39127) );
  NAND2HSV0 U43864 ( .A1(n39446), .A2(n39487), .ZN(n39126) );
  XOR2HSV0 U43865 ( .A1(n39127), .A2(n39126), .Z(n39128) );
  XNOR2HSV1 U43866 ( .A1(n39129), .A2(n39128), .ZN(n39146) );
  NAND2HSV0 U43867 ( .A1(n59642), .A2(n39130), .ZN(n39132) );
  NAND2HSV0 U43868 ( .A1(n39455), .A2(n48760), .ZN(n39131) );
  XOR2HSV0 U43869 ( .A1(n39132), .A2(n39131), .Z(n39136) );
  CLKNAND2HSV0 U43870 ( .A1(n39499), .A2(n39914), .ZN(n39134) );
  CLKNHSV0 U43871 ( .I(n48175), .ZN(n48829) );
  CLKNAND2HSV0 U43872 ( .A1(n48829), .A2(n39615), .ZN(n39133) );
  XOR2HSV0 U43873 ( .A1(n39134), .A2(n39133), .Z(n39135) );
  XOR2HSV0 U43874 ( .A1(n39136), .A2(n39135), .Z(n39142) );
  NAND2HSV0 U43875 ( .A1(n44335), .A2(\pe5/pvq [26]), .ZN(n39137) );
  XOR2HSV0 U43876 ( .A1(n39137), .A2(\pe5/phq [26]), .Z(n39140) );
  NAND2HSV2 U43877 ( .A1(n59941), .A2(n52610), .ZN(n39589) );
  NAND2HSV2 U43878 ( .A1(\pe5/aot [23]), .A2(n52595), .ZN(n39440) );
  OAI22HSV0 U43879 ( .A1(n40043), .A2(n39796), .B1(n45451), .B2(n45821), .ZN(
        n39138) );
  OAI21HSV1 U43880 ( .A1(n39589), .A2(n39440), .B(n39138), .ZN(n39139) );
  XOR2HSV0 U43881 ( .A1(n39140), .A2(n39139), .Z(n39141) );
  XNOR2HSV1 U43882 ( .A1(n39142), .A2(n39141), .ZN(n39145) );
  INHSV2 U43883 ( .I(n45901), .ZN(n47144) );
  NAND2HSV0 U43884 ( .A1(n30377), .A2(n47144), .ZN(n39144) );
  XOR3HSV2 U43885 ( .A1(n39146), .A2(n39145), .A3(n39144), .Z(n39148) );
  CLKNHSV0 U43886 ( .I(n30887), .ZN(n48751) );
  CLKNAND2HSV1 U43887 ( .A1(n48751), .A2(n51210), .ZN(n39147) );
  XNOR2HSV1 U43888 ( .A1(n39148), .A2(n39147), .ZN(n39184) );
  INHSV2 U43889 ( .I(n48204), .ZN(n48205) );
  NAND2HSV0 U43890 ( .A1(n48205), .A2(n45470), .ZN(n39150) );
  NAND2HSV0 U43891 ( .A1(n39887), .A2(n39495), .ZN(n39149) );
  XOR2HSV0 U43892 ( .A1(n39150), .A2(n39149), .Z(n39154) );
  NAND2HSV0 U43893 ( .A1(n59640), .A2(n31160), .ZN(n39152) );
  CLKNHSV0 U43894 ( .I(n48822), .ZN(n39921) );
  CLKNAND2HSV0 U43895 ( .A1(n48242), .A2(n39921), .ZN(n39151) );
  XOR2HSV0 U43896 ( .A1(n39152), .A2(n39151), .Z(n39153) );
  XOR2HSV0 U43897 ( .A1(n39154), .A2(n39153), .Z(n39162) );
  CLKNAND2HSV0 U43898 ( .A1(\pe5/aot [13]), .A2(n52594), .ZN(n39156) );
  NAND2HSV0 U43899 ( .A1(n40234), .A2(n39592), .ZN(n39155) );
  XOR2HSV0 U43900 ( .A1(n39156), .A2(n39155), .Z(n39160) );
  CLKNAND2HSV1 U43901 ( .A1(n59879), .A2(n50668), .ZN(n39158) );
  CLKNHSV0 U43902 ( .I(n30150), .ZN(n48634) );
  NAND2HSV0 U43903 ( .A1(n48634), .A2(n40221), .ZN(n39157) );
  XOR2HSV0 U43904 ( .A1(n39158), .A2(n39157), .Z(n39159) );
  XOR2HSV0 U43905 ( .A1(n39160), .A2(n39159), .Z(n39161) );
  XOR2HSV0 U43906 ( .A1(n39162), .A2(n39161), .Z(n39180) );
  INHSV2 U43907 ( .I(n48823), .ZN(n47278) );
  CLKNAND2HSV1 U43908 ( .A1(n47278), .A2(n30692), .ZN(n39165) );
  CLKNAND2HSV1 U43909 ( .A1(n52675), .A2(n39436), .ZN(n39164) );
  XOR2HSV0 U43910 ( .A1(n39165), .A2(n39164), .Z(n39170) );
  CLKNAND2HSV0 U43911 ( .A1(n51247), .A2(n30789), .ZN(n39168) );
  CLKNAND2HSV0 U43912 ( .A1(\pe5/aot [18]), .A2(n46933), .ZN(n39167) );
  XOR2HSV0 U43913 ( .A1(n39168), .A2(n39167), .Z(n39169) );
  XOR2HSV0 U43914 ( .A1(n39170), .A2(n39169), .Z(n39178) );
  NOR2HSV0 U43915 ( .A1(n50518), .A2(n45844), .ZN(n39172) );
  CLKNHSV0 U43916 ( .I(n30163), .ZN(n48663) );
  CLKNAND2HSV0 U43917 ( .A1(n48663), .A2(n48170), .ZN(n39171) );
  XOR2HSV0 U43918 ( .A1(n39172), .A2(n39171), .Z(n39176) );
  NAND2HSV0 U43919 ( .A1(n48658), .A2(n39449), .ZN(n39174) );
  CLKNHSV0 U43920 ( .I(n46978), .ZN(n52573) );
  NAND2HSV0 U43921 ( .A1(n52573), .A2(n30918), .ZN(n39173) );
  XOR2HSV0 U43922 ( .A1(n39174), .A2(n39173), .Z(n39175) );
  XOR2HSV0 U43923 ( .A1(n39176), .A2(n39175), .Z(n39177) );
  XOR2HSV0 U43924 ( .A1(n39178), .A2(n39177), .Z(n39179) );
  XOR2HSV0 U43925 ( .A1(n39180), .A2(n39179), .Z(n39182) );
  CLKNAND2HSV0 U43926 ( .A1(n48014), .A2(n52641), .ZN(n39181) );
  XNOR2HSV1 U43927 ( .A1(n39182), .A2(n39181), .ZN(n39183) );
  XNOR2HSV1 U43928 ( .A1(n39184), .A2(n39183), .ZN(n39185) );
  XOR2HSV0 U43929 ( .A1(n39186), .A2(n39185), .Z(n39187) );
  XNOR2HSV1 U43930 ( .A1(n39188), .A2(n39187), .ZN(n39191) );
  CLKNHSV0 U43931 ( .I(n45817), .ZN(n39655) );
  CLKNAND2HSV0 U43932 ( .A1(n39654), .A2(n39655), .ZN(n39190) );
  BUFHSV2 U43933 ( .I(n48848), .Z(n39954) );
  CLKNAND2HSV1 U43934 ( .A1(n39954), .A2(n39582), .ZN(n39189) );
  XOR3HSV2 U43935 ( .A1(n39191), .A2(n39190), .A3(n39189), .Z(n39192) );
  XNOR2HSV1 U43936 ( .A1(n39193), .A2(n39192), .ZN(n39194) );
  XNOR2HSV1 U43937 ( .A1(n39195), .A2(n39194), .ZN(n39196) );
  XOR2HSV0 U43938 ( .A1(n39197), .A2(n39196), .Z(n39198) );
  XNOR2HSV1 U43939 ( .A1(n39199), .A2(n39198), .ZN(n39200) );
  XOR2HSV0 U43940 ( .A1(n39201), .A2(n39200), .Z(n39202) );
  XNOR2HSV1 U43941 ( .A1(n39203), .A2(n39202), .ZN(n39205) );
  INHSV2 U43942 ( .I(n30516), .ZN(n51228) );
  CLKNAND2HSV0 U43943 ( .A1(n44694), .A2(n51228), .ZN(n39204) );
  XOR2HSV0 U43944 ( .A1(n39205), .A2(n39204), .Z(n39206) );
  XNOR2HSV1 U43945 ( .A1(n39207), .A2(n39206), .ZN(n39209) );
  BUFHSV2 U43946 ( .I(n39341), .Z(n51205) );
  NAND2HSV0 U43947 ( .A1(n51205), .A2(n30840), .ZN(n39208) );
  XNOR2HSV1 U43948 ( .A1(n39209), .A2(n39208), .ZN(n39210) );
  BUFHSV2 U43949 ( .I(n39542), .Z(n48746) );
  NAND2HSV2 U43950 ( .A1(n48746), .A2(n37630), .ZN(n39213) );
  INHSV3 U43951 ( .I(n39255), .ZN(n40116) );
  CLKNAND2HSV1 U43952 ( .A1(n40116), .A2(n48742), .ZN(n39212) );
  NOR2HSV0 U43953 ( .A1(n39215), .A2(n39222), .ZN(n39217) );
  NAND2HSV2 U43954 ( .A1(n39217), .A2(n39216), .ZN(n39221) );
  CLKNHSV1 U43955 ( .I(n39218), .ZN(n39219) );
  OAI21HSV2 U43956 ( .A1(n39221), .A2(n39223), .B(n39219), .ZN(n39220) );
  INHSV2 U43957 ( .I(n39220), .ZN(n39225) );
  NAND3HSV2 U43958 ( .A1(n39221), .A2(n39223), .A3(n40006), .ZN(n39224) );
  CLKNAND2HSV2 U43959 ( .A1(n39225), .A2(n39224), .ZN(n39356) );
  CLKNHSV2 U43960 ( .I(n39356), .ZN(n39226) );
  INHSV2 U43961 ( .I(n39416), .ZN(n39670) );
  NOR2HSV0 U43962 ( .A1(n39418), .A2(n40130), .ZN(n39229) );
  OAI21HSV1 U43963 ( .A1(n39416), .A2(n39230), .B(n39229), .ZN(n39233) );
  CLKNHSV0 U43964 ( .I(n40133), .ZN(n39683) );
  NOR2HSV0 U43965 ( .A1(n39354), .A2(n39683), .ZN(n39231) );
  CLKNAND2HSV1 U43966 ( .A1(n39364), .A2(n39231), .ZN(n39232) );
  CLKNAND2HSV1 U43967 ( .A1(n39233), .A2(n39232), .ZN(n39236) );
  CLKNHSV0 U43968 ( .I(n39413), .ZN(n39359) );
  MUX2NHSV1 U43969 ( .I0(n39359), .I1(n39234), .S(n39416), .ZN(n39235) );
  NAND2HSV2 U43970 ( .A1(n39236), .A2(n39235), .ZN(n39237) );
  XNOR2HSV4 U43971 ( .A1(n39238), .A2(n39237), .ZN(n39575) );
  NAND2HSV2 U43972 ( .A1(\pe5/ti_7t [23]), .A2(n39239), .ZN(n39742) );
  CLKNHSV1 U43973 ( .I(n39742), .ZN(n39688) );
  AOI21HSV1 U43974 ( .A1(n39742), .A2(n39241), .B(n39240), .ZN(n39242) );
  INHSV2 U43975 ( .I(n39575), .ZN(n39244) );
  INHSV1 U43976 ( .I(n39247), .ZN(n39248) );
  AOI22HSV4 U43977 ( .A1(n39249), .A2(n29722), .B1(n60025), .B2(n39248), .ZN(
        n39353) );
  CLKNHSV0 U43978 ( .I(n39251), .ZN(n39252) );
  INHSV2 U43979 ( .I(n39879), .ZN(n48164) );
  NOR2HSV2 U43980 ( .A1(n39255), .A2(n48164), .ZN(n39349) );
  NAND2HSV2 U43981 ( .A1(n39256), .A2(n48742), .ZN(n39345) );
  CLKNAND2HSV1 U43982 ( .A1(n45417), .A2(n45500), .ZN(n39340) );
  CLKNAND2HSV1 U43983 ( .A1(n39257), .A2(n39532), .ZN(n39336) );
  CLKNAND2HSV0 U43984 ( .A1(n45820), .A2(n37656), .ZN(n39334) );
  CLKNAND2HSV1 U43985 ( .A1(n48748), .A2(n45816), .ZN(n39332) );
  CLKNAND2HSV1 U43986 ( .A1(n40171), .A2(n39432), .ZN(n39330) );
  CLKNAND2HSV0 U43987 ( .A1(n40172), .A2(n39433), .ZN(n39328) );
  NAND2HSV0 U43988 ( .A1(n39258), .A2(n46974), .ZN(n39326) );
  CLKNAND2HSV1 U43989 ( .A1(n48168), .A2(n39259), .ZN(n39321) );
  CLKNAND2HSV0 U43990 ( .A1(n59639), .A2(n39655), .ZN(n39319) );
  CLKNAND2HSV0 U43991 ( .A1(\pe5/aot [23]), .A2(n39443), .ZN(n39261) );
  NAND2HSV0 U43992 ( .A1(n30788), .A2(n39445), .ZN(n39260) );
  XOR2HSV0 U43993 ( .A1(n39261), .A2(n39260), .Z(n39265) );
  NAND2HSV0 U43994 ( .A1(n59938), .A2(n52619), .ZN(n39262) );
  XOR2HSV0 U43995 ( .A1(n39263), .A2(n39262), .Z(n39264) );
  XOR2HSV0 U43996 ( .A1(n39265), .A2(n39264), .Z(n39281) );
  CLKNAND2HSV0 U43997 ( .A1(n39266), .A2(n39471), .ZN(n39268) );
  CLKNAND2HSV0 U43998 ( .A1(n39455), .A2(n48170), .ZN(n39267) );
  XOR2HSV0 U43999 ( .A1(n39268), .A2(n39267), .Z(n39273) );
  NAND2HSV0 U44000 ( .A1(n39269), .A2(n52610), .ZN(n39271) );
  CLKNHSV0 U44001 ( .I(n48175), .ZN(n39902) );
  NAND2HSV0 U44002 ( .A1(n39902), .A2(n39472), .ZN(n39270) );
  XOR2HSV0 U44003 ( .A1(n39271), .A2(n39270), .Z(n39272) );
  XOR2HSV0 U44004 ( .A1(n39273), .A2(n39272), .Z(n39277) );
  NAND2HSV0 U44005 ( .A1(n44335), .A2(\pe5/pvq [24]), .ZN(n39274) );
  XNOR2HSV1 U44006 ( .A1(n39274), .A2(\pe5/phq [24]), .ZN(n39275) );
  XNOR2HSV1 U44007 ( .A1(n39275), .A2(n40227), .ZN(n39276) );
  XNOR2HSV1 U44008 ( .A1(n39277), .A2(n39276), .ZN(n39280) );
  NAND2HSV0 U44009 ( .A1(n39278), .A2(n53289), .ZN(n39279) );
  XOR3HSV2 U44010 ( .A1(n39281), .A2(n39280), .A3(n39279), .Z(n39283) );
  NAND2HSV0 U44011 ( .A1(n39466), .A2(\pe5/got [12]), .ZN(n39282) );
  XNOR2HSV1 U44012 ( .A1(n39283), .A2(n39282), .ZN(n39317) );
  CLKNAND2HSV0 U44013 ( .A1(n39473), .A2(\pe5/bq[15] ), .ZN(n39285) );
  NAND2HSV0 U44014 ( .A1(n39616), .A2(n30692), .ZN(n39284) );
  XOR2HSV0 U44015 ( .A1(n39285), .A2(n39284), .Z(n39289) );
  NAND2HSV0 U44016 ( .A1(n50653), .A2(n52594), .ZN(n39287) );
  NAND2HSV0 U44017 ( .A1(\pe5/aot [16]), .A2(n52585), .ZN(n39286) );
  XOR2HSV0 U44018 ( .A1(n39287), .A2(n39286), .Z(n39288) );
  XOR2HSV0 U44019 ( .A1(n39289), .A2(n39288), .Z(n39297) );
  NOR2HSV1 U44020 ( .A1(n31029), .A2(n45844), .ZN(n39291) );
  NAND2HSV0 U44021 ( .A1(\pe5/aot [18]), .A2(n31160), .ZN(n39290) );
  XOR2HSV0 U44022 ( .A1(n39291), .A2(n39290), .Z(n39295) );
  CLKNAND2HSV0 U44023 ( .A1(n39499), .A2(n52595), .ZN(n39293) );
  NAND2HSV0 U44024 ( .A1(n39490), .A2(n39449), .ZN(n39292) );
  XOR2HSV0 U44025 ( .A1(n39293), .A2(n39292), .Z(n39294) );
  XOR2HSV0 U44026 ( .A1(n39295), .A2(n39294), .Z(n39296) );
  XOR2HSV0 U44027 ( .A1(n39297), .A2(n39296), .Z(n39313) );
  CLKNAND2HSV0 U44028 ( .A1(\pe5/aot [9]), .A2(n31192), .ZN(n39299) );
  NAND2HSV0 U44029 ( .A1(\pe5/got [9]), .A2(n37584), .ZN(n39298) );
  XOR2HSV0 U44030 ( .A1(n39299), .A2(n39298), .Z(n39303) );
  NAND2HSV0 U44031 ( .A1(n59427), .A2(\pe5/bq[11] ), .ZN(n39301) );
  NAND2HSV0 U44032 ( .A1(n48205), .A2(n39495), .ZN(n39300) );
  XOR2HSV0 U44033 ( .A1(n39301), .A2(n39300), .Z(n39302) );
  XOR2HSV0 U44034 ( .A1(n39303), .A2(n39302), .Z(n39311) );
  CLKNAND2HSV1 U44035 ( .A1(n51187), .A2(n39487), .ZN(n39305) );
  NAND2HSV0 U44036 ( .A1(\pe5/aot [13]), .A2(n45470), .ZN(n39304) );
  XOR2HSV0 U44037 ( .A1(n39305), .A2(n39304), .Z(n39309) );
  NAND2HSV0 U44038 ( .A1(n59896), .A2(n30230), .ZN(n39307) );
  NAND2HSV0 U44039 ( .A1(n59642), .A2(n39436), .ZN(n39306) );
  XOR2HSV0 U44040 ( .A1(n39307), .A2(n39306), .Z(n39308) );
  XOR2HSV0 U44041 ( .A1(n39309), .A2(n39308), .Z(n39310) );
  XOR2HSV0 U44042 ( .A1(n39311), .A2(n39310), .Z(n39312) );
  XOR2HSV0 U44043 ( .A1(n39313), .A2(n39312), .Z(n39315) );
  NAND2HSV0 U44044 ( .A1(n48014), .A2(n51305), .ZN(n39314) );
  XNOR2HSV1 U44045 ( .A1(n39315), .A2(n39314), .ZN(n39316) );
  XNOR2HSV1 U44046 ( .A1(n39317), .A2(n39316), .ZN(n39318) );
  XOR2HSV0 U44047 ( .A1(n39319), .A2(n39318), .Z(n39320) );
  XNOR2HSV1 U44048 ( .A1(n39321), .A2(n39320), .ZN(n39324) );
  CLKNAND2HSV1 U44049 ( .A1(n39654), .A2(n39516), .ZN(n39323) );
  CLKNAND2HSV0 U44050 ( .A1(n48848), .A2(n39434), .ZN(n39322) );
  XOR3HSV2 U44051 ( .A1(n39324), .A2(n39323), .A3(n39322), .Z(n39325) );
  XNOR2HSV1 U44052 ( .A1(n39326), .A2(n39325), .ZN(n39327) );
  XNOR2HSV1 U44053 ( .A1(n39328), .A2(n39327), .ZN(n39329) );
  XOR2HSV0 U44054 ( .A1(n39330), .A2(n39329), .Z(n39331) );
  XNOR2HSV1 U44055 ( .A1(n39332), .A2(n39331), .ZN(n39333) );
  XOR2HSV0 U44056 ( .A1(n39334), .A2(n39333), .Z(n39335) );
  CLKNAND2HSV0 U44057 ( .A1(n44694), .A2(n31148), .ZN(n39337) );
  XOR2HSV0 U44058 ( .A1(n39338), .A2(n39337), .Z(n39339) );
  CLKNAND2HSV0 U44059 ( .A1(n39341), .A2(n48739), .ZN(n39342) );
  XNOR2HSV4 U44060 ( .A1(n39345), .A2(n39344), .ZN(n39347) );
  NAND2HSV2 U44061 ( .A1(n39542), .A2(n30254), .ZN(n39346) );
  XOR2HSV2 U44062 ( .A1(n39347), .A2(n39346), .Z(n39348) );
  XNOR2HSV4 U44063 ( .A1(n39349), .A2(n39348), .ZN(n39350) );
  XNOR2HSV4 U44064 ( .A1(n39351), .A2(n39350), .ZN(n39352) );
  XNOR2HSV4 U44065 ( .A1(n39353), .A2(n39352), .ZN(n39377) );
  INHSV3 U44066 ( .I(n39377), .ZN(n39374) );
  INHSV2 U44067 ( .I(n39354), .ZN(n39414) );
  CLKNAND2HSV1 U44068 ( .A1(n39360), .A2(n39414), .ZN(n39358) );
  NOR3HSV2 U44069 ( .A1(n39367), .A2(n40009), .A3(n39356), .ZN(n39357) );
  CLKNAND2HSV2 U44070 ( .A1(n39362), .A2(n39361), .ZN(n39375) );
  AND2HSV2 U44071 ( .A1(n39365), .A2(n39414), .Z(n39363) );
  NAND2HSV0 U44072 ( .A1(n39368), .A2(n39413), .ZN(n39369) );
  INHSV2 U44073 ( .I(n39369), .ZN(n39371) );
  OR2HSV1 U44074 ( .A1(n39418), .A2(n40169), .Z(n39370) );
  AOI21HSV4 U44075 ( .A1(n39372), .A2(n39371), .B(n39370), .ZN(n39376) );
  CLKNAND2HSV2 U44076 ( .A1(n39375), .A2(n39376), .ZN(n39373) );
  CLKNAND2HSV3 U44077 ( .A1(n39374), .A2(n39373), .ZN(n39378) );
  NOR2HSV2 U44078 ( .A1(n51115), .A2(n39379), .ZN(n39380) );
  AND2HSV2 U44079 ( .A1(n39383), .A2(\pe5/ti_7t [24]), .Z(n39384) );
  AOI21HSV4 U44080 ( .A1(n29689), .A2(n59573), .B(n39384), .ZN(n39577) );
  INHSV2 U44081 ( .I(n39722), .ZN(n44329) );
  CLKNHSV2 U44082 ( .I(n39869), .ZN(n39386) );
  CLKNAND2HSV1 U44083 ( .A1(n40009), .A2(\pe5/ti_7t [26]), .ZN(n40143) );
  INHSV2 U44084 ( .I(n40143), .ZN(n39877) );
  NOR2HSV2 U44085 ( .A1(n39386), .A2(n39877), .ZN(n39573) );
  NAND2HSV4 U44086 ( .A1(n39577), .A2(n39576), .ZN(n39716) );
  INHSV4 U44087 ( .I(n39716), .ZN(n39554) );
  NOR2HSV4 U44088 ( .A1(n39554), .A2(n30421), .ZN(n39867) );
  CLKNHSV0 U44089 ( .I(n39867), .ZN(n39563) );
  OR2HSV2 U44090 ( .A1(n39570), .A2(n39877), .Z(n39562) );
  NAND3HSV2 U44091 ( .A1(n39677), .A2(n39390), .A3(n39389), .ZN(n39391) );
  CLKNHSV2 U44092 ( .I(n39401), .ZN(n39394) );
  NOR2HSV4 U44093 ( .A1(n39395), .A2(n39394), .ZN(n39396) );
  NAND2HSV0 U44094 ( .A1(n39399), .A2(n39398), .ZN(n39400) );
  CLKNHSV0 U44095 ( .I(n39400), .ZN(n39402) );
  CLKNAND2HSV0 U44096 ( .A1(n39402), .A2(n39678), .ZN(n39410) );
  NOR2HSV0 U44097 ( .A1(n39404), .A2(n47387), .ZN(n39407) );
  OAI21HSV0 U44098 ( .A1(n39405), .A2(\pe5/ti_7t [23]), .B(n52799), .ZN(n39406) );
  AOI31HSV2 U44099 ( .A1(n39677), .A2(n39408), .A3(n39407), .B(n39406), .ZN(
        n39409) );
  NAND3HSV2 U44100 ( .A1(n39681), .A2(n39718), .A3(n39680), .ZN(n39411) );
  CLKNHSV0 U44101 ( .I(n39418), .ZN(n39419) );
  AND2HSV2 U44102 ( .A1(n39419), .A2(n48885), .Z(n39420) );
  CLKNHSV0 U44103 ( .I(n39420), .ZN(n39422) );
  INAND2HSV2 U44104 ( .A1(n39669), .B1(n39420), .ZN(n39421) );
  CLKNAND2HSV2 U44105 ( .A1(n39670), .A2(n39671), .ZN(n47948) );
  NAND2HSV2 U44106 ( .A1(n39429), .A2(n39428), .ZN(n45416) );
  NAND2HSV2 U44107 ( .A1(n45416), .A2(n39430), .ZN(n39547) );
  NAND2HSV2 U44108 ( .A1(n51158), .A2(\pe5/got [25]), .ZN(n39541) );
  CLKNAND2HSV1 U44109 ( .A1(n45417), .A2(n30840), .ZN(n39536) );
  NAND2HSV2 U44110 ( .A1(n51019), .A2(n40170), .ZN(n39531) );
  CLKNAND2HSV0 U44111 ( .A1(n45820), .A2(n45816), .ZN(n39529) );
  NAND2HSV2 U44112 ( .A1(n48748), .A2(n39432), .ZN(n39527) );
  CLKNAND2HSV1 U44113 ( .A1(n59513), .A2(n39433), .ZN(n39525) );
  NAND2HSV0 U44114 ( .A1(n52578), .A2(n46974), .ZN(n39523) );
  NAND2HSV0 U44115 ( .A1(n39882), .A2(n39434), .ZN(n39521) );
  CLKNAND2HSV1 U44116 ( .A1(n48168), .A2(n39435), .ZN(n39515) );
  CLKNAND2HSV0 U44117 ( .A1(n39583), .A2(n48167), .ZN(n39513) );
  NAND2HSV0 U44118 ( .A1(n39616), .A2(n47305), .ZN(n39438) );
  NAND2HSV0 U44119 ( .A1(n39887), .A2(n39436), .ZN(n39437) );
  XOR2HSV0 U44120 ( .A1(n39438), .A2(n39437), .Z(n39442) );
  NAND2HSV0 U44121 ( .A1(n59896), .A2(n30357), .ZN(n39439) );
  XOR2HSV0 U44122 ( .A1(n39440), .A2(n39439), .Z(n39441) );
  XOR2HSV0 U44123 ( .A1(n39442), .A2(n39441), .Z(n39465) );
  CLKNAND2HSV1 U44124 ( .A1(n39278), .A2(n40257), .ZN(n39464) );
  NAND2HSV0 U44125 ( .A1(n39444), .A2(n39443), .ZN(n39448) );
  NAND2HSV0 U44126 ( .A1(n39446), .A2(n39445), .ZN(n39447) );
  XOR2HSV0 U44127 ( .A1(n39448), .A2(n39447), .Z(n39453) );
  CLKNAND2HSV0 U44128 ( .A1(\pe5/got [8]), .A2(n30693), .ZN(n39451) );
  NAND2HSV0 U44129 ( .A1(\pe5/aot [13]), .A2(n39449), .ZN(n39450) );
  XOR2HSV0 U44130 ( .A1(n39451), .A2(n39450), .Z(n39452) );
  XOR2HSV0 U44131 ( .A1(n39453), .A2(n39452), .Z(n39462) );
  CLKNAND2HSV0 U44132 ( .A1(n51187), .A2(n39454), .ZN(n39457) );
  CLKNAND2HSV0 U44133 ( .A1(n39455), .A2(n50533), .ZN(n39456) );
  XOR2HSV0 U44134 ( .A1(n39457), .A2(n39456), .Z(n39460) );
  NAND2HSV0 U44135 ( .A1(n48039), .A2(\pe5/pvq [25]), .ZN(n39458) );
  XOR2HSV0 U44136 ( .A1(n39458), .A2(\pe5/phq [25]), .Z(n39459) );
  XOR2HSV0 U44137 ( .A1(n39460), .A2(n39459), .Z(n39461) );
  XOR2HSV0 U44138 ( .A1(n39462), .A2(n39461), .Z(n39463) );
  XOR3HSV2 U44139 ( .A1(n39465), .A2(n39464), .A3(n39463), .Z(n39468) );
  CLKNAND2HSV0 U44140 ( .A1(n39466), .A2(n48749), .ZN(n39467) );
  XNOR2HSV1 U44141 ( .A1(n39468), .A2(n39467), .ZN(n39511) );
  CLKNAND2HSV1 U44142 ( .A1(n50511), .A2(n30789), .ZN(n39470) );
  CLKNAND2HSV1 U44143 ( .A1(n48634), .A2(n39914), .ZN(n39469) );
  XOR2HSV0 U44144 ( .A1(n39470), .A2(n39469), .Z(n39477) );
  CLKNAND2HSV1 U44145 ( .A1(n39902), .A2(n39471), .ZN(n39475) );
  NAND2HSV0 U44146 ( .A1(n39473), .A2(n39472), .ZN(n39474) );
  XOR2HSV0 U44147 ( .A1(n39475), .A2(n39474), .Z(n39476) );
  XOR2HSV0 U44148 ( .A1(n39477), .A2(n39476), .Z(n39486) );
  CLKNAND2HSV1 U44149 ( .A1(n59640), .A2(n30891), .ZN(n39479) );
  NAND2HSV0 U44150 ( .A1(n50653), .A2(n46622), .ZN(n39478) );
  XOR2HSV0 U44151 ( .A1(n39479), .A2(n39478), .Z(n39484) );
  CLKNAND2HSV0 U44152 ( .A1(\pe5/aot [18]), .A2(n39480), .ZN(n39482) );
  NAND2HSV0 U44153 ( .A1(n39629), .A2(n48170), .ZN(n39481) );
  XOR2HSV0 U44154 ( .A1(n39482), .A2(n39481), .Z(n39483) );
  XOR2HSV0 U44155 ( .A1(n39484), .A2(n39483), .Z(n39485) );
  XOR2HSV0 U44156 ( .A1(n39486), .A2(n39485), .Z(n39507) );
  NAND2HSV0 U44157 ( .A1(n52591), .A2(n39487), .ZN(n39489) );
  CLKNAND2HSV0 U44158 ( .A1(n48663), .A2(n39592), .ZN(n39488) );
  XOR2HSV0 U44159 ( .A1(n39489), .A2(n39488), .Z(n39494) );
  CLKNAND2HSV0 U44160 ( .A1(n39490), .A2(n30222), .ZN(n39492) );
  NAND2HSV0 U44161 ( .A1(n48205), .A2(n39130), .ZN(n39491) );
  XOR2HSV0 U44162 ( .A1(n39492), .A2(n39491), .Z(n39493) );
  XOR2HSV0 U44163 ( .A1(n39494), .A2(n39493), .Z(n39505) );
  NAND2HSV0 U44164 ( .A1(n59642), .A2(n39495), .ZN(n39498) );
  NAND2HSV0 U44165 ( .A1(n39496), .A2(\pe5/bq[8] ), .ZN(n39497) );
  XOR2HSV0 U44166 ( .A1(n39498), .A2(n39497), .Z(n39503) );
  CLKNAND2HSV1 U44167 ( .A1(n40234), .A2(n39615), .ZN(n39501) );
  CLKNAND2HSV1 U44168 ( .A1(n39499), .A2(n52610), .ZN(n39500) );
  XOR2HSV0 U44169 ( .A1(n39501), .A2(n39500), .Z(n39502) );
  XOR2HSV0 U44170 ( .A1(n39503), .A2(n39502), .Z(n39504) );
  XOR2HSV0 U44171 ( .A1(n39505), .A2(n39504), .Z(n39506) );
  XOR2HSV0 U44172 ( .A1(n39507), .A2(n39506), .Z(n39509) );
  CLKNAND2HSV1 U44173 ( .A1(n48014), .A2(n51210), .ZN(n39508) );
  XNOR2HSV1 U44174 ( .A1(n39509), .A2(n39508), .ZN(n39510) );
  XNOR2HSV1 U44175 ( .A1(n39511), .A2(n39510), .ZN(n39512) );
  XNOR2HSV1 U44176 ( .A1(n39513), .A2(n39512), .ZN(n39514) );
  XNOR2HSV1 U44177 ( .A1(n39515), .A2(n39514), .ZN(n39519) );
  CLKNAND2HSV1 U44178 ( .A1(n39654), .A2(n39582), .ZN(n39518) );
  NAND2HSV2 U44179 ( .A1(n39954), .A2(n39516), .ZN(n39517) );
  XOR3HSV2 U44180 ( .A1(n39519), .A2(n39518), .A3(n39517), .Z(n39520) );
  XNOR2HSV1 U44181 ( .A1(n39521), .A2(n39520), .ZN(n39522) );
  XNOR2HSV1 U44182 ( .A1(n39523), .A2(n39522), .ZN(n39524) );
  XOR2HSV0 U44183 ( .A1(n39525), .A2(n39524), .Z(n39526) );
  XOR2HSV0 U44184 ( .A1(n39527), .A2(n39526), .Z(n39528) );
  XOR2HSV0 U44185 ( .A1(n39529), .A2(n39528), .Z(n39530) );
  XNOR2HSV1 U44186 ( .A1(n39531), .A2(n39530), .ZN(n39534) );
  CLKNAND2HSV1 U44187 ( .A1(n44694), .A2(n39532), .ZN(n39533) );
  XOR2HSV0 U44188 ( .A1(n39534), .A2(n39533), .Z(n39535) );
  XNOR2HSV1 U44189 ( .A1(n39536), .A2(n39535), .ZN(n39539) );
  NAND2HSV0 U44190 ( .A1(n39537), .A2(n45500), .ZN(n39538) );
  XNOR2HSV1 U44191 ( .A1(n39539), .A2(n39538), .ZN(n39540) );
  XNOR2HSV1 U44192 ( .A1(n39541), .A2(n39540), .ZN(n39545) );
  CLKNAND2HSV1 U44193 ( .A1(n48746), .A2(n48742), .ZN(n39544) );
  NAND2HSV2 U44194 ( .A1(n40116), .A2(n31225), .ZN(n39543) );
  XOR3HSV2 U44195 ( .A1(n39545), .A2(n39544), .A3(n39543), .Z(n39546) );
  XNOR2HSV1 U44196 ( .A1(n39547), .A2(n39546), .ZN(n39552) );
  CLKNHSV2 U44197 ( .I(n39549), .ZN(n39550) );
  OAI21HSV1 U44198 ( .A1(n60025), .A2(n29722), .B(n39550), .ZN(n39551) );
  XNOR2HSV1 U44199 ( .A1(n39552), .A2(n39551), .ZN(n39556) );
  XNOR2HSV4 U44200 ( .A1(n39557), .A2(n39556), .ZN(n39725) );
  NOR2HSV4 U44201 ( .A1(n39725), .A2(n39239), .ZN(n39553) );
  INHSV2 U44202 ( .I(n39569), .ZN(n39581) );
  NOR2HSV2 U44203 ( .A1(n39705), .A2(\pe5/ti_7t [25]), .ZN(n39996) );
  NOR2HSV0 U44204 ( .A1(n39996), .A2(n39733), .ZN(n39567) );
  CLKNHSV0 U44205 ( .I(n39567), .ZN(n39555) );
  NOR2HSV0 U44206 ( .A1(n39877), .A2(n39555), .ZN(n39559) );
  AND2HSV2 U44207 ( .A1(n39559), .A2(n39568), .Z(n39560) );
  NAND2HSV2 U44208 ( .A1(n39581), .A2(n39560), .ZN(n39561) );
  OAI21HSV4 U44209 ( .A1(n39563), .A2(n39562), .B(n39561), .ZN(n39572) );
  INHSV2 U44210 ( .I(n39379), .ZN(n45414) );
  OAI21HSV2 U44211 ( .A1(n39570), .A2(n59946), .B(n45414), .ZN(n39564) );
  INHSV2 U44212 ( .I(n39564), .ZN(n39566) );
  NAND2HSV4 U44213 ( .A1(n39566), .A2(n39565), .ZN(n40139) );
  CLKNAND2HSV4 U44214 ( .A1(n39867), .A2(n26683), .ZN(n40141) );
  CLKNAND2HSV1 U44215 ( .A1(n40138), .A2(n40141), .ZN(n39571) );
  OAI22HSV4 U44216 ( .A1(n39573), .A2(n39572), .B1(n40139), .B2(n39571), .ZN(
        n47041) );
  BUFHSV2 U44217 ( .I(n47041), .Z(n59535) );
  INHSV2 U44218 ( .I(n39874), .ZN(n39580) );
  CLKNAND2HSV0 U44219 ( .A1(n39576), .A2(n39577), .ZN(n39579) );
  BUFHSV2 U44220 ( .I(n51158), .Z(n59882) );
  INHSV2 U44221 ( .I(\pe5/got [18]), .ZN(n46583) );
  CLKNAND2HSV1 U44222 ( .A1(n40171), .A2(n39881), .ZN(n39663) );
  INHSV2 U44223 ( .I(n48722), .ZN(n51157) );
  NAND2HSV0 U44224 ( .A1(n48624), .A2(n51157), .ZN(n39662) );
  NAND2HSV0 U44225 ( .A1(n39882), .A2(n39582), .ZN(n39660) );
  CLKNHSV0 U44226 ( .I(n47143), .ZN(n48749) );
  NAND2HSV2 U44227 ( .A1(n48168), .A2(n48749), .ZN(n39653) );
  BUFHSV2 U44228 ( .I(n39583), .Z(n48169) );
  CLKNAND2HSV1 U44229 ( .A1(n48169), .A2(n51210), .ZN(n39651) );
  CLKNAND2HSV0 U44230 ( .A1(n37707), .A2(\pe5/pvq [27]), .ZN(n39584) );
  XOR2HSV0 U44231 ( .A1(n39584), .A2(\pe5/phq [27]), .Z(n39588) );
  CLKNAND2HSV0 U44232 ( .A1(\pe5/aot [23]), .A2(n51191), .ZN(n47323) );
  OAI22HSV0 U44233 ( .A1(n31044), .A2(n46136), .B1(n40043), .B2(n51057), .ZN(
        n39585) );
  OAI21HSV0 U44234 ( .A1(n39586), .A2(n47323), .B(n39585), .ZN(n39587) );
  XNOR2HSV1 U44235 ( .A1(n39588), .A2(n39587), .ZN(n39591) );
  NAND2HSV0 U44236 ( .A1(n39887), .A2(n48755), .ZN(n45462) );
  XOR2HSV0 U44237 ( .A1(n39589), .A2(n45462), .Z(n39590) );
  XNOR2HSV1 U44238 ( .A1(n39591), .A2(n39590), .ZN(n39610) );
  CLKNHSV0 U44239 ( .I(n46978), .ZN(n51359) );
  NAND2HSV0 U44240 ( .A1(n30377), .A2(n51359), .ZN(n39609) );
  NAND2HSV0 U44241 ( .A1(n48829), .A2(n39592), .ZN(n39594) );
  BUFHSV2 U44242 ( .I(\pe5/aot [6]), .Z(n52682) );
  NAND2HSV0 U44243 ( .A1(n52682), .A2(n31192), .ZN(n39593) );
  XOR2HSV0 U44244 ( .A1(n39594), .A2(n39593), .Z(n39598) );
  NAND2HSV0 U44245 ( .A1(n39490), .A2(n30341), .ZN(n39596) );
  INHSV2 U44246 ( .I(n47230), .ZN(n53304) );
  CLKNAND2HSV0 U44247 ( .A1(n53304), .A2(n30698), .ZN(n39595) );
  XOR2HSV0 U44248 ( .A1(n39596), .A2(n39595), .Z(n39597) );
  XOR2HSV0 U44249 ( .A1(n39598), .A2(n39597), .Z(n39607) );
  NOR2HSV0 U44250 ( .A1(n31029), .A2(n46134), .ZN(n39600) );
  CLKNAND2HSV1 U44251 ( .A1(n51187), .A2(n48236), .ZN(n39599) );
  XOR2HSV0 U44252 ( .A1(n39600), .A2(n39599), .Z(n39605) );
  NAND2HSV0 U44253 ( .A1(n39601), .A2(\pe5/bq[7] ), .ZN(n39603) );
  NAND2HSV0 U44254 ( .A1(n48658), .A2(n30222), .ZN(n39602) );
  XOR2HSV0 U44255 ( .A1(n39603), .A2(n39602), .Z(n39604) );
  XOR2HSV0 U44256 ( .A1(n39605), .A2(n39604), .Z(n39606) );
  XOR2HSV0 U44257 ( .A1(n39607), .A2(n39606), .Z(n39608) );
  XOR3HSV2 U44258 ( .A1(n39610), .A2(n39609), .A3(n39608), .Z(n39612) );
  CLKNAND2HSV1 U44259 ( .A1(n48751), .A2(n40257), .ZN(n39611) );
  XNOR2HSV1 U44260 ( .A1(n39612), .A2(n39611), .ZN(n39649) );
  NAND2HSV0 U44261 ( .A1(\pe5/aot [18]), .A2(n51048), .ZN(n39614) );
  CLKNAND2HSV0 U44262 ( .A1(n30788), .A2(n39921), .ZN(n39613) );
  XOR2HSV0 U44263 ( .A1(n39614), .A2(n39613), .Z(n39620) );
  CLKNAND2HSV1 U44264 ( .A1(n31175), .A2(n39615), .ZN(n39618) );
  NAND2HSV0 U44265 ( .A1(n39616), .A2(n46933), .ZN(n39617) );
  XOR2HSV0 U44266 ( .A1(n39618), .A2(n39617), .Z(n39619) );
  XOR2HSV0 U44267 ( .A1(n39620), .A2(n39619), .Z(n39628) );
  CLKNAND2HSV0 U44268 ( .A1(n48663), .A2(n50533), .ZN(n39622) );
  NAND2HSV0 U44269 ( .A1(\pe5/got [6]), .A2(n37584), .ZN(n39621) );
  XOR2HSV0 U44270 ( .A1(n39622), .A2(n39621), .Z(n39626) );
  CLKNAND2HSV1 U44271 ( .A1(\pe5/aot [16]), .A2(n47059), .ZN(n39624) );
  NAND2HSV0 U44272 ( .A1(n48205), .A2(n30256), .ZN(n39623) );
  XOR2HSV0 U44273 ( .A1(n39624), .A2(n39623), .Z(n39625) );
  XOR2HSV0 U44274 ( .A1(n39626), .A2(n39625), .Z(n39627) );
  XOR2HSV0 U44275 ( .A1(n39628), .A2(n39627), .Z(n39645) );
  NAND2HSV0 U44276 ( .A1(n59642), .A2(n48802), .ZN(n39631) );
  NAND2HSV0 U44277 ( .A1(n39629), .A2(n48760), .ZN(n39630) );
  XOR2HSV0 U44278 ( .A1(n39631), .A2(n39630), .Z(n39635) );
  NAND2HSV0 U44279 ( .A1(n50511), .A2(n40074), .ZN(n39633) );
  NAND2HSV0 U44280 ( .A1(n40234), .A2(n48170), .ZN(n39632) );
  XOR2HSV0 U44281 ( .A1(n39633), .A2(n39632), .Z(n39634) );
  XOR2HSV0 U44282 ( .A1(n39635), .A2(n39634), .Z(n39643) );
  NOR2HSV0 U44283 ( .A1(n30150), .A2(n48050), .ZN(n39637) );
  NAND2HSV0 U44284 ( .A1(n39499), .A2(n40221), .ZN(n39636) );
  XOR2HSV0 U44285 ( .A1(n39637), .A2(n39636), .Z(n39641) );
  NAND2HSV0 U44286 ( .A1(\pe5/aot [13]), .A2(n46622), .ZN(n39639) );
  NAND2HSV0 U44287 ( .A1(n47278), .A2(n30607), .ZN(n39638) );
  XOR2HSV0 U44288 ( .A1(n39639), .A2(n39638), .Z(n39640) );
  XOR2HSV0 U44289 ( .A1(n39641), .A2(n39640), .Z(n39642) );
  XOR2HSV0 U44290 ( .A1(n39643), .A2(n39642), .Z(n39644) );
  XOR2HSV0 U44291 ( .A1(n39645), .A2(n39644), .Z(n39647) );
  CLKNAND2HSV0 U44292 ( .A1(n30785), .A2(\pe5/got [8]), .ZN(n39646) );
  XNOR2HSV1 U44293 ( .A1(n39647), .A2(n39646), .ZN(n39648) );
  XNOR2HSV1 U44294 ( .A1(n39649), .A2(n39648), .ZN(n39650) );
  XOR2HSV0 U44295 ( .A1(n39651), .A2(n39650), .Z(n39652) );
  XNOR2HSV1 U44296 ( .A1(n39653), .A2(n39652), .ZN(n39658) );
  CLKNAND2HSV0 U44297 ( .A1(n39654), .A2(n48167), .ZN(n39657) );
  CLKNAND2HSV1 U44298 ( .A1(n39954), .A2(n39655), .ZN(n39656) );
  XOR3HSV2 U44299 ( .A1(n39658), .A2(n39657), .A3(n39656), .Z(n39659) );
  XNOR2HSV1 U44300 ( .A1(n39660), .A2(n39659), .ZN(n39661) );
  CLKNHSV0 U44301 ( .I(n39664), .ZN(n59517) );
  XNOR2HSV4 U44302 ( .A1(n39668), .A2(n39667), .ZN(n39674) );
  CLKNHSV0 U44303 ( .I(n44520), .ZN(n47387) );
  NAND2HSV2 U44304 ( .A1(n45489), .A2(n39879), .ZN(n39673) );
  NAND3HSV2 U44305 ( .A1(n29706), .A2(n40133), .A3(n39679), .ZN(n39691) );
  CLKNHSV0 U44306 ( .I(n39680), .ZN(n39685) );
  NAND2HSV0 U44307 ( .A1(n39681), .A2(n39682), .ZN(n39684) );
  NOR3HSV2 U44308 ( .A1(n39685), .A2(n39684), .A3(n39683), .ZN(n39687) );
  CLKNAND2HSV1 U44309 ( .A1(n39687), .A2(n39686), .ZN(n39690) );
  CLKNAND2HSV1 U44310 ( .A1(n39688), .A2(n30142), .ZN(n39689) );
  NAND2HSV2 U44311 ( .A1(n25904), .A2(n39693), .ZN(n39694) );
  CLKNHSV2 U44312 ( .I(n39694), .ZN(n39695) );
  OR2HSV1 U44313 ( .A1(n39733), .A2(n39702), .Z(n39703) );
  NOR2HSV4 U44314 ( .A1(n39732), .A2(n39703), .ZN(n39710) );
  NAND2HSV2 U44315 ( .A1(n25904), .A2(n31133), .ZN(n39708) );
  OAI21HSV0 U44316 ( .A1(\pe5/ti_7t [27]), .A2(n39705), .B(n39704), .ZN(n39706) );
  INHSV2 U44317 ( .I(n39706), .ZN(n39707) );
  NAND2HSV2 U44318 ( .A1(n39708), .A2(n39707), .ZN(n39709) );
  AOI21HSV4 U44319 ( .A1(n59423), .A2(n39710), .B(n39709), .ZN(n39711) );
  NOR2HSV0 U44320 ( .A1(n39725), .A2(n47927), .ZN(n39723) );
  NOR2HSV2 U44321 ( .A1(n39724), .A2(n39723), .ZN(n39729) );
  CLKNHSV0 U44322 ( .I(n39726), .ZN(n39727) );
  NAND2HSV2 U44323 ( .A1(n39717), .A2(n39727), .ZN(n39728) );
  NAND2HSV2 U44324 ( .A1(\pe5/ti_7t [25]), .A2(n39730), .ZN(n40131) );
  NAND2HSV2 U44325 ( .A1(n40290), .A2(n30046), .ZN(n39865) );
  INAND2HSV2 U44326 ( .A1(n30431), .B1(n45415), .ZN(n39864) );
  BUFHSV2 U44327 ( .I(n39880), .Z(n48165) );
  NAND2HSV2 U44328 ( .A1(n48165), .A2(\pe5/got [25]), .ZN(n39859) );
  BUFHSV2 U44329 ( .I(n45489), .Z(n59926) );
  INHSV2 U44330 ( .I(n59926), .ZN(n50692) );
  NOR2HSV2 U44331 ( .A1(n50692), .A2(n40020), .ZN(n39857) );
  CLKNHSV2 U44332 ( .I(n40278), .ZN(n47145) );
  BUFHSV2 U44333 ( .I(n47145), .Z(n51217) );
  NAND2HSV2 U44334 ( .A1(n48745), .A2(\pe5/got [23]), .ZN(n39855) );
  NOR2HSV2 U44335 ( .A1(n48166), .A2(n47140), .ZN(n39853) );
  NAND2HSV2 U44336 ( .A1(n52570), .A2(n51103), .ZN(n39848) );
  INHSV1 U44337 ( .I(n50422), .ZN(n51156) );
  CLKNAND2HSV0 U44338 ( .A1(n52572), .A2(n51156), .ZN(n39844) );
  INHSV2 U44339 ( .I(n48722), .ZN(n51015) );
  NAND2HSV0 U44340 ( .A1(n51160), .A2(n51015), .ZN(n39839) );
  BUFHSV2 U44341 ( .I(n39744), .Z(n59392) );
  CLKNHSV0 U44342 ( .I(n31199), .ZN(n52652) );
  NAND2HSV0 U44343 ( .A1(n52574), .A2(n52652), .ZN(n39837) );
  CLKNHSV0 U44344 ( .I(n45817), .ZN(n52568) );
  NAND2HSV0 U44345 ( .A1(n59871), .A2(n52568), .ZN(n39835) );
  CLKNAND2HSV1 U44346 ( .A1(n39745), .A2(n48167), .ZN(n39833) );
  NAND2HSV0 U44347 ( .A1(n48624), .A2(n48749), .ZN(n39831) );
  BUFHSV2 U44348 ( .I(n59381), .Z(n52580) );
  NAND2HSV0 U44349 ( .A1(n52580), .A2(n51210), .ZN(n39829) );
  NAND2HSV0 U44350 ( .A1(n37558), .A2(n51359), .ZN(n39823) );
  NAND2HSV0 U44351 ( .A1(n48751), .A2(n48841), .ZN(n39819) );
  INHSV2 U44352 ( .I(n50507), .ZN(n52584) );
  NAND2HSV0 U44353 ( .A1(n52584), .A2(n47059), .ZN(n39747) );
  INHSV2 U44354 ( .I(n48204), .ZN(n52611) );
  NAND2HSV0 U44355 ( .A1(n52611), .A2(n47305), .ZN(n39746) );
  XOR2HSV0 U44356 ( .A1(n39747), .A2(n39746), .Z(n39751) );
  CLKNHSV0 U44357 ( .I(n51021), .ZN(n48686) );
  NAND2HSV0 U44358 ( .A1(n48663), .A2(n48686), .ZN(n39749) );
  NAND2HSV0 U44359 ( .A1(\pe5/aot [6]), .A2(n48802), .ZN(n39748) );
  XOR2HSV0 U44360 ( .A1(n39749), .A2(n39748), .Z(n39750) );
  XOR2HSV0 U44361 ( .A1(n39751), .A2(n39750), .Z(n39759) );
  NAND2HSV0 U44362 ( .A1(n51313), .A2(n30891), .ZN(n39753) );
  NAND2HSV0 U44363 ( .A1(n40190), .A2(n50500), .ZN(n39752) );
  XOR2HSV0 U44364 ( .A1(n39753), .A2(n39752), .Z(n39757) );
  NAND2HSV2 U44365 ( .A1(\pe5/aot [13]), .A2(n39445), .ZN(n39755) );
  NAND2HSV0 U44366 ( .A1(n59944), .A2(n48787), .ZN(n39754) );
  XOR2HSV0 U44367 ( .A1(n39755), .A2(n39754), .Z(n39756) );
  XOR2HSV0 U44368 ( .A1(n39757), .A2(n39756), .Z(n39758) );
  XOR2HSV0 U44369 ( .A1(n39759), .A2(n39758), .Z(n39761) );
  INHSV2 U44370 ( .I(n51231), .ZN(n59355) );
  NAND2HSV0 U44371 ( .A1(n30377), .A2(n59355), .ZN(n39760) );
  XNOR2HSV1 U44372 ( .A1(n39761), .A2(n39760), .ZN(n39763) );
  NAND2HSV0 U44373 ( .A1(n30270), .A2(n51302), .ZN(n39762) );
  XNOR2HSV1 U44374 ( .A1(n39763), .A2(n39762), .ZN(n39818) );
  NAND2HSV0 U44375 ( .A1(\pe5/aot [23]), .A2(\pe5/bq[11] ), .ZN(n39765) );
  NAND2HSV0 U44376 ( .A1(\pe5/aot [4]), .A2(n48198), .ZN(n39764) );
  XOR2HSV0 U44377 ( .A1(n39765), .A2(n39764), .Z(n39769) );
  NAND2HSV0 U44378 ( .A1(n40210), .A2(n48236), .ZN(n39767) );
  CLKNHSV0 U44379 ( .I(n45451), .ZN(n48171) );
  NAND2HSV0 U44380 ( .A1(n48171), .A2(n31045), .ZN(n39766) );
  XOR2HSV0 U44381 ( .A1(n39767), .A2(n39766), .Z(n39768) );
  XOR2HSV0 U44382 ( .A1(n39769), .A2(n39768), .Z(n39778) );
  NAND2HSV0 U44383 ( .A1(n39473), .A2(n48760), .ZN(n39771) );
  NAND2HSV0 U44384 ( .A1(n52600), .A2(n30698), .ZN(n39770) );
  XOR2HSV0 U44385 ( .A1(n39771), .A2(n39770), .Z(n39776) );
  CLKNHSV0 U44386 ( .I(n30150), .ZN(n48761) );
  NAND2HSV0 U44387 ( .A1(n48761), .A2(n48775), .ZN(n39774) );
  NAND2HSV0 U44388 ( .A1(n59880), .A2(n30222), .ZN(n39773) );
  XOR2HSV0 U44389 ( .A1(n39774), .A2(n39773), .Z(n39775) );
  XOR2HSV0 U44390 ( .A1(n39776), .A2(n39775), .Z(n39777) );
  XOR2HSV0 U44391 ( .A1(n39778), .A2(n39777), .Z(n39793) );
  INHSV2 U44392 ( .I(\pe5/got [2]), .ZN(n51306) );
  INHSV2 U44393 ( .I(n51306), .ZN(n59357) );
  NAND2HSV0 U44394 ( .A1(n59357), .A2(n30918), .ZN(n39781) );
  CLKNHSV0 U44395 ( .I(n39779), .ZN(n48172) );
  CLKNHSV0 U44396 ( .I(n48031), .ZN(n40226) );
  NAND2HSV0 U44397 ( .A1(n48172), .A2(n40226), .ZN(n39780) );
  XOR2HSV0 U44398 ( .A1(n39781), .A2(n39780), .Z(n39785) );
  CLKNHSV0 U44399 ( .I(n48822), .ZN(n51167) );
  NAND2HSV2 U44400 ( .A1(\pe5/aot [16]), .A2(n51167), .ZN(n39783) );
  CLKNHSV0 U44401 ( .I(n44704), .ZN(n48243) );
  BUFHSV2 U44402 ( .I(\pe5/bq[10] ), .Z(n53216) );
  NAND2HSV0 U44403 ( .A1(n48243), .A2(n53216), .ZN(n39782) );
  XOR2HSV0 U44404 ( .A1(n39783), .A2(n39782), .Z(n39784) );
  XOR2HSV0 U44405 ( .A1(n39785), .A2(n39784), .Z(n39791) );
  NAND2HSV0 U44406 ( .A1(n46628), .A2(\pe5/pvq [31]), .ZN(n39786) );
  XOR2HSV0 U44407 ( .A1(n39786), .A2(\pe5/phq [31]), .Z(n39789) );
  NAND2HSV0 U44408 ( .A1(n48681), .A2(\pe5/bq[19] ), .ZN(n48827) );
  INHSV2 U44409 ( .I(n48823), .ZN(n50505) );
  NAND2HSV2 U44410 ( .A1(n50505), .A2(n48237), .ZN(n40232) );
  OAI22HSV0 U44411 ( .A1(n46134), .A2(n48823), .B1(n59641), .B2(n45426), .ZN(
        n39787) );
  OAI21HSV0 U44412 ( .A1(n48827), .A2(n40232), .B(n39787), .ZN(n39788) );
  XOR2HSV0 U44413 ( .A1(n39789), .A2(n39788), .Z(n39790) );
  XNOR2HSV1 U44414 ( .A1(n39791), .A2(n39790), .ZN(n39792) );
  XNOR2HSV1 U44415 ( .A1(n39793), .A2(n39792), .ZN(n39816) );
  BUFHSV2 U44416 ( .I(\pe5/aot [21]), .Z(n48242) );
  NAND2HSV0 U44417 ( .A1(n48242), .A2(n50668), .ZN(n39795) );
  NAND2HSV0 U44418 ( .A1(n52591), .A2(n40221), .ZN(n39794) );
  XOR2HSV0 U44419 ( .A1(n39795), .A2(n39794), .Z(n39814) );
  CLKNHSV0 U44420 ( .I(n51232), .ZN(n51419) );
  NAND2HSV0 U44421 ( .A1(n51419), .A2(n48181), .ZN(n50585) );
  OAI22HSV0 U44422 ( .A1(n39166), .A2(n51232), .B1(n45858), .B2(n39796), .ZN(
        n39798) );
  OAI21HSV0 U44423 ( .A1(n39799), .A2(n50585), .B(n39798), .ZN(n39805) );
  NAND2HSV0 U44424 ( .A1(n39902), .A2(\pe5/bq[2] ), .ZN(n47322) );
  NOR2HSV0 U44425 ( .A1(n39800), .A2(n47322), .ZN(n39803) );
  AOI22HSV0 U44426 ( .A1(n59366), .A2(\pe5/bq[2] ), .B1(n39801), .B2(
        \pe5/bq[7] ), .ZN(n39802) );
  NOR2HSV2 U44427 ( .A1(n39803), .A2(n39802), .ZN(n39804) );
  XNOR2HSV1 U44428 ( .A1(n39805), .A2(n39804), .ZN(n39813) );
  NAND2HSV0 U44429 ( .A1(\pe5/aot [9]), .A2(n46622), .ZN(n39807) );
  NAND2HSV0 U44430 ( .A1(n39266), .A2(n50526), .ZN(n39806) );
  XOR2HSV0 U44431 ( .A1(n39807), .A2(n39806), .Z(n39811) );
  CLKNHSV0 U44432 ( .I(n47409), .ZN(n51363) );
  NAND2HSV0 U44433 ( .A1(n51363), .A2(n30230), .ZN(n39809) );
  NAND2HSV0 U44434 ( .A1(n59427), .A2(\pe5/bq[4] ), .ZN(n39808) );
  XOR2HSV0 U44435 ( .A1(n39809), .A2(n39808), .Z(n39810) );
  XOR2HSV0 U44436 ( .A1(n39811), .A2(n39810), .Z(n39812) );
  XOR3HSV2 U44437 ( .A1(n39814), .A2(n39813), .A3(n39812), .Z(n39815) );
  XNOR2HSV1 U44438 ( .A1(n39816), .A2(n39815), .ZN(n39817) );
  XOR3HSV2 U44439 ( .A1(n39819), .A2(n39818), .A3(n39817), .Z(n39821) );
  NAND2HSV0 U44440 ( .A1(n48169), .A2(\pe5/got [6]), .ZN(n39820) );
  XOR2HSV0 U44441 ( .A1(n39821), .A2(n39820), .Z(n39822) );
  XNOR2HSV1 U44442 ( .A1(n39823), .A2(n39822), .ZN(n39827) );
  INHSV2 U44443 ( .I(n44332), .ZN(n48750) );
  NAND2HSV0 U44444 ( .A1(n48750), .A2(n50698), .ZN(n39826) );
  NAND2HSV0 U44445 ( .A1(n39954), .A2(n40257), .ZN(n39825) );
  XOR3HSV2 U44446 ( .A1(n39827), .A2(n39826), .A3(n39825), .Z(n39828) );
  XNOR2HSV1 U44447 ( .A1(n39829), .A2(n39828), .ZN(n39830) );
  XNOR2HSV1 U44448 ( .A1(n39831), .A2(n39830), .ZN(n39832) );
  XOR2HSV0 U44449 ( .A1(n39833), .A2(n39832), .Z(n39834) );
  XNOR2HSV1 U44450 ( .A1(n39835), .A2(n39834), .ZN(n39836) );
  XOR2HSV0 U44451 ( .A1(n39837), .A2(n39836), .Z(n39838) );
  XNOR2HSV1 U44452 ( .A1(n39839), .A2(n39838), .ZN(n39842) );
  INHSV2 U44453 ( .I(n30888), .ZN(n51224) );
  CLKNAND2HSV1 U44454 ( .A1(n44694), .A2(n51224), .ZN(n39841) );
  XOR2HSV0 U44455 ( .A1(n39842), .A2(n39841), .Z(n39843) );
  XNOR2HSV1 U44456 ( .A1(n39844), .A2(n39843), .ZN(n39846) );
  NAND2HSV0 U44457 ( .A1(n59517), .A2(n50495), .ZN(n39845) );
  XNOR2HSV1 U44458 ( .A1(n39846), .A2(n39845), .ZN(n39847) );
  XOR2HSV0 U44459 ( .A1(n39848), .A2(n39847), .Z(n39851) );
  NAND2HSV0 U44460 ( .A1(n48746), .A2(n40185), .ZN(n39850) );
  CLKNHSV1 U44461 ( .I(n40116), .ZN(n46960) );
  CLKNAND2HSV0 U44462 ( .A1(n40116), .A2(n40170), .ZN(n39849) );
  XOR3HSV2 U44463 ( .A1(n39851), .A2(n39850), .A3(n39849), .Z(n39852) );
  XOR2HSV0 U44464 ( .A1(n39853), .A2(n39852), .Z(n39854) );
  XNOR2HSV1 U44465 ( .A1(n39855), .A2(n39854), .ZN(n39856) );
  XNOR2HSV1 U44466 ( .A1(n39857), .A2(n39856), .ZN(n39858) );
  NAND2HSV2 U44467 ( .A1(n39860), .A2(n48742), .ZN(n39861) );
  XNOR2HSV1 U44468 ( .A1(n39862), .A2(n39861), .ZN(n39863) );
  BUFHSV8 U44469 ( .I(n47041), .Z(n45499) );
  CLKNAND2HSV2 U44470 ( .A1(n39867), .A2(n39866), .ZN(n40136) );
  INHSV2 U44471 ( .I(n40136), .ZN(n39868) );
  NOR2HSV2 U44472 ( .A1(n39868), .A2(n40169), .ZN(n39870) );
  INHSV2 U44473 ( .I(n40139), .ZN(n39876) );
  CLKNAND2HSV1 U44474 ( .A1(n39872), .A2(n39871), .ZN(n39873) );
  NOR2HSV0 U44475 ( .A1(n39874), .A2(n39873), .ZN(n39875) );
  CLKNAND2HSV1 U44476 ( .A1(n39877), .A2(n59946), .ZN(n39878) );
  CLKNHSV0 U44477 ( .I(n45489), .ZN(n40018) );
  NOR2HSV1 U44478 ( .A1(n40018), .A2(n37635), .ZN(n39985) );
  CLKBUFHSV2 U44479 ( .I(n40278), .Z(n40019) );
  CLKNAND2HSV1 U44480 ( .A1(n40019), .A2(n48742), .ZN(n39984) );
  BUFHSV2 U44481 ( .I(n51158), .Z(n48747) );
  NAND2HSV2 U44482 ( .A1(n48747), .A2(n47267), .ZN(n39977) );
  CLKNAND2HSV1 U44483 ( .A1(n40021), .A2(n45816), .ZN(n39973) );
  CLKNAND2HSV0 U44484 ( .A1(n51160), .A2(n50495), .ZN(n39969) );
  CLKNAND2HSV1 U44485 ( .A1(n59392), .A2(n46974), .ZN(n39967) );
  NAND2HSV0 U44486 ( .A1(n59871), .A2(n39881), .ZN(n39965) );
  CLKNAND2HSV0 U44487 ( .A1(n30781), .A2(n51157), .ZN(n39963) );
  NAND2HSV0 U44488 ( .A1(n48624), .A2(n40186), .ZN(n39961) );
  CLKNHSV0 U44489 ( .I(n45817), .ZN(n50497) );
  NAND2HSV0 U44490 ( .A1(n39258), .A2(n50497), .ZN(n39959) );
  CLKNAND2HSV0 U44491 ( .A1(n37558), .A2(\pe5/got [10]), .ZN(n39953) );
  CLKNAND2HSV0 U44492 ( .A1(n48169), .A2(n40257), .ZN(n39951) );
  NAND2HSV0 U44493 ( .A1(n44335), .A2(\pe5/pvq [28]), .ZN(n39883) );
  XOR2HSV0 U44494 ( .A1(n39883), .A2(\pe5/phq [28]), .Z(n39886) );
  NAND2HSV0 U44495 ( .A1(n48658), .A2(n31160), .ZN(n40233) );
  OAI22HSV0 U44496 ( .A1(n30287), .A2(n50507), .B1(n59641), .B2(n37564), .ZN(
        n39884) );
  OAI21HSV0 U44497 ( .A1(n48680), .A2(n40233), .B(n39884), .ZN(n39885) );
  XNOR2HSV1 U44498 ( .A1(n39886), .A2(n39885), .ZN(n39893) );
  CLKNAND2HSV0 U44499 ( .A1(n39887), .A2(\pe5/bq[7] ), .ZN(n50678) );
  OAI21HSV0 U44500 ( .A1(n48246), .A2(n30116), .B(n40238), .ZN(n39888) );
  OAI21HSV0 U44501 ( .A1(n39889), .A2(n50678), .B(n39888), .ZN(n39891) );
  CLKNHSV0 U44502 ( .I(n47409), .ZN(n50588) );
  NAND2HSV0 U44503 ( .A1(n50588), .A2(n30789), .ZN(n39890) );
  XNOR2HSV1 U44504 ( .A1(n39891), .A2(n39890), .ZN(n39892) );
  XNOR2HSV1 U44505 ( .A1(n39893), .A2(n39892), .ZN(n39911) );
  NAND2HSV0 U44506 ( .A1(n59393), .A2(n51200), .ZN(n39910) );
  NAND2HSV0 U44507 ( .A1(n40210), .A2(n51048), .ZN(n39895) );
  CLKNAND2HSV0 U44508 ( .A1(n48172), .A2(n51191), .ZN(n39894) );
  XOR2HSV0 U44509 ( .A1(n39895), .A2(n39894), .Z(n39899) );
  NAND2HSV0 U44510 ( .A1(n40234), .A2(\pe5/bq[9] ), .ZN(n39897) );
  CLKNHSV0 U44511 ( .I(n51021), .ZN(n50504) );
  NAND2HSV0 U44512 ( .A1(n39496), .A2(n50504), .ZN(n39896) );
  XOR2HSV0 U44513 ( .A1(n39897), .A2(n39896), .Z(n39898) );
  XOR2HSV0 U44514 ( .A1(n39899), .A2(n39898), .Z(n39908) );
  CLKNAND2HSV0 U44515 ( .A1(n39499), .A2(n50668), .ZN(n39901) );
  NAND2HSV0 U44516 ( .A1(\pe5/got [5]), .A2(n37584), .ZN(n39900) );
  XOR2HSV0 U44517 ( .A1(n39901), .A2(n39900), .Z(n39906) );
  NAND2HSV0 U44518 ( .A1(n47278), .A2(n47059), .ZN(n39904) );
  BUFHSV2 U44519 ( .I(\pe5/bq[10] ), .Z(n48778) );
  NAND2HSV0 U44520 ( .A1(n39902), .A2(n48778), .ZN(n39903) );
  XOR2HSV0 U44521 ( .A1(n39904), .A2(n39903), .Z(n39905) );
  XOR2HSV0 U44522 ( .A1(n39906), .A2(n39905), .Z(n39907) );
  XOR2HSV0 U44523 ( .A1(n39908), .A2(n39907), .Z(n39909) );
  XOR3HSV2 U44524 ( .A1(n39911), .A2(n39910), .A3(n39909), .Z(n39913) );
  NAND2HSV0 U44525 ( .A1(n48751), .A2(n50698), .ZN(n39912) );
  XNOR2HSV1 U44526 ( .A1(n39913), .A2(n39912), .ZN(n39949) );
  NAND2HSV0 U44527 ( .A1(\pe5/aot [13]), .A2(n30692), .ZN(n39916) );
  NAND2HSV0 U44528 ( .A1(n48171), .A2(n39914), .ZN(n39915) );
  XOR2HSV0 U44529 ( .A1(n39916), .A2(n39915), .Z(n39920) );
  NAND2HSV0 U44530 ( .A1(n48634), .A2(n39615), .ZN(n39918) );
  NAND2HSV0 U44531 ( .A1(n31175), .A2(\pe5/bq[11] ), .ZN(n39917) );
  XOR2HSV0 U44532 ( .A1(n39918), .A2(n39917), .Z(n39919) );
  XOR2HSV0 U44533 ( .A1(n39920), .A2(n39919), .Z(n39929) );
  NAND2HSV0 U44534 ( .A1(n48663), .A2(n48760), .ZN(n39923) );
  NAND2HSV0 U44535 ( .A1(n40190), .A2(n39921), .ZN(n39922) );
  XOR2HSV0 U44536 ( .A1(n39923), .A2(n39922), .Z(n39927) );
  NAND2HSV0 U44537 ( .A1(n50511), .A2(n30230), .ZN(n39925) );
  CLKNAND2HSV0 U44538 ( .A1(n59640), .A2(n46933), .ZN(n39924) );
  XOR2HSV0 U44539 ( .A1(n39925), .A2(n39924), .Z(n39926) );
  XOR2HSV0 U44540 ( .A1(n39927), .A2(n39926), .Z(n39928) );
  XOR2HSV0 U44541 ( .A1(n39929), .A2(n39928), .Z(n39945) );
  NAND2HSV0 U44542 ( .A1(n59642), .A2(n30256), .ZN(n39931) );
  NAND2HSV0 U44543 ( .A1(\pe5/aot [18]), .A2(n39454), .ZN(n39930) );
  XOR2HSV0 U44544 ( .A1(n39931), .A2(n39930), .Z(n39935) );
  NAND2HSV0 U44545 ( .A1(\pe5/aot [23]), .A2(n40221), .ZN(n39933) );
  NAND2HSV0 U44546 ( .A1(n48205), .A2(n40207), .ZN(n39932) );
  XOR2HSV0 U44547 ( .A1(n39933), .A2(n39932), .Z(n39934) );
  XOR2HSV0 U44548 ( .A1(n39935), .A2(n39934), .Z(n39943) );
  CLKNAND2HSV0 U44549 ( .A1(n52591), .A2(n48236), .ZN(n39937) );
  NAND2HSV0 U44550 ( .A1(n51187), .A2(n52610), .ZN(n39936) );
  XOR2HSV0 U44551 ( .A1(n39937), .A2(n39936), .Z(n39941) );
  NAND2HSV0 U44552 ( .A1(n53304), .A2(n40074), .ZN(n39939) );
  NAND2HSV0 U44553 ( .A1(\pe5/aot [6]), .A2(n39436), .ZN(n39938) );
  XOR2HSV0 U44554 ( .A1(n39939), .A2(n39938), .Z(n39940) );
  XOR2HSV0 U44555 ( .A1(n39941), .A2(n39940), .Z(n39942) );
  XOR2HSV0 U44556 ( .A1(n39943), .A2(n39942), .Z(n39944) );
  XOR2HSV0 U44557 ( .A1(n39945), .A2(n39944), .Z(n39947) );
  CLKNHSV0 U44558 ( .I(n46978), .ZN(n51159) );
  NAND2HSV0 U44559 ( .A1(n48014), .A2(n51159), .ZN(n39946) );
  XNOR2HSV1 U44560 ( .A1(n39947), .A2(n39946), .ZN(n39948) );
  XNOR2HSV1 U44561 ( .A1(n39949), .A2(n39948), .ZN(n39950) );
  XNOR2HSV1 U44562 ( .A1(n39951), .A2(n39950), .ZN(n39952) );
  XNOR2HSV1 U44563 ( .A1(n39953), .A2(n39952), .ZN(n39957) );
  CLKNAND2HSV0 U44564 ( .A1(n48750), .A2(n59643), .ZN(n39956) );
  NAND2HSV0 U44565 ( .A1(n39954), .A2(n48167), .ZN(n39955) );
  XOR3HSV2 U44566 ( .A1(n39957), .A2(n39956), .A3(n39955), .Z(n39958) );
  XNOR2HSV1 U44567 ( .A1(n39959), .A2(n39958), .ZN(n39960) );
  XNOR2HSV1 U44568 ( .A1(n39961), .A2(n39960), .ZN(n39962) );
  XOR2HSV0 U44569 ( .A1(n39963), .A2(n39962), .Z(n39964) );
  XNOR2HSV1 U44570 ( .A1(n39965), .A2(n39964), .ZN(n39966) );
  XOR2HSV0 U44571 ( .A1(n39967), .A2(n39966), .Z(n39968) );
  XNOR2HSV1 U44572 ( .A1(n39969), .A2(n39968), .ZN(n39971) );
  NAND2HSV0 U44573 ( .A1(n44694), .A2(n51103), .ZN(n39970) );
  XOR2HSV0 U44574 ( .A1(n39971), .A2(n39970), .Z(n39972) );
  XNOR2HSV1 U44575 ( .A1(n39973), .A2(n39972), .ZN(n39975) );
  NAND2HSV0 U44576 ( .A1(n51205), .A2(n37656), .ZN(n39974) );
  XNOR2HSV1 U44577 ( .A1(n39975), .A2(n39974), .ZN(n39976) );
  XNOR2HSV1 U44578 ( .A1(n39977), .A2(n39976), .ZN(n39980) );
  BUFHSV4 U44579 ( .I(n48746), .Z(n45818) );
  NAND2HSV2 U44580 ( .A1(n45818), .A2(n59948), .ZN(n39979) );
  CLKNAND2HSV0 U44581 ( .A1(n40116), .A2(n48743), .ZN(n39978) );
  XNOR3HSV1 U44582 ( .A1(n39980), .A2(n39979), .A3(n39978), .ZN(n39981) );
  XOR2HSV0 U44583 ( .A1(n39982), .A2(n39981), .Z(n39983) );
  CLKNAND2HSV1 U44584 ( .A1(n39985), .A2(n39987), .ZN(n39986) );
  INHSV2 U44585 ( .I(n39986), .ZN(n39989) );
  AOI21HSV2 U44586 ( .A1(n59926), .A2(n31225), .B(n39987), .ZN(n39988) );
  NOR2HSV2 U44587 ( .A1(n39989), .A2(n39988), .ZN(n39990) );
  NAND2HSV2 U44588 ( .A1(n39860), .A2(n30142), .ZN(n39993) );
  NOR2HSV2 U44589 ( .A1(n39996), .A2(n39995), .ZN(n39997) );
  OAI21HSV4 U44590 ( .A1(n60068), .A2(n39230), .B(n39997), .ZN(n39998) );
  INHSV2 U44591 ( .I(n39998), .ZN(n39999) );
  NOR2HSV4 U44592 ( .A1(n52836), .A2(n39383), .ZN(n40001) );
  XNOR2HSV4 U44593 ( .A1(n40005), .A2(n40004), .ZN(n40010) );
  INHSV3 U44594 ( .I(n40166), .ZN(n40165) );
  NOR2HSV4 U44595 ( .A1(n40010), .A2(n40009), .ZN(n40011) );
  OAI21HSV1 U44596 ( .A1(n40012), .A2(\pe5/ti_7t [28]), .B(n52694), .ZN(n40157) );
  NOR2HSV1 U44597 ( .A1(n40157), .A2(n39730), .ZN(n40013) );
  NAND2HSV2 U44598 ( .A1(n40159), .A2(n40013), .ZN(n40016) );
  AOI21HSV4 U44599 ( .A1(n39739), .A2(n40017), .B(n39246), .ZN(n40149) );
  NOR2HSV2 U44600 ( .A1(n40018), .A2(n31081), .ZN(n40125) );
  CLKNAND2HSV0 U44601 ( .A1(n40278), .A2(n37630), .ZN(n40123) );
  NAND2HSV0 U44602 ( .A1(n52570), .A2(n40170), .ZN(n40115) );
  CLKNAND2HSV0 U44603 ( .A1(n40021), .A2(n47056), .ZN(n40111) );
  CLKNAND2HSV0 U44604 ( .A1(n51019), .A2(n46974), .ZN(n40107) );
  NAND2HSV0 U44605 ( .A1(n59392), .A2(n51224), .ZN(n40105) );
  NAND2HSV0 U44606 ( .A1(n52575), .A2(n51157), .ZN(n40103) );
  NAND2HSV0 U44607 ( .A1(n40171), .A2(n40186), .ZN(n40101) );
  NAND2HSV0 U44608 ( .A1(n48624), .A2(n50497), .ZN(n40099) );
  NAND2HSV0 U44609 ( .A1(n39882), .A2(n48167), .ZN(n40097) );
  NAND2HSV0 U44610 ( .A1(n37558), .A2(n59891), .ZN(n40092) );
  NAND2HSV0 U44611 ( .A1(n48751), .A2(n52573), .ZN(n40088) );
  NAND2HSV0 U44612 ( .A1(n47278), .A2(n46933), .ZN(n40023) );
  NAND2HSV0 U44613 ( .A1(n48761), .A2(\pe5/bq[11] ), .ZN(n40022) );
  XOR2HSV0 U44614 ( .A1(n40023), .A2(n40022), .Z(n40027) );
  NAND2HSV0 U44615 ( .A1(n31175), .A2(n48778), .ZN(n40025) );
  CLKNHSV0 U44616 ( .I(n48822), .ZN(n50444) );
  NAND2HSV0 U44617 ( .A1(\pe5/aot [18]), .A2(n50444), .ZN(n40024) );
  XOR2HSV0 U44618 ( .A1(n40025), .A2(n40024), .Z(n40026) );
  XOR2HSV0 U44619 ( .A1(n40027), .A2(n40026), .Z(n40035) );
  NAND2HSV0 U44620 ( .A1(n39490), .A2(n47059), .ZN(n40029) );
  NAND2HSV0 U44621 ( .A1(\pe5/aot [13]), .A2(n31160), .ZN(n40028) );
  XOR2HSV0 U44622 ( .A1(n40029), .A2(n40028), .Z(n40033) );
  NAND2HSV0 U44623 ( .A1(n53304), .A2(n30230), .ZN(n40031) );
  NAND2HSV0 U44624 ( .A1(n51313), .A2(n30222), .ZN(n40030) );
  XOR2HSV0 U44625 ( .A1(n40031), .A2(n40030), .Z(n40032) );
  XOR2HSV0 U44626 ( .A1(n40033), .A2(n40032), .Z(n40034) );
  XOR2HSV0 U44627 ( .A1(n40035), .A2(n40034), .Z(n40051) );
  NAND2HSV0 U44628 ( .A1(\pe5/got [4]), .A2(n37584), .ZN(n40037) );
  NAND2HSV0 U44629 ( .A1(n40234), .A2(n48760), .ZN(n40036) );
  XOR2HSV0 U44630 ( .A1(n40037), .A2(n40036), .Z(n40041) );
  NAND2HSV0 U44631 ( .A1(n39499), .A2(n31045), .ZN(n40039) );
  NAND2HSV0 U44632 ( .A1(n48663), .A2(\pe5/bq[7] ), .ZN(n40038) );
  XOR2HSV0 U44633 ( .A1(n40039), .A2(n40038), .Z(n40040) );
  XOR2HSV0 U44634 ( .A1(n40041), .A2(n40040), .Z(n40049) );
  NAND2HSV0 U44635 ( .A1(\pe5/pvq [29]), .A2(n48029), .ZN(n40042) );
  XOR2HSV0 U44636 ( .A1(n40042), .A2(\pe5/phq [29]), .Z(n40047) );
  NAND2HSV0 U44637 ( .A1(\pe5/aot [23]), .A2(\pe5/bq[5] ), .ZN(n47241) );
  OAI22HSV0 U44638 ( .A1(n39779), .A2(n51021), .B1(n40043), .B2(n48050), .ZN(
        n40044) );
  OAI21HSV0 U44639 ( .A1(n40045), .A2(n47241), .B(n40044), .ZN(n40046) );
  XOR2HSV0 U44640 ( .A1(n40047), .A2(n40046), .Z(n40048) );
  XNOR2HSV1 U44641 ( .A1(n40049), .A2(n40048), .ZN(n40050) );
  XNOR2HSV1 U44642 ( .A1(n40051), .A2(n40050), .ZN(n40053) );
  NAND2HSV0 U44643 ( .A1(n39278), .A2(n48841), .ZN(n40052) );
  XNOR2HSV1 U44644 ( .A1(n40053), .A2(n40052), .ZN(n40087) );
  NAND2HSV0 U44645 ( .A1(n52584), .A2(n30891), .ZN(n40055) );
  NAND2HSV0 U44646 ( .A1(n48829), .A2(n51307), .ZN(n40054) );
  XOR2HSV0 U44647 ( .A1(n40055), .A2(n40054), .Z(n40059) );
  NAND2HSV0 U44648 ( .A1(n39496), .A2(\pe5/bq[4] ), .ZN(n40057) );
  NAND2HSV0 U44649 ( .A1(n51187), .A2(n39914), .ZN(n40056) );
  XOR2HSV0 U44650 ( .A1(n40057), .A2(n40056), .Z(n40058) );
  XOR2HSV0 U44651 ( .A1(n40059), .A2(n40058), .Z(n40067) );
  NAND2HSV0 U44652 ( .A1(n40190), .A2(n48236), .ZN(n40061) );
  NAND2HSV0 U44653 ( .A1(\pe5/aot [16]), .A2(n48237), .ZN(n40060) );
  XOR2HSV0 U44654 ( .A1(n40061), .A2(n40060), .Z(n40065) );
  NAND2HSV0 U44655 ( .A1(n50501), .A2(n30789), .ZN(n40063) );
  NAND2HSV0 U44656 ( .A1(n51188), .A2(n40221), .ZN(n40062) );
  XOR2HSV0 U44657 ( .A1(n40063), .A2(n40062), .Z(n40064) );
  XOR2HSV0 U44658 ( .A1(n40065), .A2(n40064), .Z(n40066) );
  XOR2HSV0 U44659 ( .A1(n40067), .A2(n40066), .Z(n40083) );
  NAND2HSV0 U44660 ( .A1(\pe5/aot [9]), .A2(n30256), .ZN(n40069) );
  NAND2HSV0 U44661 ( .A1(n50511), .A2(n48802), .ZN(n40068) );
  XOR2HSV0 U44662 ( .A1(n40069), .A2(n40068), .Z(n40073) );
  NAND2HSV0 U44663 ( .A1(n48205), .A2(n46622), .ZN(n40071) );
  NAND2HSV0 U44664 ( .A1(n59427), .A2(n50526), .ZN(n40070) );
  XOR2HSV0 U44665 ( .A1(n40071), .A2(n40070), .Z(n40072) );
  XOR2HSV0 U44666 ( .A1(n40073), .A2(n40072), .Z(n40081) );
  NOR2HSV0 U44667 ( .A1(n45815), .A2(n39796), .ZN(n40076) );
  NAND2HSV0 U44668 ( .A1(\pe5/aot [6]), .A2(n40074), .ZN(n40075) );
  XOR2HSV0 U44669 ( .A1(n40076), .A2(n40075), .Z(n40079) );
  NAND2HSV0 U44670 ( .A1(n40210), .A2(n39454), .ZN(n51170) );
  NAND2HSV0 U44671 ( .A1(n51363), .A2(n30698), .ZN(n40077) );
  XOR2HSV0 U44672 ( .A1(n51170), .A2(n40077), .Z(n40078) );
  XOR2HSV0 U44673 ( .A1(n40079), .A2(n40078), .Z(n40080) );
  XOR2HSV0 U44674 ( .A1(n40081), .A2(n40080), .Z(n40082) );
  XOR2HSV0 U44675 ( .A1(n40083), .A2(n40082), .Z(n40085) );
  NAND2HSV0 U44676 ( .A1(n48014), .A2(n51200), .ZN(n40084) );
  XNOR2HSV1 U44677 ( .A1(n40085), .A2(n40084), .ZN(n40086) );
  XOR3HSV2 U44678 ( .A1(n40088), .A2(n40087), .A3(n40086), .Z(n40090) );
  NAND2HSV0 U44679 ( .A1(n48169), .A2(n47144), .ZN(n40089) );
  XOR2HSV0 U44680 ( .A1(n40090), .A2(n40089), .Z(n40091) );
  XNOR2HSV1 U44681 ( .A1(n40092), .A2(n40091), .ZN(n40095) );
  NAND2HSV0 U44682 ( .A1(n48750), .A2(n51210), .ZN(n40094) );
  NAND2HSV0 U44683 ( .A1(n39954), .A2(n59643), .ZN(n40093) );
  XOR3HSV2 U44684 ( .A1(n40095), .A2(n40094), .A3(n40093), .Z(n40096) );
  XNOR2HSV1 U44685 ( .A1(n40097), .A2(n40096), .ZN(n40098) );
  XNOR2HSV1 U44686 ( .A1(n40099), .A2(n40098), .ZN(n40100) );
  XOR2HSV0 U44687 ( .A1(n40101), .A2(n40100), .Z(n40102) );
  XNOR2HSV1 U44688 ( .A1(n40103), .A2(n40102), .ZN(n40104) );
  XOR2HSV0 U44689 ( .A1(n40105), .A2(n40104), .Z(n40106) );
  XNOR2HSV1 U44690 ( .A1(n40107), .A2(n40106), .ZN(n40109) );
  NAND2HSV0 U44691 ( .A1(n44694), .A2(n52566), .ZN(n40108) );
  XOR2HSV0 U44692 ( .A1(n40109), .A2(n40108), .Z(n40110) );
  XNOR2HSV1 U44693 ( .A1(n40111), .A2(n40110), .ZN(n40113) );
  NAND2HSV0 U44694 ( .A1(n59517), .A2(n40185), .ZN(n40112) );
  XNOR2HSV1 U44695 ( .A1(n40113), .A2(n40112), .ZN(n40114) );
  XNOR2HSV1 U44696 ( .A1(n40115), .A2(n40114), .ZN(n40119) );
  NAND2HSV2 U44697 ( .A1(n45818), .A2(n47267), .ZN(n40118) );
  NAND2HSV0 U44698 ( .A1(n40116), .A2(n59948), .ZN(n40117) );
  XOR3HSV2 U44699 ( .A1(n40119), .A2(n40118), .A3(n40117), .Z(n40120) );
  XOR2HSV0 U44700 ( .A1(n40121), .A2(n40120), .Z(n40122) );
  XNOR2HSV1 U44701 ( .A1(n40123), .A2(n40122), .ZN(n40124) );
  XNOR2HSV1 U44702 ( .A1(n40125), .A2(n40124), .ZN(n40126) );
  NOR2HSV2 U44703 ( .A1(n44329), .A2(n48164), .ZN(n40128) );
  XOR2HSV0 U44704 ( .A1(n40129), .A2(n40128), .Z(n40135) );
  NOR2HSV1 U44705 ( .A1(n40131), .A2(n40130), .ZN(n40132) );
  AOI21HSV2 U44706 ( .A1(n60068), .A2(n40133), .B(n40132), .ZN(n40134) );
  NAND3HSV2 U44707 ( .A1(n40137), .A2(n59395), .A3(n40136), .ZN(n40146) );
  CLKNHSV0 U44708 ( .I(n40138), .ZN(n40140) );
  NOR2HSV2 U44709 ( .A1(n40143), .A2(n31003), .ZN(n40144) );
  XNOR2HSV4 U44710 ( .A1(n40148), .A2(n40147), .ZN(n40150) );
  NAND2HSV2 U44711 ( .A1(n40149), .A2(n40150), .ZN(n40154) );
  CLKAND2HSV2 U44712 ( .A1(n47387), .A2(\pe5/ti_7t [29]), .Z(n40155) );
  AOI21HSV4 U44713 ( .A1(n40156), .A2(n52838), .B(n40155), .ZN(n44662) );
  INHSV2 U44714 ( .I(n40157), .ZN(n40158) );
  INHSV2 U44715 ( .I(n40160), .ZN(n40161) );
  NAND2HSV4 U44716 ( .A1(n25829), .A2(n40161), .ZN(n52839) );
  NOR2HSV4 U44717 ( .A1(n52838), .A2(n40162), .ZN(n40163) );
  CLKNAND2HSV4 U44718 ( .A1(n40163), .A2(n52839), .ZN(n44663) );
  CLKNAND2HSV3 U44719 ( .A1(n40168), .A2(n40167), .ZN(n40314) );
  INHSV2 U44720 ( .I(n40314), .ZN(n47392) );
  NOR2HSV2 U44721 ( .A1(n40302), .A2(n40169), .ZN(n40292) );
  NAND2HSV2 U44722 ( .A1(n45818), .A2(n40170), .ZN(n40180) );
  NAND2HSV2 U44723 ( .A1(n40021), .A2(n50495), .ZN(n40176) );
  CLKNAND2HSV1 U44724 ( .A1(n29770), .A2(n50497), .ZN(n40174) );
  NAND2HSV0 U44725 ( .A1(n40172), .A2(n48167), .ZN(n40173) );
  XOR2HSV0 U44726 ( .A1(n40174), .A2(n40173), .Z(n40175) );
  XNOR2HSV1 U44727 ( .A1(n40176), .A2(n40175), .ZN(n40178) );
  NAND2HSV0 U44728 ( .A1(n51205), .A2(n47056), .ZN(n40177) );
  XNOR2HSV1 U44729 ( .A1(n40178), .A2(n40177), .ZN(n40179) );
  XOR2HSV0 U44730 ( .A1(n40180), .A2(n40179), .Z(n40182) );
  NAND2HSV2 U44731 ( .A1(n51211), .A2(n39532), .ZN(n40181) );
  XNOR2HSV1 U44732 ( .A1(n40182), .A2(n40181), .ZN(n40184) );
  OAI21HSV2 U44733 ( .A1(n51361), .A2(n39743), .B(n40184), .ZN(n40183) );
  OAI31HSV2 U44734 ( .A1(n48166), .A2(n39743), .A3(n40184), .B(n40183), .ZN(
        n40274) );
  NAND2HSV2 U44735 ( .A1(n48747), .A2(n40185), .ZN(n40272) );
  CLKNAND2HSV0 U44736 ( .A1(n39257), .A2(n52658), .ZN(n40268) );
  NAND2HSV2 U44737 ( .A1(n59392), .A2(n51015), .ZN(n40266) );
  NAND2HSV2 U44738 ( .A1(n59871), .A2(n40186), .ZN(n40264) );
  NAND2HSV2 U44739 ( .A1(n30885), .A2(n59643), .ZN(n40262) );
  CLKNAND2HSV1 U44740 ( .A1(n30515), .A2(n47144), .ZN(n40256) );
  NAND2HSV0 U44741 ( .A1(n40187), .A2(n51200), .ZN(n40252) );
  NAND2HSV0 U44742 ( .A1(\pe5/aot [16]), .A2(\pe5/bq[19] ), .ZN(n40189) );
  CLKNAND2HSV1 U44743 ( .A1(\pe5/aot [18]), .A2(n48236), .ZN(n40188) );
  XOR2HSV0 U44744 ( .A1(n40189), .A2(n40188), .Z(n40194) );
  NAND2HSV2 U44745 ( .A1(n40190), .A2(n48181), .ZN(n40192) );
  NAND2HSV0 U44746 ( .A1(n51313), .A2(n46622), .ZN(n40191) );
  XOR2HSV0 U44747 ( .A1(n40192), .A2(n40191), .Z(n40193) );
  XOR2HSV0 U44748 ( .A1(n40194), .A2(n40193), .Z(n40202) );
  NAND2HSV0 U44749 ( .A1(n53295), .A2(n48755), .ZN(n40196) );
  CLKNAND2HSV0 U44750 ( .A1(n48829), .A2(n48760), .ZN(n40195) );
  XOR2HSV0 U44751 ( .A1(n40196), .A2(n40195), .Z(n40200) );
  NAND2HSV2 U44752 ( .A1(n48761), .A2(n48778), .ZN(n40198) );
  NAND2HSV0 U44753 ( .A1(n53304), .A2(n30357), .ZN(n40197) );
  XOR2HSV0 U44754 ( .A1(n40198), .A2(n40197), .Z(n40199) );
  XOR2HSV0 U44755 ( .A1(n40200), .A2(n40199), .Z(n40201) );
  XOR2HSV0 U44756 ( .A1(n40202), .A2(n40201), .Z(n40204) );
  NAND2HSV0 U44757 ( .A1(n30806), .A2(n52577), .ZN(n40203) );
  XNOR2HSV1 U44758 ( .A1(n40204), .A2(n40203), .ZN(n40206) );
  NAND2HSV0 U44759 ( .A1(n48014), .A2(n48841), .ZN(n40205) );
  XNOR2HSV1 U44760 ( .A1(n40206), .A2(n40205), .ZN(n40251) );
  NAND2HSV0 U44761 ( .A1(\pe5/aot [14]), .A2(n31190), .ZN(n40209) );
  NAND2HSV0 U44762 ( .A1(\pe5/aot [9]), .A2(n40207), .ZN(n40208) );
  XOR2HSV0 U44763 ( .A1(n40209), .A2(n40208), .Z(n40212) );
  XOR2HSV0 U44764 ( .A1(n40212), .A2(n40211), .Z(n40218) );
  NAND2HSV0 U44765 ( .A1(n30529), .A2(n50526), .ZN(n40214) );
  NAND2HSV0 U44766 ( .A1(\pe5/aot [4]), .A2(n30698), .ZN(n40213) );
  XOR2HSV0 U44767 ( .A1(n40214), .A2(n40213), .Z(n40216) );
  XOR2HSV0 U44768 ( .A1(n40216), .A2(n40215), .Z(n40217) );
  XOR2HSV0 U44769 ( .A1(n40218), .A2(n40217), .Z(n40231) );
  NAND2HSV2 U44770 ( .A1(n52591), .A2(n39914), .ZN(n40220) );
  NAND2HSV0 U44771 ( .A1(n59355), .A2(n30693), .ZN(n40219) );
  XOR2HSV0 U44772 ( .A1(n40220), .A2(n40219), .Z(n40225) );
  NAND2HSV0 U44773 ( .A1(\pe5/aot [3]), .A2(n30789), .ZN(n40223) );
  NAND2HSV0 U44774 ( .A1(n48242), .A2(n40221), .ZN(n40222) );
  XOR2HSV0 U44775 ( .A1(n40223), .A2(n40222), .Z(n40224) );
  XOR2HSV0 U44776 ( .A1(n40225), .A2(n40224), .Z(n40229) );
  CLKNAND2HSV1 U44777 ( .A1(n39473), .A2(n40226), .ZN(n47325) );
  XNOR2HSV1 U44778 ( .A1(n40229), .A2(n40228), .ZN(n40230) );
  XNOR2HSV1 U44779 ( .A1(n40231), .A2(n40230), .ZN(n40249) );
  XOR2HSV0 U44780 ( .A1(n40233), .A2(n40232), .Z(n40247) );
  CLKNAND2HSV0 U44781 ( .A1(n40234), .A2(n51373), .ZN(n48828) );
  OAI22HSV0 U44782 ( .A1(n40236), .A2(n51021), .B1(n40235), .B2(n47207), .ZN(
        n40237) );
  OAI21HSV2 U44783 ( .A1(n40238), .A2(n48828), .B(n40237), .ZN(n40239) );
  NAND2HSV2 U44784 ( .A1(\pe5/aot [13]), .A2(n47059), .ZN(n51164) );
  XNOR2HSV1 U44785 ( .A1(n40239), .A2(n51164), .ZN(n40246) );
  NAND2HSV0 U44786 ( .A1(n59945), .A2(n48198), .ZN(n40241) );
  NAND2HSV0 U44787 ( .A1(n52675), .A2(n48787), .ZN(n40240) );
  XOR2HSV0 U44788 ( .A1(n40241), .A2(n40240), .Z(n40244) );
  NAND2HSV2 U44789 ( .A1(n48172), .A2(\pe5/bq[4] ), .ZN(n48815) );
  CLKNAND2HSV0 U44790 ( .A1(n48205), .A2(n30341), .ZN(n40242) );
  XOR2HSV0 U44791 ( .A1(n48815), .A2(n40242), .Z(n40243) );
  XOR2HSV0 U44792 ( .A1(n40244), .A2(n40243), .Z(n40245) );
  XOR3HSV2 U44793 ( .A1(n40247), .A2(n40246), .A3(n40245), .Z(n40248) );
  XNOR2HSV1 U44794 ( .A1(n40249), .A2(n40248), .ZN(n40250) );
  XOR3HSV2 U44795 ( .A1(n40252), .A2(n40251), .A3(n40250), .Z(n40254) );
  CLKNAND2HSV1 U44796 ( .A1(n48169), .A2(n51159), .ZN(n40253) );
  XOR2HSV0 U44797 ( .A1(n40254), .A2(n40253), .Z(n40255) );
  XNOR2HSV1 U44798 ( .A1(n40256), .A2(n40255), .ZN(n40260) );
  NAND2HSV2 U44799 ( .A1(n48750), .A2(n40257), .ZN(n40259) );
  NAND2HSV2 U44800 ( .A1(n47058), .A2(n51210), .ZN(n40258) );
  XOR3HSV2 U44801 ( .A1(n40260), .A2(n40259), .A3(n40258), .Z(n40261) );
  XNOR2HSV1 U44802 ( .A1(n40262), .A2(n40261), .ZN(n40263) );
  XNOR2HSV1 U44803 ( .A1(n40264), .A2(n40263), .ZN(n40265) );
  XOR2HSV0 U44804 ( .A1(n40266), .A2(n40265), .Z(n40267) );
  XNOR2HSV1 U44805 ( .A1(n40268), .A2(n40267), .ZN(n40270) );
  CLKNAND2HSV0 U44806 ( .A1(n44694), .A2(\pe5/got [17]), .ZN(n40269) );
  XOR2HSV0 U44807 ( .A1(n40270), .A2(n40269), .Z(n40271) );
  XNOR2HSV1 U44808 ( .A1(n40272), .A2(n40271), .ZN(n40273) );
  XOR2HSV0 U44809 ( .A1(n40274), .A2(n40273), .Z(n40277) );
  NOR2HSV2 U44810 ( .A1(n50692), .A2(n30210), .ZN(n40276) );
  XNOR3HSV1 U44811 ( .A1(n40277), .A2(n40276), .A3(n40275), .ZN(n40284) );
  CLKNAND2HSV1 U44812 ( .A1(n40019), .A2(n48743), .ZN(n40279) );
  AOI21HSV2 U44813 ( .A1(n53344), .A2(n31225), .B(n40279), .ZN(n40282) );
  CLKNAND2HSV0 U44814 ( .A1(n40279), .A2(n31225), .ZN(n40280) );
  NOR2HSV1 U44815 ( .A1(n39554), .A2(n40280), .ZN(n40281) );
  NOR2HSV2 U44816 ( .A1(n40282), .A2(n40281), .ZN(n40283) );
  XOR2HSV2 U44817 ( .A1(n40284), .A2(n40283), .Z(n40286) );
  CLKNHSV2 U44818 ( .I(n40287), .ZN(n40289) );
  CLKNHSV2 U44819 ( .I(n30046), .ZN(n40288) );
  INHSV3 U44820 ( .I(n40318), .ZN(n40301) );
  INHSV2 U44821 ( .I(n40301), .ZN(n40291) );
  MUX2NHSV2 U44822 ( .I0(n40293), .I1(n40292), .S(n40291), .ZN(n40299) );
  CLKNHSV0 U44823 ( .I(n40320), .ZN(n40298) );
  NAND3HSV3 U44824 ( .A1(n40296), .A2(n40295), .A3(n40294), .ZN(n45902) );
  INHSV4 U44825 ( .I(n45902), .ZN(n47139) );
  AOI21HSV2 U44826 ( .A1(n47139), .A2(n40301), .B(n37551), .ZN(n40297) );
  CLKNAND2HSV0 U44827 ( .A1(n40302), .A2(n40301), .ZN(n40303) );
  CLKNAND2HSV1 U44828 ( .A1(n40304), .A2(n40303), .ZN(n40308) );
  CLKNAND2HSV2 U44829 ( .A1(n40318), .A2(n30048), .ZN(n40306) );
  CLKAND2HSV2 U44830 ( .A1(n40306), .A2(n40305), .Z(n40307) );
  CLKNHSV0 U44831 ( .I(\pe5/ti_7t [30]), .ZN(n40311) );
  AOI21HSV1 U44832 ( .A1(n40311), .A2(n40310), .B(n40309), .ZN(n40312) );
  NOR2HSV4 U44833 ( .A1(n40316), .A2(n40315), .ZN(n47391) );
  CLKXOR2HSV4 U44834 ( .A1(n40319), .A2(n40318), .Z(n40322) );
  CLKNAND2HSV4 U44835 ( .A1(n40320), .A2(n52694), .ZN(n40321) );
  XNOR2HSV4 U44836 ( .A1(n40322), .A2(n40321), .ZN(n60067) );
  INHSV4 U44837 ( .I(\pe1/bq[31] ), .ZN(n40328) );
  BUFHSV8 U44838 ( .I(n40328), .Z(n40736) );
  CLKNHSV6 U44839 ( .I(ctro1), .ZN(n40343) );
  INHSV6 U44840 ( .I(n40343), .ZN(n40969) );
  INHSV4 U44841 ( .I(n40558), .ZN(n40332) );
  INHSV2 U44842 ( .I(n40649), .ZN(n53518) );
  NAND2HSV2 U44843 ( .A1(n41880), .A2(n53518), .ZN(n40325) );
  XNOR2HSV4 U44844 ( .A1(n40326), .A2(n40325), .ZN(n40337) );
  INHSV2 U44845 ( .I(n40445), .ZN(n59376) );
  INHSV4 U44846 ( .I(n40445), .ZN(n40568) );
  CLKNHSV6 U44847 ( .I(ctro1), .ZN(n40338) );
  CLKBUFHSV4 U44848 ( .I(n40338), .Z(n40598) );
  INHSV2 U44849 ( .I(\pe1/ti_7t [2]), .ZN(n40327) );
  INHSV2 U44850 ( .I(n40328), .ZN(n40385) );
  NAND2HSV4 U44851 ( .A1(n40385), .A2(\pe1/aot [32]), .ZN(n51112) );
  NAND2HSV0 U44852 ( .A1(n40568), .A2(\pe1/aot [32]), .ZN(n40330) );
  INHSV2 U44853 ( .I(n40330), .ZN(n40367) );
  NOR2HSV2 U44854 ( .A1(n40569), .A2(n40558), .ZN(n60110) );
  BUFHSV8 U44855 ( .I(n40338), .Z(n40547) );
  BUFHSV2 U44856 ( .I(n40335), .Z(n40525) );
  INHSV2 U44857 ( .I(n53787), .ZN(n40393) );
  XNOR2HSV4 U44858 ( .A1(n40337), .A2(n40336), .ZN(n40358) );
  INHSV4 U44859 ( .I(n40358), .ZN(n40355) );
  NOR2HSV4 U44860 ( .A1(n40339), .A2(n40335), .ZN(n40341) );
  NAND2HSV2 U44861 ( .A1(n40568), .A2(n40385), .ZN(n40348) );
  BUFHSV8 U44862 ( .I(n40343), .Z(n40437) );
  INHSV2 U44863 ( .I(n42335), .ZN(n41238) );
  INHSV2 U44864 ( .I(\pe1/got [32]), .ZN(n40520) );
  CLKNHSV1 U44865 ( .I(n40520), .ZN(n42339) );
  OA21HSV2 U44866 ( .A1(n40437), .A2(\pe1/ti_7t [3]), .B(n42339), .Z(n40344)
         );
  INHSV2 U44867 ( .I(n40654), .ZN(n59999) );
  XOR2HSV0 U44868 ( .A1(n40351), .A2(n25857), .Z(n40352) );
  CLKNAND2HSV2 U44869 ( .A1(n40353), .A2(n40352), .ZN(n40356) );
  NAND3HSV4 U44870 ( .A1(n40358), .A2(n40357), .A3(n40356), .ZN(n40359) );
  INHSV2 U44871 ( .I(n40396), .ZN(n60108) );
  NOR2HSV0 U44872 ( .A1(n40363), .A2(n40362), .ZN(n40370) );
  CLKNHSV0 U44873 ( .I(n51112), .ZN(n40364) );
  CLKNHSV0 U44874 ( .I(n40364), .ZN(n40369) );
  NOR2HSV1 U44875 ( .A1(n40367), .A2(n40366), .ZN(n40368) );
  NAND3HSV2 U44876 ( .A1(n40370), .A2(n40369), .A3(n40368), .ZN(n40373) );
  INHSV2 U44877 ( .I(n40520), .ZN(n53367) );
  NAND2HSV2 U44878 ( .A1(n40371), .A2(n53367), .ZN(n40372) );
  CLKNAND2HSV2 U44879 ( .A1(n40373), .A2(n40372), .ZN(n40374) );
  XNOR2HSV4 U44880 ( .A1(n40377), .A2(n40376), .ZN(n60009) );
  INHSV2 U44881 ( .I(\pe1/ti_7t [3]), .ZN(n40378) );
  BUFHSV4 U44882 ( .I(n40493), .Z(n42212) );
  INHSV2 U44883 ( .I(\pe1/bq[28] ), .ZN(n40446) );
  NOR2HSV2 U44884 ( .A1(n42212), .A2(n40416), .ZN(n40382) );
  INHSV2 U44885 ( .I(n40455), .ZN(n41339) );
  NAND2HSV2 U44886 ( .A1(n41339), .A2(n40879), .ZN(n40381) );
  CLKXOR2HSV4 U44887 ( .A1(n40382), .A2(n40381), .Z(n40384) );
  INHSV2 U44888 ( .I(n41228), .ZN(n54033) );
  CLKNAND2HSV2 U44889 ( .A1(n41880), .A2(n54033), .ZN(n40383) );
  NAND2HSV2 U44890 ( .A1(\pe1/aot [28]), .A2(n40385), .ZN(n40419) );
  BUFHSV6 U44891 ( .I(n40736), .Z(n41952) );
  INHSV4 U44892 ( .I(n40558), .ZN(n40501) );
  OAI22HSV4 U44893 ( .A1(n41952), .A2(n40412), .B1(n53447), .B2(n41334), .ZN(
        n40386) );
  NAND2HSV2 U44894 ( .A1(n40876), .A2(n53411), .ZN(n40387) );
  XNOR2HSV4 U44895 ( .A1(n40388), .A2(n40387), .ZN(n40389) );
  XNOR2HSV4 U44896 ( .A1(n40390), .A2(n40389), .ZN(n40392) );
  BUFHSV2 U44897 ( .I(n40649), .Z(n41331) );
  INHSV2 U44898 ( .I(n41331), .ZN(n40427) );
  INHSV2 U44899 ( .I(n40957), .ZN(n40394) );
  INHSV2 U44900 ( .I(n40404), .ZN(n40401) );
  INHSV2 U44901 ( .I(\pe1/ti_7t [4]), .ZN(n40395) );
  CLKNAND2HSV1 U44902 ( .A1(n40467), .A2(n41712), .ZN(n40408) );
  CLKAND2HSV2 U44903 ( .A1(n40408), .A2(n53367), .Z(n40397) );
  CLKNAND2HSV4 U44904 ( .A1(n40410), .A2(n40397), .ZN(n40402) );
  BUFHSV8 U44905 ( .I(n40786), .Z(n41930) );
  INHSV2 U44906 ( .I(n40398), .ZN(n40399) );
  NOR2HSV4 U44907 ( .A1(n41930), .A2(n40399), .ZN(n40403) );
  NOR2HSV4 U44908 ( .A1(n40402), .A2(n40403), .ZN(n40400) );
  CLKNAND2HSV3 U44909 ( .A1(n40400), .A2(n40401), .ZN(n40406) );
  NAND2HSV4 U44910 ( .A1(n40406), .A2(n40405), .ZN(n40477) );
  INHSV4 U44911 ( .I(n40477), .ZN(n40484) );
  CLKAND2HSV2 U44912 ( .A1(n40408), .A2(n40407), .Z(n40409) );
  CLKNAND2HSV2 U44913 ( .A1(n40410), .A2(n40409), .ZN(n40432) );
  INHSV2 U44914 ( .I(\pe1/got [28]), .ZN(n48450) );
  NAND2HSV2 U44915 ( .A1(n41880), .A2(\pe1/got [28]), .ZN(n40415) );
  NAND2HSV2 U44916 ( .A1(n40898), .A2(n40501), .ZN(n41162) );
  NOR2HSV2 U44917 ( .A1(n40445), .A2(n40416), .ZN(n40418) );
  INAND2HSV2 U44918 ( .A1(n40493), .B1(n40494), .ZN(n40417) );
  INHSV2 U44919 ( .I(n40455), .ZN(n42223) );
  XNOR2HSV4 U44920 ( .A1(n40421), .A2(n40420), .ZN(n40422) );
  XNOR2HSV4 U44921 ( .A1(n40423), .A2(n40422), .ZN(n40426) );
  XNOR2HSV4 U44922 ( .A1(n40426), .A2(n40425), .ZN(n40430) );
  CLKNHSV1 U44923 ( .I(n40427), .ZN(n40428) );
  NOR2HSV4 U44924 ( .A1(n40430), .A2(n40428), .ZN(n40429) );
  AOI22HSV4 U44925 ( .A1(n40431), .A2(n40430), .B1(n40429), .B2(n41930), .ZN(
        n40433) );
  INHSV2 U44926 ( .I(n40432), .ZN(n40435) );
  INHSV2 U44927 ( .I(n40433), .ZN(n40434) );
  CLKNAND2HSV3 U44928 ( .A1(n40435), .A2(n40434), .ZN(n40436) );
  INHSV2 U44929 ( .I(n40329), .ZN(n41328) );
  NAND2HSV2 U44930 ( .A1(n41225), .A2(n41328), .ZN(n40973) );
  NAND3HSV4 U44931 ( .A1(n59498), .A2(n40579), .A3(n40438), .ZN(n40442) );
  NOR2HSV4 U44932 ( .A1(n40479), .A2(n41230), .ZN(n40441) );
  CLKNAND2HSV2 U44933 ( .A1(n40477), .A2(n53650), .ZN(n40440) );
  NAND2HSV4 U44934 ( .A1(n40441), .A2(n40440), .ZN(n40634) );
  NAND2HSV2 U44935 ( .A1(n41230), .A2(\pe1/ti_7t [6]), .ZN(n40633) );
  NAND3HSV4 U44936 ( .A1(n40442), .A2(n40634), .A3(n40633), .ZN(n40474) );
  CLKNAND2HSV2 U44937 ( .A1(n40474), .A2(\pe1/got [31]), .ZN(n40471) );
  NOR2HSV2 U44938 ( .A1(n41333), .A2(n44337), .ZN(n40452) );
  NAND2HSV2 U44939 ( .A1(n40898), .A2(n53411), .ZN(n40444) );
  CLKNHSV0 U44940 ( .I(n40443), .ZN(n42139) );
  INHSV2 U44941 ( .I(n42264), .ZN(n53718) );
  NAND2HSV2 U44942 ( .A1(n42139), .A2(n53718), .ZN(n41253) );
  XOR2HSV0 U44943 ( .A1(n40444), .A2(n41253), .Z(n40450) );
  INHSV2 U44944 ( .I(n40445), .ZN(n40879) );
  CLKNAND2HSV1 U44945 ( .A1(n40879), .A2(n40557), .ZN(n40448) );
  INHSV2 U44946 ( .I(n48347), .ZN(n40608) );
  CLKNAND2HSV0 U44947 ( .A1(n40608), .A2(n40488), .ZN(n40447) );
  XOR2HSV0 U44948 ( .A1(n40448), .A2(n40447), .Z(n40449) );
  XNOR2HSV1 U44949 ( .A1(n40450), .A2(n40449), .ZN(n40451) );
  NAND2HSV2 U44950 ( .A1(n40876), .A2(n40494), .ZN(n40454) );
  CLKNAND2HSV0 U44951 ( .A1(\pe1/aot [25]), .A2(n40501), .ZN(n40453) );
  XOR2HSV0 U44952 ( .A1(n40454), .A2(n40453), .Z(n40459) );
  INHSV2 U44953 ( .I(n46629), .ZN(n53931) );
  INHSV2 U44954 ( .I(n40736), .ZN(n53526) );
  CLKNAND2HSV1 U44955 ( .A1(n53931), .A2(n53526), .ZN(n40457) );
  INHSV2 U44956 ( .I(n40455), .ZN(n40733) );
  CLKNAND2HSV0 U44957 ( .A1(n40683), .A2(n40733), .ZN(n40456) );
  XOR2HSV0 U44958 ( .A1(n40457), .A2(n40456), .Z(n40458) );
  XOR2HSV0 U44959 ( .A1(n40459), .A2(n40458), .Z(n40461) );
  BUFHSV2 U44960 ( .I(n41880), .Z(n40741) );
  INHSV4 U44961 ( .I(\pe1/got [26]), .ZN(n42086) );
  CLKNAND2HSV1 U44962 ( .A1(n40741), .A2(n40605), .ZN(n40460) );
  XNOR2HSV1 U44963 ( .A1(n40461), .A2(n40460), .ZN(n40462) );
  CLKXOR2HSV2 U44964 ( .A1(n40463), .A2(n40462), .Z(n40465) );
  INHSV2 U44965 ( .I(n48450), .ZN(n41731) );
  NAND2HSV2 U44966 ( .A1(n41422), .A2(n41731), .ZN(n40464) );
  XNOR2HSV4 U44967 ( .A1(n40465), .A2(n40464), .ZN(n40470) );
  INHSV2 U44968 ( .I(n40719), .ZN(n40636) );
  INHSV4 U44969 ( .I(n40466), .ZN(n40962) );
  INHSV2 U44970 ( .I(n40962), .ZN(n41410) );
  XNOR2HSV2 U44971 ( .A1(n40470), .A2(n40469), .ZN(n40472) );
  CLKNAND2HSV2 U44972 ( .A1(n40471), .A2(n40472), .ZN(n40476) );
  NOR2HSV4 U44973 ( .A1(n40472), .A2(n42070), .ZN(n40473) );
  INHSV2 U44974 ( .I(n59999), .ZN(n41234) );
  NAND2HSV4 U44975 ( .A1(n40477), .A2(n41234), .ZN(n40510) );
  NAND2HSV2 U44976 ( .A1(n41230), .A2(\pe1/ti_7t [5]), .ZN(n40509) );
  NAND2HSV4 U44977 ( .A1(n40510), .A2(n40509), .ZN(n40514) );
  INHSV4 U44978 ( .I(n40514), .ZN(n40678) );
  INHSV4 U44979 ( .I(n40678), .ZN(n53524) );
  XNOR2HSV4 U44980 ( .A1(n40478), .A2(n29639), .ZN(n40599) );
  INHSV2 U44981 ( .I(n40973), .ZN(n40580) );
  NAND2HSV2 U44982 ( .A1(n40479), .A2(n40580), .ZN(n40480) );
  INHSV2 U44983 ( .I(n40480), .ZN(n40481) );
  NAND2HSV4 U44984 ( .A1(n59498), .A2(n40481), .ZN(n40635) );
  INHSV2 U44985 ( .I(n41414), .ZN(n40482) );
  INHSV2 U44986 ( .I(n40483), .ZN(n40487) );
  CLKNHSV2 U44987 ( .I(n40579), .ZN(n46610) );
  INHSV2 U44988 ( .I(n40484), .ZN(n40485) );
  INHSV2 U44989 ( .I(n40580), .ZN(n44521) );
  INHSV2 U44990 ( .I(n48468), .ZN(n42328) );
  NOR2HSV4 U44991 ( .A1(n40485), .A2(n42328), .ZN(n40486) );
  CLKNAND2HSV4 U44992 ( .A1(n46610), .A2(n40486), .ZN(n40523) );
  INHSV1 U44993 ( .I(n40719), .ZN(n40822) );
  INHSV2 U44994 ( .I(n41074), .ZN(n59986) );
  NAND2HSV2 U44995 ( .A1(n53526), .A2(n59986), .ZN(n40490) );
  INHSV2 U44996 ( .I(n40455), .ZN(n40553) );
  XNOR2HSV4 U44997 ( .A1(n40490), .A2(n40489), .ZN(n40492) );
  BUFHSV2 U44998 ( .I(n41256), .Z(n41460) );
  NOR2HSV2 U44999 ( .A1(n41460), .A2(n40446), .ZN(n40788) );
  XNOR2HSV4 U45000 ( .A1(n40492), .A2(n40788), .ZN(n40498) );
  CLKNHSV0 U45001 ( .I(n40493), .ZN(n59591) );
  NAND2HSV2 U45002 ( .A1(n59591), .A2(n40557), .ZN(n40496) );
  CLKNAND2HSV0 U45003 ( .A1(n40568), .A2(n40494), .ZN(n40495) );
  XOR2HSV0 U45004 ( .A1(n40496), .A2(n40495), .Z(n40497) );
  XNOR2HSV4 U45005 ( .A1(n40498), .A2(n40497), .ZN(n40500) );
  NAND2HSV2 U45006 ( .A1(n40741), .A2(\pe1/got [27]), .ZN(n40499) );
  XNOR2HSV4 U45007 ( .A1(n40500), .A2(n40499), .ZN(n40502) );
  INHSV2 U45008 ( .I(n46629), .ZN(n54293) );
  NAND2HSV2 U45009 ( .A1(n54293), .A2(n40501), .ZN(n41270) );
  BUFHSV4 U45010 ( .I(n40786), .Z(n41422) );
  NAND2HSV4 U45011 ( .A1(n40700), .A2(n40781), .ZN(n40527) );
  INHSV2 U45012 ( .I(n42488), .ZN(n42344) );
  BUFHSV2 U45013 ( .I(n47935), .Z(n44522) );
  NAND2HSV2 U45014 ( .A1(n41238), .A2(\pe1/ti_7t [7]), .ZN(n40512) );
  INHSV2 U45015 ( .I(n40512), .ZN(n40542) );
  INHSV2 U45016 ( .I(n40542), .ZN(n40646) );
  OAI22HSV2 U45017 ( .A1(n40504), .A2(n40641), .B1(n44522), .B2(n40646), .ZN(
        n40519) );
  INHSV2 U45018 ( .I(n42196), .ZN(n59394) );
  NAND2HSV2 U45019 ( .A1(n29688), .A2(n40785), .ZN(n40544) );
  INHSV2 U45020 ( .I(n40544), .ZN(n40517) );
  AND2HSV2 U45021 ( .A1(n40512), .A2(n40668), .Z(n40513) );
  CLKNAND2HSV0 U45022 ( .A1(n40534), .A2(n40513), .ZN(n40515) );
  INHSV4 U45023 ( .I(n40514), .ZN(n46609) );
  NOR2HSV2 U45024 ( .A1(n40515), .A2(n46609), .ZN(n40516) );
  NOR2HSV2 U45025 ( .A1(n40517), .A2(n40516), .ZN(n40518) );
  OR2HSV1 U45026 ( .A1(n40633), .A2(n40520), .Z(n40521) );
  CLKNAND2HSV3 U45027 ( .A1(n40635), .A2(n40521), .ZN(n40522) );
  INHSV3 U45028 ( .I(n40522), .ZN(n40524) );
  NAND2HSV4 U45029 ( .A1(n40524), .A2(n40523), .ZN(n48007) );
  NOR2HSV2 U45030 ( .A1(n40526), .A2(n40668), .ZN(n40531) );
  NAND3HSV2 U45031 ( .A1(n40528), .A2(n42067), .A3(n40527), .ZN(n40529) );
  INHSV2 U45032 ( .I(n59999), .ZN(n41727) );
  CLKNAND2HSV1 U45033 ( .A1(n40529), .A2(n41727), .ZN(n40530) );
  NOR2HSV2 U45034 ( .A1(n40531), .A2(n40530), .ZN(n40532) );
  INHSV1 U45035 ( .I(n46609), .ZN(n40535) );
  INOR2HSV2 U45036 ( .A1(n40668), .B1(n40534), .ZN(n40546) );
  CLKNAND2HSV2 U45037 ( .A1(n40535), .A2(n40546), .ZN(n40536) );
  NAND2HSV4 U45038 ( .A1(n40538), .A2(n40648), .ZN(n40600) );
  INHSV2 U45039 ( .I(n40973), .ZN(n40972) );
  INHSV4 U45040 ( .I(n48007), .ZN(n40645) );
  NOR2HSV4 U45041 ( .A1(n40678), .A2(n42037), .ZN(n48006) );
  INHSV2 U45042 ( .I(n48006), .ZN(n40540) );
  INAND2HSV2 U45043 ( .A1(n40639), .B1(n40646), .ZN(n40539) );
  OAI22HSV2 U45044 ( .A1(n40645), .A2(n40542), .B1(n40540), .B2(n40539), .ZN(
        n40551) );
  NOR2HSV2 U45045 ( .A1(n29715), .A2(n48320), .ZN(n40543) );
  NAND2HSV2 U45046 ( .A1(n40544), .A2(n40543), .ZN(n40550) );
  NAND2HSV0 U45047 ( .A1(n40639), .A2(n40785), .ZN(n40545) );
  OA21HSV2 U45048 ( .A1(n40546), .A2(n40785), .B(n40545), .Z(n40549) );
  NOR2HSV2 U45049 ( .A1(n42070), .A2(n40962), .ZN(n40604) );
  NAND2HSV2 U45050 ( .A1(n48007), .A2(n40604), .ZN(n40548) );
  OAI22HSV4 U45051 ( .A1(n40551), .A2(n40550), .B1(n40549), .B2(n40548), .ZN(
        n40666) );
  BUFHSV2 U45052 ( .I(n40700), .Z(n41472) );
  BUFHSV2 U45053 ( .I(n41930), .Z(n40720) );
  CLKNAND2HSV3 U45054 ( .A1(n40720), .A2(n40923), .ZN(n40578) );
  NAND2HSV2 U45055 ( .A1(n53931), .A2(n53411), .ZN(n40555) );
  CLKNAND2HSV1 U45056 ( .A1(n40898), .A2(n40553), .ZN(n40554) );
  XOR2HSV0 U45057 ( .A1(n40555), .A2(n40554), .Z(n40562) );
  INHSV2 U45058 ( .I(n41870), .ZN(n40876) );
  CLKNAND2HSV1 U45059 ( .A1(n40876), .A2(n40557), .ZN(n40560) );
  NAND2HSV2 U45060 ( .A1(n54307), .A2(n40684), .ZN(n40559) );
  XOR2HSV0 U45061 ( .A1(n40560), .A2(n40559), .Z(n40561) );
  XOR2HSV0 U45062 ( .A1(n40562), .A2(n40561), .Z(n40576) );
  INHSV2 U45063 ( .I(\pe1/got [25]), .ZN(n41848) );
  INHSV2 U45064 ( .I(n41848), .ZN(n41201) );
  CLKNAND2HSV1 U45065 ( .A1(n40741), .A2(n41201), .ZN(n40566) );
  NOR2HSV2 U45066 ( .A1(n53447), .A2(n40446), .ZN(n40564) );
  CLKNAND2HSV1 U45067 ( .A1(n59385), .A2(n41771), .ZN(n40563) );
  XOR2HSV0 U45068 ( .A1(n40564), .A2(n40563), .Z(n40565) );
  XNOR2HSV1 U45069 ( .A1(n40566), .A2(n40565), .ZN(n40575) );
  INHSV2 U45070 ( .I(n40567), .ZN(n59590) );
  NAND2HSV2 U45071 ( .A1(n59590), .A2(n40605), .ZN(n40574) );
  INHSV2 U45072 ( .I(n54185), .ZN(n54318) );
  CLKNAND2HSV0 U45073 ( .A1(n54318), .A2(n40568), .ZN(n40613) );
  INHSV2 U45074 ( .I(n40569), .ZN(n44566) );
  OAI21HSV2 U45075 ( .A1(n41253), .A2(n40613), .B(n40570), .ZN(n40572) );
  CLKNAND2HSV1 U45076 ( .A1(n59589), .A2(n25179), .ZN(n40571) );
  XNOR2HSV1 U45077 ( .A1(n40572), .A2(n40571), .ZN(n40573) );
  XOR3HSV2 U45078 ( .A1(n40576), .A2(n40575), .A3(n29679), .Z(n40577) );
  NAND2HSV2 U45079 ( .A1(n40485), .A2(n40579), .ZN(n40582) );
  CLKNAND2HSV0 U45080 ( .A1(n40580), .A2(n40933), .ZN(n40581) );
  OAI22HSV2 U45081 ( .A1(n40582), .A2(n40581), .B1(n40936), .B2(n40633), .ZN(
        n40583) );
  INHSV2 U45082 ( .I(n40583), .ZN(n40586) );
  CLKNHSV2 U45083 ( .I(n40634), .ZN(n40584) );
  CLKNAND2HSV1 U45084 ( .A1(n40584), .A2(n59394), .ZN(n40585) );
  NAND2HSV2 U45085 ( .A1(n40586), .A2(n40585), .ZN(n40588) );
  INHSV2 U45086 ( .I(n40588), .ZN(n40589) );
  CLKNAND2HSV3 U45087 ( .A1(n40590), .A2(n40589), .ZN(n40591) );
  CLKNAND2HSV3 U45088 ( .A1(n40592), .A2(n40591), .ZN(n40665) );
  XNOR2HSV4 U45089 ( .A1(n40666), .A2(n40665), .ZN(n40657) );
  NOR2HSV4 U45090 ( .A1(n40673), .A2(n40657), .ZN(n40658) );
  AND2HSV2 U45091 ( .A1(n40671), .A2(n53367), .Z(n40593) );
  NOR2HSV4 U45092 ( .A1(n40658), .A2(n40593), .ZN(n40596) );
  NAND3HSV2 U45093 ( .A1(n40594), .A2(n40657), .A3(n40972), .ZN(n40595) );
  NAND2HSV4 U45094 ( .A1(n40596), .A2(n40595), .ZN(n40664) );
  INHSV2 U45095 ( .I(\pe1/ti_7t [8]), .ZN(n40597) );
  NOR2HSV4 U45096 ( .A1(n40598), .A2(n40597), .ZN(n40716) );
  CLKNAND2HSV2 U45097 ( .A1(n40599), .A2(n40600), .ZN(n40603) );
  CLKNAND2HSV4 U45098 ( .A1(n40602), .A2(n40603), .ZN(n40677) );
  INHSV2 U45099 ( .I(n40604), .ZN(n48324) );
  INHSV2 U45100 ( .I(n48324), .ZN(n42059) );
  AOI22HSV4 U45101 ( .A1(n53787), .A2(n40716), .B1(n40677), .B2(n42059), .ZN(
        n40653) );
  NAND2HSV2 U45102 ( .A1(n40720), .A2(n40605), .ZN(n40628) );
  CLKNAND2HSV1 U45103 ( .A1(n41145), .A2(n41644), .ZN(n40607) );
  CLKNAND2HSV0 U45104 ( .A1(n53931), .A2(n40733), .ZN(n40606) );
  XOR2HSV0 U45105 ( .A1(n40607), .A2(n40606), .Z(n40612) );
  CLKNAND2HSV1 U45106 ( .A1(n40898), .A2(n40608), .ZN(n40610) );
  INHSV2 U45107 ( .I(n46142), .ZN(n54288) );
  CLKNAND2HSV1 U45108 ( .A1(n54288), .A2(n40684), .ZN(n40609) );
  XOR2HSV0 U45109 ( .A1(n40610), .A2(n40609), .Z(n40611) );
  XOR2HSV0 U45110 ( .A1(n40612), .A2(n40611), .Z(n40619) );
  CLKNAND2HSV0 U45111 ( .A1(n59589), .A2(n53411), .ZN(n40789) );
  XOR2HSV0 U45112 ( .A1(n40613), .A2(n40789), .Z(n40617) );
  NAND2HSV0 U45113 ( .A1(n40683), .A2(n41771), .ZN(n40615) );
  INHSV2 U45114 ( .I(n42264), .ZN(n54319) );
  CLKNAND2HSV1 U45115 ( .A1(n40876), .A2(n54319), .ZN(n40614) );
  XOR2HSV0 U45116 ( .A1(n40615), .A2(n40614), .Z(n40616) );
  XOR2HSV0 U45117 ( .A1(n40617), .A2(n40616), .Z(n40618) );
  XOR2HSV0 U45118 ( .A1(n40619), .A2(n40618), .Z(n40626) );
  INHSV2 U45119 ( .I(\pe1/got [24]), .ZN(n41392) );
  INHSV2 U45120 ( .I(n41392), .ZN(n41143) );
  CLKNAND2HSV1 U45121 ( .A1(n40741), .A2(n41143), .ZN(n40622) );
  INHSV2 U45122 ( .I(\pe1/bq[23] ), .ZN(n41461) );
  INHSV2 U45123 ( .I(n41461), .ZN(n54048) );
  NAND2HSV2 U45124 ( .A1(\pe1/aot [24]), .A2(n54048), .ZN(n41082) );
  CLKNAND2HSV2 U45125 ( .A1(n25226), .A2(\pe1/bq[23] ), .ZN(n42214) );
  OAI21HSV1 U45126 ( .A1(n41952), .A2(n41974), .B(n42214), .ZN(n40620) );
  OAI21HSV0 U45127 ( .A1(n41082), .A2(n51112), .B(n40620), .ZN(n40621) );
  XOR2HSV0 U45128 ( .A1(n40622), .A2(n40621), .Z(n40624) );
  CLKNAND2HSV1 U45129 ( .A1(n59590), .A2(n41201), .ZN(n40623) );
  XOR2HSV0 U45130 ( .A1(n40624), .A2(n40623), .Z(n40625) );
  XNOR2HSV1 U45131 ( .A1(n40626), .A2(n40625), .ZN(n40627) );
  XNOR2HSV2 U45132 ( .A1(n40628), .A2(n40627), .ZN(n40630) );
  BUFHSV2 U45133 ( .I(n40700), .Z(n40910) );
  INHSV2 U45134 ( .I(n44337), .ZN(n40823) );
  XNOR2HSV4 U45135 ( .A1(n40632), .A2(n40631), .ZN(n40638) );
  NAND3HSV2 U45136 ( .A1(n40635), .A2(n40634), .A3(n40633), .ZN(n41017) );
  CLKBUFHSV4 U45137 ( .I(n41017), .Z(n40801) );
  NAND2HSV2 U45138 ( .A1(n40801), .A2(n40636), .ZN(n40637) );
  XNOR2HSV4 U45139 ( .A1(n40638), .A2(n40637), .ZN(n40651) );
  INHSV2 U45140 ( .I(n40639), .ZN(n48005) );
  CLKNAND2HSV2 U45141 ( .A1(n48006), .A2(n48005), .ZN(n40644) );
  NOR2HSV4 U45142 ( .A1(n40642), .A2(n40641), .ZN(n40643) );
  NAND3HSV3 U45143 ( .A1(n40645), .A2(n40644), .A3(n40643), .ZN(n40647) );
  NAND3HSV4 U45144 ( .A1(n40648), .A2(n40647), .A3(n40646), .ZN(n40757) );
  INHSV2 U45145 ( .I(n40649), .ZN(n40933) );
  XNOR2HSV4 U45146 ( .A1(n40651), .A2(n40650), .ZN(n40652) );
  XNOR2HSV4 U45147 ( .A1(n40653), .A2(n40652), .ZN(n40663) );
  XNOR2HSV4 U45148 ( .A1(n40664), .A2(n40663), .ZN(n40803) );
  INHSV2 U45149 ( .I(n40654), .ZN(n41242) );
  NAND2HSV2 U45150 ( .A1(n48331), .A2(\pe1/ti_7t [10]), .ZN(n40655) );
  OAI21HSV4 U45151 ( .A1(n40803), .A2(n41242), .B(n40655), .ZN(n40656) );
  INHSV4 U45152 ( .I(n40656), .ZN(n40821) );
  CLKNHSV6 U45153 ( .I(n40821), .ZN(n40928) );
  BUFHSV2 U45154 ( .I(n48450), .Z(n44528) );
  NAND2HSV0 U45155 ( .A1(n40928), .A2(n40873), .ZN(n40662) );
  INHSV2 U45156 ( .I(n25398), .ZN(n52736) );
  INHSV2 U45157 ( .I(n44649), .ZN(n41056) );
  NOR2HSV2 U45158 ( .A1(n40962), .A2(n53650), .ZN(n42478) );
  NOR2HSV2 U45159 ( .A1(n40669), .A2(n42478), .ZN(n40660) );
  NOR2HSV2 U45160 ( .A1(n40658), .A2(n40671), .ZN(n40659) );
  OAI21HSV4 U45161 ( .A1(n52736), .A2(n40660), .B(n40659), .ZN(n40874) );
  CLKNAND2HSV1 U45162 ( .A1(n29762), .A2(n40823), .ZN(n40661) );
  XNOR2HSV1 U45163 ( .A1(n40662), .A2(n40661), .ZN(n40819) );
  XNOR2HSV4 U45164 ( .A1(n40664), .A2(n40663), .ZN(n40771) );
  NOR2HSV4 U45165 ( .A1(n40771), .A2(n42328), .ZN(n40713) );
  NOR2HSV0 U45166 ( .A1(n40671), .A2(n42478), .ZN(n40667) );
  NAND2HSV2 U45167 ( .A1(n40672), .A2(n40667), .ZN(n40670) );
  OAI21HSV2 U45168 ( .A1(n40670), .A2(n40669), .B(n40668), .ZN(n40675) );
  NOR2HSV4 U45169 ( .A1(n40675), .A2(n40674), .ZN(n40807) );
  INHSV2 U45170 ( .I(n41331), .ZN(n53786) );
  NOR2HSV0 U45171 ( .A1(n40936), .A2(n41056), .ZN(n40676) );
  AOI22HSV2 U45172 ( .A1(n40716), .A2(n53786), .B1(n40677), .B2(n40676), .ZN(
        n40709) );
  AND2HSV2 U45173 ( .A1(n40757), .A2(n40822), .Z(n40707) );
  INHSV2 U45174 ( .I(n40678), .ZN(n40914) );
  CLKNAND2HSV3 U45175 ( .A1(n40914), .A2(n40923), .ZN(n40703) );
  NAND2HSV2 U45176 ( .A1(n40720), .A2(n41201), .ZN(n40699) );
  CLKNAND2HSV0 U45177 ( .A1(n59589), .A2(n40733), .ZN(n40680) );
  CLKNAND2HSV0 U45178 ( .A1(n40876), .A2(n54318), .ZN(n40679) );
  XOR2HSV0 U45179 ( .A1(n40680), .A2(n40679), .Z(n40693) );
  CLKNAND2HSV1 U45180 ( .A1(n54288), .A2(n54302), .ZN(n41364) );
  INHSV2 U45181 ( .I(n41947), .ZN(n40889) );
  CLKNAND2HSV1 U45182 ( .A1(n59591), .A2(n40889), .ZN(n41155) );
  OAI21HSV0 U45183 ( .A1(n46142), .A2(n41952), .B(n41155), .ZN(n40681) );
  OAI21HSV0 U45184 ( .A1(n41364), .A2(n51112), .B(n40681), .ZN(n40682) );
  NOR2HSV1 U45185 ( .A1(n40445), .A2(n41461), .ZN(n41738) );
  XNOR2HSV1 U45186 ( .A1(n40682), .A2(n41738), .ZN(n40692) );
  NAND2HSV0 U45187 ( .A1(n40683), .A2(n41644), .ZN(n40686) );
  CLKNAND2HSV0 U45188 ( .A1(\pe1/aot [22]), .A2(n40684), .ZN(n40685) );
  XOR2HSV0 U45189 ( .A1(n40686), .A2(n40685), .Z(n40690) );
  CLKNHSV2 U45190 ( .I(n40446), .ZN(n53922) );
  CLKNAND2HSV0 U45191 ( .A1(n53931), .A2(n53922), .ZN(n40688) );
  NAND2HSV0 U45192 ( .A1(n54307), .A2(n53411), .ZN(n40687) );
  XOR2HSV0 U45193 ( .A1(n40688), .A2(n40687), .Z(n40689) );
  XOR2HSV0 U45194 ( .A1(n40690), .A2(n40689), .Z(n40691) );
  XOR3HSV2 U45195 ( .A1(n40693), .A2(n40692), .A3(n40691), .Z(n40697) );
  INHSV2 U45196 ( .I(\pe1/got [23]), .ZN(n41926) );
  INHSV2 U45197 ( .I(n41926), .ZN(n41298) );
  CLKNAND2HSV0 U45198 ( .A1(n59590), .A2(n41143), .ZN(n40694) );
  XNOR2HSV1 U45199 ( .A1(n40695), .A2(n40694), .ZN(n40696) );
  XNOR2HSV1 U45200 ( .A1(n40697), .A2(n40696), .ZN(n40698) );
  XNOR2HSV1 U45201 ( .A1(n40699), .A2(n40698), .ZN(n40702) );
  BUFHSV2 U45202 ( .I(n40700), .Z(n59674) );
  NAND2HSV2 U45203 ( .A1(n40801), .A2(n40873), .ZN(n40704) );
  XNOR2HSV4 U45204 ( .A1(n40707), .A2(n40706), .ZN(n40708) );
  XNOR2HSV4 U45205 ( .A1(n40709), .A2(n40708), .ZN(n40806) );
  NAND2HSV2 U45206 ( .A1(n40807), .A2(n40806), .ZN(n40712) );
  INHSV4 U45207 ( .I(n40807), .ZN(n40808) );
  INHSV2 U45208 ( .I(n40806), .ZN(n40710) );
  CLKNAND2HSV3 U45209 ( .A1(n40710), .A2(n40808), .ZN(n40711) );
  BUFHSV2 U45210 ( .I(n41134), .Z(n41217) );
  INHSV1 U45211 ( .I(n40809), .ZN(n40714) );
  CLKNAND2HSV3 U45212 ( .A1(n40715), .A2(n51114), .ZN(n40764) );
  INHSV2 U45213 ( .I(n40716), .ZN(n40717) );
  NAND2HSV4 U45214 ( .A1(n40718), .A2(n40717), .ZN(n47999) );
  INAND2HSV2 U45215 ( .A1(n40719), .B1(n47999), .ZN(n40761) );
  NAND2HSV2 U45216 ( .A1(n40914), .A2(n41689), .ZN(n40754) );
  NAND2HSV2 U45217 ( .A1(n40720), .A2(n41143), .ZN(n40750) );
  NAND2HSV2 U45218 ( .A1(n41160), .A2(n41298), .ZN(n40724) );
  NAND2HSV0 U45219 ( .A1(n54288), .A2(n53411), .ZN(n40722) );
  INHSV2 U45220 ( .I(n41944), .ZN(n54663) );
  NAND2HSV2 U45221 ( .A1(n54663), .A2(n40890), .ZN(n40721) );
  XOR2HSV0 U45222 ( .A1(n40722), .A2(n40721), .Z(n40723) );
  XNOR2HSV1 U45223 ( .A1(n40724), .A2(n40723), .ZN(n40732) );
  BUFHSV2 U45224 ( .I(n41461), .Z(n53819) );
  NOR2HSV2 U45225 ( .A1(n41256), .A2(n53819), .ZN(n40726) );
  NAND2HSV0 U45226 ( .A1(n54293), .A2(n41771), .ZN(n40725) );
  XOR2HSV0 U45227 ( .A1(n40726), .A2(n40725), .Z(n40730) );
  CLKNAND2HSV0 U45228 ( .A1(n59589), .A2(n53922), .ZN(n40728) );
  NAND2HSV0 U45229 ( .A1(n40683), .A2(n53718), .ZN(n40727) );
  XOR2HSV0 U45230 ( .A1(n40728), .A2(n40727), .Z(n40729) );
  XOR2HSV0 U45231 ( .A1(n40730), .A2(n40729), .Z(n40731) );
  XNOR2HSV1 U45232 ( .A1(n40732), .A2(n40731), .ZN(n40748) );
  NAND2HSV0 U45233 ( .A1(n54307), .A2(n40733), .ZN(n40735) );
  CLKNAND2HSV0 U45234 ( .A1(n59385), .A2(n54318), .ZN(n40734) );
  XOR2HSV0 U45235 ( .A1(n40735), .A2(n40734), .Z(n40740) );
  CLKBUFHSV2 U45236 ( .I(n41952), .Z(n41453) );
  INHSV2 U45237 ( .I(n41453), .ZN(n40897) );
  NAND2HSV2 U45238 ( .A1(n54078), .A2(n40897), .ZN(n40738) );
  NAND2HSV0 U45239 ( .A1(n40898), .A2(n41644), .ZN(n40737) );
  XOR2HSV0 U45240 ( .A1(n40738), .A2(n40737), .Z(n40739) );
  XOR2HSV0 U45241 ( .A1(n40740), .A2(n40739), .Z(n40746) );
  INHSV2 U45242 ( .I(n42209), .ZN(n40875) );
  CLKNAND2HSV0 U45243 ( .A1(n40741), .A2(n40875), .ZN(n40744) );
  INHSV2 U45244 ( .I(\pe1/bq[21] ), .ZN(n44703) );
  CLKNAND2HSV0 U45245 ( .A1(n40879), .A2(\pe1/bq[21] ), .ZN(n40828) );
  BUFHSV2 U45246 ( .I(n41947), .Z(n48393) );
  NAND2HSV0 U45247 ( .A1(n59591), .A2(\pe1/bq[21] ), .ZN(n41077) );
  OAI21HSV0 U45248 ( .A1(n48393), .A2(n40445), .B(n41077), .ZN(n40742) );
  OAI21HSV1 U45249 ( .A1(n40828), .A2(n41155), .B(n40742), .ZN(n40743) );
  XOR2HSV0 U45250 ( .A1(n40744), .A2(n40743), .Z(n40745) );
  XOR2HSV0 U45251 ( .A1(n40746), .A2(n40745), .Z(n40747) );
  XNOR2HSV1 U45252 ( .A1(n40748), .A2(n40747), .ZN(n40749) );
  XNOR2HSV2 U45253 ( .A1(n40750), .A2(n40749), .ZN(n40752) );
  BUFHSV2 U45254 ( .I(n41472), .Z(n41287) );
  NAND2HSV2 U45255 ( .A1(n41287), .A2(\pe1/got [25]), .ZN(n40751) );
  XNOR2HSV1 U45256 ( .A1(n40752), .A2(n40751), .ZN(n40753) );
  XNOR2HSV2 U45257 ( .A1(n40754), .A2(n40753), .ZN(n40756) );
  NAND2HSV2 U45258 ( .A1(n40917), .A2(n40923), .ZN(n40755) );
  INHSV2 U45259 ( .I(n40757), .ZN(n41893) );
  INHSV2 U45260 ( .I(n41893), .ZN(n40920) );
  CLKNAND2HSV1 U45261 ( .A1(n40920), .A2(n40873), .ZN(n40758) );
  XNOR2HSV4 U45262 ( .A1(n40761), .A2(n40760), .ZN(n40763) );
  CLKNAND2HSV2 U45263 ( .A1(n40874), .A2(n40933), .ZN(n40762) );
  XNOR2HSV4 U45264 ( .A1(n40763), .A2(n40762), .ZN(n47987) );
  XNOR2HSV4 U45265 ( .A1(n40764), .A2(n47987), .ZN(n40860) );
  INHSV2 U45266 ( .I(n40767), .ZN(n40858) );
  INHSV4 U45267 ( .I(n40928), .ZN(n40766) );
  OR2HSV1 U45268 ( .A1(n41056), .A2(n48320), .Z(n40765) );
  NOR2HSV4 U45269 ( .A1(n40766), .A2(n40765), .ZN(n40859) );
  NOR2HSV4 U45270 ( .A1(n40859), .A2(n40767), .ZN(n40943) );
  CLKNHSV2 U45271 ( .I(n40943), .ZN(n40768) );
  CLKNAND2HSV2 U45272 ( .A1(n40768), .A2(n40781), .ZN(n40769) );
  AOI21HSV4 U45273 ( .A1(n40941), .A2(n40858), .B(n40769), .ZN(n40784) );
  NAND2HSV0 U45274 ( .A1(n40809), .A2(n53650), .ZN(n40770) );
  CLKAND2HSV2 U45275 ( .A1(n40810), .A2(n40770), .Z(n40778) );
  NOR2HSV2 U45276 ( .A1(n40805), .A2(n44521), .ZN(n40773) );
  CLKNHSV0 U45277 ( .I(n40771), .ZN(n60008) );
  INHSV2 U45278 ( .I(n60008), .ZN(n40772) );
  CLKNAND2HSV1 U45279 ( .A1(n40773), .A2(n40772), .ZN(n40776) );
  NAND3HSV2 U45280 ( .A1(n40778), .A2(n40777), .A3(n40776), .ZN(n40779) );
  NAND2HSV4 U45281 ( .A1(n40780), .A2(n40779), .ZN(n40942) );
  NAND3HSV3 U45282 ( .A1(n40942), .A2(n29653), .A3(n40781), .ZN(n40782) );
  INHSV4 U45283 ( .I(n40782), .ZN(n40783) );
  NOR2HSV4 U45284 ( .A1(n40784), .A2(n40783), .ZN(n40818) );
  BUFHSV2 U45285 ( .I(n47999), .Z(n41929) );
  INHSV2 U45286 ( .I(\pe1/got [21]), .ZN(n48337) );
  INHSV2 U45287 ( .I(n48337), .ZN(n40886) );
  NOR2HSV2 U45288 ( .A1(n53957), .A2(n44703), .ZN(n40827) );
  INHSV2 U45289 ( .I(\pe1/bq[18] ), .ZN(n41512) );
  NAND2HSV0 U45290 ( .A1(n40898), .A2(\pe1/bq[18] ), .ZN(n41363) );
  NAND2HSV0 U45291 ( .A1(n40879), .A2(n42092), .ZN(n53671) );
  INHSV2 U45292 ( .I(n44705), .ZN(n42099) );
  NOR2HSV2 U45293 ( .A1(n41885), .A2(n48060), .ZN(n41763) );
  CLKNAND2HSV0 U45294 ( .A1(n54669), .A2(n41173), .ZN(n41352) );
  NAND2HSV0 U45295 ( .A1(\pe1/aot [25]), .A2(n41173), .ZN(n40984) );
  INHSV2 U45296 ( .I(n41333), .ZN(n41248) );
  NOR2HSV0 U45297 ( .A1(n53447), .A2(n48393), .ZN(n40793) );
  INHSV2 U45298 ( .I(n54185), .ZN(n40982) );
  NAND2HSV0 U45299 ( .A1(\pe1/aot [26]), .A2(n40982), .ZN(n40792) );
  XOR2HSV0 U45300 ( .A1(n40793), .A2(n40792), .Z(n40796) );
  CLKNAND2HSV1 U45301 ( .A1(n40733), .A2(n59987), .ZN(n40795) );
  CLKNHSV0 U45302 ( .I(n46142), .ZN(n40996) );
  CLKNAND2HSV0 U45303 ( .A1(n40996), .A2(n41771), .ZN(n40794) );
  CLKNAND2HSV0 U45304 ( .A1(\pe1/aot [24]), .A2(n41644), .ZN(n40798) );
  INHSV2 U45305 ( .I(n41931), .ZN(n54916) );
  CLKNAND2HSV1 U45306 ( .A1(n54916), .A2(n41083), .ZN(n40797) );
  XOR2HSV0 U45307 ( .A1(n40798), .A2(n40797), .Z(n40800) );
  BUFHSV2 U45308 ( .I(n41880), .Z(n41752) );
  CLKBUFHSV2 U45309 ( .I(n41752), .Z(n41152) );
  INHSV2 U45310 ( .I(n41928), .ZN(n41188) );
  CLKNAND2HSV1 U45311 ( .A1(n41152), .A2(n41188), .ZN(n40799) );
  INHSV2 U45312 ( .I(n42209), .ZN(n41387) );
  BUFHSV2 U45313 ( .I(n40801), .Z(n40917) );
  INHSV2 U45314 ( .I(n41392), .ZN(n40913) );
  INHSV2 U45315 ( .I(n41893), .ZN(n42431) );
  CLKNHSV0 U45316 ( .I(n40814), .ZN(n40802) );
  NOR2HSV2 U45317 ( .A1(n40802), .A2(n40719), .ZN(n40816) );
  CLKNAND2HSV1 U45318 ( .A1(n40803), .A2(n41129), .ZN(n40804) );
  MUX2NHSV1 U45319 ( .I0(n40808), .I1(n40807), .S(n40806), .ZN(n52743) );
  BUFHSV2 U45320 ( .I(n42478), .Z(n48471) );
  AOI21HSV2 U45321 ( .A1(n52743), .A2(n48471), .B(n40809), .ZN(n40811) );
  INHSV6 U45322 ( .I(n41391), .ZN(n40820) );
  INHSV6 U45323 ( .I(n40820), .ZN(n54683) );
  AOI21HSV2 U45324 ( .A1(n59934), .A2(n42084), .B(n40814), .ZN(n40815) );
  XOR3HSV2 U45325 ( .A1(n40819), .A2(n40818), .A3(n40817), .Z(n40872) );
  CLKNHSV6 U45326 ( .I(n40820), .ZN(n54732) );
  INHSV4 U45327 ( .I(n40821), .ZN(n41026) );
  INHSV1 U45328 ( .I(n40936), .ZN(n41319) );
  CLKNAND2HSV4 U45329 ( .A1(n41026), .A2(n41319), .ZN(n40856) );
  NAND2HSV2 U45330 ( .A1(n40874), .A2(n40822), .ZN(n40855) );
  CLKNAND2HSV1 U45331 ( .A1(n40920), .A2(n40823), .ZN(n40853) );
  NAND2HSV2 U45332 ( .A1(n40914), .A2(\pe1/got [25]), .ZN(n40848) );
  NAND2HSV2 U45333 ( .A1(n41549), .A2(\pe1/got [23]), .ZN(n40844) );
  NAND2HSV2 U45334 ( .A1(n41169), .A2(n53411), .ZN(n41761) );
  NAND2HSV0 U45335 ( .A1(n59589), .A2(n41771), .ZN(n54084) );
  XOR2HSV0 U45336 ( .A1(n41761), .A2(n54084), .Z(n40826) );
  CLKNHSV1 U45337 ( .I(n41870), .ZN(n41358) );
  NAND2HSV2 U45338 ( .A1(n41358), .A2(n40889), .ZN(n41258) );
  NAND2HSV0 U45339 ( .A1(n40898), .A2(n53718), .ZN(n40824) );
  XOR2HSV0 U45340 ( .A1(n41258), .A2(n40824), .Z(n40825) );
  XOR2HSV0 U45341 ( .A1(n40826), .A2(n40825), .Z(n40842) );
  CLKNAND2HSV1 U45342 ( .A1(n40683), .A2(n40982), .ZN(n41260) );
  CLKNHSV0 U45343 ( .I(\pe1/bq[28] ), .ZN(n48347) );
  NOR2HSV2 U45344 ( .A1(n41974), .A2(n48347), .ZN(n40830) );
  CLKNAND2HSV0 U45345 ( .A1(\pe1/aot [26]), .A2(n41644), .ZN(n40829) );
  XOR2HSV0 U45346 ( .A1(n40830), .A2(n40829), .Z(n40834) );
  NAND2HSV2 U45347 ( .A1(n40733), .A2(n40996), .ZN(n40832) );
  CLKNAND2HSV1 U45348 ( .A1(n54669), .A2(n40890), .ZN(n40831) );
  XOR2HSV0 U45349 ( .A1(n40832), .A2(n40831), .Z(n40833) );
  XOR2HSV0 U45350 ( .A1(n40834), .A2(n40833), .Z(n40839) );
  NAND2HSV2 U45351 ( .A1(n41152), .A2(n40886), .ZN(n40837) );
  CLKNAND2HSV1 U45352 ( .A1(n59987), .A2(n41760), .ZN(n41874) );
  NAND2HSV0 U45353 ( .A1(n42139), .A2(\pe1/bq[20] ), .ZN(n41617) );
  OAI21HSV0 U45354 ( .A1(n41952), .A2(n41944), .B(n41617), .ZN(n40835) );
  OAI21HSV0 U45355 ( .A1(n51112), .A2(n41874), .B(n40835), .ZN(n40836) );
  XOR2HSV0 U45356 ( .A1(n40837), .A2(n40836), .Z(n40838) );
  XOR2HSV0 U45357 ( .A1(n40839), .A2(n40838), .Z(n40840) );
  XOR3HSV2 U45358 ( .A1(n40842), .A2(n40841), .A3(n40840), .Z(n40843) );
  XNOR2HSV1 U45359 ( .A1(n40844), .A2(n40843), .ZN(n40846) );
  NAND2HSV2 U45360 ( .A1(n40910), .A2(n40913), .ZN(n40845) );
  XNOR2HSV1 U45361 ( .A1(n40846), .A2(n40845), .ZN(n40847) );
  CLKNAND2HSV1 U45362 ( .A1(n40917), .A2(n41689), .ZN(n40849) );
  XOR2HSV0 U45363 ( .A1(n40850), .A2(n40849), .Z(n40852) );
  CLKNAND2HSV2 U45364 ( .A1(n47999), .A2(n40873), .ZN(n40851) );
  XOR3HSV2 U45365 ( .A1(n40853), .A2(n40852), .A3(n40851), .Z(n40854) );
  XOR2HSV4 U45366 ( .A1(n40856), .A2(n29692), .Z(n40857) );
  AOI21HSV4 U45367 ( .A1(n54732), .A2(n40957), .B(n40857), .ZN(n40865) );
  INHSV4 U45368 ( .I(n40865), .ZN(n40949) );
  BUFHSV2 U45369 ( .I(n53649), .Z(n40975) );
  NAND3HSV3 U45370 ( .A1(n40857), .A2(n54732), .A3(n40975), .ZN(n40948) );
  NAND2HSV4 U45371 ( .A1(n40949), .A2(n40948), .ZN(n40955) );
  CLKNHSV2 U45372 ( .I(n40955), .ZN(n40870) );
  INHSV2 U45373 ( .I(n40858), .ZN(n40939) );
  AOI21HSV4 U45374 ( .A1(n40860), .A2(n40859), .B(n40939), .ZN(n40862) );
  CLKNAND2HSV4 U45375 ( .A1(n40862), .A2(n40861), .ZN(n41061) );
  CLKNHSV0 U45376 ( .I(n40973), .ZN(n42484) );
  CLKBUFHSV4 U45377 ( .I(n41061), .Z(n41142) );
  CLKNAND2HSV1 U45378 ( .A1(n41229), .A2(n42471), .ZN(n40864) );
  INHSV2 U45379 ( .I(n40864), .ZN(n40863) );
  CLKNAND2HSV2 U45380 ( .A1(n40948), .A2(n40863), .ZN(n40866) );
  AOI21HSV4 U45381 ( .A1(n40870), .A2(n29648), .B(n40869), .ZN(n40871) );
  XNOR2HSV4 U45382 ( .A1(n40872), .A2(n40871), .ZN(n52762) );
  INHSV4 U45383 ( .I(n54683), .ZN(n47984) );
  CLKAND2HSV2 U45384 ( .A1(n40874), .A2(n40873), .Z(n40927) );
  CLKNAND2HSV1 U45385 ( .A1(n41549), .A2(n40875), .ZN(n40909) );
  CLKNAND2HSV0 U45386 ( .A1(n40876), .A2(\pe1/bq[21] ), .ZN(n40878) );
  CLKNAND2HSV1 U45387 ( .A1(n59987), .A2(n53411), .ZN(n40877) );
  XOR2HSV0 U45388 ( .A1(n40878), .A2(n40877), .Z(n40882) );
  CLKNAND2HSV0 U45389 ( .A1(n40879), .A2(n42238), .ZN(n41075) );
  CLKNAND2HSV0 U45390 ( .A1(n40683), .A2(n54048), .ZN(n40880) );
  XOR2HSV0 U45391 ( .A1(n41075), .A2(n40880), .Z(n40881) );
  XOR2HSV0 U45392 ( .A1(n40882), .A2(n40881), .Z(n40907) );
  CLKNAND2HSV1 U45393 ( .A1(n41752), .A2(\pe1/got [20]), .ZN(n40885) );
  CLKNAND2HSV0 U45394 ( .A1(\pe1/aot [26]), .A2(\pe1/bq[19] ), .ZN(n41351) );
  OAI22HSV2 U45395 ( .A1(n41076), .A2(n41963), .B1(n46629), .B2(n42264), .ZN(
        n40883) );
  OAI21HSV0 U45396 ( .A1(n41351), .A2(n41253), .B(n40883), .ZN(n40884) );
  XOR2HSV0 U45397 ( .A1(n40885), .A2(n40884), .Z(n40888) );
  CLKNAND2HSV1 U45398 ( .A1(n41248), .A2(n40886), .ZN(n40887) );
  INHSV2 U45399 ( .I(n44705), .ZN(n54824) );
  NAND2HSV0 U45400 ( .A1(\pe1/aot [24]), .A2(n41771), .ZN(n40892) );
  CLKNAND2HSV0 U45401 ( .A1(n41169), .A2(n42125), .ZN(n40891) );
  XOR2HSV0 U45402 ( .A1(n40892), .A2(n40891), .Z(n40893) );
  XOR2HSV0 U45403 ( .A1(n40894), .A2(n40893), .Z(n40904) );
  NOR2HSV0 U45404 ( .A1(n46142), .A2(n48347), .ZN(n40896) );
  NAND2HSV0 U45405 ( .A1(n59589), .A2(n41644), .ZN(n40895) );
  XOR2HSV0 U45406 ( .A1(n40896), .A2(n40895), .Z(n40902) );
  CLKNAND2HSV1 U45407 ( .A1(n54669), .A2(n40897), .ZN(n40900) );
  NAND2HSV0 U45408 ( .A1(n40898), .A2(n54318), .ZN(n40899) );
  XOR2HSV0 U45409 ( .A1(n40900), .A2(n40899), .Z(n40901) );
  XOR2HSV0 U45410 ( .A1(n40902), .A2(n40901), .Z(n40903) );
  XOR2HSV0 U45411 ( .A1(n40904), .A2(n40903), .Z(n40905) );
  XOR3HSV2 U45412 ( .A1(n40907), .A2(n40906), .A3(n40905), .Z(n40908) );
  XNOR2HSV1 U45413 ( .A1(n40909), .A2(n40908), .ZN(n40912) );
  NAND2HSV2 U45414 ( .A1(n40910), .A2(n41298), .ZN(n40911) );
  XNOR2HSV1 U45415 ( .A1(n40912), .A2(n40911), .ZN(n40916) );
  NAND2HSV2 U45416 ( .A1(n40914), .A2(n40913), .ZN(n40915) );
  XNOR2HSV1 U45417 ( .A1(n40916), .A2(n40915), .ZN(n40919) );
  CLKNAND2HSV1 U45418 ( .A1(n40917), .A2(\pe1/got [25]), .ZN(n40918) );
  XNOR2HSV1 U45419 ( .A1(n40919), .A2(n40918), .ZN(n40922) );
  CLKNAND2HSV1 U45420 ( .A1(n40920), .A2(n41689), .ZN(n40921) );
  XNOR2HSV1 U45421 ( .A1(n40922), .A2(n40921), .ZN(n40925) );
  CLKNAND2HSV2 U45422 ( .A1(n47999), .A2(n40923), .ZN(n40924) );
  XNOR2HSV4 U45423 ( .A1(n40925), .A2(n40924), .ZN(n40926) );
  XNOR2HSV4 U45424 ( .A1(n40927), .A2(n40926), .ZN(n40930) );
  NOR2HSV2 U45425 ( .A1(n40930), .A2(n40719), .ZN(n40929) );
  AOI22HSV2 U45426 ( .A1(n40930), .A2(n40719), .B1(n40929), .B2(n40928), .ZN(
        n40932) );
  INAND2HSV1 U45427 ( .A1(n41026), .B1(n40930), .ZN(n40931) );
  NAND2HSV2 U45428 ( .A1(n40932), .A2(n40931), .ZN(n40934) );
  INHSV2 U45429 ( .I(n40934), .ZN(n40935) );
  OAI21HSV4 U45430 ( .A1(n47984), .A2(n40936), .B(n40935), .ZN(n40937) );
  OAI21HSV4 U45431 ( .A1(n47984), .A2(n40938), .B(n40937), .ZN(n40960) );
  NOR2HSV4 U45432 ( .A1(n29653), .A2(n40939), .ZN(n40940) );
  INHSV4 U45433 ( .I(n40942), .ZN(n40944) );
  NAND2HSV4 U45434 ( .A1(n40944), .A2(n40943), .ZN(n40947) );
  INHSV2 U45435 ( .I(n41701), .ZN(n53649) );
  NAND3HSV3 U45436 ( .A1(n40946), .A2(n40947), .A3(n53649), .ZN(n40945) );
  NOR2HSV4 U45437 ( .A1(n40954), .A2(n40366), .ZN(n40951) );
  NAND2HSV2 U45438 ( .A1(n40949), .A2(n40948), .ZN(n40950) );
  XNOR2HSV4 U45439 ( .A1(n40951), .A2(n40950), .ZN(n59576) );
  NAND3HSV4 U45440 ( .A1(n52763), .A2(n59576), .A3(n40972), .ZN(n41115) );
  CLKNAND2HSV0 U45441 ( .A1(n41115), .A2(n40952), .ZN(n40953) );
  NOR2HSV4 U45442 ( .A1(n52762), .A2(n40953), .ZN(n40966) );
  XNOR2HSV4 U45443 ( .A1(n40955), .A2(n40954), .ZN(n41111) );
  CLKNAND2HSV2 U45444 ( .A1(n41111), .A2(n40438), .ZN(n40967) );
  INHSV2 U45445 ( .I(n42478), .ZN(n41919) );
  NOR2HSV4 U45446 ( .A1(n41142), .A2(n41919), .ZN(n40956) );
  INHSV2 U45447 ( .I(n40960), .ZN(n40964) );
  NAND2HSV0 U45448 ( .A1(n48471), .A2(n40957), .ZN(n42315) );
  CLKNHSV0 U45449 ( .I(n42315), .ZN(n40958) );
  AND2HSV2 U45450 ( .A1(n42478), .A2(n42070), .Z(n40963) );
  INHSV2 U45451 ( .I(n47935), .ZN(n51114) );
  INHSV2 U45452 ( .I(n52760), .ZN(n40965) );
  NAND2HSV4 U45453 ( .A1(n40966), .A2(n40965), .ZN(n41051) );
  INHSV2 U45454 ( .I(n41115), .ZN(n52761) );
  NAND2HSV2 U45455 ( .A1(n52762), .A2(n52761), .ZN(n41050) );
  NOR2HSV0 U45456 ( .A1(n26381), .A2(n40967), .ZN(n40968) );
  NAND2HSV2 U45457 ( .A1(n52762), .A2(n40968), .ZN(n41053) );
  NAND2HSV2 U45458 ( .A1(n41720), .A2(\pe1/ti_7t [15]), .ZN(n41052) );
  CLKNAND2HSV4 U45459 ( .A1(n41053), .A2(n41052), .ZN(n40970) );
  NOR2HSV8 U45460 ( .A1(n40971), .A2(n40970), .ZN(n41421) );
  INHSV2 U45461 ( .I(\pe1/got [31]), .ZN(n42037) );
  NOR2HSV0 U45462 ( .A1(n40973), .A2(n42037), .ZN(n48312) );
  NAND3HSV2 U45463 ( .A1(n52763), .A2(n59576), .A3(n48312), .ZN(n40974) );
  INHSV2 U45464 ( .I(n40974), .ZN(n41043) );
  CLKNAND2HSV2 U45465 ( .A1(n41111), .A2(n42059), .ZN(n41034) );
  NOR2HSV0 U45466 ( .A1(n41034), .A2(n52763), .ZN(n41033) );
  NAND2HSV4 U45467 ( .A1(n41117), .A2(n40975), .ZN(n41038) );
  CLKNAND2HSV0 U45468 ( .A1(n41929), .A2(n41201), .ZN(n41023) );
  CLKNAND2HSV0 U45469 ( .A1(n41144), .A2(n41387), .ZN(n41016) );
  NAND2HSV0 U45470 ( .A1(n41549), .A2(n44530), .ZN(n41012) );
  NOR2HSV0 U45471 ( .A1(n41944), .A2(n48347), .ZN(n40977) );
  INHSV2 U45472 ( .I(n44705), .ZN(n41736) );
  NAND2HSV0 U45473 ( .A1(n41736), .A2(n53411), .ZN(n40976) );
  XOR2HSV0 U45474 ( .A1(n40977), .A2(n40976), .Z(n40981) );
  NAND2HSV0 U45475 ( .A1(n42139), .A2(\pe1/bq[17] ), .ZN(n40979) );
  CLKNHSV0 U45476 ( .I(n40445), .ZN(n42412) );
  CLKNAND2HSV0 U45477 ( .A1(n42412), .A2(\pe1/bq[18] ), .ZN(n40978) );
  XOR2HSV0 U45478 ( .A1(n40979), .A2(n40978), .Z(n40980) );
  XOR2HSV0 U45479 ( .A1(n40981), .A2(n40980), .Z(n40988) );
  CLKNAND2HSV0 U45480 ( .A1(n41152), .A2(\pe1/got [18]), .ZN(n40986) );
  NAND2HSV0 U45481 ( .A1(\pe1/aot [24]), .A2(n40982), .ZN(n41163) );
  CLKNHSV0 U45482 ( .I(n54185), .ZN(n41355) );
  CLKNAND2HSV1 U45483 ( .A1(\pe1/aot [25]), .A2(n41355), .ZN(n54187) );
  OAI21HSV0 U45484 ( .A1(n41974), .A2(n42264), .B(n54187), .ZN(n40983) );
  OAI21HSV0 U45485 ( .A1(n40984), .A2(n41163), .B(n40983), .ZN(n40985) );
  XOR2HSV0 U45486 ( .A1(n40986), .A2(n40985), .Z(n40987) );
  XNOR2HSV1 U45487 ( .A1(n40988), .A2(n40987), .ZN(n40993) );
  CLKNAND2HSV0 U45488 ( .A1(n41160), .A2(n41188), .ZN(n40991) );
  NAND2HSV2 U45489 ( .A1(n41145), .A2(n41760), .ZN(n53663) );
  CLKNAND2HSV1 U45490 ( .A1(n40898), .A2(n54302), .ZN(n40989) );
  XOR2HSV0 U45491 ( .A1(n53663), .A2(n40989), .Z(n40990) );
  XOR2HSV0 U45492 ( .A1(n40991), .A2(n40990), .Z(n40992) );
  XNOR2HSV1 U45493 ( .A1(n40993), .A2(n40992), .ZN(n41010) );
  NAND2HSV0 U45494 ( .A1(n41169), .A2(n41771), .ZN(n40995) );
  NAND2HSV0 U45495 ( .A1(\pe1/aot [20]), .A2(n42223), .ZN(n40994) );
  XOR2HSV0 U45496 ( .A1(n40995), .A2(n40994), .Z(n41000) );
  CLKNAND2HSV0 U45497 ( .A1(n41153), .A2(\pe1/bq[23] ), .ZN(n40998) );
  NAND2HSV0 U45498 ( .A1(n40996), .A2(n41644), .ZN(n40997) );
  XOR2HSV0 U45499 ( .A1(n40998), .A2(n40997), .Z(n40999) );
  XOR2HSV0 U45500 ( .A1(n41000), .A2(n40999), .Z(n41008) );
  NOR2HSV0 U45501 ( .A1(n41870), .A2(n41963), .ZN(n41002) );
  CLKNHSV0 U45502 ( .I(n41453), .ZN(n41170) );
  CLKNAND2HSV0 U45503 ( .A1(n54916), .A2(n41170), .ZN(n41001) );
  XOR2HSV0 U45504 ( .A1(n41002), .A2(n41001), .Z(n41006) );
  NAND2HSV0 U45505 ( .A1(n40683), .A2(\pe1/bq[21] ), .ZN(n41004) );
  CLKNAND2HSV0 U45506 ( .A1(\pe1/aot [17]), .A2(n41083), .ZN(n41003) );
  XOR2HSV0 U45507 ( .A1(n41004), .A2(n41003), .Z(n41005) );
  XOR2HSV0 U45508 ( .A1(n41006), .A2(n41005), .Z(n41007) );
  XOR2HSV0 U45509 ( .A1(n41008), .A2(n41007), .Z(n41009) );
  XNOR2HSV1 U45510 ( .A1(n41010), .A2(n41009), .ZN(n41011) );
  XNOR2HSV1 U45511 ( .A1(n41012), .A2(n41011), .ZN(n41014) );
  NAND2HSV2 U45512 ( .A1(n41472), .A2(n54724), .ZN(n41013) );
  XNOR2HSV1 U45513 ( .A1(n41014), .A2(n41013), .ZN(n41015) );
  XNOR2HSV1 U45514 ( .A1(n41016), .A2(n41015), .ZN(n41019) );
  BUFHSV2 U45515 ( .I(n41017), .Z(n59686) );
  BUFHSV2 U45516 ( .I(n59686), .Z(n41557) );
  CLKNAND2HSV1 U45517 ( .A1(n41557), .A2(\pe1/got [23]), .ZN(n41018) );
  XOR2HSV0 U45518 ( .A1(n41019), .A2(n41018), .Z(n41021) );
  NAND2HSV0 U45519 ( .A1(n42431), .A2(n41143), .ZN(n41020) );
  XOR2HSV0 U45520 ( .A1(n41021), .A2(n41020), .Z(n41022) );
  XNOR2HSV1 U45521 ( .A1(n41023), .A2(n41022), .ZN(n41025) );
  CLKNAND2HSV0 U45522 ( .A1(n41677), .A2(n41689), .ZN(n41024) );
  XOR2HSV0 U45523 ( .A1(n41025), .A2(n41024), .Z(n41028) );
  BUFHSV6 U45524 ( .I(n41026), .Z(n41390) );
  INAND2HSV2 U45525 ( .A1(n44337), .B1(n41390), .ZN(n41027) );
  XOR2HSV4 U45526 ( .A1(n41028), .A2(n41027), .Z(n41030) );
  NAND2HSV0 U45527 ( .A1(n54683), .A2(n40873), .ZN(n41029) );
  XNOR2HSV4 U45528 ( .A1(n41030), .A2(n41029), .ZN(n41032) );
  NAND2HSV2 U45529 ( .A1(n41061), .A2(n53512), .ZN(n41031) );
  XNOR2HSV4 U45530 ( .A1(n41032), .A2(n41031), .ZN(n41040) );
  CLKNHSV6 U45531 ( .I(n41040), .ZN(n41036) );
  INAND3HSV4 U45532 ( .A1(n41033), .B1(n41038), .B2(n41036), .ZN(n41042) );
  INHSV2 U45533 ( .I(n41034), .ZN(n41035) );
  AOI21HSV4 U45534 ( .A1(n41038), .A2(n41037), .B(n41036), .ZN(n41039) );
  AOI21HSV4 U45535 ( .A1(n41043), .A2(n41040), .B(n41039), .ZN(n41041) );
  OAI21HSV4 U45536 ( .A1(n41043), .A2(n41042), .B(n41041), .ZN(n41047) );
  INHSV2 U45537 ( .I(n41238), .ZN(n44649) );
  NAND2HSV2 U45538 ( .A1(n41238), .A2(\pe1/ti_7t [13]), .ZN(n41044) );
  CLKNAND2HSV3 U45539 ( .A1(n41045), .A2(n41044), .ZN(n44696) );
  BUFHSV8 U45540 ( .I(n44696), .Z(n41243) );
  INHSV2 U45541 ( .I(n41331), .ZN(n41212) );
  XNOR2HSV4 U45542 ( .A1(n41047), .A2(n41046), .ZN(n41240) );
  NOR2HSV2 U45543 ( .A1(n41217), .A2(\pe1/ti_7t [16]), .ZN(n41140) );
  NOR2HSV2 U45544 ( .A1(n41140), .A2(n42067), .ZN(n41048) );
  NAND2HSV2 U45545 ( .A1(n41051), .A2(n41050), .ZN(n41055) );
  CLKNAND2HSV2 U45546 ( .A1(n41053), .A2(n41052), .ZN(n41054) );
  NOR2HSV4 U45547 ( .A1(n41055), .A2(n41054), .ZN(n41312) );
  CLKNHSV2 U45548 ( .I(n41919), .ZN(n41057) );
  AOI21HSV4 U45549 ( .A1(n41312), .A2(n41129), .B(n41057), .ZN(n41058) );
  NOR2HSV4 U45550 ( .A1(n41241), .A2(n41058), .ZN(n41059) );
  NOR2HSV4 U45551 ( .A1(n41060), .A2(n41059), .ZN(n41131) );
  INHSV4 U45552 ( .I(n41131), .ZN(n41136) );
  CLKNAND2HSV2 U45553 ( .A1(n41239), .A2(n41212), .ZN(n41124) );
  BUFHSV2 U45554 ( .I(n41061), .Z(n54162) );
  NAND2HSV2 U45555 ( .A1(n54162), .A2(n40823), .ZN(n41110) );
  BUFHSV2 U45556 ( .I(n41929), .Z(n41332) );
  NAND2HSV2 U45557 ( .A1(n41332), .A2(n41298), .ZN(n41103) );
  CLKNAND2HSV0 U45558 ( .A1(n41144), .A2(n41676), .ZN(n41097) );
  CLKNHSV0 U45559 ( .I(n46142), .ZN(n41735) );
  CLKNAND2HSV1 U45560 ( .A1(n41735), .A2(n41355), .ZN(n41063) );
  NAND2HSV0 U45561 ( .A1(n41736), .A2(n53922), .ZN(n41062) );
  XOR2HSV0 U45562 ( .A1(n41063), .A2(n41062), .Z(n41067) );
  NAND2HSV0 U45563 ( .A1(n59987), .A2(n41644), .ZN(n41065) );
  CLKNAND2HSV0 U45564 ( .A1(n59989), .A2(n41170), .ZN(n41064) );
  XOR2HSV0 U45565 ( .A1(n41065), .A2(n41064), .Z(n41066) );
  XOR2HSV0 U45566 ( .A1(n41067), .A2(n41066), .Z(n41073) );
  NAND2HSV0 U45567 ( .A1(n41358), .A2(\pe1/bq[17] ), .ZN(n41069) );
  CLKNAND2HSV0 U45568 ( .A1(n41145), .A2(\pe1/bq[18] ), .ZN(n41068) );
  XOR2HSV0 U45569 ( .A1(n41069), .A2(n41068), .Z(n41071) );
  INHSV2 U45570 ( .I(n53793), .ZN(n41374) );
  NAND2HSV0 U45571 ( .A1(n41152), .A2(n41374), .ZN(n41070) );
  XOR2HSV0 U45572 ( .A1(n41071), .A2(n41070), .Z(n41072) );
  XNOR2HSV1 U45573 ( .A1(n41073), .A2(n41072), .ZN(n41079) );
  NAND2HSV0 U45574 ( .A1(n40898), .A2(\pe1/bq[16] ), .ZN(n41630) );
  BUFHSV2 U45575 ( .I(n41074), .Z(n53833) );
  INHSV2 U45576 ( .I(n54973), .ZN(n41424) );
  CLKNAND2HSV0 U45577 ( .A1(n41153), .A2(n41424), .ZN(n54074) );
  INHSV2 U45578 ( .I(n53911), .ZN(n41284) );
  XNOR2HSV1 U45579 ( .A1(n41079), .A2(n41078), .ZN(n41091) );
  NOR2HSV0 U45580 ( .A1(n53447), .A2(n41963), .ZN(n53832) );
  CLKNAND2HSV1 U45581 ( .A1(\pe1/aot [20]), .A2(\pe1/bq[27] ), .ZN(n41251) );
  XOR2HSV0 U45582 ( .A1(n53832), .A2(n41251), .Z(n41081) );
  INHSV2 U45583 ( .I(n41931), .ZN(n59733) );
  NAND2HSV0 U45584 ( .A1(n59733), .A2(n41339), .ZN(n41759) );
  CLKNHSV0 U45585 ( .I(n42264), .ZN(n42366) );
  NAND2HSV2 U45586 ( .A1(n41169), .A2(n42366), .ZN(n53822) );
  XOR2HSV0 U45587 ( .A1(n41759), .A2(n53822), .Z(n41080) );
  XOR2HSV0 U45588 ( .A1(n41081), .A2(n41080), .Z(n41089) );
  CLKNAND2HSV1 U45589 ( .A1(\pe1/aot [25]), .A2(n54302), .ZN(n44540) );
  XOR2HSV0 U45590 ( .A1(n41082), .A2(n44540), .Z(n41087) );
  INHSV2 U45591 ( .I(n54829), .ZN(n59988) );
  NAND2HSV2 U45592 ( .A1(n59988), .A2(n25428), .ZN(n41085) );
  CLKNAND2HSV0 U45593 ( .A1(n55186), .A2(n41083), .ZN(n41084) );
  XOR2HSV0 U45594 ( .A1(n41085), .A2(n41084), .Z(n41086) );
  XOR2HSV0 U45595 ( .A1(n41087), .A2(n41086), .Z(n41088) );
  XOR2HSV0 U45596 ( .A1(n41089), .A2(n41088), .Z(n41090) );
  XNOR2HSV1 U45597 ( .A1(n41091), .A2(n41090), .ZN(n41093) );
  CLKNAND2HSV1 U45598 ( .A1(n42210), .A2(n54716), .ZN(n41092) );
  XOR2HSV0 U45599 ( .A1(n41093), .A2(n41092), .Z(n41095) );
  NAND2HSV2 U45600 ( .A1(n41287), .A2(n41188), .ZN(n41094) );
  XNOR2HSV1 U45601 ( .A1(n41095), .A2(n41094), .ZN(n41096) );
  XNOR2HSV1 U45602 ( .A1(n41097), .A2(n41096), .ZN(n41099) );
  CLKNAND2HSV1 U45603 ( .A1(n41557), .A2(n54724), .ZN(n41098) );
  XOR2HSV0 U45604 ( .A1(n41099), .A2(n41098), .Z(n41101) );
  NAND2HSV0 U45605 ( .A1(n42431), .A2(n41387), .ZN(n41100) );
  XOR2HSV0 U45606 ( .A1(n41101), .A2(n41100), .Z(n41102) );
  XNOR2HSV1 U45607 ( .A1(n41103), .A2(n41102), .ZN(n41105) );
  NAND2HSV0 U45608 ( .A1(n29763), .A2(n41143), .ZN(n41104) );
  XOR2HSV0 U45609 ( .A1(n41105), .A2(n41104), .Z(n41108) );
  INHSV2 U45610 ( .I(n41390), .ZN(n41301) );
  NOR2HSV2 U45611 ( .A1(n41301), .A2(n41848), .ZN(n41107) );
  BUFHSV2 U45612 ( .I(n41391), .Z(n42439) );
  NAND2HSV2 U45613 ( .A1(n42439), .A2(n41689), .ZN(n41106) );
  XOR3HSV2 U45614 ( .A1(n41108), .A2(n41107), .A3(n41106), .Z(n41109) );
  XOR2HSV0 U45615 ( .A1(n41110), .A2(n41109), .Z(n41123) );
  INHSV2 U45616 ( .I(n41112), .ZN(n41113) );
  NAND2HSV2 U45617 ( .A1(n41114), .A2(n41113), .ZN(n41116) );
  INHSV2 U45618 ( .I(n41118), .ZN(n41119) );
  NOR2HSV4 U45619 ( .A1(n41120), .A2(n41119), .ZN(n41309) );
  NOR2HSV4 U45620 ( .A1(n41309), .A2(n41507), .ZN(n41122) );
  CLKAND2HSV2 U45621 ( .A1(n41243), .A2(n40873), .Z(n41121) );
  XOR3HSV2 U45622 ( .A1(n41123), .A2(n41122), .A3(n41121), .Z(n41125) );
  NAND2HSV2 U45623 ( .A1(n41124), .A2(n41125), .ZN(n41128) );
  CLKNHSV2 U45624 ( .I(n41125), .ZN(n41126) );
  INHSV4 U45625 ( .I(n41130), .ZN(n41137) );
  INHSV2 U45626 ( .I(n41238), .ZN(n41129) );
  CLKNAND2HSV2 U45627 ( .A1(n41220), .A2(n41129), .ZN(n41133) );
  CLKNAND2HSV2 U45628 ( .A1(n41131), .A2(n41130), .ZN(n41219) );
  INHSV2 U45629 ( .I(n41219), .ZN(n41132) );
  NOR2HSV4 U45630 ( .A1(n41133), .A2(n41132), .ZN(n41216) );
  CLKNAND2HSV3 U45631 ( .A1(n41136), .A2(n41135), .ZN(n41139) );
  CLKNHSV2 U45632 ( .I(n41137), .ZN(n41138) );
  OAI22HSV4 U45633 ( .A1(n41219), .A2(n41218), .B1(n41139), .B2(n41138), .ZN(
        n41215) );
  XNOR2HSV4 U45634 ( .A1(n41240), .A2(n41421), .ZN(n41235) );
  NAND2HSV4 U45635 ( .A1(n41235), .A2(n41234), .ZN(n41141) );
  CLKNAND2HSV4 U45636 ( .A1(n41141), .A2(n41236), .ZN(n41237) );
  BUFHSV8 U45637 ( .I(n41142), .Z(n59534) );
  CLKAND2HSV2 U45638 ( .A1(n59534), .A2(n40873), .Z(n41208) );
  CLKNAND2HSV0 U45639 ( .A1(n41929), .A2(n41143), .ZN(n41200) );
  CLKNAND2HSV0 U45640 ( .A1(n41144), .A2(n54724), .ZN(n41194) );
  CLKNAND2HSV0 U45641 ( .A1(n41145), .A2(\pe1/bq[19] ), .ZN(n41147) );
  CLKNAND2HSV0 U45642 ( .A1(n42412), .A2(\pe1/bq[17] ), .ZN(n41146) );
  XOR2HSV0 U45643 ( .A1(n41147), .A2(n41146), .Z(n41151) );
  CLKNAND2HSV1 U45644 ( .A1(n59733), .A2(n25428), .ZN(n41149) );
  NAND2HSV0 U45645 ( .A1(n41736), .A2(n42223), .ZN(n41148) );
  XOR2HSV0 U45646 ( .A1(n41149), .A2(n41148), .Z(n41150) );
  XOR2HSV0 U45647 ( .A1(n41151), .A2(n41150), .Z(n41159) );
  CLKNAND2HSV0 U45648 ( .A1(n41152), .A2(n41284), .ZN(n41157) );
  CLKNAND2HSV1 U45649 ( .A1(n41153), .A2(n54836), .ZN(n41777) );
  NAND2HSV0 U45650 ( .A1(n41153), .A2(n54302), .ZN(n53443) );
  OAI21HSV0 U45651 ( .A1(n45814), .A2(n41076), .B(n53443), .ZN(n41154) );
  OAI21HSV0 U45652 ( .A1(n41155), .A2(n41777), .B(n41154), .ZN(n41156) );
  XOR2HSV0 U45653 ( .A1(n41157), .A2(n41156), .Z(n41158) );
  XOR2HSV0 U45654 ( .A1(n41159), .A2(n41158), .Z(n41168) );
  NAND2HSV0 U45655 ( .A1(n41160), .A2(n42359), .ZN(n41166) );
  NAND2HSV0 U45656 ( .A1(\pe1/aot [16]), .A2(\pe1/bq[21] ), .ZN(n42372) );
  NAND2HSV0 U45657 ( .A1(n40898), .A2(\pe1/bq[21] ), .ZN(n41632) );
  OAI21HSV2 U45658 ( .A1(n54673), .A2(n41967), .B(n41632), .ZN(n41161) );
  OAI21HSV0 U45659 ( .A1(n42372), .A2(n41162), .B(n41161), .ZN(n41164) );
  XNOR2HSV1 U45660 ( .A1(n41164), .A2(n41163), .ZN(n41165) );
  XNOR2HSV1 U45661 ( .A1(n41166), .A2(n41165), .ZN(n41167) );
  XNOR2HSV1 U45662 ( .A1(n41168), .A2(n41167), .ZN(n41187) );
  NAND2HSV0 U45663 ( .A1(n41169), .A2(n41644), .ZN(n41172) );
  INHSV2 U45664 ( .I(n54829), .ZN(n42220) );
  CLKNAND2HSV0 U45665 ( .A1(n42220), .A2(n41170), .ZN(n41171) );
  XOR2HSV0 U45666 ( .A1(n41172), .A2(n41171), .Z(n41177) );
  NAND2HSV0 U45667 ( .A1(n41735), .A2(n41173), .ZN(n41175) );
  NAND2HSV0 U45668 ( .A1(n41358), .A2(\pe1/bq[18] ), .ZN(n41174) );
  XOR2HSV0 U45669 ( .A1(n41175), .A2(n41174), .Z(n41176) );
  XOR2HSV0 U45670 ( .A1(n41177), .A2(n41176), .Z(n41185) );
  NAND2HSV0 U45671 ( .A1(n59987), .A2(n41771), .ZN(n41179) );
  NAND2HSV0 U45672 ( .A1(\pe1/aot [25]), .A2(\pe1/bq[23] ), .ZN(n41178) );
  XOR2HSV0 U45673 ( .A1(n41179), .A2(n41178), .Z(n41183) );
  CLKNAND2HSV1 U45674 ( .A1(\pe1/aot [28]), .A2(n54565), .ZN(n41181) );
  NAND2HSV0 U45675 ( .A1(\pe1/aot [20]), .A2(n53922), .ZN(n41180) );
  XOR2HSV0 U45676 ( .A1(n41181), .A2(n41180), .Z(n41182) );
  XOR2HSV0 U45677 ( .A1(n41183), .A2(n41182), .Z(n41184) );
  XOR2HSV0 U45678 ( .A1(n41185), .A2(n41184), .Z(n41186) );
  XNOR2HSV1 U45679 ( .A1(n41187), .A2(n41186), .ZN(n41190) );
  CLKNAND2HSV1 U45680 ( .A1(n42210), .A2(n41188), .ZN(n41189) );
  XOR2HSV0 U45681 ( .A1(n41190), .A2(n41189), .Z(n41192) );
  NAND2HSV2 U45682 ( .A1(n41287), .A2(n41676), .ZN(n41191) );
  XNOR2HSV1 U45683 ( .A1(n41192), .A2(n41191), .ZN(n41193) );
  XNOR2HSV1 U45684 ( .A1(n41194), .A2(n41193), .ZN(n41196) );
  CLKNAND2HSV0 U45685 ( .A1(n41557), .A2(n41387), .ZN(n41195) );
  XOR2HSV0 U45686 ( .A1(n41196), .A2(n41195), .Z(n41198) );
  NAND2HSV0 U45687 ( .A1(n42431), .A2(n41298), .ZN(n41197) );
  XOR2HSV0 U45688 ( .A1(n41198), .A2(n41197), .Z(n41199) );
  XNOR2HSV1 U45689 ( .A1(n41200), .A2(n41199), .ZN(n41203) );
  NAND2HSV0 U45690 ( .A1(n29773), .A2(n41201), .ZN(n41202) );
  XOR2HSV0 U45691 ( .A1(n41203), .A2(n41202), .Z(n41207) );
  INAND2HSV2 U45692 ( .A1(n42086), .B1(n41390), .ZN(n41204) );
  INHSV2 U45693 ( .I(n41204), .ZN(n41206) );
  NAND2HSV0 U45694 ( .A1(n54732), .A2(n40823), .ZN(n41205) );
  XOR3HSV2 U45695 ( .A1(n41207), .A2(n41206), .A3(n41205), .Z(n41209) );
  CLKNAND2HSV1 U45696 ( .A1(n41208), .A2(n41209), .ZN(n41211) );
  AOI21HSV2 U45697 ( .A1(n59534), .A2(n40873), .B(n41209), .ZN(n41210) );
  INOR2HSV4 U45698 ( .A1(n41211), .B1(n41210), .ZN(n41232) );
  INAND2HSV2 U45699 ( .A1(n41309), .B1(n41212), .ZN(n41231) );
  INHSV2 U45700 ( .I(n42037), .ZN(n59365) );
  NAND2HSV4 U45701 ( .A1(n41239), .A2(n59365), .ZN(n41233) );
  NOR2HSV1 U45702 ( .A1(n41218), .A2(n41217), .ZN(n41222) );
  NAND2HSV2 U45703 ( .A1(n41220), .A2(n41219), .ZN(n41221) );
  MUX2NHSV2 U45704 ( .I0(n41218), .I1(n41222), .S(n41221), .ZN(n41223) );
  CLKNAND2HSV3 U45705 ( .A1(n41224), .A2(n41223), .ZN(n60106) );
  NAND2HSV2 U45706 ( .A1(n41712), .A2(\pe1/ti_7t [18]), .ZN(n41226) );
  BUFHSV8 U45707 ( .I(n41412), .Z(n54730) );
  INHSV2 U45708 ( .I(n41228), .ZN(n53512) );
  NAND2HSV2 U45709 ( .A1(n41238), .A2(\pe1/ti_7t [17]), .ZN(n41329) );
  NAND2HSV4 U45710 ( .A1(n41330), .A2(n41329), .ZN(n41847) );
  CLKNAND2HSV0 U45711 ( .A1(n48331), .A2(\pe1/ti_7t [16]), .ZN(n41505) );
  NAND2HSV2 U45712 ( .A1(n41734), .A2(n40823), .ZN(n41308) );
  CLKNAND2HSV0 U45713 ( .A1(n54162), .A2(n40605), .ZN(n41306) );
  CLKNAND2HSV1 U45714 ( .A1(n41332), .A2(n41387), .ZN(n41297) );
  CLKNAND2HSV1 U45715 ( .A1(n41609), .A2(n41188), .ZN(n41291) );
  NOR2HSV0 U45716 ( .A1(n40445), .A2(n54973), .ZN(n41245) );
  CLKNAND2HSV0 U45717 ( .A1(n53538), .A2(n54995), .ZN(n41244) );
  XOR2HSV0 U45718 ( .A1(n41245), .A2(n41244), .Z(n41247) );
  BUFHSV2 U45719 ( .I(n41752), .Z(n41522) );
  CLKNAND2HSV1 U45720 ( .A1(n41522), .A2(n41550), .ZN(n41246) );
  XOR2HSV0 U45721 ( .A1(n41247), .A2(n41246), .Z(n41250) );
  NAND2HSV0 U45722 ( .A1(n41248), .A2(n41374), .ZN(n41249) );
  XNOR2HSV1 U45723 ( .A1(n41250), .A2(n41249), .ZN(n41266) );
  CLKNAND2HSV0 U45724 ( .A1(n41736), .A2(\pe1/bq[26] ), .ZN(n41350) );
  NAND2HSV0 U45725 ( .A1(n59987), .A2(\pe1/bq[14] ), .ZN(n44537) );
  OAI22HSV0 U45726 ( .A1(n41076), .A2(n54281), .B1(n41944), .B2(n42264), .ZN(
        n41252) );
  OAI21HSV0 U45727 ( .A1(n41253), .A2(n44537), .B(n41252), .ZN(n41254) );
  XOR2HSV0 U45728 ( .A1(n41255), .A2(n41254), .Z(n41264) );
  NAND2HSV0 U45729 ( .A1(n54307), .A2(n55100), .ZN(n41423) );
  OAI22HSV0 U45730 ( .A1(n45814), .A2(n41256), .B1(n41974), .B2(n41947), .ZN(
        n41257) );
  OAI21HSV0 U45731 ( .A1(n41258), .A2(n41423), .B(n41257), .ZN(n41262) );
  NAND2HSV0 U45732 ( .A1(n41169), .A2(\pe1/bq[18] ), .ZN(n41886) );
  CLKNAND2HSV0 U45733 ( .A1(\pe1/aot [28]), .A2(\pe1/bq[18] ), .ZN(n41634) );
  OAI21HSV0 U45734 ( .A1(n41885), .A2(n54185), .B(n41634), .ZN(n41259) );
  OAI21HSV0 U45735 ( .A1(n41260), .A2(n41886), .B(n41259), .ZN(n41261) );
  XOR2HSV0 U45736 ( .A1(n41262), .A2(n41261), .Z(n41263) );
  XOR2HSV0 U45737 ( .A1(n41264), .A2(n41263), .Z(n41265) );
  XOR2HSV0 U45738 ( .A1(n41266), .A2(n41265), .Z(n41283) );
  NAND2HSV0 U45739 ( .A1(n59989), .A2(n53411), .ZN(n41268) );
  NAND2HSV0 U45740 ( .A1(n59733), .A2(n53922), .ZN(n41267) );
  XOR2HSV0 U45741 ( .A1(n41268), .A2(n41267), .Z(n41281) );
  INHSV2 U45742 ( .I(\pe1/aot [14]), .ZN(n54843) );
  NAND2HSV0 U45743 ( .A1(\pe1/aot [14]), .A2(\pe1/bq[20] ), .ZN(n48344) );
  OAI22HSV0 U45744 ( .A1(n41967), .A2(n54843), .B1(n46629), .B2(n48060), .ZN(
        n41269) );
  OAI21HSV0 U45745 ( .A1(n41270), .A2(n48344), .B(n41269), .ZN(n41272) );
  NAND2HSV0 U45746 ( .A1(n59988), .A2(n41339), .ZN(n41271) );
  XNOR2HSV1 U45747 ( .A1(n41272), .A2(n41271), .ZN(n41280) );
  NAND2HSV0 U45748 ( .A1(n40898), .A2(n42092), .ZN(n41274) );
  NAND2HSV0 U45749 ( .A1(\pe1/aot [25]), .A2(\pe1/bq[21] ), .ZN(n41273) );
  XOR2HSV0 U45750 ( .A1(n41274), .A2(n41273), .Z(n41278) );
  NAND2HSV0 U45751 ( .A1(n41735), .A2(\pe1/bq[23] ), .ZN(n41276) );
  CLKNAND2HSV0 U45752 ( .A1(n42132), .A2(n48055), .ZN(n41275) );
  XOR2HSV0 U45753 ( .A1(n41276), .A2(n41275), .Z(n41277) );
  XOR2HSV0 U45754 ( .A1(n41278), .A2(n41277), .Z(n41279) );
  XOR3HSV2 U45755 ( .A1(n41281), .A2(n41280), .A3(n41279), .Z(n41282) );
  XNOR2HSV1 U45756 ( .A1(n41283), .A2(n41282), .ZN(n41286) );
  CLKNAND2HSV0 U45757 ( .A1(n42210), .A2(n41284), .ZN(n41285) );
  XOR2HSV0 U45758 ( .A1(n41286), .A2(n41285), .Z(n41289) );
  CLKNAND2HSV1 U45759 ( .A1(n42275), .A2(n54716), .ZN(n41288) );
  XNOR2HSV1 U45760 ( .A1(n41289), .A2(n41288), .ZN(n41290) );
  XNOR2HSV1 U45761 ( .A1(n41291), .A2(n41290), .ZN(n41293) );
  NAND2HSV0 U45762 ( .A1(n41557), .A2(n41676), .ZN(n41292) );
  XOR2HSV0 U45763 ( .A1(n41293), .A2(n41292), .Z(n41295) );
  NAND2HSV0 U45764 ( .A1(n42431), .A2(n54724), .ZN(n41294) );
  XOR2HSV0 U45765 ( .A1(n41295), .A2(n41294), .Z(n41296) );
  XNOR2HSV1 U45766 ( .A1(n41297), .A2(n41296), .ZN(n41300) );
  NAND2HSV0 U45767 ( .A1(n29762), .A2(n41298), .ZN(n41299) );
  XOR2HSV0 U45768 ( .A1(n41300), .A2(n41299), .Z(n41304) );
  NOR2HSV2 U45769 ( .A1(n41301), .A2(n41392), .ZN(n41303) );
  NAND2HSV2 U45770 ( .A1(n41894), .A2(\pe1/got [25]), .ZN(n41302) );
  XOR3HSV2 U45771 ( .A1(n41304), .A2(n41303), .A3(n41302), .Z(n41305) );
  XNOR2HSV1 U45772 ( .A1(n41306), .A2(n41305), .ZN(n41307) );
  CLKXOR2HSV4 U45773 ( .A1(n41308), .A2(n41307), .Z(n41311) );
  BUFHSV2 U45774 ( .I(n41309), .Z(n53393) );
  INHSV2 U45775 ( .I(n53393), .ZN(n41733) );
  NAND2HSV2 U45776 ( .A1(n41733), .A2(n40873), .ZN(n41310) );
  XNOR2HSV4 U45777 ( .A1(n41311), .A2(n41310), .ZN(n41314) );
  INHSV4 U45778 ( .I(n41312), .ZN(n41575) );
  NAND2HSV2 U45779 ( .A1(n41575), .A2(n59994), .ZN(n41313) );
  XNOR2HSV4 U45780 ( .A1(n41314), .A2(n41313), .ZN(n41317) );
  CLKNHSV1 U45781 ( .I(n41319), .ZN(n41315) );
  NOR2HSV4 U45782 ( .A1(n41317), .A2(n41315), .ZN(n41316) );
  NAND2HSV2 U45783 ( .A1(n41420), .A2(n41316), .ZN(n41322) );
  CLKNHSV2 U45784 ( .I(n41317), .ZN(n41318) );
  AOI21HSV2 U45785 ( .A1(n41420), .A2(n41319), .B(n41318), .ZN(n41324) );
  CLKNHSV2 U45786 ( .I(n41322), .ZN(n41325) );
  OAI21HSV4 U45787 ( .A1(n41325), .A2(n41324), .B(n41323), .ZN(n41326) );
  XNOR2HSV4 U45788 ( .A1(n54730), .A2(n41699), .ZN(n41592) );
  INHSV2 U45789 ( .I(n41331), .ZN(n53514) );
  CLKNAND2HSV4 U45790 ( .A1(n41508), .A2(n53514), .ZN(n41406) );
  CLKNAND2HSV1 U45791 ( .A1(n41733), .A2(n40823), .ZN(n41402) );
  CLKNAND2HSV2 U45792 ( .A1(n41575), .A2(n40873), .ZN(n41401) );
  NAND2HSV2 U45793 ( .A1(n42088), .A2(\pe1/got [26]), .ZN(n41399) );
  BUFHSV2 U45794 ( .I(n54162), .Z(n54362) );
  CLKBUFHSV4 U45795 ( .I(n54362), .Z(n54264) );
  NAND2HSV2 U45796 ( .A1(n54264), .A2(\pe1/got [25]), .ZN(n41397) );
  CLKNAND2HSV0 U45797 ( .A1(n41332), .A2(n54724), .ZN(n41386) );
  CLKNAND2HSV0 U45798 ( .A1(n41609), .A2(n54716), .ZN(n41380) );
  CLKNAND2HSV1 U45799 ( .A1(n59590), .A2(n41550), .ZN(n41336) );
  NAND2HSV2 U45800 ( .A1(n41743), .A2(n41760), .ZN(n53965) );
  INHSV2 U45801 ( .I(n53672), .ZN(n54912) );
  NAND2HSV2 U45802 ( .A1(n54912), .A2(n41083), .ZN(n42266) );
  XOR2HSV0 U45803 ( .A1(n53965), .A2(n42266), .Z(n41335) );
  XNOR2HSV1 U45804 ( .A1(n41336), .A2(n41335), .ZN(n41373) );
  NOR2HSV0 U45805 ( .A1(n41885), .A2(n53819), .ZN(n41338) );
  NAND2HSV0 U45806 ( .A1(\pe1/aot [28]), .A2(n54995), .ZN(n41337) );
  XOR2HSV0 U45807 ( .A1(n41338), .A2(n41337), .Z(n41343) );
  NAND2HSV0 U45808 ( .A1(n54916), .A2(n40494), .ZN(n41341) );
  NAND2HSV0 U45809 ( .A1(n59989), .A2(n41339), .ZN(n41340) );
  XOR2HSV0 U45810 ( .A1(n41341), .A2(n41340), .Z(n41342) );
  XOR2HSV0 U45811 ( .A1(n41343), .A2(n41342), .Z(n41349) );
  NAND2HSV0 U45812 ( .A1(n42412), .A2(n41641), .ZN(n41345) );
  NAND2HSV0 U45813 ( .A1(n42139), .A2(n41645), .ZN(n41344) );
  XOR2HSV0 U45814 ( .A1(n41345), .A2(n41344), .Z(n41347) );
  CLKNAND2HSV0 U45815 ( .A1(n41522), .A2(\pe1/got [14]), .ZN(n41346) );
  XOR2HSV0 U45816 ( .A1(n41347), .A2(n41346), .Z(n41348) );
  XOR2HSV0 U45817 ( .A1(n41349), .A2(n41348), .Z(n41372) );
  NOR2HSV2 U45818 ( .A1(n42361), .A2(n41622), .ZN(n41625) );
  XOR2HSV0 U45819 ( .A1(n41625), .A2(n41350), .Z(n41354) );
  XOR2HSV0 U45820 ( .A1(n41352), .A2(n41351), .Z(n41353) );
  XOR2HSV0 U45821 ( .A1(n41354), .A2(n41353), .Z(n41371) );
  NAND2HSV0 U45822 ( .A1(n59987), .A2(n41355), .ZN(n41357) );
  NAND2HSV0 U45823 ( .A1(n42220), .A2(n53922), .ZN(n41356) );
  XOR2HSV0 U45824 ( .A1(n41357), .A2(n41356), .Z(n41362) );
  NAND2HSV0 U45825 ( .A1(n54307), .A2(\pe1/bq[21] ), .ZN(n41360) );
  NAND2HSV0 U45826 ( .A1(n41358), .A2(n41424), .ZN(n41359) );
  XOR2HSV0 U45827 ( .A1(n41360), .A2(n41359), .Z(n41361) );
  XOR2HSV0 U45828 ( .A1(n41362), .A2(n41361), .Z(n41369) );
  XOR2HSV0 U45829 ( .A1(n41364), .A2(n41363), .Z(n41367) );
  CLKNAND2HSV1 U45830 ( .A1(n53538), .A2(n55100), .ZN(n53958) );
  CLKNAND2HSV0 U45831 ( .A1(\pe1/aot [14]), .A2(n42231), .ZN(n41365) );
  XOR2HSV0 U45832 ( .A1(n53958), .A2(n41365), .Z(n41366) );
  XOR2HSV0 U45833 ( .A1(n41367), .A2(n41366), .Z(n41368) );
  XOR2HSV0 U45834 ( .A1(n41369), .A2(n41368), .Z(n41370) );
  XOR4HSV1 U45835 ( .A1(n41373), .A2(n41372), .A3(n41371), .A4(n41370), .Z(
        n41376) );
  NAND2HSV0 U45836 ( .A1(n42210), .A2(n41374), .ZN(n41375) );
  XNOR2HSV1 U45837 ( .A1(n41376), .A2(n41375), .ZN(n41378) );
  INHSV2 U45838 ( .I(n53911), .ZN(n41851) );
  CLKNAND2HSV1 U45839 ( .A1(n59674), .A2(n41851), .ZN(n41377) );
  XNOR2HSV1 U45840 ( .A1(n41378), .A2(n41377), .ZN(n41379) );
  XNOR2HSV1 U45841 ( .A1(n41380), .A2(n41379), .ZN(n41382) );
  NAND2HSV0 U45842 ( .A1(n41557), .A2(n41188), .ZN(n41381) );
  XOR2HSV0 U45843 ( .A1(n41382), .A2(n41381), .Z(n41384) );
  NAND2HSV0 U45844 ( .A1(n42431), .A2(n41676), .ZN(n41383) );
  XOR2HSV0 U45845 ( .A1(n41384), .A2(n41383), .Z(n41385) );
  XNOR2HSV1 U45846 ( .A1(n41386), .A2(n41385), .ZN(n41389) );
  NAND2HSV0 U45847 ( .A1(n29763), .A2(n41387), .ZN(n41388) );
  XOR2HSV0 U45848 ( .A1(n41389), .A2(n41388), .Z(n41395) );
  BUFHSV2 U45849 ( .I(n41390), .Z(n44532) );
  INHSV2 U45850 ( .I(n44532), .ZN(n41566) );
  NOR2HSV2 U45851 ( .A1(n41566), .A2(n41926), .ZN(n41394) );
  NAND2HSV2 U45852 ( .A1(n54115), .A2(n40913), .ZN(n41393) );
  XOR3HSV2 U45853 ( .A1(n41395), .A2(n41394), .A3(n41393), .Z(n41396) );
  XNOR2HSV1 U45854 ( .A1(n41397), .A2(n41396), .ZN(n41398) );
  XOR2HSV0 U45855 ( .A1(n41399), .A2(n41398), .Z(n41400) );
  XOR3HSV2 U45856 ( .A1(n41402), .A2(n41401), .A3(n41400), .Z(n41404) );
  NAND2HSV2 U45857 ( .A1(n41420), .A2(n59994), .ZN(n41403) );
  XNOR2HSV4 U45858 ( .A1(n41404), .A2(n41403), .ZN(n41405) );
  XNOR2HSV4 U45859 ( .A1(n41406), .A2(n41405), .ZN(n41409) );
  INHSV4 U45860 ( .I(n41409), .ZN(n41407) );
  NAND2HSV4 U45861 ( .A1(n41593), .A2(n41595), .ZN(n41590) );
  NAND2HSV2 U45862 ( .A1(\pe1/ti_7t [20]), .A2(n41242), .ZN(n41411) );
  BUFHSV4 U45863 ( .I(n41699), .Z(n41413) );
  OAI21HSV4 U45864 ( .A1(n44529), .A2(n41414), .B(n41413), .ZN(n41417) );
  NOR2HSV2 U45865 ( .A1(n41699), .A2(n41414), .ZN(n41415) );
  INHSV2 U45866 ( .I(n41418), .ZN(n41924) );
  MUX2NHSV2 U45867 ( .I0(pov1[19]), .I1(\pe1/ti_7t [19]), .S(n41924), .ZN(
        n41419) );
  INHSV4 U45868 ( .I(n41419), .ZN(n41925) );
  INHSV4 U45869 ( .I(n41925), .ZN(n42356) );
  NOR2HSV2 U45870 ( .A1(n42356), .A2(n44337), .ZN(n41504) );
  BUFHSV2 U45871 ( .I(n26839), .Z(n41927) );
  CLKNAND2HSV1 U45872 ( .A1(n41927), .A2(n41689), .ZN(n41502) );
  BUFHSV8 U45873 ( .I(n41508), .Z(n59592) );
  NAND2HSV2 U45874 ( .A1(n59592), .A2(\pe1/got [25]), .ZN(n41500) );
  CLKBUFHSV4 U45875 ( .I(n41420), .Z(n44531) );
  NOR2HSV2 U45876 ( .A1(n41849), .A2(n41392), .ZN(n41498) );
  CLKNHSV0 U45877 ( .I(n53393), .ZN(n59518) );
  INHSV2 U45878 ( .I(n42209), .ZN(n54452) );
  NAND2HSV0 U45879 ( .A1(n59518), .A2(n54452), .ZN(n41496) );
  BUFHSV4 U45880 ( .I(n41421), .Z(n54691) );
  CLKNAND2HSV0 U45881 ( .A1(n41850), .A2(\pe1/got [23]), .ZN(n41495) );
  NAND2HSV0 U45882 ( .A1(n53913), .A2(n54724), .ZN(n41493) );
  NAND2HSV0 U45883 ( .A1(n54041), .A2(n44530), .ZN(n41491) );
  BUFHSV2 U45884 ( .I(n41929), .Z(n42089) );
  INHSV2 U45885 ( .I(n53793), .ZN(n42162) );
  NAND2HSV0 U45886 ( .A1(n42089), .A2(n42162), .ZN(n41483) );
  CLKNAND2HSV0 U45887 ( .A1(n41609), .A2(n42155), .ZN(n41477) );
  BUFHSV8 U45888 ( .I(n41422), .Z(n59529) );
  NAND2HSV2 U45889 ( .A1(n59529), .A2(n55214), .ZN(n41475) );
  XOR2HSV0 U45890 ( .A1(n41423), .A2(n41886), .Z(n41427) );
  CLKNAND2HSV0 U45891 ( .A1(n41743), .A2(n41424), .ZN(n41633) );
  NAND2HSV0 U45892 ( .A1(n55103), .A2(n41771), .ZN(n41889) );
  XOR2HSV0 U45893 ( .A1(n41633), .A2(n41889), .Z(n41426) );
  XOR2HSV0 U45894 ( .A1(n41427), .A2(n41426), .Z(n41435) );
  BUFHSV2 U45895 ( .I(\pe1/aot [11]), .Z(n59593) );
  CLKNHSV0 U45896 ( .I(n40455), .ZN(n42125) );
  NAND2HSV0 U45897 ( .A1(n59593), .A2(n42125), .ZN(n41429) );
  NAND2HSV0 U45898 ( .A1(n42255), .A2(n54995), .ZN(n41428) );
  XOR2HSV0 U45899 ( .A1(n41429), .A2(n41428), .Z(n41433) );
  NAND2HSV0 U45900 ( .A1(\pe1/aot [14]), .A2(n40557), .ZN(n41431) );
  CLKNHSV0 U45901 ( .I(n41947), .ZN(n42106) );
  NAND2HSV0 U45902 ( .A1(n54916), .A2(n42106), .ZN(n41430) );
  XOR2HSV0 U45903 ( .A1(n41431), .A2(n41430), .Z(n41432) );
  XOR2HSV0 U45904 ( .A1(n41433), .A2(n41432), .Z(n41434) );
  XOR2HSV0 U45905 ( .A1(n41435), .A2(n41434), .Z(n41452) );
  CLKNHSV0 U45906 ( .I(n54185), .ZN(n54479) );
  NAND2HSV0 U45907 ( .A1(n59989), .A2(n54479), .ZN(n41437) );
  NAND2HSV0 U45908 ( .A1(n54663), .A2(n42092), .ZN(n41436) );
  XOR2HSV0 U45909 ( .A1(n41437), .A2(n41436), .Z(n41441) );
  NAND2HSV0 U45910 ( .A1(n42099), .A2(\pe1/bq[21] ), .ZN(n41439) );
  NAND2HSV0 U45911 ( .A1(n54293), .A2(n41641), .ZN(n41438) );
  XOR2HSV0 U45912 ( .A1(n41439), .A2(n41438), .Z(n41440) );
  XOR2HSV0 U45913 ( .A1(n41441), .A2(n41440), .Z(n41450) );
  INHSV2 U45914 ( .I(\pe1/aot [12]), .ZN(n41653) );
  INHSV2 U45915 ( .I(n41653), .ZN(n53812) );
  NAND2HSV0 U45916 ( .A1(n53812), .A2(n53922), .ZN(n41444) );
  NAND2HSV0 U45917 ( .A1(\pe1/aot [27]), .A2(n41645), .ZN(n41443) );
  XOR2HSV0 U45918 ( .A1(n41444), .A2(n41443), .Z(n41448) );
  NAND2HSV0 U45919 ( .A1(n41768), .A2(n42238), .ZN(n41446) );
  NAND2HSV0 U45920 ( .A1(n55452), .A2(n40890), .ZN(n41445) );
  XOR2HSV0 U45921 ( .A1(n41446), .A2(n41445), .Z(n41447) );
  XOR2HSV0 U45922 ( .A1(n41448), .A2(n41447), .Z(n41449) );
  XOR2HSV0 U45923 ( .A1(n41450), .A2(n41449), .Z(n41451) );
  XOR2HSV0 U45924 ( .A1(n41452), .A2(n41451), .Z(n41471) );
  INHSV2 U45925 ( .I(n54472), .ZN(n55380) );
  NAND2HSV0 U45926 ( .A1(n55380), .A2(n42231), .ZN(n41455) );
  CLKNHSV0 U45927 ( .I(n40445), .ZN(n41877) );
  NAND2HSV0 U45928 ( .A1(n41877), .A2(\pe1/bq[9] ), .ZN(n41454) );
  XOR2HSV0 U45929 ( .A1(n41455), .A2(n41454), .Z(n41457) );
  NAND2HSV0 U45930 ( .A1(n41752), .A2(n44605), .ZN(n41456) );
  XOR2HSV0 U45931 ( .A1(n41457), .A2(n41456), .Z(n41459) );
  XNOR2HSV1 U45932 ( .A1(n41459), .A2(n41458), .ZN(n41469) );
  CLKNAND2HSV0 U45933 ( .A1(n40683), .A2(n55379), .ZN(n42217) );
  CLKNAND2HSV0 U45934 ( .A1(n41964), .A2(n42373), .ZN(n41776) );
  NAND2HSV0 U45935 ( .A1(n42132), .A2(\pe1/bq[23] ), .ZN(n42211) );
  NAND2HSV0 U45936 ( .A1(n42220), .A2(n42366), .ZN(n41739) );
  XOR2HSV0 U45937 ( .A1(n41463), .A2(n41462), .Z(n41467) );
  CLKNAND2HSV0 U45938 ( .A1(n44569), .A2(n53708), .ZN(n42375) );
  CLKNAND2HSV1 U45939 ( .A1(n44566), .A2(n54311), .ZN(n41615) );
  NAND2HSV0 U45940 ( .A1(n44566), .A2(n53708), .ZN(n53529) );
  OAI21HSV0 U45941 ( .A1(n48030), .A2(n53957), .B(n53529), .ZN(n41464) );
  OAI21HSV1 U45942 ( .A1(n42375), .A2(n41615), .B(n41464), .ZN(n41465) );
  NOR2HSV0 U45943 ( .A1(n54846), .A2(n41622), .ZN(n42364) );
  XNOR2HSV1 U45944 ( .A1(n41465), .A2(n42364), .ZN(n41466) );
  XNOR2HSV1 U45945 ( .A1(n41467), .A2(n41466), .ZN(n41468) );
  XNOR2HSV1 U45946 ( .A1(n41469), .A2(n41468), .ZN(n41470) );
  XNOR2HSV1 U45947 ( .A1(n41471), .A2(n41470), .ZN(n41474) );
  BUFHSV2 U45948 ( .I(n41472), .Z(n42275) );
  NAND2HSV0 U45949 ( .A1(n42275), .A2(n55337), .ZN(n41473) );
  XOR3HSV2 U45950 ( .A1(n41475), .A2(n41474), .A3(n41473), .Z(n41476) );
  XNOR2HSV1 U45951 ( .A1(n41477), .A2(n41476), .ZN(n41479) );
  NAND2HSV0 U45952 ( .A1(n59686), .A2(n54969), .ZN(n41478) );
  XOR2HSV0 U45953 ( .A1(n41479), .A2(n41478), .Z(n41481) );
  CLKNHSV0 U45954 ( .I(n41893), .ZN(n54265) );
  NAND2HSV0 U45955 ( .A1(n54265), .A2(n54241), .ZN(n41480) );
  XOR2HSV0 U45956 ( .A1(n41481), .A2(n41480), .Z(n41482) );
  XNOR2HSV1 U45957 ( .A1(n41483), .A2(n41482), .ZN(n41486) );
  NAND2HSV0 U45958 ( .A1(n29762), .A2(n41851), .ZN(n41485) );
  XOR2HSV0 U45959 ( .A1(n41486), .A2(n41485), .Z(n41489) );
  NOR2HSV2 U45960 ( .A1(n41802), .A2(n54248), .ZN(n41488) );
  NAND2HSV0 U45961 ( .A1(n41894), .A2(n59995), .ZN(n41487) );
  XOR3HSV2 U45962 ( .A1(n41489), .A2(n41488), .A3(n41487), .Z(n41490) );
  XNOR2HSV1 U45963 ( .A1(n41491), .A2(n41490), .ZN(n41492) );
  XOR2HSV0 U45964 ( .A1(n41493), .A2(n41492), .Z(n41494) );
  XOR3HSV2 U45965 ( .A1(n41496), .A2(n41495), .A3(n41494), .Z(n41497) );
  XOR2HSV0 U45966 ( .A1(n41498), .A2(n41497), .Z(n41499) );
  XNOR2HSV1 U45967 ( .A1(n41500), .A2(n41499), .ZN(n41501) );
  XNOR2HSV1 U45968 ( .A1(n41502), .A2(n41501), .ZN(n41503) );
  NAND2HSV4 U45969 ( .A1(n53657), .A2(n40873), .ZN(n41511) );
  INHSV4 U45970 ( .I(n41511), .ZN(n41510) );
  NOR2HSV3 U45971 ( .A1(n41510), .A2(n41507), .ZN(n41509) );
  NAND2HSV2 U45972 ( .A1(n41509), .A2(n41508), .ZN(n41582) );
  NAND2HSV2 U45973 ( .A1(n41510), .A2(n41507), .ZN(n41580) );
  CLKNAND2HSV1 U45974 ( .A1(n41582), .A2(n41580), .ZN(n41579) );
  NAND2HSV0 U45975 ( .A1(n54162), .A2(\pe1/got [24]), .ZN(n41571) );
  NAND2HSV2 U45976 ( .A1(n42089), .A2(n41676), .ZN(n41563) );
  CLKNAND2HSV0 U45977 ( .A1(n41609), .A2(n41851), .ZN(n41556) );
  CLKNAND2HSV1 U45978 ( .A1(n41160), .A2(n54969), .ZN(n41515) );
  NOR2HSV0 U45979 ( .A1(n44705), .A2(n42264), .ZN(n41627) );
  XNOR2HSV1 U45980 ( .A1(n41513), .A2(n41627), .ZN(n41514) );
  XNOR2HSV1 U45981 ( .A1(n41515), .A2(n41514), .ZN(n41548) );
  NOR2HSV0 U45982 ( .A1(n53957), .A2(n54973), .ZN(n41517) );
  INHSV2 U45983 ( .I(\pe1/aot [12]), .ZN(n54672) );
  CLKNAND2HSV0 U45984 ( .A1(n55113), .A2(n41083), .ZN(n41516) );
  XOR2HSV0 U45985 ( .A1(n41517), .A2(n41516), .Z(n41521) );
  NAND2HSV0 U45986 ( .A1(n54916), .A2(n41644), .ZN(n41519) );
  CLKNAND2HSV1 U45987 ( .A1(n41768), .A2(n54479), .ZN(n41518) );
  XOR2HSV0 U45988 ( .A1(n41519), .A2(n41518), .Z(n41520) );
  XOR2HSV0 U45989 ( .A1(n41521), .A2(n41520), .Z(n41524) );
  XOR2HSV0 U45990 ( .A1(n41524), .A2(n41523), .Z(n41547) );
  NOR2HSV0 U45991 ( .A1(n54673), .A2(n48347), .ZN(n41526) );
  NAND2HSV0 U45992 ( .A1(\pe1/aot [14]), .A2(n53411), .ZN(n41525) );
  XOR2HSV0 U45993 ( .A1(n41526), .A2(n41525), .Z(n41530) );
  NAND2HSV2 U45994 ( .A1(n42132), .A2(n42125), .ZN(n41528) );
  CLKNAND2HSV0 U45995 ( .A1(n59990), .A2(n42231), .ZN(n41527) );
  XOR2HSV0 U45996 ( .A1(n41528), .A2(n41527), .Z(n41529) );
  XOR2HSV0 U45997 ( .A1(n41530), .A2(n41529), .Z(n41546) );
  NAND2HSV0 U45998 ( .A1(n41169), .A2(n42106), .ZN(n41532) );
  NAND2HSV0 U45999 ( .A1(n42220), .A2(n41771), .ZN(n41531) );
  XOR2HSV0 U46000 ( .A1(n41532), .A2(n41531), .Z(n41536) );
  NAND2HSV0 U46001 ( .A1(n41735), .A2(\pe1/bq[21] ), .ZN(n41534) );
  CLKNAND2HSV1 U46002 ( .A1(n41964), .A2(n41641), .ZN(n41533) );
  XOR2HSV0 U46003 ( .A1(n41534), .A2(n41533), .Z(n41535) );
  XOR2HSV0 U46004 ( .A1(n41536), .A2(n41535), .Z(n41544) );
  CLKNAND2HSV0 U46005 ( .A1(n41743), .A2(n42092), .ZN(n41538) );
  CLKNAND2HSV0 U46006 ( .A1(n54663), .A2(\pe1/bq[23] ), .ZN(n41537) );
  XOR2HSV0 U46007 ( .A1(n41538), .A2(n41537), .Z(n41542) );
  NAND2HSV0 U46008 ( .A1(n54307), .A2(n41760), .ZN(n41540) );
  CLKNAND2HSV1 U46009 ( .A1(n40898), .A2(n42098), .ZN(n41539) );
  XOR2HSV0 U46010 ( .A1(n41540), .A2(n41539), .Z(n41541) );
  XOR2HSV0 U46011 ( .A1(n41542), .A2(n41541), .Z(n41543) );
  XOR2HSV0 U46012 ( .A1(n41544), .A2(n41543), .Z(n41545) );
  XOR4HSV1 U46013 ( .A1(n41548), .A2(n41547), .A3(n41546), .A4(n41545), .Z(
        n41552) );
  NAND2HSV2 U46014 ( .A1(n42210), .A2(n41550), .ZN(n41551) );
  XNOR2HSV1 U46015 ( .A1(n41552), .A2(n41551), .ZN(n41554) );
  CLKNAND2HSV1 U46016 ( .A1(n59674), .A2(n42162), .ZN(n41553) );
  XNOR2HSV1 U46017 ( .A1(n41554), .A2(n41553), .ZN(n41555) );
  XNOR2HSV1 U46018 ( .A1(n41556), .A2(n41555), .ZN(n41559) );
  NAND2HSV0 U46019 ( .A1(n41557), .A2(n54716), .ZN(n41558) );
  XOR2HSV0 U46020 ( .A1(n41559), .A2(n41558), .Z(n41561) );
  NAND2HSV0 U46021 ( .A1(n42431), .A2(n41188), .ZN(n41560) );
  XOR2HSV0 U46022 ( .A1(n41561), .A2(n41560), .Z(n41562) );
  XNOR2HSV1 U46023 ( .A1(n41563), .A2(n41562), .ZN(n41565) );
  NAND2HSV0 U46024 ( .A1(n29762), .A2(n54724), .ZN(n41564) );
  XOR2HSV0 U46025 ( .A1(n41565), .A2(n41564), .Z(n41569) );
  NOR2HSV2 U46026 ( .A1(n41566), .A2(n42209), .ZN(n41568) );
  BUFHSV2 U46027 ( .I(n42439), .Z(n53996) );
  NAND2HSV2 U46028 ( .A1(n53996), .A2(\pe1/got [23]), .ZN(n41567) );
  XOR3HSV2 U46029 ( .A1(n41569), .A2(n41568), .A3(n41567), .Z(n41570) );
  XNOR2HSV1 U46030 ( .A1(n41571), .A2(n41570), .ZN(n41574) );
  NAND2HSV2 U46031 ( .A1(n42088), .A2(\pe1/got [25]), .ZN(n41573) );
  CLKNAND2HSV0 U46032 ( .A1(n41733), .A2(n41689), .ZN(n41572) );
  XOR3HSV2 U46033 ( .A1(n41574), .A2(n41573), .A3(n41572), .Z(n41577) );
  NAND2HSV2 U46034 ( .A1(n41575), .A2(n59374), .ZN(n41576) );
  XNOR2HSV1 U46035 ( .A1(n41577), .A2(n41576), .ZN(n41581) );
  INHSV2 U46036 ( .I(n41581), .ZN(n41578) );
  OAI21HSV2 U46037 ( .A1(n41579), .A2(n41583), .B(n41578), .ZN(n41585) );
  NAND2HSV2 U46038 ( .A1(n41585), .A2(n41584), .ZN(n41587) );
  XNOR2HSV4 U46039 ( .A1(n47957), .A2(n41588), .ZN(n41604) );
  CLKNHSV0 U46040 ( .I(n41592), .ZN(n41599) );
  INHSV2 U46041 ( .I(n41594), .ZN(n41598) );
  NOR2HSV2 U46042 ( .A1(n41596), .A2(n42344), .ZN(n41597) );
  OAI21HSV0 U46043 ( .A1(n42335), .A2(\pe1/ti_7t [20]), .B(n51114), .ZN(n41600) );
  CLKNHSV0 U46044 ( .I(n41600), .ZN(n41601) );
  INHSV3 U46045 ( .I(n41604), .ZN(n41606) );
  CLKNAND2HSV3 U46046 ( .A1(n41606), .A2(n41605), .ZN(n41607) );
  INHSV2 U46047 ( .I(n41924), .ZN(n42202) );
  CLKNAND2HSV1 U46048 ( .A1(n41720), .A2(\pe1/ti_7t [21]), .ZN(n41825) );
  INHSV2 U46049 ( .I(n41825), .ZN(n41827) );
  INHSV2 U46050 ( .I(n41827), .ZN(n41704) );
  CLKNAND2HSV4 U46051 ( .A1(n59592), .A2(n41731), .ZN(n41695) );
  INHSV4 U46052 ( .I(n44531), .ZN(n41732) );
  NOR2HSV4 U46053 ( .A1(n41732), .A2(n44337), .ZN(n41693) );
  NAND2HSV2 U46054 ( .A1(n41734), .A2(\pe1/got [24]), .ZN(n41686) );
  CLKNAND2HSV1 U46055 ( .A1(n54362), .A2(\pe1/got [23]), .ZN(n41684) );
  NAND2HSV0 U46056 ( .A1(n41929), .A2(n59995), .ZN(n41675) );
  NAND2HSV0 U46057 ( .A1(n41609), .A2(n42162), .ZN(n41669) );
  CLKNAND2HSV1 U46058 ( .A1(n54663), .A2(n42106), .ZN(n41611) );
  CLKNAND2HSV0 U46059 ( .A1(\pe1/aot [14]), .A2(n42125), .ZN(n41610) );
  XOR2HSV0 U46060 ( .A1(n41611), .A2(n41610), .Z(n41614) );
  NAND2HSV0 U46061 ( .A1(\pe1/aot [24]), .A2(n42092), .ZN(n54198) );
  NAND2HSV0 U46062 ( .A1(n59989), .A2(n40494), .ZN(n41612) );
  XOR2HSV0 U46063 ( .A1(n54198), .A2(n41612), .Z(n41613) );
  XOR2HSV0 U46064 ( .A1(n41614), .A2(n41613), .Z(n41663) );
  NAND2HSV0 U46065 ( .A1(n41752), .A2(\pe1/got [12]), .ZN(n41619) );
  NAND2HSV0 U46066 ( .A1(n41735), .A2(n55166), .ZN(n48343) );
  OAI21HSV0 U46067 ( .A1(n48060), .A2(n46142), .B(n41615), .ZN(n41616) );
  OAI21HSV0 U46068 ( .A1(n48343), .A2(n41617), .B(n41616), .ZN(n41618) );
  XOR2HSV0 U46069 ( .A1(n41619), .A2(n41618), .Z(n41621) );
  NAND2HSV0 U46070 ( .A1(n59590), .A2(n42155), .ZN(n41620) );
  XOR2HSV0 U46071 ( .A1(n41621), .A2(n41620), .Z(n41662) );
  NOR2HSV0 U46072 ( .A1(n53672), .A2(n48347), .ZN(n41888) );
  AOI22HSV0 U46073 ( .A1(n55186), .A2(n41623), .B1(n25428), .B2(n44541), .ZN(
        n41624) );
  AOI21HSV2 U46074 ( .A1(n41888), .A2(n41625), .B(n41624), .ZN(n41629) );
  NOR2HSV0 U46075 ( .A1(n41931), .A2(n54185), .ZN(n41757) );
  AOI22HSV0 U46076 ( .A1(n54916), .A2(n42366), .B1(n54318), .B2(n41736), .ZN(
        n41626) );
  AOI21HSV0 U46077 ( .A1(n41757), .A2(n41627), .B(n41626), .ZN(n41628) );
  XOR2HSV0 U46078 ( .A1(n41629), .A2(n41628), .Z(n41640) );
  NAND2HSV0 U46079 ( .A1(n54078), .A2(n55100), .ZN(n54077) );
  OAI21HSV0 U46080 ( .A1(n44703), .A2(n41885), .B(n41630), .ZN(n41631) );
  OAI21HSV0 U46081 ( .A1(n41632), .A2(n54077), .B(n41631), .ZN(n41638) );
  NOR2HSV0 U46082 ( .A1(n41634), .A2(n41633), .ZN(n41636) );
  AOI22HSV0 U46083 ( .A1(n40683), .A2(n41424), .B1(n41743), .B2(\pe1/bq[18] ), 
        .ZN(n41635) );
  NOR2HSV1 U46084 ( .A1(n41636), .A2(n41635), .ZN(n41637) );
  XOR2HSV0 U46085 ( .A1(n41638), .A2(n41637), .Z(n41639) );
  XOR2HSV0 U46086 ( .A1(n41640), .A2(n41639), .Z(n41661) );
  CLKNAND2HSV0 U46087 ( .A1(n41877), .A2(\pe1/bq[12] ), .ZN(n41643) );
  NAND2HSV0 U46088 ( .A1(n44569), .A2(n41641), .ZN(n41642) );
  XOR2HSV0 U46089 ( .A1(n41643), .A2(n41642), .Z(n41649) );
  NAND2HSV0 U46090 ( .A1(n42220), .A2(n41644), .ZN(n41647) );
  CLKNAND2HSV0 U46091 ( .A1(n41964), .A2(n41645), .ZN(n41646) );
  XOR2HSV0 U46092 ( .A1(n41647), .A2(n41646), .Z(n41648) );
  XOR2HSV0 U46093 ( .A1(n41649), .A2(n41648), .Z(n41659) );
  NOR2HSV0 U46094 ( .A1(n41650), .A2(n53819), .ZN(n41652) );
  CLKNAND2HSV1 U46095 ( .A1(n41153), .A2(n42098), .ZN(n41651) );
  XOR2HSV0 U46096 ( .A1(n41652), .A2(n41651), .Z(n41657) );
  NAND2HSV2 U46097 ( .A1(n44533), .A2(n42231), .ZN(n41655) );
  CLKBUFHSV2 U46098 ( .I(\pe1/aot [11]), .Z(n55393) );
  NAND2HSV0 U46099 ( .A1(n55393), .A2(n40890), .ZN(n41654) );
  XOR2HSV0 U46100 ( .A1(n41655), .A2(n41654), .Z(n41656) );
  XOR2HSV0 U46101 ( .A1(n41657), .A2(n41656), .Z(n41658) );
  XOR2HSV0 U46102 ( .A1(n41659), .A2(n41658), .Z(n41660) );
  XOR4HSV1 U46103 ( .A1(n41663), .A2(n41662), .A3(n41661), .A4(n41660), .Z(
        n41665) );
  CLKNAND2HSV1 U46104 ( .A1(n59529), .A2(n54969), .ZN(n41664) );
  XNOR2HSV1 U46105 ( .A1(n41665), .A2(n41664), .ZN(n41667) );
  NAND2HSV2 U46106 ( .A1(n42275), .A2(n41550), .ZN(n41666) );
  XNOR2HSV1 U46107 ( .A1(n41667), .A2(n41666), .ZN(n41668) );
  XNOR2HSV1 U46108 ( .A1(n41669), .A2(n41668), .ZN(n41671) );
  CLKNAND2HSV1 U46109 ( .A1(n53602), .A2(n41851), .ZN(n41670) );
  XOR2HSV0 U46110 ( .A1(n41671), .A2(n41670), .Z(n41673) );
  NAND2HSV0 U46111 ( .A1(n42431), .A2(n42359), .ZN(n41672) );
  XOR2HSV0 U46112 ( .A1(n41673), .A2(n41672), .Z(n41674) );
  XNOR2HSV1 U46113 ( .A1(n41675), .A2(n41674), .ZN(n41679) );
  NAND2HSV0 U46114 ( .A1(n29773), .A2(n41676), .ZN(n41678) );
  XOR2HSV0 U46115 ( .A1(n41679), .A2(n41678), .Z(n41682) );
  NOR2HSV2 U46116 ( .A1(n41802), .A2(n48337), .ZN(n41681) );
  CLKNAND2HSV0 U46117 ( .A1(n41894), .A2(n54452), .ZN(n41680) );
  XOR3HSV2 U46118 ( .A1(n41682), .A2(n41681), .A3(n41680), .Z(n41683) );
  XNOR2HSV1 U46119 ( .A1(n41684), .A2(n41683), .ZN(n41685) );
  XOR2HSV0 U46120 ( .A1(n41686), .A2(n41685), .Z(n41688) );
  NAND2HSV0 U46121 ( .A1(n41733), .A2(\pe1/got [25]), .ZN(n41687) );
  XNOR2HSV1 U46122 ( .A1(n41688), .A2(n41687), .ZN(n41691) );
  CLKNAND2HSV1 U46123 ( .A1(n41850), .A2(n41689), .ZN(n41690) );
  XOR2HSV0 U46124 ( .A1(n41691), .A2(n41690), .Z(n41692) );
  XNOR2HSV4 U46125 ( .A1(n41693), .A2(n41692), .ZN(n41694) );
  NAND2HSV2 U46126 ( .A1(n26851), .A2(n54033), .ZN(n41696) );
  INHSV2 U46127 ( .I(n42196), .ZN(n42200) );
  CLKNAND2HSV1 U46128 ( .A1(n41697), .A2(n42200), .ZN(n41698) );
  INHSV4 U46129 ( .I(n41707), .ZN(n42029) );
  BUFHSV2 U46130 ( .I(n41708), .Z(n41700) );
  INHSV4 U46131 ( .I(n41707), .ZN(n41706) );
  NOR2HSV2 U46132 ( .A1(n41908), .A2(n41706), .ZN(n41726) );
  NAND2HSV0 U46133 ( .A1(n41707), .A2(n41701), .ZN(n41723) );
  CLKNAND2HSV0 U46134 ( .A1(n41723), .A2(n40541), .ZN(n41702) );
  NOR3HSV4 U46135 ( .A1(n41725), .A2(n41726), .A3(n41702), .ZN(n41703) );
  NAND2HSV2 U46136 ( .A1(n41707), .A2(n40407), .ZN(n41709) );
  NOR2HSV2 U46137 ( .A1(n41709), .A2(n41708), .ZN(n41715) );
  NAND2HSV4 U46138 ( .A1(n42029), .A2(n48320), .ZN(n41713) );
  NAND2HSV2 U46139 ( .A1(n41713), .A2(n41418), .ZN(n41710) );
  NOR3HSV2 U46140 ( .A1(n41716), .A2(n41715), .A3(n41710), .ZN(n41711) );
  NAND2HSV2 U46141 ( .A1(n42352), .A2(n59365), .ZN(n41841) );
  BUFHSV2 U46142 ( .I(n41841), .Z(n41835) );
  INHSV4 U46143 ( .I(n41713), .ZN(n41714) );
  NOR2HSV4 U46144 ( .A1(n41715), .A2(n41714), .ZN(n41718) );
  CLKNAND2HSV2 U46145 ( .A1(n41718), .A2(n41717), .ZN(n41719) );
  INHSV4 U46146 ( .I(n41914), .ZN(n41913) );
  CLKNHSV0 U46147 ( .I(\pe1/ti_7t [22]), .ZN(n41721) );
  AO21HSV1 U46148 ( .A1(n41721), .A2(n41720), .B(n41414), .Z(n41722) );
  CLKNHSV1 U46149 ( .I(n41723), .ZN(n41724) );
  NOR2HSV4 U46150 ( .A1(n41725), .A2(n41724), .ZN(n41729) );
  INHSV2 U46151 ( .I(n41726), .ZN(n41728) );
  INHSV4 U46152 ( .I(n41915), .ZN(n41730) );
  INHSV4 U46153 ( .I(n41730), .ZN(n41839) );
  CLKNAND2HSV2 U46154 ( .A1(n41840), .A2(n41839), .ZN(n41833) );
  NAND2HSV2 U46155 ( .A1(n41925), .A2(n59994), .ZN(n41820) );
  NAND2HSV2 U46156 ( .A1(n41927), .A2(n41731), .ZN(n41818) );
  NAND2HSV2 U46157 ( .A1(n59592), .A2(n59374), .ZN(n41816) );
  NOR2HSV2 U46158 ( .A1(n41732), .A2(n42086), .ZN(n41814) );
  NAND2HSV0 U46159 ( .A1(n41733), .A2(\pe1/got [24]), .ZN(n41812) );
  CLKNAND2HSV1 U46160 ( .A1(n41850), .A2(\pe1/got [25]), .ZN(n41811) );
  NAND2HSV2 U46161 ( .A1(n41734), .A2(\pe1/got [23]), .ZN(n41809) );
  CLKNAND2HSV0 U46162 ( .A1(n54041), .A2(n54452), .ZN(n41807) );
  CLKNAND2HSV0 U46163 ( .A1(n42089), .A2(n42359), .ZN(n41799) );
  CLKNAND2HSV1 U46164 ( .A1(n41609), .A2(n48339), .ZN(n41793) );
  NAND2HSV0 U46165 ( .A1(n41735), .A2(n42092), .ZN(n41887) );
  NOR2HSV0 U46166 ( .A1(n44705), .A2(n48030), .ZN(n53938) );
  AOI22HSV0 U46167 ( .A1(n59376), .A2(n54311), .B1(\pe1/bq[23] ), .B2(n41736), 
        .ZN(n41737) );
  AOI21HSV0 U46168 ( .A1(n41738), .A2(n53938), .B(n41737), .ZN(n41742) );
  NAND2HSV0 U46169 ( .A1(\pe1/aot [14]), .A2(n53922), .ZN(n41890) );
  INHSV2 U46170 ( .I(n41890), .ZN(n41740) );
  XOR2HSV0 U46171 ( .A1(n41740), .A2(n41739), .Z(n41741) );
  XOR3HSV1 U46172 ( .A1(n41887), .A2(n41742), .A3(n41741), .Z(n41787) );
  NOR2HSV0 U46173 ( .A1(n53833), .A2(n54973), .ZN(n41745) );
  NAND2HSV0 U46174 ( .A1(n41743), .A2(n42098), .ZN(n41744) );
  XOR2HSV0 U46175 ( .A1(n41745), .A2(n41744), .Z(n41749) );
  CLKNAND2HSV0 U46176 ( .A1(n59593), .A2(n42231), .ZN(n41747) );
  NAND2HSV0 U46177 ( .A1(\pe1/aot [10]), .A2(n41083), .ZN(n41746) );
  XOR2HSV0 U46178 ( .A1(n41747), .A2(n41746), .Z(n41748) );
  XOR2HSV0 U46179 ( .A1(n41749), .A2(n41748), .Z(n41756) );
  CLKNAND2HSV1 U46180 ( .A1(n44569), .A2(n54179), .ZN(n41751) );
  NAND2HSV0 U46181 ( .A1(n44566), .A2(\pe1/bq[10] ), .ZN(n41750) );
  XOR2HSV0 U46182 ( .A1(n41751), .A2(n41750), .Z(n41754) );
  NAND2HSV0 U46183 ( .A1(n41752), .A2(\pe1/got [11]), .ZN(n41753) );
  XOR2HSV0 U46184 ( .A1(n41754), .A2(n41753), .Z(n41755) );
  XOR2HSV0 U46185 ( .A1(n41756), .A2(n41755), .Z(n41786) );
  NAND2HSV0 U46186 ( .A1(n59990), .A2(n54479), .ZN(n42371) );
  BUFHSV2 U46187 ( .I(n40455), .Z(n53410) );
  OAI21HSV0 U46188 ( .A1(n42371), .A2(n41759), .B(n41758), .ZN(n41765) );
  NOR2HSV0 U46189 ( .A1(n54672), .A2(n41622), .ZN(n41762) );
  NAND2HSV0 U46190 ( .A1(n53812), .A2(n41760), .ZN(n53666) );
  OAI22HSV0 U46191 ( .A1(n41763), .A2(n41762), .B1(n41761), .B2(n53666), .ZN(
        n41764) );
  XOR2HSV0 U46192 ( .A1(n41765), .A2(n41764), .Z(n41766) );
  XNOR2HSV1 U46193 ( .A1(n41767), .A2(n41766), .ZN(n41785) );
  NAND2HSV0 U46194 ( .A1(n41768), .A2(n42106), .ZN(n41770) );
  NAND2HSV0 U46195 ( .A1(n54307), .A2(\pe1/bq[18] ), .ZN(n41769) );
  XOR2HSV0 U46196 ( .A1(n41770), .A2(n41769), .Z(n41775) );
  NAND2HSV0 U46197 ( .A1(n54663), .A2(\pe1/bq[21] ), .ZN(n41773) );
  NAND2HSV0 U46198 ( .A1(n42132), .A2(n41771), .ZN(n41772) );
  XOR2HSV0 U46199 ( .A1(n41773), .A2(n41772), .Z(n41774) );
  XOR2HSV0 U46200 ( .A1(n41775), .A2(n41774), .Z(n41783) );
  XOR2HSV0 U46201 ( .A1(n41777), .A2(n41776), .Z(n41781) );
  NAND2HSV0 U46202 ( .A1(n59989), .A2(\pe1/bq[26] ), .ZN(n41779) );
  NAND2HSV0 U46203 ( .A1(n40683), .A2(n53571), .ZN(n41778) );
  XOR2HSV0 U46204 ( .A1(n41779), .A2(n41778), .Z(n41780) );
  XOR2HSV0 U46205 ( .A1(n41781), .A2(n41780), .Z(n41782) );
  XOR2HSV0 U46206 ( .A1(n41783), .A2(n41782), .Z(n41784) );
  XOR4HSV1 U46207 ( .A1(n41787), .A2(n41786), .A3(n41785), .A4(n41784), .Z(
        n41789) );
  NAND2HSV0 U46208 ( .A1(n42210), .A2(n42155), .ZN(n41788) );
  XNOR2HSV1 U46209 ( .A1(n41789), .A2(n41788), .ZN(n41791) );
  CLKNAND2HSV0 U46210 ( .A1(n42275), .A2(n54969), .ZN(n41790) );
  XNOR2HSV1 U46211 ( .A1(n41791), .A2(n41790), .ZN(n41792) );
  XNOR2HSV1 U46212 ( .A1(n41793), .A2(n41792), .ZN(n41795) );
  CLKNAND2HSV0 U46213 ( .A1(n53602), .A2(n42162), .ZN(n41794) );
  XOR2HSV0 U46214 ( .A1(n41795), .A2(n41794), .Z(n41797) );
  NAND2HSV0 U46215 ( .A1(n54265), .A2(n41851), .ZN(n41796) );
  XOR2HSV0 U46216 ( .A1(n41797), .A2(n41796), .Z(n41798) );
  XNOR2HSV1 U46217 ( .A1(n41799), .A2(n41798), .ZN(n41801) );
  NAND2HSV0 U46218 ( .A1(n29773), .A2(n54728), .ZN(n41800) );
  XOR2HSV0 U46219 ( .A1(n41801), .A2(n41800), .Z(n41805) );
  NOR2HSV1 U46220 ( .A1(n41802), .A2(n48338), .ZN(n41804) );
  NAND2HSV0 U46221 ( .A1(n41894), .A2(\pe1/got [21]), .ZN(n41803) );
  XOR3HSV2 U46222 ( .A1(n41805), .A2(n41804), .A3(n41803), .Z(n41806) );
  XNOR2HSV1 U46223 ( .A1(n41807), .A2(n41806), .ZN(n41808) );
  XOR2HSV0 U46224 ( .A1(n41809), .A2(n41808), .Z(n41810) );
  XOR3HSV2 U46225 ( .A1(n41812), .A2(n41811), .A3(n41810), .Z(n41813) );
  XOR2HSV0 U46226 ( .A1(n41814), .A2(n41813), .Z(n41815) );
  XNOR2HSV1 U46227 ( .A1(n41816), .A2(n41815), .ZN(n41817) );
  XNOR2HSV4 U46228 ( .A1(n41820), .A2(n41819), .ZN(n41821) );
  XNOR2HSV4 U46229 ( .A1(n41822), .A2(n41821), .ZN(n41830) );
  AOI21HSV2 U46230 ( .A1(n41825), .A2(n25448), .B(n42070), .ZN(n41826) );
  OAI21HSV4 U46231 ( .A1(n41828), .A2(n41827), .B(n41826), .ZN(n41829) );
  NOR2HSV4 U46232 ( .A1(n41833), .A2(n41832), .ZN(n41834) );
  INOR2HSV4 U46233 ( .A1(n29726), .B1(n41834), .ZN(n41837) );
  NAND3HSV4 U46234 ( .A1(n41921), .A2(n41922), .A3(n41831), .ZN(n41836) );
  NOR2HSV4 U46235 ( .A1(n26888), .A2(n42082), .ZN(n41842) );
  NOR2HSV8 U46236 ( .A1(n41842), .A2(n41841), .ZN(n41845) );
  NAND2HSV2 U46237 ( .A1(n42316), .A2(n29735), .ZN(n52829) );
  NAND2HSV2 U46238 ( .A1(n52829), .A2(n42484), .ZN(n42347) );
  NAND2HSV2 U46239 ( .A1(n42355), .A2(n59365), .ZN(n41912) );
  NAND2HSV2 U46240 ( .A1(n41846), .A2(n53518), .ZN(n41911) );
  CLKNAND2HSV1 U46241 ( .A1(n41927), .A2(\pe1/got [27]), .ZN(n41905) );
  BUFHSV2 U46242 ( .I(n41848), .Z(n42207) );
  NOR2HSV2 U46243 ( .A1(n41849), .A2(n42207), .ZN(n41901) );
  NAND2HSV0 U46244 ( .A1(n59518), .A2(\pe1/got [23]), .ZN(n41899) );
  CLKNAND2HSV0 U46245 ( .A1(n41850), .A2(n41143), .ZN(n41898) );
  BUFHSV2 U46246 ( .I(n44696), .Z(n42088) );
  NAND2HSV2 U46247 ( .A1(n42088), .A2(n53390), .ZN(n41896) );
  INHSV2 U46248 ( .I(n41931), .ZN(n42399) );
  NAND2HSV2 U46249 ( .A1(n42399), .A2(\pe1/bq[23] ), .ZN(n41853) );
  CLKNAND2HSV0 U46250 ( .A1(n44569), .A2(n42373), .ZN(n41852) );
  XOR2HSV0 U46251 ( .A1(n41853), .A2(n41852), .Z(n41857) );
  NAND2HSV0 U46252 ( .A1(n42132), .A2(n40557), .ZN(n41855) );
  INHSV2 U46253 ( .I(n54846), .ZN(n53717) );
  NAND2HSV0 U46254 ( .A1(n53717), .A2(n42231), .ZN(n41854) );
  XOR2HSV0 U46255 ( .A1(n41855), .A2(n41854), .Z(n41856) );
  NAND2HSV0 U46256 ( .A1(n40898), .A2(n41641), .ZN(n41859) );
  CLKNAND2HSV1 U46257 ( .A1(n53848), .A2(n55100), .ZN(n41858) );
  XOR2HSV0 U46258 ( .A1(n41859), .A2(n41858), .Z(n41863) );
  NAND2HSV0 U46259 ( .A1(n59989), .A2(n42366), .ZN(n41861) );
  NAND2HSV0 U46260 ( .A1(n42093), .A2(\pe1/bq[21] ), .ZN(n41860) );
  XOR2HSV0 U46261 ( .A1(n41861), .A2(n41860), .Z(n41862) );
  NAND2HSV0 U46262 ( .A1(n53936), .A2(n53411), .ZN(n41865) );
  CLKNAND2HSV0 U46263 ( .A1(n40683), .A2(n54179), .ZN(n41864) );
  XOR2HSV0 U46264 ( .A1(n41865), .A2(n41864), .Z(n41869) );
  NAND2HSV0 U46265 ( .A1(\pe1/aot [24]), .A2(n54995), .ZN(n41867) );
  INHSV2 U46266 ( .I(n54472), .ZN(n54188) );
  NAND2HSV0 U46267 ( .A1(n54188), .A2(n41083), .ZN(n41866) );
  XOR2HSV0 U46268 ( .A1(n41867), .A2(n41866), .Z(n41868) );
  CLKNAND2HSV0 U46269 ( .A1(n41964), .A2(n54311), .ZN(n41872) );
  NAND2HSV0 U46270 ( .A1(n42220), .A2(n54479), .ZN(n41871) );
  XOR2HSV0 U46271 ( .A1(n41872), .A2(n41871), .Z(n41876) );
  NAND2HSV0 U46272 ( .A1(n42099), .A2(n42106), .ZN(n41873) );
  XOR2HSV0 U46273 ( .A1(n41874), .A2(n41873), .Z(n41875) );
  INHSV2 U46274 ( .I(n53723), .ZN(n55250) );
  NAND2HSV0 U46275 ( .A1(n41877), .A2(n55250), .ZN(n41879) );
  NAND2HSV0 U46276 ( .A1(n44566), .A2(\pe1/bq[9] ), .ZN(n41878) );
  XOR2HSV0 U46277 ( .A1(n41879), .A2(n41878), .Z(n41882) );
  BUFHSV2 U46278 ( .I(n41752), .Z(n59675) );
  CLKNAND2HSV0 U46279 ( .A1(n59675), .A2(n53473), .ZN(n41881) );
  XOR2HSV0 U46280 ( .A1(n41882), .A2(n41881), .Z(n41884) );
  NAND2HSV0 U46281 ( .A1(n53812), .A2(n42125), .ZN(n42365) );
  XOR2HSV0 U46282 ( .A1(n54074), .A2(n42365), .Z(n41891) );
  CLKNHSV0 U46283 ( .I(n41893), .ZN(n59919) );
  XOR2HSV0 U46284 ( .A1(n41896), .A2(n41895), .Z(n41897) );
  XOR3HSV2 U46285 ( .A1(n41899), .A2(n41898), .A3(n41897), .Z(n41900) );
  XOR2HSV0 U46286 ( .A1(n41901), .A2(n41900), .Z(n41902) );
  XNOR2HSV1 U46287 ( .A1(n41905), .A2(n41904), .ZN(n41906) );
  XOR2HSV0 U46288 ( .A1(n41907), .A2(n41906), .Z(n41910) );
  XNOR2HSV4 U46289 ( .A1(n41912), .A2(n42060), .ZN(n41918) );
  NAND2HSV2 U46290 ( .A1(n42352), .A2(n44523), .ZN(n41916) );
  XNOR2HSV4 U46291 ( .A1(n41918), .A2(n29754), .ZN(n60104) );
  INAND2HSV2 U46292 ( .A1(n41919), .B1(n29735), .ZN(n41920) );
  NAND2HSV2 U46293 ( .A1(n25448), .A2(\pe1/ti_7t [25]), .ZN(n42318) );
  CLKNAND2HSV0 U46294 ( .A1(n41922), .A2(n41921), .ZN(n41923) );
  NAND2HSV0 U46295 ( .A1(n41924), .A2(\pe1/ti_7t [23]), .ZN(n42203) );
  INHSV2 U46296 ( .I(n42203), .ZN(n42205) );
  INHSV2 U46297 ( .I(n42205), .ZN(n53655) );
  CLKNHSV0 U46298 ( .I(n42355), .ZN(n54037) );
  NAND2HSV0 U46299 ( .A1(n42085), .A2(n53520), .ZN(n42028) );
  BUFHSV4 U46300 ( .I(n41925), .Z(n59360) );
  INHSV2 U46301 ( .I(n59360), .ZN(n53391) );
  BUFHSV2 U46302 ( .I(n41926), .Z(n42087) );
  NOR2HSV2 U46303 ( .A1(n53391), .A2(n42087), .ZN(n42026) );
  BUFHSV2 U46304 ( .I(n41927), .Z(n42357) );
  NAND2HSV0 U46305 ( .A1(n42357), .A2(n53390), .ZN(n42024) );
  NAND2HSV2 U46306 ( .A1(n53392), .A2(n40886), .ZN(n42022) );
  NOR2HSV0 U46307 ( .A1(n41849), .A2(n48338), .ZN(n42020) );
  NAND2HSV0 U46308 ( .A1(n59518), .A2(\pe1/got [18]), .ZN(n42018) );
  NAND2HSV2 U46309 ( .A1(n54600), .A2(n54728), .ZN(n42017) );
  INHSV2 U46310 ( .I(n53911), .ZN(n54965) );
  NAND2HSV0 U46311 ( .A1(n53913), .A2(n54965), .ZN(n42015) );
  INHSV2 U46312 ( .I(n53793), .ZN(n54161) );
  NAND2HSV2 U46313 ( .A1(n54041), .A2(n54161), .ZN(n42013) );
  CLKNAND2HSV0 U46314 ( .A1(n41929), .A2(n55337), .ZN(n42006) );
  NAND2HSV0 U46315 ( .A1(n42360), .A2(n44605), .ZN(n42000) );
  BUFHSV2 U46316 ( .I(n41422), .Z(n53979) );
  CLKNHSV0 U46317 ( .I(n55019), .ZN(n42417) );
  CLKNAND2HSV1 U46318 ( .A1(n53979), .A2(n42417), .ZN(n41998) );
  BUFHSV2 U46319 ( .I(n59674), .Z(n53795) );
  NAND2HSV2 U46320 ( .A1(n53795), .A2(n55339), .ZN(n41997) );
  CLKNAND2HSV0 U46321 ( .A1(n41248), .A2(n53523), .ZN(n41935) );
  CLKNAND2HSV1 U46322 ( .A1(n54500), .A2(n54836), .ZN(n48365) );
  NAND2HSV0 U46323 ( .A1(n42093), .A2(\pe1/bq[18] ), .ZN(n42215) );
  OAI22HSV0 U46324 ( .A1(n41650), .A2(n45814), .B1(n41931), .B2(n41512), .ZN(
        n41932) );
  OAI21HSV1 U46325 ( .A1(n48365), .A2(n42215), .B(n41932), .ZN(n41933) );
  INHSV2 U46326 ( .I(n54472), .ZN(n54818) );
  CLKNAND2HSV0 U46327 ( .A1(n54818), .A2(n40494), .ZN(n53839) );
  XNOR2HSV1 U46328 ( .A1(n41933), .A2(n53839), .ZN(n41934) );
  XNOR2HSV1 U46329 ( .A1(n41935), .A2(n41934), .ZN(n41943) );
  NAND2HSV0 U46330 ( .A1(n54912), .A2(\pe1/bq[23] ), .ZN(n41937) );
  CLKNHSV0 U46331 ( .I(n54185), .ZN(n53578) );
  NAND2HSV0 U46332 ( .A1(n44533), .A2(n53578), .ZN(n41936) );
  XOR2HSV0 U46333 ( .A1(n41937), .A2(n41936), .Z(n41941) );
  CLKNAND2HSV1 U46334 ( .A1(n42132), .A2(\pe1/bq[21] ), .ZN(n41939) );
  NAND2HSV0 U46335 ( .A1(n53848), .A2(\pe1/bq[11] ), .ZN(n41938) );
  XOR2HSV0 U46336 ( .A1(n41939), .A2(n41938), .Z(n41940) );
  XOR2HSV0 U46337 ( .A1(n41941), .A2(n41940), .Z(n41942) );
  XNOR2HSV1 U46338 ( .A1(n41943), .A2(n41942), .ZN(n41962) );
  NAND2HSV0 U46339 ( .A1(n59987), .A2(n48380), .ZN(n41946) );
  INHSV2 U46340 ( .I(\pe1/aot [7]), .ZN(n42230) );
  NAND2HSV0 U46341 ( .A1(n54578), .A2(n42125), .ZN(n41945) );
  XOR2HSV0 U46342 ( .A1(n41946), .A2(n41945), .Z(n41951) );
  NAND2HSV0 U46343 ( .A1(n54904), .A2(n41623), .ZN(n41949) );
  CLKNAND2HSV0 U46344 ( .A1(\pe1/aot [14]), .A2(n42106), .ZN(n41948) );
  XOR2HSV0 U46345 ( .A1(n41949), .A2(n41948), .Z(n41950) );
  XOR2HSV0 U46346 ( .A1(n41951), .A2(n41950), .Z(n41960) );
  NAND2HSV0 U46347 ( .A1(n53717), .A2(n41644), .ZN(n41954) );
  CLKNHSV0 U46348 ( .I(n41952), .ZN(n48055) );
  NAND2HSV0 U46349 ( .A1(n59993), .A2(n48055), .ZN(n41953) );
  XOR2HSV0 U46350 ( .A1(n41954), .A2(n41953), .Z(n41958) );
  CLKNHSV0 U46351 ( .I(n44705), .ZN(n44556) );
  NAND2HSV0 U46352 ( .A1(n44556), .A2(n42098), .ZN(n41956) );
  NAND2HSV0 U46353 ( .A1(n54293), .A2(n55352), .ZN(n41955) );
  XOR2HSV0 U46354 ( .A1(n41956), .A2(n41955), .Z(n41957) );
  XOR2HSV0 U46355 ( .A1(n41958), .A2(n41957), .Z(n41959) );
  XOR2HSV0 U46356 ( .A1(n41960), .A2(n41959), .Z(n41961) );
  XOR2HSV0 U46357 ( .A1(n41962), .A2(n41961), .Z(n41995) );
  CLKNHSV0 U46358 ( .I(n54829), .ZN(n48396) );
  NAND2HSV0 U46359 ( .A1(n48396), .A2(n42092), .ZN(n41966) );
  NAND2HSV0 U46360 ( .A1(n41964), .A2(n55231), .ZN(n41965) );
  XOR2HSV0 U46361 ( .A1(n41966), .A2(n41965), .Z(n41971) );
  INHSV2 U46362 ( .I(n54901), .ZN(n59992) );
  NAND2HSV0 U46363 ( .A1(n59992), .A2(n53411), .ZN(n41969) );
  NAND2HSV0 U46364 ( .A1(\pe1/aot [4]), .A2(n40684), .ZN(n41968) );
  XOR2HSV0 U46365 ( .A1(n41969), .A2(n41968), .Z(n41970) );
  XOR2HSV0 U46366 ( .A1(n41971), .A2(n41970), .Z(n41980) );
  NOR2HSV0 U46367 ( .A1(n54673), .A2(n48060), .ZN(n41973) );
  NAND2HSV0 U46368 ( .A1(n40683), .A2(n53708), .ZN(n41972) );
  XOR2HSV0 U46369 ( .A1(n41973), .A2(n41972), .Z(n41978) );
  NAND2HSV0 U46370 ( .A1(n54307), .A2(n42373), .ZN(n41976) );
  NAND2HSV0 U46371 ( .A1(n54078), .A2(n53571), .ZN(n41975) );
  XOR2HSV0 U46372 ( .A1(n41976), .A2(n41975), .Z(n41977) );
  XOR2HSV0 U46373 ( .A1(n41978), .A2(n41977), .Z(n41979) );
  XOR2HSV0 U46374 ( .A1(n41980), .A2(n41979), .Z(n41993) );
  CLKNHSV0 U46375 ( .I(n40445), .ZN(n53673) );
  NAND2HSV0 U46376 ( .A1(n53673), .A2(\pe1/bq[5] ), .ZN(n41982) );
  BUFHSV2 U46377 ( .I(\pe1/bq[4] ), .Z(n54371) );
  NAND2HSV0 U46378 ( .A1(n44566), .A2(n54371), .ZN(n41981) );
  XOR2HSV0 U46379 ( .A1(n41982), .A2(n41981), .Z(n41986) );
  BUFHSV2 U46380 ( .I(\pe1/aot [11]), .Z(n53936) );
  NAND2HSV0 U46381 ( .A1(n53936), .A2(n42366), .ZN(n41984) );
  CLKNAND2HSV1 U46382 ( .A1(n53954), .A2(n54179), .ZN(n41983) );
  XOR2HSV0 U46383 ( .A1(n41984), .A2(n41983), .Z(n41985) );
  XOR2HSV0 U46384 ( .A1(n41986), .A2(n41985), .Z(n41991) );
  CLKNAND2HSV0 U46385 ( .A1(n41522), .A2(\pe1/got [5]), .ZN(n41989) );
  NAND2HSV0 U46386 ( .A1(n44569), .A2(\pe1/bq[9] ), .ZN(n42225) );
  INHSV2 U46387 ( .I(n54093), .ZN(n55394) );
  NAND2HSV0 U46388 ( .A1(n40898), .A2(n55394), .ZN(n48366) );
  OAI22HSV0 U46389 ( .A1(n53957), .A2(n54093), .B1(n53833), .B2(n55385), .ZN(
        n41987) );
  OAI21HSV0 U46390 ( .A1(n42225), .A2(n48366), .B(n41987), .ZN(n41988) );
  XOR2HSV0 U46391 ( .A1(n41989), .A2(n41988), .Z(n41990) );
  XOR2HSV0 U46392 ( .A1(n41991), .A2(n41990), .Z(n41992) );
  XOR2HSV0 U46393 ( .A1(n41993), .A2(n41992), .Z(n41994) );
  XOR2HSV0 U46394 ( .A1(n41995), .A2(n41994), .Z(n41996) );
  XOR3HSV2 U46395 ( .A1(n41998), .A2(n41997), .A3(n41996), .Z(n41999) );
  XNOR2HSV1 U46396 ( .A1(n42000), .A2(n41999), .ZN(n42002) );
  NAND2HSV0 U46397 ( .A1(n40917), .A2(n55088), .ZN(n42001) );
  XOR2HSV0 U46398 ( .A1(n42002), .A2(n42001), .Z(n42004) );
  NAND2HSV0 U46399 ( .A1(n54265), .A2(\pe1/got [11]), .ZN(n42003) );
  XOR2HSV0 U46400 ( .A1(n42004), .A2(n42003), .Z(n42005) );
  XNOR2HSV1 U46401 ( .A1(n42006), .A2(n42005), .ZN(n42008) );
  NAND2HSV0 U46402 ( .A1(n29762), .A2(n54812), .ZN(n42007) );
  XOR2HSV0 U46403 ( .A1(n42008), .A2(n42007), .Z(n42011) );
  CLKNHSV0 U46404 ( .I(n44532), .ZN(n42438) );
  NOR2HSV1 U46405 ( .A1(n42438), .A2(n54884), .ZN(n42010) );
  NAND2HSV0 U46406 ( .A1(n42439), .A2(n48339), .ZN(n42009) );
  XOR3HSV2 U46407 ( .A1(n42011), .A2(n42010), .A3(n42009), .Z(n42012) );
  XNOR2HSV1 U46408 ( .A1(n42013), .A2(n42012), .ZN(n42014) );
  XOR2HSV0 U46409 ( .A1(n42015), .A2(n42014), .Z(n42016) );
  XOR3HSV2 U46410 ( .A1(n42018), .A2(n42017), .A3(n42016), .Z(n42019) );
  XOR2HSV0 U46411 ( .A1(n42020), .A2(n42019), .Z(n42021) );
  XNOR2HSV1 U46412 ( .A1(n42022), .A2(n42021), .ZN(n42023) );
  XNOR2HSV1 U46413 ( .A1(n42024), .A2(n42023), .ZN(n42025) );
  XOR2HSV0 U46414 ( .A1(n42026), .A2(n42025), .Z(n42027) );
  INHSV3 U46415 ( .I(n25826), .ZN(n59377) );
  CLKNHSV1 U46416 ( .I(n59377), .ZN(n55018) );
  CLKNAND2HSV2 U46417 ( .A1(n42033), .A2(n53650), .ZN(n42030) );
  INAND2HSV2 U46418 ( .A1(n42031), .B1(n40482), .ZN(n42032) );
  INHSV2 U46419 ( .I(n42032), .ZN(n42034) );
  NAND2HSV2 U46420 ( .A1(n42034), .A2(n42033), .ZN(n42035) );
  CLKNAND2HSV0 U46421 ( .A1(n41720), .A2(\pe1/ti_7t [24]), .ZN(n42068) );
  CLKNAND2HSV1 U46422 ( .A1(n42069), .A2(n42068), .ZN(n42039) );
  INHSV2 U46423 ( .I(n42060), .ZN(n42072) );
  CLKNHSV0 U46424 ( .I(n42068), .ZN(n42038) );
  OAI22HSV1 U46425 ( .A1(n42049), .A2(n42039), .B1(n42072), .B2(n42038), .ZN(
        n42040) );
  INHSV2 U46426 ( .I(n42040), .ZN(n42048) );
  INHSV4 U46427 ( .I(n42069), .ZN(n42050) );
  INHSV2 U46428 ( .I(n42041), .ZN(n42054) );
  CLKNAND2HSV2 U46429 ( .A1(n42050), .A2(n42054), .ZN(n42046) );
  INOR2HSV1 U46430 ( .A1(n42471), .B1(n41242), .ZN(n42043) );
  CLKNHSV0 U46431 ( .I(n42043), .ZN(n42044) );
  CLKNAND2HSV0 U46432 ( .A1(n42060), .A2(n41129), .ZN(n42053) );
  NOR2HSV2 U46433 ( .A1(n42062), .A2(n42053), .ZN(n42055) );
  NAND2HSV2 U46434 ( .A1(n42054), .A2(n42069), .ZN(n42064) );
  INHSV3 U46435 ( .I(n42466), .ZN(n55144) );
  CLKNAND2HSV0 U46436 ( .A1(n42060), .A2(n42059), .ZN(n42061) );
  NOR2HSV2 U46437 ( .A1(n42062), .A2(n42061), .ZN(n42063) );
  INHSV2 U46438 ( .I(n42063), .ZN(n42066) );
  NOR2HSV1 U46439 ( .A1(n42068), .A2(n42067), .ZN(n42071) );
  INHSV2 U46440 ( .I(n42071), .ZN(n42076) );
  CLKAND2HSV1 U46441 ( .A1(n42069), .A2(n42076), .Z(n42074) );
  AOI21HSV2 U46442 ( .A1(n42072), .A2(n42471), .B(n42071), .ZN(n42073) );
  AOI21HSV2 U46443 ( .A1(n42075), .A2(n42074), .B(n42073), .ZN(n42079) );
  CLKNAND2HSV1 U46444 ( .A1(n42077), .A2(n42076), .ZN(n42078) );
  AOI22HSV4 U46445 ( .A1(n42081), .A2(n42080), .B1(n42078), .B2(n42079), .ZN(
        n42325) );
  NAND2HSV1 U46446 ( .A1(n42352), .A2(n53518), .ZN(n42083) );
  CLKNAND2HSV1 U46447 ( .A1(n42355), .A2(n42084), .ZN(n42185) );
  NOR2HSV2 U46448 ( .A1(n42356), .A2(n42086), .ZN(n42182) );
  NAND2HSV2 U46449 ( .A1(n42357), .A2(n41201), .ZN(n42180) );
  CLKNAND2HSV1 U46450 ( .A1(n42358), .A2(n53520), .ZN(n42178) );
  NOR2HSV2 U46451 ( .A1(n41849), .A2(n42087), .ZN(n42176) );
  NAND2HSV0 U46452 ( .A1(n59518), .A2(\pe1/got [21]), .ZN(n42174) );
  NAND2HSV2 U46453 ( .A1(n54600), .A2(n53390), .ZN(n42173) );
  NAND2HSV0 U46454 ( .A1(n42088), .A2(n44530), .ZN(n42171) );
  NAND2HSV0 U46455 ( .A1(n54264), .A2(n59995), .ZN(n42169) );
  NAND2HSV0 U46456 ( .A1(n42089), .A2(n41550), .ZN(n42161) );
  CLKNAND2HSV1 U46457 ( .A1(n42360), .A2(n55337), .ZN(n42154) );
  CLKNAND2HSV1 U46458 ( .A1(n59529), .A2(n53473), .ZN(n42152) );
  CLKNAND2HSV0 U46459 ( .A1(\pe1/aot [16]), .A2(\pe1/bq[23] ), .ZN(n42091) );
  NAND2HSV0 U46460 ( .A1(n59987), .A2(\pe1/bq[18] ), .ZN(n42090) );
  XOR2HSV0 U46461 ( .A1(n42091), .A2(n42090), .Z(n42097) );
  NAND2HSV0 U46462 ( .A1(n42093), .A2(n42092), .ZN(n42095) );
  NAND2HSV0 U46463 ( .A1(n54307), .A2(n41424), .ZN(n42094) );
  XOR2HSV0 U46464 ( .A1(n42095), .A2(n42094), .Z(n42096) );
  XOR2HSV0 U46465 ( .A1(n42097), .A2(n42096), .Z(n42105) );
  CLKNAND2HSV1 U46466 ( .A1(n41964), .A2(\pe1/bq[9] ), .ZN(n53413) );
  NAND2HSV0 U46467 ( .A1(n54078), .A2(n42098), .ZN(n54189) );
  XOR2HSV0 U46468 ( .A1(n53413), .A2(n54189), .Z(n42103) );
  CLKNAND2HSV1 U46469 ( .A1(n54912), .A2(n41644), .ZN(n42101) );
  NAND2HSV0 U46470 ( .A1(n42099), .A2(n42238), .ZN(n42100) );
  XOR2HSV0 U46471 ( .A1(n42101), .A2(n42100), .Z(n42102) );
  XOR2HSV0 U46472 ( .A1(n42103), .A2(n42102), .Z(n42104) );
  XOR2HSV0 U46473 ( .A1(n42105), .A2(n42104), .Z(n42122) );
  NAND2HSV0 U46474 ( .A1(n42220), .A2(n42106), .ZN(n42108) );
  NAND2HSV0 U46475 ( .A1(n53812), .A2(n41771), .ZN(n42107) );
  XOR2HSV0 U46476 ( .A1(n42108), .A2(n42107), .Z(n42112) );
  CLKNAND2HSV0 U46477 ( .A1(n59593), .A2(n53805), .ZN(n42110) );
  NAND2HSV0 U46478 ( .A1(n40898), .A2(n42373), .ZN(n42109) );
  XOR2HSV0 U46479 ( .A1(n42110), .A2(n42109), .Z(n42111) );
  XOR2HSV0 U46480 ( .A1(n42112), .A2(n42111), .Z(n42120) );
  NAND2HSV0 U46481 ( .A1(n41153), .A2(\pe1/bq[13] ), .ZN(n42114) );
  NAND2HSV0 U46482 ( .A1(\pe1/aot [8]), .A2(n42231), .ZN(n42113) );
  XOR2HSV0 U46483 ( .A1(n42114), .A2(n42113), .Z(n42118) );
  CLKNAND2HSV1 U46484 ( .A1(n53848), .A2(n53571), .ZN(n42116) );
  INHSV2 U46485 ( .I(\pe1/aot [7]), .ZN(n42362) );
  INHSV2 U46486 ( .I(n42362), .ZN(n55547) );
  NAND2HSV0 U46487 ( .A1(n55547), .A2(n40890), .ZN(n42115) );
  XOR2HSV0 U46488 ( .A1(n42116), .A2(n42115), .Z(n42117) );
  XOR2HSV0 U46489 ( .A1(n42118), .A2(n42117), .Z(n42119) );
  XOR2HSV0 U46490 ( .A1(n42120), .A2(n42119), .Z(n42121) );
  XOR2HSV0 U46491 ( .A1(n42122), .A2(n42121), .Z(n42149) );
  CLKNAND2HSV0 U46492 ( .A1(n42255), .A2(n55100), .ZN(n42124) );
  NAND2HSV0 U46493 ( .A1(n44569), .A2(n55250), .ZN(n42123) );
  XOR2HSV0 U46494 ( .A1(n42124), .A2(n42123), .Z(n42129) );
  INHSV2 U46495 ( .I(n54846), .ZN(n59991) );
  NAND2HSV0 U46496 ( .A1(n59991), .A2(n42125), .ZN(n42127) );
  NAND2HSV0 U46497 ( .A1(n54818), .A2(n53411), .ZN(n42126) );
  XOR2HSV0 U46498 ( .A1(n42127), .A2(n42126), .Z(n42128) );
  XOR2HSV0 U46499 ( .A1(n42129), .A2(n42128), .Z(n42138) );
  NAND2HSV0 U46500 ( .A1(n40683), .A2(n54311), .ZN(n42131) );
  NAND2HSV0 U46501 ( .A1(\pe1/aot [14]), .A2(n54319), .ZN(n42130) );
  XOR2HSV0 U46502 ( .A1(n42131), .A2(n42130), .Z(n42136) );
  NAND2HSV0 U46503 ( .A1(n42132), .A2(n54479), .ZN(n42134) );
  NAND2HSV0 U46504 ( .A1(n42399), .A2(\pe1/bq[21] ), .ZN(n42133) );
  XOR2HSV0 U46505 ( .A1(n42134), .A2(n42133), .Z(n42135) );
  XOR2HSV0 U46506 ( .A1(n42136), .A2(n42135), .Z(n42137) );
  XOR2HSV0 U46507 ( .A1(n42138), .A2(n42137), .Z(n42147) );
  NAND2HSV0 U46508 ( .A1(n42139), .A2(n55394), .ZN(n42141) );
  CLKNAND2HSV0 U46509 ( .A1(n53673), .A2(n53708), .ZN(n42140) );
  XOR2HSV0 U46510 ( .A1(n42141), .A2(n42140), .Z(n42143) );
  NAND2HSV0 U46511 ( .A1(n59675), .A2(\pe1/got [8]), .ZN(n42142) );
  XOR2HSV0 U46512 ( .A1(n42143), .A2(n42142), .Z(n42145) );
  XNOR2HSV1 U46513 ( .A1(n42145), .A2(n42144), .ZN(n42146) );
  XNOR2HSV1 U46514 ( .A1(n42147), .A2(n42146), .ZN(n42148) );
  XNOR2HSV1 U46515 ( .A1(n42149), .A2(n42148), .ZN(n42151) );
  NAND2HSV0 U46516 ( .A1(n42275), .A2(n55214), .ZN(n42150) );
  XOR3HSV2 U46517 ( .A1(n42152), .A2(n42151), .A3(n42150), .Z(n42153) );
  XNOR2HSV1 U46518 ( .A1(n42154), .A2(n42153), .ZN(n42157) );
  NAND2HSV0 U46519 ( .A1(n53602), .A2(n42155), .ZN(n42156) );
  XOR2HSV0 U46520 ( .A1(n42157), .A2(n42156), .Z(n42159) );
  NAND2HSV0 U46521 ( .A1(n59919), .A2(n54969), .ZN(n42158) );
  XOR2HSV0 U46522 ( .A1(n42159), .A2(n42158), .Z(n42160) );
  XNOR2HSV1 U46523 ( .A1(n42161), .A2(n42160), .ZN(n42164) );
  NAND2HSV0 U46524 ( .A1(n29763), .A2(n42162), .ZN(n42163) );
  XOR2HSV0 U46525 ( .A1(n42164), .A2(n42163), .Z(n42167) );
  NOR2HSV2 U46526 ( .A1(n42438), .A2(n53911), .ZN(n42166) );
  NAND2HSV0 U46527 ( .A1(n42439), .A2(n42359), .ZN(n42165) );
  XOR3HSV2 U46528 ( .A1(n42167), .A2(n42166), .A3(n42165), .Z(n42168) );
  XNOR2HSV1 U46529 ( .A1(n42169), .A2(n42168), .ZN(n42170) );
  XOR2HSV0 U46530 ( .A1(n42171), .A2(n42170), .Z(n42172) );
  XOR3HSV2 U46531 ( .A1(n42174), .A2(n42173), .A3(n42172), .Z(n42175) );
  XOR2HSV0 U46532 ( .A1(n42176), .A2(n42175), .Z(n42177) );
  XNOR2HSV1 U46533 ( .A1(n42178), .A2(n42177), .ZN(n42179) );
  XNOR2HSV1 U46534 ( .A1(n42180), .A2(n42179), .ZN(n42181) );
  XOR2HSV0 U46535 ( .A1(n42182), .A2(n42181), .Z(n42183) );
  OAI22HSV4 U46536 ( .A1(n42186), .A2(n29760), .B1(n44522), .B2(n42318), .ZN(
        n42322) );
  CLKAND2HSV2 U46537 ( .A1(n41056), .A2(\pe1/ti_7t [26]), .Z(n42191) );
  NOR2HSV1 U46538 ( .A1(n42322), .A2(n42191), .ZN(n42190) );
  CLKNHSV0 U46539 ( .I(n42323), .ZN(n42189) );
  NOR2HSV2 U46540 ( .A1(n42191), .A2(n41134), .ZN(n42188) );
  AOI31HSV2 U46541 ( .A1(n42320), .A2(n42190), .A3(n42189), .B(n42188), .ZN(
        n42195) );
  NOR2HSV4 U46542 ( .A1(n42322), .A2(n42323), .ZN(n42329) );
  CLKNHSV2 U46543 ( .I(n42329), .ZN(n42193) );
  CLKNAND2HSV3 U46544 ( .A1(n42195), .A2(n42194), .ZN(n48451) );
  INHSV2 U46545 ( .I(n42198), .ZN(n42199) );
  AOI21HSV2 U46546 ( .A1(n42203), .A2(n41924), .B(n41507), .ZN(n42204) );
  OAI21HSV2 U46547 ( .A1(pov1[23]), .A2(n42205), .B(n42204), .ZN(n42314) );
  CLKNAND2HSV0 U46548 ( .A1(n42355), .A2(\pe1/got [28]), .ZN(n42312) );
  CLKNHSV2 U46549 ( .I(n42206), .ZN(n59391) );
  CLKNAND2HSV1 U46550 ( .A1(n42085), .A2(n40605), .ZN(n42308) );
  INHSV2 U46551 ( .I(n59360), .ZN(n42208) );
  NOR2HSV2 U46552 ( .A1(n42208), .A2(n42207), .ZN(n42306) );
  CLKNAND2HSV1 U46553 ( .A1(n42357), .A2(n53520), .ZN(n42304) );
  CLKNAND2HSV0 U46554 ( .A1(n42358), .A2(\pe1/got [23]), .ZN(n42302) );
  NOR2HSV2 U46555 ( .A1(n41849), .A2(n42209), .ZN(n42300) );
  NAND2HSV0 U46556 ( .A1(n59518), .A2(n44530), .ZN(n42298) );
  CLKNAND2HSV1 U46557 ( .A1(n54600), .A2(n40886), .ZN(n42297) );
  INHSV4 U46558 ( .I(n41928), .ZN(n54728) );
  NAND2HSV0 U46559 ( .A1(n53913), .A2(n54728), .ZN(n42295) );
  NAND2HSV0 U46560 ( .A1(n54264), .A2(n42359), .ZN(n42293) );
  CLKNAND2HSV1 U46561 ( .A1(n42089), .A2(n54969), .ZN(n42286) );
  CLKNAND2HSV0 U46562 ( .A1(n42360), .A2(n55214), .ZN(n42280) );
  NAND2HSV0 U46563 ( .A1(n42210), .A2(n44605), .ZN(n42278) );
  NAND2HSV2 U46564 ( .A1(n42132), .A2(n54911), .ZN(n54558) );
  OAI21HSV0 U46565 ( .A1(n41076), .A2(n54735), .B(n42211), .ZN(n42213) );
  OAI21HSV0 U46566 ( .A1(n42214), .A2(n54558), .B(n42213), .ZN(n42216) );
  XNOR2HSV1 U46567 ( .A1(n42216), .A2(n42215), .ZN(n42219) );
  XOR2HSV0 U46568 ( .A1(n54077), .A2(n42217), .Z(n42218) );
  XNOR2HSV1 U46569 ( .A1(n42219), .A2(n42218), .ZN(n42229) );
  NAND2HSV0 U46570 ( .A1(n42220), .A2(\pe1/bq[21] ), .ZN(n42222) );
  NAND2HSV0 U46571 ( .A1(n53717), .A2(n53805), .ZN(n42221) );
  XOR2HSV0 U46572 ( .A1(n42222), .A2(n42221), .Z(n42227) );
  NAND2HSV0 U46573 ( .A1(n54188), .A2(n42223), .ZN(n42224) );
  XOR2HSV0 U46574 ( .A1(n42225), .A2(n42224), .Z(n42226) );
  XOR2HSV0 U46575 ( .A1(n42227), .A2(n42226), .Z(n42228) );
  XOR2HSV0 U46576 ( .A1(n42229), .A2(n42228), .Z(n42248) );
  NAND2HSV0 U46577 ( .A1(n54578), .A2(n42231), .ZN(n42233) );
  CLKNAND2HSV0 U46578 ( .A1(n44556), .A2(n42092), .ZN(n42232) );
  XOR2HSV0 U46579 ( .A1(n42233), .A2(n42232), .Z(n42237) );
  NAND2HSV0 U46580 ( .A1(n59985), .A2(n53708), .ZN(n42235) );
  NAND2HSV0 U46581 ( .A1(n44533), .A2(n40557), .ZN(n42234) );
  XOR2HSV0 U46582 ( .A1(n42235), .A2(n42234), .Z(n42236) );
  XOR2HSV0 U46583 ( .A1(n42237), .A2(n42236), .Z(n42246) );
  NAND2HSV0 U46584 ( .A1(n42399), .A2(n42238), .ZN(n42240) );
  NAND2HSV0 U46585 ( .A1(\pe1/aot [27]), .A2(n54311), .ZN(n42239) );
  XOR2HSV0 U46586 ( .A1(n42240), .A2(n42239), .Z(n42244) );
  CLKNAND2HSV1 U46587 ( .A1(n59989), .A2(n54465), .ZN(n42242) );
  NAND2HSV0 U46588 ( .A1(\pe1/aot [14]), .A2(n53578), .ZN(n42241) );
  XOR2HSV0 U46589 ( .A1(n42242), .A2(n42241), .Z(n42243) );
  XOR2HSV0 U46590 ( .A1(n42244), .A2(n42243), .Z(n42245) );
  XOR2HSV0 U46591 ( .A1(n42246), .A2(n42245), .Z(n42247) );
  XOR2HSV0 U46592 ( .A1(n42248), .A2(n42247), .Z(n42274) );
  NAND2HSV0 U46593 ( .A1(\pe1/aot [8]), .A2(n25428), .ZN(n42250) );
  INHSV2 U46594 ( .I(n54093), .ZN(n55045) );
  CLKNAND2HSV0 U46595 ( .A1(n53673), .A2(n55045), .ZN(n42249) );
  XOR2HSV0 U46596 ( .A1(n42250), .A2(n42249), .Z(n42254) );
  NAND2HSV0 U46597 ( .A1(n54293), .A2(n42373), .ZN(n42252) );
  NAND2HSV0 U46598 ( .A1(n54307), .A2(n53571), .ZN(n42251) );
  XOR2HSV0 U46599 ( .A1(n42252), .A2(n42251), .Z(n42253) );
  XOR2HSV0 U46600 ( .A1(n42254), .A2(n42253), .Z(n42263) );
  CLKNAND2HSV1 U46601 ( .A1(n53848), .A2(n41645), .ZN(n42257) );
  NAND2HSV0 U46602 ( .A1(n42255), .A2(n41424), .ZN(n42256) );
  XOR2HSV0 U46603 ( .A1(n42257), .A2(n42256), .Z(n42261) );
  NAND2HSV0 U46604 ( .A1(n59593), .A2(n41771), .ZN(n42259) );
  CLKNAND2HSV0 U46605 ( .A1(n59987), .A2(n42098), .ZN(n42258) );
  XOR2HSV0 U46606 ( .A1(n42259), .A2(n42258), .Z(n42260) );
  XOR2HSV0 U46607 ( .A1(n42261), .A2(n42260), .Z(n42262) );
  XOR2HSV0 U46608 ( .A1(n42263), .A2(n42262), .Z(n42272) );
  CLKNAND2HSV1 U46609 ( .A1(n41522), .A2(n42417), .ZN(n42268) );
  INHSV2 U46610 ( .I(n54901), .ZN(n55492) );
  NAND2HSV0 U46611 ( .A1(n55492), .A2(n54319), .ZN(n53409) );
  OAI22HSV0 U46612 ( .A1(n41967), .A2(n54901), .B1(n53672), .B2(n42264), .ZN(
        n42265) );
  OAI21HSV0 U46613 ( .A1(n42266), .A2(n53409), .B(n42265), .ZN(n42267) );
  XOR2HSV0 U46614 ( .A1(n42268), .A2(n42267), .Z(n42270) );
  NAND2HSV0 U46615 ( .A1(n41160), .A2(n55339), .ZN(n42269) );
  XOR2HSV0 U46616 ( .A1(n42270), .A2(n42269), .Z(n42271) );
  XNOR2HSV1 U46617 ( .A1(n42272), .A2(n42271), .ZN(n42273) );
  XNOR2HSV1 U46618 ( .A1(n42274), .A2(n42273), .ZN(n42277) );
  NAND2HSV0 U46619 ( .A1(n42275), .A2(n53473), .ZN(n42276) );
  XOR3HSV2 U46620 ( .A1(n42278), .A2(n42277), .A3(n42276), .Z(n42279) );
  XNOR2HSV1 U46621 ( .A1(n42280), .A2(n42279), .ZN(n42282) );
  NAND2HSV0 U46622 ( .A1(n53602), .A2(n55337), .ZN(n42281) );
  XOR2HSV0 U46623 ( .A1(n42282), .A2(n42281), .Z(n42284) );
  NAND2HSV0 U46624 ( .A1(n54265), .A2(\pe1/got [13]), .ZN(n42283) );
  XOR2HSV0 U46625 ( .A1(n42284), .A2(n42283), .Z(n42285) );
  XNOR2HSV1 U46626 ( .A1(n42286), .A2(n42285), .ZN(n42288) );
  NAND2HSV0 U46627 ( .A1(n29763), .A2(\pe1/got [15]), .ZN(n42287) );
  XOR2HSV0 U46628 ( .A1(n42288), .A2(n42287), .Z(n42291) );
  NOR2HSV1 U46629 ( .A1(n42438), .A2(n53793), .ZN(n42290) );
  INHSV2 U46630 ( .I(n53911), .ZN(n54135) );
  NAND2HSV0 U46631 ( .A1(n42439), .A2(n54135), .ZN(n42289) );
  XOR3HSV2 U46632 ( .A1(n42291), .A2(n42290), .A3(n42289), .Z(n42292) );
  XNOR2HSV1 U46633 ( .A1(n42293), .A2(n42292), .ZN(n42294) );
  XOR2HSV0 U46634 ( .A1(n42295), .A2(n42294), .Z(n42296) );
  XOR3HSV2 U46635 ( .A1(n42298), .A2(n42297), .A3(n42296), .Z(n42299) );
  XOR2HSV0 U46636 ( .A1(n42300), .A2(n42299), .Z(n42301) );
  XNOR2HSV1 U46637 ( .A1(n42302), .A2(n42301), .ZN(n42303) );
  XNOR2HSV1 U46638 ( .A1(n42304), .A2(n42303), .ZN(n42305) );
  XOR2HSV0 U46639 ( .A1(n42306), .A2(n42305), .Z(n42307) );
  XNOR2HSV1 U46640 ( .A1(n42308), .A2(n42307), .ZN(n42310) );
  CLKNAND2HSV1 U46641 ( .A1(n59377), .A2(\pe1/got [27]), .ZN(n42309) );
  XOR2HSV0 U46642 ( .A1(n42310), .A2(n42309), .Z(n42311) );
  NOR2HSV1 U46643 ( .A1(n42318), .A2(n42037), .ZN(n42319) );
  XNOR2HSV4 U46644 ( .A1(n42337), .A2(n42336), .ZN(n42343) );
  NOR2HSV2 U46645 ( .A1(n42323), .A2(n42322), .ZN(n42326) );
  XNOR2HSV4 U46646 ( .A1(n42325), .A2(n42324), .ZN(n42330) );
  AND2HSV2 U46647 ( .A1(n42471), .A2(n42488), .Z(n42327) );
  NOR2HSV4 U46648 ( .A1(n42330), .A2(n42329), .ZN(n44651) );
  CLKNAND2HSV1 U46649 ( .A1(n41056), .A2(\pe1/ti_7t [27]), .ZN(n42490) );
  CLKNHSV1 U46650 ( .I(n42490), .ZN(n42340) );
  INHSV2 U46651 ( .I(n44524), .ZN(n48321) );
  NAND2HSV2 U46652 ( .A1(n48325), .A2(n48321), .ZN(n42482) );
  CLKNAND2HSV1 U46653 ( .A1(n42340), .A2(n42339), .ZN(n42341) );
  NAND2HSV2 U46654 ( .A1(n42489), .A2(n48468), .ZN(n42342) );
  NOR2HSV4 U46655 ( .A1(n48329), .A2(n42344), .ZN(n45782) );
  CLKNAND2HSV1 U46656 ( .A1(n29760), .A2(n59394), .ZN(n42348) );
  NOR2HSV2 U46657 ( .A1(n42347), .A2(n42348), .ZN(n42349) );
  INHSV2 U46658 ( .I(n42349), .ZN(n42350) );
  NAND2HSV0 U46659 ( .A1(n42352), .A2(n40873), .ZN(n42353) );
  NOR2HSV2 U46660 ( .A1(n42354), .A2(n42353), .ZN(n42465) );
  NAND2HSV0 U46661 ( .A1(n42355), .A2(n59374), .ZN(n42463) );
  NAND2HSV2 U46662 ( .A1(n42085), .A2(\pe1/got [25]), .ZN(n42459) );
  NOR2HSV1 U46663 ( .A1(n42356), .A2(n41392), .ZN(n42457) );
  CLKNAND2HSV0 U46664 ( .A1(n42357), .A2(\pe1/got [23]), .ZN(n42455) );
  CLKNAND2HSV0 U46665 ( .A1(n42358), .A2(n54160), .ZN(n42453) );
  NOR2HSV1 U46666 ( .A1(n54040), .A2(n48337), .ZN(n42451) );
  NAND2HSV0 U46667 ( .A1(n59518), .A2(n59995), .ZN(n42449) );
  CLKNAND2HSV0 U46668 ( .A1(n54600), .A2(n44530), .ZN(n42448) );
  CLKNAND2HSV1 U46669 ( .A1(n53913), .A2(n42359), .ZN(n42446) );
  CLKNHSV2 U46670 ( .I(n53911), .ZN(n59996) );
  NAND2HSV0 U46671 ( .A1(n54264), .A2(n59996), .ZN(n42444) );
  CLKNAND2HSV0 U46672 ( .A1(n42089), .A2(\pe1/got [13]), .ZN(n42435) );
  NAND2HSV0 U46673 ( .A1(n42360), .A2(n55088), .ZN(n42428) );
  NAND2HSV0 U46674 ( .A1(n41549), .A2(n55339), .ZN(n42426) );
  NOR2HSV0 U46675 ( .A1(n42361), .A2(n48393), .ZN(n54384) );
  CLKNAND2HSV1 U46676 ( .A1(n44556), .A2(\pe1/bq[18] ), .ZN(n54823) );
  XOR2HSV0 U46677 ( .A1(n54384), .A2(n54823), .Z(n42380) );
  NOR2HSV0 U46678 ( .A1(n55307), .A2(n41425), .ZN(n48342) );
  AOI22HSV0 U46679 ( .A1(n59991), .A2(n41771), .B1(n53411), .B2(n55547), .ZN(
        n42363) );
  AOI21HSV0 U46680 ( .A1(n42364), .A2(n48342), .B(n42363), .ZN(n42370) );
  NAND2HSV0 U46681 ( .A1(\pe1/aot [8]), .A2(n53718), .ZN(n53535) );
  NOR2HSV0 U46682 ( .A1(n42365), .A2(n53535), .ZN(n42368) );
  AOI22HSV0 U46683 ( .A1(\pe1/aot [12]), .A2(n42366), .B1(n42125), .B2(
        \pe1/aot [8]), .ZN(n42367) );
  NOR2HSV1 U46684 ( .A1(n42368), .A2(n42367), .ZN(n42369) );
  XOR2HSV0 U46685 ( .A1(n42370), .A2(n42369), .Z(n42379) );
  XOR2HSV0 U46686 ( .A1(n42372), .A2(n42371), .Z(n42377) );
  CLKNAND2HSV0 U46687 ( .A1(n53848), .A2(n42373), .ZN(n42374) );
  XOR2HSV0 U46688 ( .A1(n42375), .A2(n42374), .Z(n42376) );
  XOR2HSV0 U46689 ( .A1(n42377), .A2(n42376), .Z(n42378) );
  XOR3HSV2 U46690 ( .A1(n42380), .A2(n42379), .A3(n42378), .Z(n42396) );
  NAND2HSV0 U46691 ( .A1(n59992), .A2(n48055), .ZN(n42382) );
  NAND2HSV0 U46692 ( .A1(\pe1/aot [27]), .A2(n55250), .ZN(n42381) );
  XOR2HSV0 U46693 ( .A1(n42382), .A2(n42381), .Z(n42386) );
  CLKNAND2HSV0 U46694 ( .A1(n53936), .A2(n41644), .ZN(n42384) );
  NAND2HSV0 U46695 ( .A1(n59987), .A2(n55100), .ZN(n42383) );
  XOR2HSV0 U46696 ( .A1(n42384), .A2(n42383), .Z(n42385) );
  XOR2HSV0 U46697 ( .A1(n42386), .A2(n42385), .Z(n42394) );
  NOR2HSV0 U46698 ( .A1(n46142), .A2(n54281), .ZN(n42388) );
  CLKNAND2HSV1 U46699 ( .A1(n41768), .A2(n42098), .ZN(n42387) );
  XOR2HSV0 U46700 ( .A1(n42388), .A2(n42387), .Z(n42392) );
  NAND2HSV0 U46701 ( .A1(\pe1/aot [14]), .A2(\pe1/bq[23] ), .ZN(n42390) );
  NAND2HSV0 U46702 ( .A1(n41169), .A2(n41424), .ZN(n42389) );
  XOR2HSV0 U46703 ( .A1(n42390), .A2(n42389), .Z(n42391) );
  XOR2HSV0 U46704 ( .A1(n42392), .A2(n42391), .Z(n42393) );
  XOR2HSV0 U46705 ( .A1(n42394), .A2(n42393), .Z(n42395) );
  XOR2HSV0 U46706 ( .A1(n42396), .A2(n42395), .Z(n42423) );
  CLKNAND2HSV0 U46707 ( .A1(n54307), .A2(n41645), .ZN(n42398) );
  NAND2HSV0 U46708 ( .A1(\pe1/aot [26]), .A2(n55166), .ZN(n42397) );
  XOR2HSV0 U46709 ( .A1(n42398), .A2(n42397), .Z(n42403) );
  CLKNAND2HSV0 U46710 ( .A1(n42399), .A2(n42092), .ZN(n42401) );
  NAND2HSV0 U46711 ( .A1(n40683), .A2(\pe1/bq[9] ), .ZN(n42400) );
  XOR2HSV0 U46712 ( .A1(n42401), .A2(n42400), .Z(n42402) );
  XOR2HSV0 U46713 ( .A1(n42403), .A2(n42402), .Z(n42411) );
  NAND2HSV2 U46714 ( .A1(n48396), .A2(n54565), .ZN(n42405) );
  NAND2HSV0 U46715 ( .A1(n55553), .A2(n40890), .ZN(n42404) );
  XOR2HSV0 U46716 ( .A1(n42405), .A2(n42404), .Z(n42409) );
  NAND2HSV0 U46717 ( .A1(n41964), .A2(n55045), .ZN(n42407) );
  NAND2HSV0 U46718 ( .A1(n54818), .A2(n53805), .ZN(n42406) );
  XOR2HSV0 U46719 ( .A1(n42407), .A2(n42406), .Z(n42408) );
  XOR2HSV0 U46720 ( .A1(n42409), .A2(n42408), .Z(n42410) );
  XOR2HSV0 U46721 ( .A1(n42411), .A2(n42410), .Z(n42421) );
  NAND2HSV0 U46722 ( .A1(n42412), .A2(n54911), .ZN(n42414) );
  NAND2HSV0 U46723 ( .A1(n44566), .A2(\pe1/bq[5] ), .ZN(n42413) );
  XOR2HSV0 U46724 ( .A1(n42414), .A2(n42413), .Z(n42416) );
  CLKNAND2HSV1 U46725 ( .A1(n41522), .A2(n53523), .ZN(n42415) );
  XOR2HSV0 U46726 ( .A1(n42416), .A2(n42415), .Z(n42419) );
  CLKNAND2HSV1 U46727 ( .A1(n41160), .A2(n42417), .ZN(n42418) );
  XNOR2HSV1 U46728 ( .A1(n42419), .A2(n42418), .ZN(n42420) );
  XNOR2HSV1 U46729 ( .A1(n42421), .A2(n42420), .ZN(n42422) );
  XNOR2HSV1 U46730 ( .A1(n42423), .A2(n42422), .ZN(n42425) );
  NAND2HSV0 U46731 ( .A1(n59674), .A2(n44605), .ZN(n42424) );
  XOR3HSV2 U46732 ( .A1(n42426), .A2(n42425), .A3(n42424), .Z(n42427) );
  XNOR2HSV1 U46733 ( .A1(n42428), .A2(n42427), .ZN(n42430) );
  NAND2HSV0 U46734 ( .A1(n40917), .A2(n55214), .ZN(n42429) );
  XOR2HSV0 U46735 ( .A1(n42430), .A2(n42429), .Z(n42433) );
  NAND2HSV0 U46736 ( .A1(n42431), .A2(\pe1/got [12]), .ZN(n42432) );
  XOR2HSV0 U46737 ( .A1(n42433), .A2(n42432), .Z(n42434) );
  XNOR2HSV1 U46738 ( .A1(n42435), .A2(n42434), .ZN(n42437) );
  NAND2HSV0 U46739 ( .A1(n29773), .A2(\pe1/got [14]), .ZN(n42436) );
  XOR2HSV0 U46740 ( .A1(n42437), .A2(n42436), .Z(n42442) );
  NOR2HSV1 U46741 ( .A1(n42438), .A2(n54263), .ZN(n42441) );
  NAND2HSV0 U46742 ( .A1(n42439), .A2(n41374), .ZN(n42440) );
  XOR3HSV2 U46743 ( .A1(n42442), .A2(n42441), .A3(n42440), .Z(n42443) );
  XNOR2HSV1 U46744 ( .A1(n42444), .A2(n42443), .ZN(n42445) );
  XOR2HSV0 U46745 ( .A1(n42446), .A2(n42445), .Z(n42447) );
  XOR3HSV2 U46746 ( .A1(n42449), .A2(n42448), .A3(n42447), .Z(n42450) );
  XOR2HSV0 U46747 ( .A1(n42451), .A2(n42450), .Z(n42452) );
  XNOR2HSV1 U46748 ( .A1(n42453), .A2(n42452), .ZN(n42454) );
  XNOR2HSV1 U46749 ( .A1(n42455), .A2(n42454), .ZN(n42456) );
  XOR2HSV0 U46750 ( .A1(n42457), .A2(n42456), .Z(n42458) );
  XNOR2HSV1 U46751 ( .A1(n42459), .A2(n42458), .ZN(n42461) );
  CLKNAND2HSV0 U46752 ( .A1(n59377), .A2(n41689), .ZN(n42460) );
  XOR2HSV0 U46753 ( .A1(n42461), .A2(n42460), .Z(n42462) );
  XNOR2HSV4 U46754 ( .A1(n42469), .A2(n42468), .ZN(n48311) );
  CLKNHSV0 U46755 ( .I(n48311), .ZN(n42470) );
  NAND2HSV2 U46756 ( .A1(n48311), .A2(n42471), .ZN(n42472) );
  INHSV2 U46757 ( .I(n42472), .ZN(n42473) );
  INHSV4 U46758 ( .I(n48451), .ZN(n54146) );
  NAND2HSV2 U46759 ( .A1(n42473), .A2(n54146), .ZN(n42474) );
  NAND3HSV2 U46760 ( .A1(n44652), .A2(n48314), .A3(n42202), .ZN(n45780) );
  NOR2HSV0 U46761 ( .A1(n44524), .A2(n42478), .ZN(n42479) );
  OAI21HSV0 U46762 ( .A1(n45780), .A2(n42483), .B(n42479), .ZN(n42480) );
  AO21HSV1 U46763 ( .A1(n45782), .A2(n25873), .B(n42480), .Z(n42481) );
  NAND2HSV2 U46764 ( .A1(n42482), .A2(n42481), .ZN(n42487) );
  INHSV2 U46765 ( .I(n53503), .ZN(n55476) );
  NOR2HSV2 U46766 ( .A1(n42493), .A2(n42492), .ZN(n42495) );
  NOR2HSV1 U46767 ( .A1(n42600), .A2(n59615), .ZN(n42494) );
  CLKNAND2HSV1 U46768 ( .A1(n42495), .A2(n42494), .ZN(n42499) );
  CLKAND2HSV2 U46769 ( .A1(n42496), .A2(n36924), .Z(n42497) );
  AOI31HSV2 U46770 ( .A1(n42599), .A2(n42600), .A3(n46107), .B(n42497), .ZN(
        n42498) );
  CLKNHSV1 U46771 ( .I(n42500), .ZN(n42704) );
  INHSV2 U46772 ( .I(n42704), .ZN(n42505) );
  NOR2HSV1 U46773 ( .A1(n42501), .A2(n43752), .ZN(n42504) );
  OAI21HSV2 U46774 ( .A1(n42584), .A2(n43743), .B(n42919), .ZN(n42502) );
  NAND2HSV2 U46775 ( .A1(n55949), .A2(n42508), .ZN(n42514) );
  CLKNAND2HSV0 U46776 ( .A1(n42514), .A2(n37107), .ZN(n42519) );
  CLKNHSV0 U46777 ( .I(n42514), .ZN(n42510) );
  NAND2HSV0 U46778 ( .A1(n42513), .A2(n43234), .ZN(n42515) );
  MUX2NHSV1 U46779 ( .I0(n56057), .I1(n42515), .S(n42514), .ZN(n42516) );
  NOR2HSV2 U46780 ( .A1(n42517), .A2(n42516), .ZN(n42518) );
  OAI21HSV2 U46781 ( .A1(n37528), .A2(n42519), .B(n42518), .ZN(n42578) );
  CLKNAND2HSV1 U46782 ( .A1(n43622), .A2(n59616), .ZN(n42577) );
  BUFHSV2 U46783 ( .I(n59626), .Z(n55707) );
  NAND2HSV2 U46784 ( .A1(n55707), .A2(n42770), .ZN(n42571) );
  NAND2HSV0 U46785 ( .A1(n42938), .A2(n42520), .ZN(n42569) );
  CLKNAND2HSV0 U46786 ( .A1(n42710), .A2(\pe3/got [18]), .ZN(n42565) );
  CLKNHSV0 U46787 ( .I(n36694), .ZN(n55735) );
  CLKNAND2HSV0 U46788 ( .A1(n42728), .A2(n55735), .ZN(n42522) );
  CLKNAND2HSV0 U46789 ( .A1(n46363), .A2(n48538), .ZN(n42521) );
  XOR2HSV0 U46790 ( .A1(n42522), .A2(n42521), .Z(n42526) );
  CLKNAND2HSV0 U46791 ( .A1(n42950), .A2(n48522), .ZN(n42524) );
  NAND2HSV0 U46792 ( .A1(n59618), .A2(\pe3/bq[26] ), .ZN(n42523) );
  XOR2HSV0 U46793 ( .A1(n42524), .A2(n42523), .Z(n42525) );
  XOR2HSV0 U46794 ( .A1(n42526), .A2(n42525), .Z(n42536) );
  NAND2HSV0 U46795 ( .A1(n42818), .A2(n42527), .ZN(n42529) );
  NAND2HSV0 U46796 ( .A1(n59368), .A2(n56213), .ZN(n42528) );
  XOR2HSV0 U46797 ( .A1(n42529), .A2(n42528), .Z(n42534) );
  NAND2HSV0 U46798 ( .A1(\pe3/aot [24]), .A2(n42530), .ZN(n42532) );
  NAND2HSV0 U46799 ( .A1(n43547), .A2(n42642), .ZN(n42531) );
  XOR2HSV0 U46800 ( .A1(n42532), .A2(n42531), .Z(n42533) );
  XOR2HSV0 U46801 ( .A1(n42534), .A2(n42533), .Z(n42535) );
  XOR2HSV0 U46802 ( .A1(n42536), .A2(n42535), .Z(n42538) );
  NAND2HSV0 U46803 ( .A1(n42725), .A2(\pe3/got [17]), .ZN(n42537) );
  XNOR2HSV1 U46804 ( .A1(n42538), .A2(n42537), .ZN(n42562) );
  NOR2HSV0 U46805 ( .A1(n42539), .A2(n45525), .ZN(n42542) );
  INHSV2 U46806 ( .I(\pe3/aot [16]), .ZN(n49265) );
  CLKNAND2HSV0 U46807 ( .A1(n56508), .A2(n42540), .ZN(n42541) );
  XOR2HSV0 U46808 ( .A1(n42542), .A2(n42541), .Z(n42546) );
  NAND2HSV0 U46809 ( .A1(n56204), .A2(n42634), .ZN(n42544) );
  NAND2HSV0 U46810 ( .A1(n42743), .A2(n43146), .ZN(n42543) );
  XOR2HSV0 U46811 ( .A1(n42544), .A2(n42543), .Z(n42545) );
  XOR2HSV0 U46812 ( .A1(n42546), .A2(n42545), .Z(n42553) );
  CLKNHSV1 U46813 ( .I(n43059), .ZN(n42831) );
  INHSV2 U46814 ( .I(n42831), .ZN(n46125) );
  NAND2HSV2 U46815 ( .A1(n46125), .A2(\pe3/pvq [17]), .ZN(n42547) );
  XOR2HSV0 U46816 ( .A1(n42547), .A2(\pe3/phq [17]), .Z(n42551) );
  NAND2HSV0 U46817 ( .A1(n59622), .A2(\pe3/bq[19] ), .ZN(n42736) );
  OAI22HSV0 U46818 ( .A1(n36989), .A2(n46131), .B1(n42843), .B2(n43039), .ZN(
        n42548) );
  OAI21HSV1 U46819 ( .A1(n42736), .A2(n42549), .B(n42548), .ZN(n42550) );
  XOR2HSV0 U46820 ( .A1(n42551), .A2(n42550), .Z(n42552) );
  XNOR2HSV1 U46821 ( .A1(n42553), .A2(n42552), .ZN(n42560) );
  CLKNAND2HSV0 U46822 ( .A1(n45554), .A2(n42971), .ZN(n42555) );
  INHSV2 U46823 ( .I(n45576), .ZN(n43437) );
  NAND2HSV0 U46824 ( .A1(n43437), .A2(n37051), .ZN(n42554) );
  XOR2HSV0 U46825 ( .A1(n42555), .A2(n42554), .Z(n42558) );
  CLKNAND2HSV1 U46826 ( .A1(n43528), .A2(n45696), .ZN(n46366) );
  NAND2HSV0 U46827 ( .A1(n43650), .A2(\pe3/bq[18] ), .ZN(n42556) );
  XOR2HSV0 U46828 ( .A1(n46366), .A2(n42556), .Z(n42557) );
  XOR2HSV0 U46829 ( .A1(n42558), .A2(n42557), .Z(n42559) );
  XNOR2HSV1 U46830 ( .A1(n42560), .A2(n42559), .ZN(n42561) );
  XNOR2HSV1 U46831 ( .A1(n42562), .A2(n42561), .ZN(n42564) );
  NAND2HSV2 U46832 ( .A1(n43516), .A2(n59965), .ZN(n42563) );
  XOR3HSV2 U46833 ( .A1(n42565), .A2(n42564), .A3(n42563), .Z(n42567) );
  CLKNAND2HSV0 U46834 ( .A1(n59621), .A2(n42996), .ZN(n42566) );
  XOR2HSV0 U46835 ( .A1(n42567), .A2(n42566), .Z(n42568) );
  XOR2HSV0 U46836 ( .A1(n42569), .A2(n42568), .Z(n42570) );
  XOR2HSV0 U46837 ( .A1(n42571), .A2(n42570), .Z(n42573) );
  NAND2HSV0 U46838 ( .A1(n42767), .A2(n42673), .ZN(n42572) );
  XOR2HSV0 U46839 ( .A1(n42573), .A2(n42572), .Z(n42575) );
  INHSV2 U46840 ( .I(n37326), .ZN(n43097) );
  CLKNAND2HSV1 U46841 ( .A1(n43097), .A2(n43452), .ZN(n42574) );
  XNOR2HSV1 U46842 ( .A1(n42575), .A2(n42574), .ZN(n42576) );
  XNOR2HSV4 U46843 ( .A1(n42578), .A2(n29683), .ZN(n42580) );
  AOI21HSV4 U46844 ( .A1(n42581), .A2(n29717), .B(n42580), .ZN(n42579) );
  CLKNHSV2 U46845 ( .I(n42579), .ZN(n42583) );
  XNOR2HSV4 U46846 ( .A1(n42586), .A2(n42585), .ZN(n42587) );
  CLKNHSV0 U46847 ( .I(\pe3/ti_7t [16]), .ZN(n42589) );
  NAND2HSV0 U46848 ( .A1(n42589), .A2(n43743), .ZN(n42786) );
  NAND2HSV0 U46849 ( .A1(n42786), .A2(n37264), .ZN(n42603) );
  OR2HSV1 U46850 ( .A1(n42603), .A2(n42689), .Z(n42798) );
  CLKNHSV1 U46851 ( .I(n42798), .ZN(n42590) );
  CLKNAND2HSV0 U46852 ( .A1(n42591), .A2(n42592), .ZN(n42593) );
  NOR2HSV2 U46853 ( .A1(n42595), .A2(n42594), .ZN(n42598) );
  INHSV2 U46854 ( .I(n42596), .ZN(n42597) );
  NOR2HSV2 U46855 ( .A1(n43226), .A2(n59998), .ZN(n42601) );
  INHSV2 U46856 ( .I(\pe3/ti_7t [17]), .ZN(n42602) );
  NOR2HSV2 U46857 ( .A1(n42698), .A2(n42602), .ZN(n42799) );
  NOR2HSV1 U46858 ( .A1(n52790), .A2(n59998), .ZN(n42604) );
  CLKNAND2HSV4 U46859 ( .A1(n42608), .A2(n42802), .ZN(n43029) );
  CLKNHSV1 U46860 ( .I(n42610), .ZN(n42611) );
  BUFHSV2 U46861 ( .I(n42612), .Z(n42614) );
  AND2HSV2 U46862 ( .A1(n42786), .A2(n36924), .Z(n42613) );
  NOR3HSV4 U46863 ( .A1(n42615), .A2(n42614), .A3(n42919), .ZN(n42791) );
  CLKNAND2HSV0 U46864 ( .A1(n59620), .A2(n59616), .ZN(n42681) );
  CLKNAND2HSV0 U46865 ( .A1(n43622), .A2(n46441), .ZN(n42679) );
  CLKNAND2HSV1 U46866 ( .A1(n55949), .A2(n59617), .ZN(n42677) );
  CLKNAND2HSV1 U46867 ( .A1(n55707), .A2(n42999), .ZN(n42670) );
  NAND2HSV0 U46868 ( .A1(n42938), .A2(n55823), .ZN(n42668) );
  NAND2HSV0 U46869 ( .A1(n42710), .A2(n56064), .ZN(n42664) );
  NAND2HSV0 U46870 ( .A1(n45695), .A2(n56213), .ZN(n42619) );
  INHSV2 U46871 ( .I(\pe3/aot [16]), .ZN(n43178) );
  NAND2HSV0 U46872 ( .A1(\pe3/aot [16]), .A2(n48538), .ZN(n42618) );
  XOR2HSV0 U46873 ( .A1(n42619), .A2(n42618), .Z(n42623) );
  CLKNHSV0 U46874 ( .I(n42833), .ZN(n42939) );
  CLKNAND2HSV1 U46875 ( .A1(n56651), .A2(n42939), .ZN(n42621) );
  INHSV2 U46876 ( .I(n46615), .ZN(n43809) );
  NAND2HSV0 U46877 ( .A1(n43528), .A2(n43809), .ZN(n42620) );
  XOR2HSV0 U46878 ( .A1(n42621), .A2(n42620), .Z(n42622) );
  XOR2HSV0 U46879 ( .A1(n42623), .A2(n42622), .Z(n42631) );
  NAND2HSV0 U46880 ( .A1(n42940), .A2(\pe3/bq[26] ), .ZN(n42625) );
  CLKNAND2HSV0 U46881 ( .A1(n42950), .A2(n55735), .ZN(n42624) );
  XOR2HSV0 U46882 ( .A1(n42625), .A2(n42624), .Z(n42629) );
  BUFHSV2 U46883 ( .I(\pe3/bq[25] ), .Z(n42949) );
  NAND2HSV0 U46884 ( .A1(n59618), .A2(n42949), .ZN(n42627) );
  INHSV2 U46885 ( .I(n45727), .ZN(n48584) );
  NAND2HSV0 U46886 ( .A1(n48584), .A2(n37007), .ZN(n42626) );
  XOR2HSV0 U46887 ( .A1(n42627), .A2(n42626), .Z(n42628) );
  XOR2HSV0 U46888 ( .A1(n42629), .A2(n42628), .Z(n42630) );
  XOR2HSV0 U46889 ( .A1(n42631), .A2(n42630), .Z(n42633) );
  NAND2HSV0 U46890 ( .A1(n42725), .A2(n43437), .ZN(n42632) );
  XNOR2HSV1 U46891 ( .A1(n42633), .A2(n42632), .ZN(n42661) );
  NAND2HSV0 U46892 ( .A1(n45648), .A2(\pe3/bq[18] ), .ZN(n42636) );
  NAND2HSV0 U46893 ( .A1(n42728), .A2(n42634), .ZN(n42635) );
  XOR2HSV0 U46894 ( .A1(n42636), .A2(n42635), .Z(n42640) );
  NAND2HSV0 U46895 ( .A1(n42818), .A2(n43052), .ZN(n42638) );
  NAND2HSV0 U46896 ( .A1(n59368), .A2(n43146), .ZN(n42637) );
  XOR2HSV0 U46897 ( .A1(n42638), .A2(n42637), .Z(n42639) );
  XOR2HSV0 U46898 ( .A1(n42640), .A2(n42639), .Z(n42648) );
  NAND2HSV0 U46899 ( .A1(n46129), .A2(\pe3/pvq [18]), .ZN(n42641) );
  XOR2HSV0 U46900 ( .A1(n42641), .A2(\pe3/phq [18]), .Z(n42646) );
  NAND2HSV0 U46901 ( .A1(n45554), .A2(n42642), .ZN(n42976) );
  OAI22HSV0 U46902 ( .A1(n43757), .A2(n55755), .B1(n45555), .B2(n46131), .ZN(
        n42644) );
  OAI21HSV0 U46903 ( .A1(n42738), .A2(n42976), .B(n42644), .ZN(n42645) );
  XOR2HSV0 U46904 ( .A1(n42646), .A2(n42645), .Z(n42647) );
  XNOR2HSV1 U46905 ( .A1(n42648), .A2(n42647), .ZN(n42659) );
  NAND2HSV0 U46906 ( .A1(\pe3/aot [17]), .A2(n43544), .ZN(n46364) );
  INHSV2 U46907 ( .I(n46138), .ZN(n56498) );
  NAND2HSV0 U46908 ( .A1(n43547), .A2(n56498), .ZN(n42963) );
  OAI21HSV0 U46909 ( .A1(n43527), .A2(n42649), .B(n42963), .ZN(n42650) );
  OAI21HSV0 U46910 ( .A1(n46364), .A2(n42651), .B(n42650), .ZN(n42652) );
  NOR2HSV0 U46911 ( .A1(n42843), .A2(n45810), .ZN(n48536) );
  XNOR2HSV1 U46912 ( .A1(n42652), .A2(n48536), .ZN(n42657) );
  NAND2HSV0 U46913 ( .A1(n56204), .A2(n42653), .ZN(n42655) );
  NAND2HSV0 U46914 ( .A1(n42743), .A2(n49439), .ZN(n42654) );
  XOR2HSV0 U46915 ( .A1(n42655), .A2(n42654), .Z(n42656) );
  XNOR2HSV1 U46916 ( .A1(n42657), .A2(n42656), .ZN(n42658) );
  XNOR2HSV1 U46917 ( .A1(n42659), .A2(n42658), .ZN(n42660) );
  XNOR2HSV1 U46918 ( .A1(n42661), .A2(n42660), .ZN(n42663) );
  CLKNAND2HSV0 U46919 ( .A1(n43516), .A2(n43374), .ZN(n42662) );
  XOR3HSV2 U46920 ( .A1(n42664), .A2(n42663), .A3(n42662), .Z(n42666) );
  NAND2HSV0 U46921 ( .A1(n59621), .A2(n42937), .ZN(n42665) );
  XNOR2HSV1 U46922 ( .A1(n42666), .A2(n42665), .ZN(n42667) );
  XOR2HSV0 U46923 ( .A1(n42668), .A2(n42667), .Z(n42669) );
  XOR2HSV0 U46924 ( .A1(n42670), .A2(n42669), .Z(n42672) );
  NAND2HSV0 U46925 ( .A1(n42767), .A2(n42770), .ZN(n42671) );
  XOR2HSV0 U46926 ( .A1(n42672), .A2(n42671), .Z(n42675) );
  CLKNAND2HSV0 U46927 ( .A1(n43097), .A2(n42673), .ZN(n42674) );
  XNOR2HSV1 U46928 ( .A1(n42675), .A2(n42674), .ZN(n42676) );
  XNOR2HSV1 U46929 ( .A1(n42677), .A2(n42676), .ZN(n42678) );
  XNOR2HSV1 U46930 ( .A1(n42679), .A2(n42678), .ZN(n42680) );
  NOR2HSV0 U46931 ( .A1(n42684), .A2(n42683), .ZN(n42685) );
  OAI21HSV2 U46932 ( .A1(n60046), .A2(n43242), .B(n42685), .ZN(n42686) );
  AND2HSV2 U46933 ( .A1(n42702), .A2(n42694), .Z(n42695) );
  XNOR2HSV4 U46934 ( .A1(n42810), .A2(n43025), .ZN(n42699) );
  NOR2HSV0 U46935 ( .A1(n42698), .A2(\pe3/ti_7t [18]), .ZN(n42907) );
  NOR2HSV2 U46936 ( .A1(n42907), .A2(n43891), .ZN(n45796) );
  AOI21HSV4 U46937 ( .A1(n42699), .A2(n45796), .B(n43912), .ZN(n42805) );
  NAND2HSV2 U46938 ( .A1(n43453), .A2(n59963), .ZN(n42783) );
  AND2HSV2 U46939 ( .A1(n42702), .A2(n59964), .Z(n42703) );
  NOR2HSV4 U46940 ( .A1(n42704), .A2(n42705), .ZN(n42708) );
  NAND2HSV2 U46941 ( .A1(n46043), .A2(n37107), .ZN(n42707) );
  XNOR2HSV4 U46942 ( .A1(n42708), .A2(n42707), .ZN(n42782) );
  MUX2NHSV1 U46943 ( .I0(n60046), .I1(\pe3/ti_7t [12]), .S(n43132), .ZN(n42709) );
  INHSV2 U46944 ( .I(n42709), .ZN(n43222) );
  NAND2HSV2 U46945 ( .A1(n43222), .A2(\pe3/got [26]), .ZN(n42780) );
  BUFHSV2 U46946 ( .I(n59620), .Z(n45517) );
  CLKBUFHSV4 U46947 ( .I(n45517), .Z(n56067) );
  NAND2HSV2 U46948 ( .A1(n45517), .A2(n46441), .ZN(n42778) );
  CLKBUFHSV4 U46949 ( .I(n43622), .Z(n59625) );
  NAND2HSV2 U46950 ( .A1(n59625), .A2(n59617), .ZN(n42776) );
  NAND2HSV2 U46951 ( .A1(n43495), .A2(n42673), .ZN(n42774) );
  NAND2HSV0 U46952 ( .A1(n55825), .A2(n42996), .ZN(n42766) );
  NAND2HSV0 U46953 ( .A1(n42938), .A2(n59965), .ZN(n42764) );
  NAND2HSV0 U46954 ( .A1(n42710), .A2(n43437), .ZN(n42760) );
  NAND2HSV0 U46955 ( .A1(n45554), .A2(\pe3/bq[18] ), .ZN(n42712) );
  CLKNAND2HSV0 U46956 ( .A1(\pe3/aot [14]), .A2(n42939), .ZN(n42711) );
  XOR2HSV0 U46957 ( .A1(n42712), .A2(n42711), .Z(n42716) );
  NAND2HSV0 U46958 ( .A1(n55864), .A2(n48538), .ZN(n42714) );
  NAND2HSV0 U46959 ( .A1(\pe3/got [14]), .A2(n37007), .ZN(n42713) );
  XOR2HSV0 U46960 ( .A1(n42714), .A2(n42713), .Z(n42715) );
  XOR2HSV0 U46961 ( .A1(n42716), .A2(n42715), .Z(n42724) );
  NAND2HSV0 U46962 ( .A1(n56182), .A2(n42949), .ZN(n42718) );
  NAND2HSV0 U46963 ( .A1(\pe3/aot [22]), .A2(\pe3/bq[24] ), .ZN(n42717) );
  XOR2HSV0 U46964 ( .A1(n42718), .A2(n42717), .Z(n42722) );
  NAND2HSV0 U46965 ( .A1(n56204), .A2(\pe3/bq[26] ), .ZN(n42720) );
  INHSV2 U46966 ( .I(n43178), .ZN(n43030) );
  NAND2HSV0 U46967 ( .A1(n43030), .A2(n43389), .ZN(n42719) );
  XOR2HSV0 U46968 ( .A1(n42720), .A2(n42719), .Z(n42721) );
  XOR2HSV0 U46969 ( .A1(n42722), .A2(n42721), .Z(n42723) );
  XOR2HSV0 U46970 ( .A1(n42724), .A2(n42723), .Z(n42727) );
  BUFHSV2 U46971 ( .I(n42725), .Z(n43424) );
  INHSV2 U46972 ( .I(n45727), .ZN(n56264) );
  CLKNAND2HSV0 U46973 ( .A1(n43424), .A2(n56264), .ZN(n42726) );
  XNOR2HSV1 U46974 ( .A1(n42727), .A2(n42726), .ZN(n42757) );
  NAND2HSV0 U46975 ( .A1(n45648), .A2(n56519), .ZN(n42730) );
  CLKNHSV0 U46976 ( .I(n45525), .ZN(n44698) );
  NAND2HSV0 U46977 ( .A1(n42728), .A2(n44698), .ZN(n42729) );
  XOR2HSV0 U46978 ( .A1(n42730), .A2(n42729), .Z(n42734) );
  CLKNHSV0 U46979 ( .I(n55714), .ZN(n43040) );
  CLKNAND2HSV0 U46980 ( .A1(n43040), .A2(n49439), .ZN(n42732) );
  NAND2HSV0 U46981 ( .A1(n42950), .A2(n55867), .ZN(n42731) );
  XOR2HSV0 U46982 ( .A1(n42732), .A2(n42731), .Z(n42733) );
  XOR2HSV0 U46983 ( .A1(n42734), .A2(n42733), .Z(n42742) );
  CLKNHSV0 U46984 ( .I(n42831), .ZN(n59537) );
  NAND2HSV2 U46985 ( .A1(n59537), .A2(\pe3/pvq [19]), .ZN(n42735) );
  XOR2HSV0 U46986 ( .A1(n42735), .A2(\pe3/phq [19]), .Z(n42740) );
  NAND2HSV0 U46987 ( .A1(n59622), .A2(n56498), .ZN(n43070) );
  OAI21HSV0 U46988 ( .A1(n46138), .A2(n43757), .B(n42736), .ZN(n42737) );
  OAI21HSV0 U46989 ( .A1(n43070), .A2(n42738), .B(n42737), .ZN(n42739) );
  XOR2HSV0 U46990 ( .A1(n42740), .A2(n42739), .Z(n42741) );
  XNOR2HSV1 U46991 ( .A1(n42742), .A2(n42741), .ZN(n42755) );
  NAND2HSV0 U46992 ( .A1(n42743), .A2(\pe3/bq[14] ), .ZN(n43182) );
  OAI22HSV0 U46993 ( .A1(n42821), .A2(n49281), .B1(n45564), .B2(n45810), .ZN(
        n42744) );
  OAI21HSV0 U46994 ( .A1(n43182), .A2(n42745), .B(n42744), .ZN(n42749) );
  CLKNHSV0 U46995 ( .I(n43527), .ZN(n43049) );
  CLKNAND2HSV0 U46996 ( .A1(n43049), .A2(n56641), .ZN(n48553) );
  CLKNAND2HSV1 U46997 ( .A1(n43265), .A2(n46323), .ZN(n43194) );
  OAI21HSV0 U46998 ( .A1(n43527), .A2(n36694), .B(n43194), .ZN(n42746) );
  OAI21HSV0 U46999 ( .A1(n42747), .A2(n48553), .B(n42746), .ZN(n42748) );
  XNOR2HSV1 U47000 ( .A1(n42749), .A2(n42748), .ZN(n42753) );
  CLKNHSV0 U47001 ( .I(n37196), .ZN(n43772) );
  CLKNAND2HSV1 U47002 ( .A1(n43034), .A2(n43772), .ZN(n42751) );
  NAND2HSV0 U47003 ( .A1(n42818), .A2(n56213), .ZN(n42750) );
  XOR2HSV0 U47004 ( .A1(n42751), .A2(n42750), .Z(n42752) );
  XNOR2HSV1 U47005 ( .A1(n42753), .A2(n42752), .ZN(n42754) );
  XNOR2HSV1 U47006 ( .A1(n42755), .A2(n42754), .ZN(n42756) );
  XNOR2HSV1 U47007 ( .A1(n42757), .A2(n42756), .ZN(n42759) );
  XOR3HSV2 U47008 ( .A1(n42760), .A2(n42759), .A3(n42758), .Z(n42762) );
  NAND2HSV0 U47009 ( .A1(n59621), .A2(n43374), .ZN(n42761) );
  XOR2HSV0 U47010 ( .A1(n42762), .A2(n42761), .Z(n42763) );
  XOR2HSV0 U47011 ( .A1(n42764), .A2(n42763), .Z(n42765) );
  XOR2HSV0 U47012 ( .A1(n42766), .A2(n42765), .Z(n42769) );
  NAND2HSV0 U47013 ( .A1(n42767), .A2(n42999), .ZN(n42768) );
  XOR2HSV0 U47014 ( .A1(n42769), .A2(n42768), .Z(n42772) );
  CLKNAND2HSV0 U47015 ( .A1(n43097), .A2(n42770), .ZN(n42771) );
  XNOR2HSV1 U47016 ( .A1(n42772), .A2(n42771), .ZN(n42773) );
  XOR2HSV0 U47017 ( .A1(n42774), .A2(n42773), .Z(n42775) );
  XOR2HSV0 U47018 ( .A1(n42776), .A2(n42775), .Z(n42777) );
  XOR2HSV0 U47019 ( .A1(n42778), .A2(n42777), .Z(n42779) );
  XNOR2HSV1 U47020 ( .A1(n42780), .A2(n42779), .ZN(n42781) );
  CLKNHSV0 U47021 ( .I(n42786), .ZN(n42787) );
  NOR2HSV1 U47022 ( .A1(n42787), .A2(n43752), .ZN(n42788) );
  CLKNAND2HSV1 U47023 ( .A1(n42789), .A2(n42788), .ZN(n42790) );
  CLKNAND2HSV1 U47024 ( .A1(n42792), .A2(n42793), .ZN(n42796) );
  INHSV2 U47025 ( .I(n42792), .ZN(n42794) );
  NAND2HSV2 U47026 ( .A1(n42796), .A2(n42795), .ZN(n42804) );
  CLKNHSV0 U47027 ( .I(n42799), .ZN(n42800) );
  OR2HSV1 U47028 ( .A1(n42800), .A2(n43361), .Z(n42801) );
  XNOR2HSV4 U47029 ( .A1(n42804), .A2(n42803), .ZN(n45799) );
  CLKNAND2HSV3 U47030 ( .A1(n42917), .A2(n42807), .ZN(n45798) );
  CLKNHSV0 U47031 ( .I(n45796), .ZN(n42808) );
  NOR2HSV1 U47032 ( .A1(n42808), .A2(n45932), .ZN(n42809) );
  CLKNAND2HSV2 U47033 ( .A1(n45798), .A2(n42809), .ZN(n42812) );
  CLKNAND2HSV2 U47034 ( .A1(n42906), .A2(n42810), .ZN(n45797) );
  NOR2HSV2 U47035 ( .A1(n42812), .A2(n42811), .ZN(n42814) );
  INHSV2 U47036 ( .I(n45799), .ZN(n42813) );
  CLKNAND2HSV3 U47037 ( .A1(n42814), .A2(n42813), .ZN(n43019) );
  INHSV2 U47038 ( .I(n42816), .ZN(n42912) );
  NOR2HSV2 U47039 ( .A1(n43448), .A2(n42817), .ZN(n42892) );
  NAND2HSV2 U47040 ( .A1(n43424), .A2(n56421), .ZN(n42825) );
  NAND2HSV2 U47041 ( .A1(n59612), .A2(n49439), .ZN(n42820) );
  INHSV2 U47042 ( .I(n50802), .ZN(n59966) );
  CLKNAND2HSV0 U47043 ( .A1(n59966), .A2(n45955), .ZN(n42819) );
  XOR2HSV0 U47044 ( .A1(n42820), .A2(n42819), .Z(n42823) );
  CLKNHSV0 U47045 ( .I(n42821), .ZN(n45962) );
  INHSV2 U47046 ( .I(\pe3/bq[12] ), .ZN(n43031) );
  INHSV2 U47047 ( .I(n43031), .ZN(n45982) );
  CLKNAND2HSV1 U47048 ( .A1(n45962), .A2(n45982), .ZN(n42822) );
  XNOR2HSV1 U47049 ( .A1(n42823), .A2(n42822), .ZN(n42824) );
  XNOR2HSV1 U47050 ( .A1(n42825), .A2(n42824), .ZN(n42828) );
  CLKNHSV0 U47051 ( .I(n42828), .ZN(n42826) );
  NOR2HSV0 U47052 ( .A1(n42826), .A2(n42827), .ZN(n42830) );
  AOI21HSV2 U47053 ( .A1(n59620), .A2(\pe3/got [23]), .B(n42828), .ZN(n42829)
         );
  AOI21HSV1 U47054 ( .A1(n42830), .A2(n59620), .B(n42829), .ZN(n42890) );
  CLKNAND2HSV0 U47055 ( .A1(n59625), .A2(n42770), .ZN(n42888) );
  NAND2HSV0 U47056 ( .A1(n55949), .A2(n43262), .ZN(n42886) );
  NAND2HSV0 U47057 ( .A1(n45949), .A2(n43374), .ZN(n42880) );
  CLKNAND2HSV1 U47058 ( .A1(n48488), .A2(n56335), .ZN(n42878) );
  INHSV2 U47059 ( .I(n42831), .ZN(n46128) );
  CLKNAND2HSV0 U47060 ( .A1(n46128), .A2(\pe3/pvq [21]), .ZN(n42832) );
  XNOR2HSV1 U47061 ( .A1(n42832), .A2(\pe3/phq [21]), .ZN(n42834) );
  INHSV2 U47062 ( .I(n53229), .ZN(n56575) );
  CLKNHSV0 U47063 ( .I(n42833), .ZN(n43499) );
  CLKNAND2HSV0 U47064 ( .A1(n56575), .A2(n43499), .ZN(n46347) );
  XNOR2HSV1 U47065 ( .A1(n42834), .A2(n46347), .ZN(n42853) );
  NAND2HSV0 U47066 ( .A1(n56464), .A2(n42949), .ZN(n42837) );
  NAND2HSV0 U47067 ( .A1(n43034), .A2(n42971), .ZN(n42836) );
  XOR2HSV0 U47068 ( .A1(n42837), .A2(n42836), .Z(n42841) );
  NAND2HSV0 U47069 ( .A1(n43040), .A2(\pe3/bq[19] ), .ZN(n42839) );
  NAND2HSV0 U47070 ( .A1(\pe3/aot [15]), .A2(n55735), .ZN(n42838) );
  XOR2HSV0 U47071 ( .A1(n42839), .A2(n42838), .Z(n42840) );
  XOR2HSV0 U47072 ( .A1(n42841), .A2(n42840), .Z(n42852) );
  NAND2HSV0 U47073 ( .A1(\pe3/aot [22]), .A2(n43772), .ZN(n49276) );
  XOR2HSV0 U47074 ( .A1(n42842), .A2(n49276), .Z(n42851) );
  CLKNHSV0 U47075 ( .I(n45555), .ZN(n45640) );
  NAND2HSV0 U47076 ( .A1(n45640), .A2(n56498), .ZN(n42845) );
  CLKNHSV0 U47077 ( .I(n42843), .ZN(n46456) );
  NAND2HSV0 U47078 ( .A1(n46456), .A2(n56519), .ZN(n42844) );
  XOR2HSV0 U47079 ( .A1(n42845), .A2(n42844), .Z(n42849) );
  NAND2HSV0 U47080 ( .A1(\pe3/aot [14]), .A2(n43389), .ZN(n42847) );
  NAND2HSV0 U47081 ( .A1(n56182), .A2(\pe3/bq[23] ), .ZN(n42846) );
  XOR2HSV0 U47082 ( .A1(n42847), .A2(n42846), .Z(n42848) );
  XOR2HSV0 U47083 ( .A1(n42849), .A2(n42848), .Z(n42850) );
  XOR4HSV1 U47084 ( .A1(n42853), .A2(n42852), .A3(n42851), .A4(n42850), .Z(
        n42869) );
  INHSV2 U47085 ( .I(\pe3/aot [13]), .ZN(n43151) );
  NAND2HSV0 U47086 ( .A1(n43280), .A2(n48538), .ZN(n42855) );
  NAND2HSV0 U47087 ( .A1(n56204), .A2(n43052), .ZN(n42854) );
  XOR2HSV0 U47088 ( .A1(n42855), .A2(n42854), .Z(n42859) );
  NAND2HSV0 U47089 ( .A1(n45648), .A2(n43809), .ZN(n42857) );
  NAND2HSV0 U47090 ( .A1(n55988), .A2(\pe3/bq[18] ), .ZN(n42856) );
  XOR2HSV0 U47091 ( .A1(n42857), .A2(n42856), .Z(n42858) );
  XOR2HSV0 U47092 ( .A1(n42859), .A2(n42858), .Z(n42867) );
  NOR2HSV0 U47093 ( .A1(n42643), .A2(n49281), .ZN(n42861) );
  NAND2HSV0 U47094 ( .A1(n42950), .A2(\pe3/bq[26] ), .ZN(n42860) );
  XOR2HSV0 U47095 ( .A1(n42861), .A2(n42860), .Z(n42865) );
  INHSV6 U47096 ( .I(\pe3/bq[13] ), .ZN(n49423) );
  INHSV2 U47097 ( .I(n49423), .ZN(n56460) );
  NAND2HSV0 U47098 ( .A1(n43265), .A2(n56460), .ZN(n42863) );
  NAND2HSV0 U47099 ( .A1(n43030), .A2(n55867), .ZN(n42862) );
  XOR2HSV0 U47100 ( .A1(n42863), .A2(n42862), .Z(n42864) );
  XOR2HSV0 U47101 ( .A1(n42865), .A2(n42864), .Z(n42866) );
  XOR2HSV0 U47102 ( .A1(n42867), .A2(n42866), .Z(n42868) );
  XNOR2HSV1 U47103 ( .A1(n42869), .A2(n42868), .ZN(n42871) );
  NAND2HSV0 U47104 ( .A1(n59797), .A2(\pe3/got [14]), .ZN(n42870) );
  XNOR2HSV1 U47105 ( .A1(n42871), .A2(n42870), .ZN(n42873) );
  CLKNHSV0 U47106 ( .I(n45727), .ZN(n59624) );
  NAND2HSV0 U47107 ( .A1(n59671), .A2(n59624), .ZN(n42872) );
  XNOR2HSV1 U47108 ( .A1(n42873), .A2(n42872), .ZN(n42876) );
  BUFHSV2 U47109 ( .I(n42874), .Z(n52727) );
  CLKNAND2HSV0 U47110 ( .A1(n52727), .A2(n43437), .ZN(n42875) );
  XOR2HSV0 U47111 ( .A1(n42876), .A2(n42875), .Z(n42877) );
  XOR2HSV0 U47112 ( .A1(n42878), .A2(n42877), .Z(n42879) );
  XOR2HSV0 U47113 ( .A1(n42880), .A2(n42879), .Z(n42882) );
  BUFHSV2 U47114 ( .I(n42767), .Z(n43211) );
  NAND2HSV0 U47115 ( .A1(n43211), .A2(n42937), .ZN(n42881) );
  XOR2HSV0 U47116 ( .A1(n42882), .A2(n42881), .Z(n42884) );
  INHSV2 U47117 ( .I(n45635), .ZN(n49404) );
  NAND2HSV0 U47118 ( .A1(n43097), .A2(n49404), .ZN(n42883) );
  XNOR2HSV1 U47119 ( .A1(n42884), .A2(n42883), .ZN(n42885) );
  XNOR2HSV1 U47120 ( .A1(n42886), .A2(n42885), .ZN(n42887) );
  XNOR2HSV1 U47121 ( .A1(n42888), .A2(n42887), .ZN(n42889) );
  XOR2HSV0 U47122 ( .A1(n42890), .A2(n42889), .Z(n42891) );
  XNOR2HSV1 U47123 ( .A1(n42892), .A2(n42891), .ZN(n42894) );
  INHSV2 U47124 ( .I(n46519), .ZN(n46043) );
  NAND2HSV2 U47125 ( .A1(n46043), .A2(n46441), .ZN(n42893) );
  XOR2HSV0 U47126 ( .A1(n42894), .A2(n42893), .Z(n42898) );
  INHSV2 U47127 ( .I(n42683), .ZN(n45633) );
  CLKNAND2HSV1 U47128 ( .A1(n43453), .A2(n45633), .ZN(n42897) );
  MUX2NHSV4 U47129 ( .I0(n60088), .I1(\pe3/ti_7t [14]), .S(n36980), .ZN(n43106) );
  CLKNHSV2 U47130 ( .I(n43106), .ZN(n43706) );
  NOR2HSV4 U47131 ( .A1(n56475), .A2(n43457), .ZN(n42896) );
  XOR3HSV2 U47132 ( .A1(n42898), .A2(n42897), .A3(n42896), .Z(n42903) );
  CLKNAND2HSV2 U47133 ( .A1(pov3[16]), .A2(n42899), .ZN(n42901) );
  NAND2HSV2 U47134 ( .A1(n43242), .A2(\pe3/ti_7t [16]), .ZN(n42900) );
  NAND2HSV4 U47135 ( .A1(n42901), .A2(n42900), .ZN(n46415) );
  XOR2HSV2 U47136 ( .A1(n42903), .A2(n42902), .Z(n42905) );
  NAND2HSV2 U47137 ( .A1(n42917), .A2(\pe3/got [29]), .ZN(n42904) );
  XNOR2HSV4 U47138 ( .A1(n42905), .A2(n42904), .ZN(n42910) );
  INHSV2 U47139 ( .I(n42907), .ZN(n42922) );
  NAND2HSV2 U47140 ( .A1(n42922), .A2(n46082), .ZN(n42908) );
  XNOR2HSV4 U47141 ( .A1(n42910), .A2(n42909), .ZN(n42911) );
  CLKNHSV0 U47142 ( .I(n43020), .ZN(n42914) );
  CLKNAND2HSV0 U47143 ( .A1(n43019), .A2(n45625), .ZN(n42913) );
  NOR2HSV4 U47144 ( .A1(n42918), .A2(n46090), .ZN(n42931) );
  CLKNHSV0 U47145 ( .I(n42926), .ZN(n42921) );
  CLKNAND2HSV0 U47146 ( .A1(n42922), .A2(n42815), .ZN(n42923) );
  NOR2HSV4 U47147 ( .A1(n42931), .A2(n42932), .ZN(n42929) );
  OAI21HSV2 U47148 ( .A1(n42933), .A2(n42932), .B(n42931), .ZN(n42934) );
  CLKNAND2HSV3 U47149 ( .A1(n42935), .A2(n42934), .ZN(n43017) );
  NOR2HSV2 U47150 ( .A1(n43106), .A2(n42683), .ZN(n43015) );
  NAND2HSV2 U47151 ( .A1(n55948), .A2(n59617), .ZN(n43007) );
  NAND2HSV2 U47152 ( .A1(n59625), .A2(n42673), .ZN(n43005) );
  NAND2HSV2 U47153 ( .A1(n43495), .A2(n42770), .ZN(n43003) );
  NAND2HSV0 U47154 ( .A1(n45949), .A2(n42937), .ZN(n42995) );
  NAND2HSV0 U47155 ( .A1(n42938), .A2(n43374), .ZN(n42993) );
  INHSV2 U47156 ( .I(n45727), .ZN(n45518) );
  NAND2HSV2 U47157 ( .A1(n59797), .A2(n45518), .ZN(n42989) );
  CLKNAND2HSV1 U47158 ( .A1(n59671), .A2(n43437), .ZN(n42988) );
  INHSV2 U47159 ( .I(n43151), .ZN(n53249) );
  CLKNAND2HSV1 U47160 ( .A1(n53249), .A2(n42939), .ZN(n42942) );
  NAND2HSV0 U47161 ( .A1(n42940), .A2(n43052), .ZN(n42941) );
  XOR2HSV0 U47162 ( .A1(n42942), .A2(n42941), .Z(n42946) );
  NAND2HSV2 U47163 ( .A1(n46456), .A2(\pe3/bq[18] ), .ZN(n42944) );
  NAND2HSV0 U47164 ( .A1(n59618), .A2(n56213), .ZN(n42943) );
  XOR2HSV0 U47165 ( .A1(n42944), .A2(n42943), .Z(n42945) );
  XOR2HSV0 U47166 ( .A1(n42946), .A2(n42945), .Z(n42956) );
  CLKNAND2HSV0 U47167 ( .A1(n43030), .A2(n55735), .ZN(n42948) );
  CLKNAND2HSV0 U47168 ( .A1(n56464), .A2(\pe3/bq[26] ), .ZN(n42947) );
  XOR2HSV0 U47169 ( .A1(n42948), .A2(n42947), .Z(n42954) );
  NAND2HSV0 U47170 ( .A1(n56204), .A2(n42949), .ZN(n42952) );
  NAND2HSV0 U47171 ( .A1(n42950), .A2(n44698), .ZN(n42951) );
  XOR2HSV0 U47172 ( .A1(n42952), .A2(n42951), .Z(n42953) );
  XOR2HSV0 U47173 ( .A1(n42954), .A2(n42953), .Z(n42955) );
  XOR2HSV0 U47174 ( .A1(n42956), .A2(n42955), .Z(n42968) );
  CLKNAND2HSV1 U47175 ( .A1(n43049), .A2(n55867), .ZN(n42958) );
  NAND2HSV0 U47176 ( .A1(\pe3/got [13]), .A2(n37051), .ZN(n42957) );
  XOR2HSV0 U47177 ( .A1(n42958), .A2(n42957), .Z(n42961) );
  NAND2HSV2 U47178 ( .A1(n46128), .A2(\pe3/pvq [20]), .ZN(n42959) );
  XNOR2HSV1 U47179 ( .A1(n42959), .A2(\pe3/phq [20]), .ZN(n42960) );
  XNOR2HSV1 U47180 ( .A1(n42961), .A2(n42960), .ZN(n42966) );
  INHSV2 U47181 ( .I(n49281), .ZN(n56379) );
  NAND2HSV0 U47182 ( .A1(n45648), .A2(n56379), .ZN(n55717) );
  BUFHSV2 U47183 ( .I(n43392), .Z(n45691) );
  OAI22HSV0 U47184 ( .A1(n45691), .A2(n49281), .B1(n36989), .B2(n46138), .ZN(
        n42962) );
  OAI21HSV2 U47185 ( .A1(n55717), .A2(n42963), .B(n42962), .ZN(n42964) );
  CLKNAND2HSV0 U47186 ( .A1(n45962), .A2(n56460), .ZN(n43068) );
  XNOR2HSV1 U47187 ( .A1(n42964), .A2(n43068), .ZN(n42965) );
  XNOR2HSV1 U47188 ( .A1(n42966), .A2(n42965), .ZN(n42967) );
  XNOR2HSV1 U47189 ( .A1(n42968), .A2(n42967), .ZN(n42986) );
  CLKNAND2HSV1 U47190 ( .A1(n43034), .A2(n49439), .ZN(n42970) );
  CLKNAND2HSV0 U47191 ( .A1(n42818), .A2(n43772), .ZN(n42969) );
  XOR2HSV0 U47192 ( .A1(n42970), .A2(n42969), .Z(n42975) );
  NAND2HSV0 U47193 ( .A1(n43040), .A2(n42971), .ZN(n42973) );
  NAND2HSV0 U47194 ( .A1(n43650), .A2(n46323), .ZN(n42972) );
  XOR2HSV0 U47195 ( .A1(n42973), .A2(n42972), .Z(n42974) );
  XOR2HSV0 U47196 ( .A1(n42975), .A2(n42974), .Z(n42982) );
  NAND2HSV2 U47197 ( .A1(n55988), .A2(\pe3/bq[19] ), .ZN(n55849) );
  XOR2HSV0 U47198 ( .A1(n42976), .A2(n55849), .Z(n42980) );
  NAND2HSV0 U47199 ( .A1(n56651), .A2(n43389), .ZN(n42978) );
  NAND2HSV2 U47200 ( .A1(n56188), .A2(n48538), .ZN(n42977) );
  XOR2HSV0 U47201 ( .A1(n42978), .A2(n42977), .Z(n42979) );
  XOR2HSV0 U47202 ( .A1(n42980), .A2(n42979), .Z(n42981) );
  XOR2HSV0 U47203 ( .A1(n42982), .A2(n42981), .Z(n42984) );
  CLKNAND2HSV1 U47204 ( .A1(n43424), .A2(n56493), .ZN(n42983) );
  XNOR2HSV1 U47205 ( .A1(n42984), .A2(n42983), .ZN(n42985) );
  XOR2HSV0 U47206 ( .A1(n42986), .A2(n42985), .Z(n42987) );
  XOR3HSV2 U47207 ( .A1(n42989), .A2(n42988), .A3(n42987), .Z(n42991) );
  NAND2HSV0 U47208 ( .A1(n59621), .A2(n56064), .ZN(n42990) );
  XNOR2HSV1 U47209 ( .A1(n42991), .A2(n42990), .ZN(n42992) );
  XOR2HSV0 U47210 ( .A1(n42993), .A2(n42992), .Z(n42994) );
  XOR2HSV0 U47211 ( .A1(n42995), .A2(n42994), .Z(n42998) );
  NAND2HSV2 U47212 ( .A1(n43211), .A2(n42996), .ZN(n42997) );
  XNOR2HSV1 U47213 ( .A1(n42998), .A2(n42997), .ZN(n43001) );
  CLKNAND2HSV0 U47214 ( .A1(n43097), .A2(n42999), .ZN(n43000) );
  XNOR2HSV1 U47215 ( .A1(n43001), .A2(n43000), .ZN(n43002) );
  XNOR2HSV1 U47216 ( .A1(n43003), .A2(n43002), .ZN(n43004) );
  XNOR2HSV1 U47217 ( .A1(n43005), .A2(n43004), .ZN(n43006) );
  XNOR2HSV1 U47218 ( .A1(n43007), .A2(n43006), .ZN(n43010) );
  NOR2HSV2 U47219 ( .A1(n43448), .A2(n43231), .ZN(n43009) );
  NOR2HSV2 U47220 ( .A1(n46519), .A2(n43457), .ZN(n43008) );
  XOR3HSV2 U47221 ( .A1(n43010), .A2(n43009), .A3(n43008), .Z(n43011) );
  NAND2HSV2 U47222 ( .A1(n46415), .A2(n37340), .ZN(n43013) );
  XNOR3HSV1 U47223 ( .A1(n43015), .A2(n43014), .A3(n43013), .ZN(n43016) );
  XNOR2HSV4 U47224 ( .A1(n43017), .A2(n43016), .ZN(n43127) );
  CLKNAND2HSV2 U47225 ( .A1(n43018), .A2(n43135), .ZN(n43023) );
  INHSV2 U47226 ( .I(\pe3/ti_7t [20]), .ZN(n43120) );
  AO21HSV1 U47227 ( .A1(n43120), .A2(n59998), .B(n45931), .Z(n43022) );
  INHSV2 U47228 ( .I(\pe3/ti_7t [21]), .ZN(n43024) );
  NOR2HSV1 U47229 ( .A1(n43604), .A2(n43024), .ZN(n43246) );
  CLKNAND2HSV1 U47230 ( .A1(n43029), .A2(n52726), .ZN(n43026) );
  CLKNAND2HSV0 U47231 ( .A1(n42689), .A2(\pe3/ti_7t [18]), .ZN(n43027) );
  CLKNAND2HSV2 U47232 ( .A1(n43621), .A2(n43868), .ZN(n43116) );
  CLKNAND2HSV0 U47233 ( .A1(n46309), .A2(n43029), .ZN(n43111) );
  BUFHSV2 U47234 ( .I(n59625), .Z(n43373) );
  NAND2HSV2 U47235 ( .A1(n43373), .A2(n43262), .ZN(n43103) );
  NAND2HSV0 U47236 ( .A1(n56180), .A2(n49404), .ZN(n43101) );
  NAND2HSV0 U47237 ( .A1(n55825), .A2(n56064), .ZN(n43094) );
  CLKNAND2HSV1 U47238 ( .A1(n48488), .A2(n43437), .ZN(n43092) );
  NAND2HSV0 U47239 ( .A1(n43030), .A2(n44698), .ZN(n43033) );
  CLKNHSV0 U47240 ( .I(n43031), .ZN(n43775) );
  NAND2HSV0 U47241 ( .A1(n43265), .A2(n43775), .ZN(n43032) );
  XOR2HSV0 U47242 ( .A1(n43033), .A2(n43032), .Z(n43038) );
  CLKNAND2HSV0 U47243 ( .A1(n43034), .A2(\pe3/bq[19] ), .ZN(n43036) );
  CLKNAND2HSV0 U47244 ( .A1(n56354), .A2(n43499), .ZN(n43035) );
  XOR2HSV0 U47245 ( .A1(n43036), .A2(n43035), .Z(n43037) );
  XOR2HSV0 U47246 ( .A1(n43038), .A2(n43037), .Z(n43048) );
  NOR2HSV0 U47247 ( .A1(n45567), .A2(n43039), .ZN(n43042) );
  NAND2HSV0 U47248 ( .A1(n43040), .A2(\pe3/bq[18] ), .ZN(n43041) );
  XOR2HSV0 U47249 ( .A1(n43042), .A2(n43041), .Z(n43046) );
  NAND2HSV0 U47250 ( .A1(n42818), .A2(n42971), .ZN(n43044) );
  NAND2HSV0 U47251 ( .A1(n42743), .A2(n55616), .ZN(n43043) );
  XOR2HSV0 U47252 ( .A1(n43044), .A2(n43043), .Z(n43045) );
  XOR2HSV0 U47253 ( .A1(n43046), .A2(n43045), .Z(n43047) );
  XOR2HSV0 U47254 ( .A1(n43048), .A2(n43047), .Z(n43066) );
  CLKNAND2HSV0 U47255 ( .A1(n43049), .A2(\pe3/bq[26] ), .ZN(n43051) );
  NAND2HSV0 U47256 ( .A1(n56204), .A2(\pe3/bq[23] ), .ZN(n43050) );
  XOR2HSV0 U47257 ( .A1(n43051), .A2(n43050), .Z(n43056) );
  NAND2HSV0 U47258 ( .A1(n56464), .A2(n43052), .ZN(n43054) );
  NAND2HSV0 U47259 ( .A1(n42950), .A2(n56071), .ZN(n43053) );
  XOR2HSV0 U47260 ( .A1(n43054), .A2(n43053), .Z(n43055) );
  XOR2HSV0 U47261 ( .A1(n43056), .A2(n43055), .Z(n43064) );
  NOR2HSV0 U47262 ( .A1(n50799), .A2(n46126), .ZN(n43058) );
  NAND2HSV0 U47263 ( .A1(n56188), .A2(n55735), .ZN(n43057) );
  XOR2HSV0 U47264 ( .A1(n43058), .A2(n43057), .Z(n43062) );
  INHSV2 U47265 ( .I(n46613), .ZN(n53221) );
  NAND2HSV2 U47266 ( .A1(n53221), .A2(\pe3/pvq [22]), .ZN(n43060) );
  XOR2HSV0 U47267 ( .A1(n43060), .A2(\pe3/phq [22]), .Z(n43061) );
  XOR2HSV0 U47268 ( .A1(n43062), .A2(n43061), .Z(n43063) );
  XOR2HSV0 U47269 ( .A1(n43064), .A2(n43063), .Z(n43065) );
  XOR2HSV0 U47270 ( .A1(n43066), .A2(n43065), .Z(n43085) );
  INHSV2 U47271 ( .I(\pe3/bq[11] ), .ZN(n56001) );
  CLKNAND2HSV1 U47272 ( .A1(n43650), .A2(\pe3/bq[11] ), .ZN(n43409) );
  OAI22HSV0 U47273 ( .A1(n59606), .A2(n56001), .B1(n43757), .B2(n49423), .ZN(
        n43067) );
  OAI21HSV0 U47274 ( .A1(n43068), .A2(n43409), .B(n43067), .ZN(n43069) );
  XNOR2HSV1 U47275 ( .A1(n43069), .A2(n55717), .ZN(n43073) );
  XOR2HSV0 U47276 ( .A1(n43071), .A2(n43070), .Z(n43072) );
  XNOR2HSV1 U47277 ( .A1(n43073), .A2(n43072), .ZN(n43081) );
  INHSV2 U47278 ( .I(n53229), .ZN(n45676) );
  CLKNAND2HSV0 U47279 ( .A1(n45676), .A2(n48538), .ZN(n43075) );
  NAND2HSV0 U47280 ( .A1(n43280), .A2(n43389), .ZN(n43074) );
  XOR2HSV0 U47281 ( .A1(n43075), .A2(n43074), .Z(n43079) );
  NAND2HSV0 U47282 ( .A1(n56651), .A2(n55867), .ZN(n43077) );
  CLKNAND2HSV0 U47283 ( .A1(n45640), .A2(n43809), .ZN(n43076) );
  XOR2HSV0 U47284 ( .A1(n43077), .A2(n43076), .Z(n43078) );
  XOR2HSV0 U47285 ( .A1(n43079), .A2(n43078), .Z(n43080) );
  XOR2HSV0 U47286 ( .A1(n43081), .A2(n43080), .Z(n43083) );
  NAND2HSV0 U47287 ( .A1(n43424), .A2(n59966), .ZN(n43082) );
  XNOR2HSV1 U47288 ( .A1(n43083), .A2(n43082), .ZN(n43084) );
  XOR2HSV0 U47289 ( .A1(n43085), .A2(n43084), .Z(n43090) );
  NAND2HSV0 U47290 ( .A1(n48511), .A2(n56493), .ZN(n43087) );
  NAND2HSV0 U47291 ( .A1(n45950), .A2(n43829), .ZN(n43086) );
  XNOR2HSV1 U47292 ( .A1(n43087), .A2(n43086), .ZN(n43089) );
  CLKNAND2HSV1 U47293 ( .A1(n52727), .A2(n59624), .ZN(n43088) );
  XOR3HSV2 U47294 ( .A1(n43090), .A2(n43089), .A3(n43088), .Z(n43091) );
  XOR2HSV0 U47295 ( .A1(n43092), .A2(n43091), .Z(n43093) );
  XOR2HSV0 U47296 ( .A1(n43094), .A2(n43093), .Z(n43096) );
  NAND2HSV0 U47297 ( .A1(n43211), .A2(n43374), .ZN(n43095) );
  XOR2HSV0 U47298 ( .A1(n43096), .A2(n43095), .Z(n43099) );
  NAND2HSV0 U47299 ( .A1(n43097), .A2(n42937), .ZN(n43098) );
  XNOR2HSV1 U47300 ( .A1(n43099), .A2(n43098), .ZN(n43100) );
  XNOR2HSV1 U47301 ( .A1(n43101), .A2(n43100), .ZN(n43102) );
  XNOR2HSV1 U47302 ( .A1(n43103), .A2(n43102), .ZN(n43104) );
  NOR2HSV2 U47303 ( .A1(n46519), .A2(n42817), .ZN(n43105) );
  CLKNAND2HSV0 U47304 ( .A1(n25893), .A2(n46311), .ZN(n43107) );
  XOR3HSV2 U47305 ( .A1(n43109), .A2(n43108), .A3(n43107), .Z(n43110) );
  CLKBUFHSV4 U47306 ( .I(n46415), .Z(n46052) );
  CLKNAND2HSV1 U47307 ( .A1(n46052), .A2(n45633), .ZN(n43112) );
  CLKNHSV2 U47308 ( .I(n43112), .ZN(n43113) );
  XNOR2HSV4 U47309 ( .A1(n43114), .A2(n43113), .ZN(n43115) );
  XNOR2HSV4 U47310 ( .A1(n43116), .A2(n43115), .ZN(n43118) );
  XNOR2HSV4 U47311 ( .A1(n43118), .A2(n43117), .ZN(n43240) );
  NOR2HSV0 U47312 ( .A1(n46559), .A2(n37264), .ZN(n43119) );
  NAND2HSV0 U47313 ( .A1(n43127), .A2(n43119), .ZN(n43122) );
  NOR2HSV0 U47314 ( .A1(n43604), .A2(n43120), .ZN(n43248) );
  INHSV2 U47315 ( .I(n43248), .ZN(n43121) );
  CLKNAND2HSV1 U47316 ( .A1(n43126), .A2(n52726), .ZN(n45616) );
  NOR2HSV2 U47317 ( .A1(n43127), .A2(n45616), .ZN(n43128) );
  NOR2HSV0 U47318 ( .A1(n43143), .A2(n43142), .ZN(n43131) );
  NOR2HSV0 U47319 ( .A1(n43912), .A2(n43361), .ZN(n45753) );
  NOR2HSV1 U47320 ( .A1(n43240), .A2(n37268), .ZN(n43138) );
  INHSV2 U47321 ( .I(n37169), .ZN(n43867) );
  CLKBUFHSV4 U47322 ( .I(n43621), .Z(n43754) );
  CLKNAND2HSV2 U47323 ( .A1(n43754), .A2(n46311), .ZN(n43230) );
  NAND2HSV0 U47324 ( .A1(n55948), .A2(n59965), .ZN(n43221) );
  CLKNAND2HSV0 U47325 ( .A1(n43373), .A2(\pe3/got [18]), .ZN(n43219) );
  BUFHSV2 U47326 ( .I(n47991), .Z(n43495) );
  CLKNAND2HSV0 U47327 ( .A1(n43495), .A2(n56335), .ZN(n43217) );
  NAND2HSV0 U47328 ( .A1(n55825), .A2(n56493), .ZN(n43210) );
  BUFHSV2 U47329 ( .I(n55951), .Z(n46314) );
  NAND2HSV0 U47330 ( .A1(n46314), .A2(\pe3/got [13]), .ZN(n43208) );
  NAND2HSV0 U47331 ( .A1(n56113), .A2(n56213), .ZN(n43145) );
  NAND2HSV0 U47332 ( .A1(n37373), .A2(\pe3/bq[11] ), .ZN(n43144) );
  XOR2HSV0 U47333 ( .A1(n43145), .A2(n43144), .Z(n43150) );
  NAND2HSV0 U47334 ( .A1(n42950), .A2(n43146), .ZN(n43148) );
  CLKNAND2HSV0 U47335 ( .A1(\pe3/aot [15]), .A2(n48520), .ZN(n43147) );
  XOR2HSV0 U47336 ( .A1(n43148), .A2(n43147), .Z(n43149) );
  XOR2HSV0 U47337 ( .A1(n43150), .A2(n43149), .Z(n43159) );
  INHSV1 U47338 ( .I(n43151), .ZN(n45952) );
  NAND2HSV0 U47339 ( .A1(n45952), .A2(n43780), .ZN(n43153) );
  NAND2HSV0 U47340 ( .A1(\pe3/aot [8]), .A2(n43499), .ZN(n43152) );
  XOR2HSV0 U47341 ( .A1(n43153), .A2(n43152), .Z(n43157) );
  NAND2HSV0 U47342 ( .A1(\pe3/aot [22]), .A2(\pe3/bq[18] ), .ZN(n43155) );
  NAND2HSV0 U47343 ( .A1(n55750), .A2(n43775), .ZN(n43154) );
  XOR2HSV0 U47344 ( .A1(n43155), .A2(n43154), .Z(n43156) );
  XOR2HSV0 U47345 ( .A1(n43157), .A2(n43156), .Z(n43158) );
  XOR2HSV0 U47346 ( .A1(n43159), .A2(n43158), .Z(n43175) );
  NAND2HSV0 U47347 ( .A1(n56204), .A2(n42971), .ZN(n43161) );
  CLKNHSV1 U47348 ( .I(n56269), .ZN(n56187) );
  NAND2HSV0 U47349 ( .A1(n48496), .A2(n56187), .ZN(n43160) );
  XOR2HSV0 U47350 ( .A1(n43161), .A2(n43160), .Z(n43165) );
  NAND2HSV0 U47351 ( .A1(n45962), .A2(n56454), .ZN(n43163) );
  NAND2HSV0 U47352 ( .A1(n45676), .A2(n43539), .ZN(n43162) );
  XOR2HSV0 U47353 ( .A1(n43163), .A2(n43162), .Z(n43164) );
  XOR2HSV0 U47354 ( .A1(n43165), .A2(n43164), .Z(n43173) );
  NOR2HSV0 U47355 ( .A1(n42539), .A2(n46131), .ZN(n43167) );
  BUFHSV2 U47356 ( .I(\pe3/aot [24]), .Z(n46332) );
  CLKNAND2HSV0 U47357 ( .A1(n46332), .A2(n43544), .ZN(n43166) );
  XOR2HSV0 U47358 ( .A1(n43167), .A2(n43166), .Z(n43171) );
  NAND2HSV0 U47359 ( .A1(\pe3/aot [23]), .A2(n56519), .ZN(n43169) );
  NAND2HSV0 U47360 ( .A1(\pe3/aot [14]), .A2(\pe3/bq[26] ), .ZN(n43168) );
  XOR2HSV0 U47361 ( .A1(n43169), .A2(n43168), .Z(n43170) );
  XOR2HSV0 U47362 ( .A1(n43171), .A2(n43170), .Z(n43172) );
  XOR2HSV0 U47363 ( .A1(n43173), .A2(n43172), .Z(n43174) );
  XOR2HSV0 U47364 ( .A1(n43175), .A2(n43174), .Z(n43177) );
  NAND2HSV0 U47365 ( .A1(n42710), .A2(n56558), .ZN(n43176) );
  XOR2HSV0 U47366 ( .A1(n43177), .A2(n43176), .Z(n43206) );
  INHSV2 U47367 ( .I(n50799), .ZN(n56557) );
  NAND2HSV0 U47368 ( .A1(n43516), .A2(n56557), .ZN(n43203) );
  CLKNAND2HSV0 U47369 ( .A1(n45645), .A2(n43052), .ZN(n43180) );
  INHSV2 U47370 ( .I(n49423), .ZN(n56644) );
  NAND2HSV0 U47371 ( .A1(n46456), .A2(n56644), .ZN(n43179) );
  XOR2HSV0 U47372 ( .A1(n43180), .A2(n43179), .Z(n43184) );
  NAND2HSV0 U47373 ( .A1(\pe3/got [8]), .A2(n37007), .ZN(n43181) );
  XOR2HSV0 U47374 ( .A1(n43182), .A2(n43181), .Z(n43183) );
  XOR2HSV0 U47375 ( .A1(n43184), .A2(n43183), .Z(n43201) );
  BUFHSV2 U47376 ( .I(n43185), .Z(n59648) );
  INHSV4 U47377 ( .I(n56680), .ZN(n56620) );
  NAND2HSV0 U47378 ( .A1(n43424), .A2(n56620), .ZN(n43200) );
  NAND2HSV0 U47379 ( .A1(n56464), .A2(n49439), .ZN(n43187) );
  NAND2HSV0 U47380 ( .A1(n59960), .A2(n45663), .ZN(n43186) );
  XOR2HSV0 U47381 ( .A1(n43187), .A2(n43186), .Z(n43191) );
  NAND2HSV0 U47382 ( .A1(n56520), .A2(n48538), .ZN(n43189) );
  BUFHSV2 U47383 ( .I(\pe3/aot [11]), .Z(n59623) );
  CLKNHSV0 U47384 ( .I(n36694), .ZN(n43793) );
  NAND2HSV0 U47385 ( .A1(n59623), .A2(n43793), .ZN(n43188) );
  XOR2HSV0 U47386 ( .A1(n43189), .A2(n43188), .Z(n43190) );
  XOR2HSV0 U47387 ( .A1(n43191), .A2(n43190), .Z(n43198) );
  CLKNAND2HSV1 U47388 ( .A1(n46124), .A2(\pe3/pvq [25]), .ZN(n43192) );
  XOR2HSV0 U47389 ( .A1(n43192), .A2(\pe3/phq [25]), .Z(n43196) );
  NAND2HSV0 U47390 ( .A1(n48530), .A2(n56785), .ZN(n46014) );
  OAI22HSV0 U47391 ( .A1(n45691), .A2(n56277), .B1(n55714), .B2(n46615), .ZN(
        n43193) );
  OAI21HSV0 U47392 ( .A1(n43194), .A2(n46014), .B(n43193), .ZN(n43195) );
  XOR2HSV0 U47393 ( .A1(n43196), .A2(n43195), .Z(n43197) );
  XNOR2HSV1 U47394 ( .A1(n43198), .A2(n43197), .ZN(n43199) );
  XOR3HSV2 U47395 ( .A1(n43201), .A2(n43200), .A3(n43199), .Z(n43202) );
  XNOR2HSV1 U47396 ( .A1(n43203), .A2(n43202), .ZN(n43205) );
  CLKNHSV0 U47397 ( .I(n50802), .ZN(n43756) );
  CLKNAND2HSV0 U47398 ( .A1(n37353), .A2(n43756), .ZN(n43204) );
  XOR3HSV2 U47399 ( .A1(n43206), .A2(n43205), .A3(n43204), .Z(n43207) );
  XOR2HSV0 U47400 ( .A1(n43208), .A2(n43207), .Z(n43209) );
  XOR2HSV0 U47401 ( .A1(n43210), .A2(n43209), .Z(n43213) );
  CLKNAND2HSV1 U47402 ( .A1(n43211), .A2(n48584), .ZN(n43212) );
  XOR2HSV0 U47403 ( .A1(n43213), .A2(n43212), .Z(n43215) );
  CLKNHSV0 U47404 ( .I(n37326), .ZN(n56127) );
  NAND2HSV0 U47405 ( .A1(n56127), .A2(n49252), .ZN(n43214) );
  XNOR2HSV1 U47406 ( .A1(n43215), .A2(n43214), .ZN(n43216) );
  XNOR2HSV1 U47407 ( .A1(n43217), .A2(n43216), .ZN(n43218) );
  XNOR2HSV1 U47408 ( .A1(n43219), .A2(n43218), .ZN(n43220) );
  XNOR2HSV1 U47409 ( .A1(n43221), .A2(n43220), .ZN(n43225) );
  NOR2HSV2 U47410 ( .A1(n45728), .A2(n45635), .ZN(n43224) );
  INHSV1 U47411 ( .I(n46519), .ZN(n56136) );
  NAND2HSV2 U47412 ( .A1(n56136), .A2(n55945), .ZN(n43223) );
  XOR3HSV2 U47413 ( .A1(n43225), .A2(n43224), .A3(n43223), .Z(n43229) );
  CLKNHSV1 U47414 ( .I(n43706), .ZN(n43577) );
  NOR2HSV1 U47415 ( .A1(n43577), .A2(n49314), .ZN(n43228) );
  BUFHSV2 U47416 ( .I(n25893), .Z(n59810) );
  NAND2HSV2 U47417 ( .A1(n45732), .A2(\pe3/got [23]), .ZN(n43227) );
  XNOR2HSV4 U47418 ( .A1(n43230), .A2(n29659), .ZN(n43239) );
  CLKBUFHSV4 U47419 ( .I(n46052), .Z(n43850) );
  CLKNAND2HSV1 U47420 ( .A1(n43850), .A2(n43452), .ZN(n43233) );
  CLKBUFHSV4 U47421 ( .I(n42918), .Z(n47430) );
  CLKNHSV0 U47422 ( .I(n43855), .ZN(n43231) );
  NOR2HSV2 U47423 ( .A1(n47430), .A2(n43231), .ZN(n43232) );
  XNOR2HSV4 U47424 ( .A1(n43233), .A2(n43232), .ZN(n43237) );
  CLKNHSV0 U47425 ( .I(\pe3/ti_7t [22]), .ZN(n43243) );
  AO21HSV1 U47426 ( .A1(n43243), .A2(n43242), .B(n45628), .Z(n43244) );
  AND2HSV2 U47427 ( .A1(n43246), .A2(n45755), .Z(n43257) );
  INHSV2 U47428 ( .I(n43257), .ZN(n43247) );
  CLKNAND2HSV0 U47429 ( .A1(n43248), .A2(n43898), .ZN(n43258) );
  CLKNHSV2 U47430 ( .I(n43258), .ZN(n43249) );
  NOR2HSV0 U47431 ( .A1(n46438), .A2(n45932), .ZN(n43261) );
  CLKNHSV0 U47432 ( .I(n43261), .ZN(n43251) );
  OAI21HSV0 U47433 ( .A1(n43257), .A2(n45625), .B(n45755), .ZN(n43250) );
  AO21HSV1 U47434 ( .A1(n43258), .A2(n43251), .B(n43250), .Z(n43252) );
  NOR2HSV2 U47435 ( .A1(n43253), .A2(n43252), .ZN(n43254) );
  INOR2HSV1 U47436 ( .A1(n43258), .B1(n43257), .ZN(n43259) );
  CLKNHSV2 U47437 ( .I(n43259), .ZN(n43260) );
  NAND2HSV2 U47438 ( .A1(n43754), .A2(n46309), .ZN(n43343) );
  NAND2HSV2 U47439 ( .A1(n59821), .A2(n45633), .ZN(n43339) );
  CLKNAND2HSV0 U47440 ( .A1(n55948), .A2(n43262), .ZN(n43331) );
  CLKNAND2HSV1 U47441 ( .A1(n43373), .A2(n49404), .ZN(n43329) );
  NAND2HSV2 U47442 ( .A1(n43495), .A2(n42937), .ZN(n43327) );
  NAND2HSV0 U47443 ( .A1(n49405), .A2(n43437), .ZN(n43321) );
  CLKNAND2HSV1 U47444 ( .A1(n48488), .A2(n59624), .ZN(n43319) );
  CLKNAND2HSV0 U47445 ( .A1(n56740), .A2(n43499), .ZN(n43264) );
  INHSV1 U47446 ( .I(n53229), .ZN(n59959) );
  NAND2HSV0 U47447 ( .A1(n59959), .A2(n43389), .ZN(n43263) );
  XOR2HSV0 U47448 ( .A1(n43264), .A2(n43263), .Z(n43269) );
  NAND2HSV0 U47449 ( .A1(n43265), .A2(\pe3/bq[11] ), .ZN(n43267) );
  NAND2HSV0 U47450 ( .A1(n56558), .A2(n37051), .ZN(n43266) );
  XOR2HSV0 U47451 ( .A1(n43267), .A2(n43266), .Z(n43268) );
  XOR2HSV0 U47452 ( .A1(n43269), .A2(n43268), .Z(n43277) );
  NAND2HSV0 U47453 ( .A1(n45962), .A2(\pe3/bq[10] ), .ZN(n43271) );
  NAND2HSV0 U47454 ( .A1(\pe3/aot [22]), .A2(n42971), .ZN(n43270) );
  XOR2HSV0 U47455 ( .A1(n43271), .A2(n43270), .Z(n43275) );
  NAND2HSV0 U47456 ( .A1(n59623), .A2(n48538), .ZN(n43273) );
  CLKNAND2HSV0 U47457 ( .A1(n45640), .A2(n56379), .ZN(n43272) );
  XOR2HSV0 U47458 ( .A1(n43273), .A2(n43272), .Z(n43274) );
  XOR2HSV0 U47459 ( .A1(n43275), .A2(n43274), .Z(n43276) );
  XOR2HSV0 U47460 ( .A1(n43277), .A2(n43276), .Z(n43294) );
  NAND2HSV0 U47461 ( .A1(n56464), .A2(\pe3/bq[23] ), .ZN(n43279) );
  CLKNAND2HSV1 U47462 ( .A1(n46363), .A2(n56071), .ZN(n43278) );
  XOR2HSV0 U47463 ( .A1(n43279), .A2(n43278), .Z(n43284) );
  CLKNAND2HSV1 U47464 ( .A1(n43650), .A2(n43775), .ZN(n43282) );
  CLKNAND2HSV0 U47465 ( .A1(n43280), .A2(n43793), .ZN(n43281) );
  XOR2HSV0 U47466 ( .A1(n43282), .A2(n43281), .Z(n43283) );
  XOR2HSV0 U47467 ( .A1(n43284), .A2(n43283), .Z(n43292) );
  NOR2HSV0 U47468 ( .A1(n42539), .A2(n43039), .ZN(n43286) );
  CLKNAND2HSV0 U47469 ( .A1(n45645), .A2(\pe3/bq[26] ), .ZN(n43285) );
  XOR2HSV0 U47470 ( .A1(n43286), .A2(n43285), .Z(n43290) );
  NAND2HSV0 U47471 ( .A1(n42950), .A2(n55872), .ZN(n43288) );
  NAND2HSV0 U47472 ( .A1(n42818), .A2(\pe3/bq[19] ), .ZN(n43287) );
  XOR2HSV0 U47473 ( .A1(n43288), .A2(n43287), .Z(n43289) );
  XOR2HSV0 U47474 ( .A1(n43290), .A2(n43289), .Z(n43291) );
  XOR2HSV0 U47475 ( .A1(n43292), .A2(n43291), .Z(n43293) );
  XOR2HSV0 U47476 ( .A1(n43294), .A2(n43293), .Z(n43296) );
  CLKNHSV0 U47477 ( .I(n50802), .ZN(n43496) );
  NAND2HSV0 U47478 ( .A1(n45950), .A2(n43496), .ZN(n43295) );
  XOR2HSV0 U47479 ( .A1(n43296), .A2(n43295), .Z(n43317) );
  NOR2HSV0 U47480 ( .A1(n45564), .A2(n46138), .ZN(n43298) );
  NAND2HSV0 U47481 ( .A1(n56204), .A2(n43772), .ZN(n43297) );
  XOR2HSV0 U47482 ( .A1(n43298), .A2(n43297), .Z(n43302) );
  NAND2HSV0 U47483 ( .A1(n56378), .A2(n43780), .ZN(n43300) );
  NAND2HSV0 U47484 ( .A1(n56188), .A2(n55867), .ZN(n43299) );
  XOR2HSV0 U47485 ( .A1(n43300), .A2(n43299), .Z(n43301) );
  XOR2HSV0 U47486 ( .A1(n43302), .A2(n43301), .Z(n43312) );
  NAND2HSV0 U47487 ( .A1(n45648), .A2(n56644), .ZN(n43304) );
  CLKNAND2HSV0 U47488 ( .A1(n46332), .A2(\pe3/bq[18] ), .ZN(n43303) );
  XOR2HSV0 U47489 ( .A1(n43304), .A2(n43303), .Z(n43307) );
  INHSV2 U47490 ( .I(n46613), .ZN(n46127) );
  NAND2HSV2 U47491 ( .A1(n46127), .A2(\pe3/pvq [23]), .ZN(n43305) );
  XNOR2HSV1 U47492 ( .A1(n43305), .A2(\pe3/phq [23]), .ZN(n43306) );
  XNOR2HSV1 U47493 ( .A1(n43307), .A2(n43306), .ZN(n43309) );
  CLKNAND2HSV0 U47494 ( .A1(n46456), .A2(n43809), .ZN(n55724) );
  NAND2HSV2 U47495 ( .A1(n48530), .A2(n56519), .ZN(n56099) );
  XOR2HSV0 U47496 ( .A1(n55724), .A2(n56099), .Z(n43308) );
  XNOR2HSV1 U47497 ( .A1(n43309), .A2(n43308), .ZN(n43311) );
  NAND2HSV0 U47498 ( .A1(n43424), .A2(n56557), .ZN(n43310) );
  XOR3HSV2 U47499 ( .A1(n43312), .A2(n43311), .A3(n43310), .Z(n43313) );
  XNOR2HSV1 U47500 ( .A1(n43314), .A2(n43313), .ZN(n43316) );
  NAND2HSV2 U47501 ( .A1(n55826), .A2(n56493), .ZN(n43315) );
  XOR3HSV2 U47502 ( .A1(n43317), .A2(n43316), .A3(n43315), .Z(n43318) );
  XOR2HSV0 U47503 ( .A1(n43319), .A2(n43318), .Z(n43320) );
  XOR2HSV0 U47504 ( .A1(n43321), .A2(n43320), .Z(n43323) );
  CLKNAND2HSV1 U47505 ( .A1(n46313), .A2(n56064), .ZN(n43322) );
  XOR2HSV0 U47506 ( .A1(n43323), .A2(n43322), .Z(n43325) );
  CLKNHSV0 U47507 ( .I(n37326), .ZN(n55895) );
  NAND2HSV0 U47508 ( .A1(n55895), .A2(n43374), .ZN(n43324) );
  XNOR2HSV1 U47509 ( .A1(n43325), .A2(n43324), .ZN(n43326) );
  XNOR2HSV1 U47510 ( .A1(n43327), .A2(n43326), .ZN(n43328) );
  XNOR2HSV1 U47511 ( .A1(n43329), .A2(n43328), .ZN(n43330) );
  XNOR2HSV1 U47512 ( .A1(n43331), .A2(n43330), .ZN(n43334) );
  NOR2HSV1 U47513 ( .A1(n43448), .A2(n49314), .ZN(n43333) );
  NAND2HSV2 U47514 ( .A1(n49468), .A2(n42673), .ZN(n43332) );
  XOR3HSV2 U47515 ( .A1(n43334), .A2(n43333), .A3(n43332), .Z(n43337) );
  NOR2HSV2 U47516 ( .A1(n43577), .A2(n42817), .ZN(n43336) );
  NAND2HSV0 U47517 ( .A1(n43453), .A2(n46441), .ZN(n43335) );
  XOR3HSV2 U47518 ( .A1(n43337), .A2(n43336), .A3(n43335), .Z(n43338) );
  XNOR2HSV1 U47519 ( .A1(n43339), .A2(n43338), .ZN(n43341) );
  NAND2HSV2 U47520 ( .A1(n43850), .A2(n46311), .ZN(n43340) );
  XOR2HSV0 U47521 ( .A1(n43341), .A2(n43340), .Z(n43342) );
  XNOR2HSV1 U47522 ( .A1(n43343), .A2(n43342), .ZN(n43346) );
  XNOR2HSV1 U47523 ( .A1(n43346), .A2(n43345), .ZN(n43351) );
  INHSV2 U47524 ( .I(n43351), .ZN(n43347) );
  NAND2HSV4 U47525 ( .A1(n43357), .A2(n43356), .ZN(n43592) );
  CLKNHSV2 U47526 ( .I(n43359), .ZN(n43363) );
  CLKNAND2HSV4 U47527 ( .A1(n43368), .A2(n43367), .ZN(n43742) );
  INHSV2 U47528 ( .I(n43479), .ZN(n43369) );
  OAI21HSV0 U47529 ( .A1(n36972), .A2(\pe3/ti_7t [24]), .B(n44669), .ZN(n43477) );
  INHSV2 U47530 ( .I(n43477), .ZN(n43482) );
  NOR2HSV4 U47531 ( .A1(n59575), .A2(n43370), .ZN(n43476) );
  INHSV2 U47532 ( .I(n45635), .ZN(n45581) );
  NAND2HSV2 U47533 ( .A1(n43755), .A2(n45581), .ZN(n43447) );
  CLKNAND2HSV0 U47534 ( .A1(n43373), .A2(n42937), .ZN(n43445) );
  CLKNAND2HSV1 U47535 ( .A1(n43495), .A2(n43374), .ZN(n43443) );
  NAND2HSV0 U47536 ( .A1(n55707), .A2(n48584), .ZN(n43436) );
  CLKNAND2HSV1 U47537 ( .A1(n46314), .A2(n56493), .ZN(n43434) );
  NAND2HSV0 U47538 ( .A1(n42950), .A2(\pe3/bq[23] ), .ZN(n43376) );
  CLKNAND2HSV0 U47539 ( .A1(n46332), .A2(n56519), .ZN(n43375) );
  XOR2HSV0 U47540 ( .A1(n43376), .A2(n43375), .Z(n43380) );
  NAND2HSV0 U47541 ( .A1(n56464), .A2(n43772), .ZN(n43378) );
  NAND2HSV0 U47542 ( .A1(n56182), .A2(n42971), .ZN(n43377) );
  XOR2HSV0 U47543 ( .A1(n43378), .A2(n43377), .Z(n43379) );
  XOR2HSV0 U47544 ( .A1(n43380), .A2(n43379), .Z(n43388) );
  CLKNAND2HSV0 U47545 ( .A1(n48530), .A2(n43544), .ZN(n43382) );
  NAND2HSV0 U47546 ( .A1(n46456), .A2(n56379), .ZN(n43381) );
  XOR2HSV0 U47547 ( .A1(n43382), .A2(n43381), .Z(n43386) );
  NAND2HSV0 U47548 ( .A1(\pe3/aot [23]), .A2(\pe3/bq[18] ), .ZN(n43384) );
  NAND2HSV0 U47549 ( .A1(n45648), .A2(n43775), .ZN(n43383) );
  XOR2HSV0 U47550 ( .A1(n43384), .A2(n43383), .Z(n43385) );
  XOR2HSV0 U47551 ( .A1(n43386), .A2(n43385), .Z(n43387) );
  XOR2HSV0 U47552 ( .A1(n43388), .A2(n43387), .Z(n43406) );
  NAND2HSV0 U47553 ( .A1(n59623), .A2(n43389), .ZN(n43391) );
  CLKNAND2HSV0 U47554 ( .A1(n46363), .A2(n55872), .ZN(n43390) );
  XOR2HSV0 U47555 ( .A1(n43391), .A2(n43390), .Z(n43396) );
  NAND2HSV0 U47556 ( .A1(\pe3/aot [14]), .A2(n43780), .ZN(n43394) );
  CLKNAND2HSV1 U47557 ( .A1(n43265), .A2(\pe3/bq[10] ), .ZN(n43393) );
  XOR2HSV0 U47558 ( .A1(n43394), .A2(n43393), .Z(n43395) );
  XOR2HSV0 U47559 ( .A1(n43396), .A2(n43395), .Z(n43404) );
  NOR2HSV0 U47560 ( .A1(n45555), .A2(n49423), .ZN(n43398) );
  INHSV2 U47561 ( .I(n56567), .ZN(n56423) );
  NAND2HSV0 U47562 ( .A1(n56423), .A2(n43499), .ZN(n43397) );
  XOR2HSV0 U47563 ( .A1(n43398), .A2(n43397), .Z(n43402) );
  CLKNAND2HSV1 U47564 ( .A1(n56651), .A2(\pe3/bq[26] ), .ZN(n43400) );
  NAND2HSV0 U47565 ( .A1(n59960), .A2(n48538), .ZN(n43399) );
  XOR2HSV0 U47566 ( .A1(n43400), .A2(n43399), .Z(n43401) );
  XOR2HSV0 U47567 ( .A1(n43402), .A2(n43401), .Z(n43403) );
  XOR2HSV0 U47568 ( .A1(n43404), .A2(n43403), .Z(n43405) );
  XOR2HSV0 U47569 ( .A1(n43406), .A2(n43405), .Z(n43408) );
  NAND2HSV0 U47570 ( .A1(n59797), .A2(n56557), .ZN(n43407) );
  XOR2HSV0 U47571 ( .A1(n43408), .A2(n43407), .Z(n43432) );
  NAND2HSV0 U47572 ( .A1(n43516), .A2(n43496), .ZN(n43429) );
  CLKNAND2HSV1 U47573 ( .A1(n45952), .A2(n43539), .ZN(n48512) );
  XOR2HSV0 U47574 ( .A1(n43409), .A2(n48512), .Z(n43413) );
  CLKNAND2HSV0 U47575 ( .A1(n45676), .A2(n43793), .ZN(n43411) );
  NAND2HSV0 U47576 ( .A1(n56620), .A2(n45955), .ZN(n43410) );
  XOR2HSV0 U47577 ( .A1(n43411), .A2(n43410), .Z(n43412) );
  XOR2HSV0 U47578 ( .A1(n43413), .A2(n43412), .Z(n43427) );
  NAND2HSV0 U47579 ( .A1(n42743), .A2(n43809), .ZN(n43415) );
  CLKNAND2HSV0 U47580 ( .A1(n45645), .A2(n48520), .ZN(n43414) );
  XOR2HSV0 U47581 ( .A1(n43415), .A2(n43414), .Z(n43418) );
  CLKNAND2HSV1 U47582 ( .A1(n53221), .A2(\pe3/pvq [24]), .ZN(n43416) );
  XNOR2HSV1 U47583 ( .A1(n43416), .A2(\pe3/phq [24]), .ZN(n43417) );
  XNOR2HSV1 U47584 ( .A1(n43418), .A2(n43417), .ZN(n43423) );
  NOR2HSV0 U47585 ( .A1(n37357), .A2(n56277), .ZN(n55829) );
  AOI22HSV0 U47586 ( .A1(n45962), .A2(n53232), .B1(n56106), .B2(\pe3/aot [20]), 
        .ZN(n43419) );
  AOI21HSV0 U47587 ( .A1(n43420), .A2(n55829), .B(n43419), .ZN(n43421) );
  NAND2HSV0 U47588 ( .A1(\pe3/aot [22]), .A2(\pe3/bq[19] ), .ZN(n55638) );
  XOR2HSV0 U47589 ( .A1(n43421), .A2(n55638), .Z(n43422) );
  XNOR2HSV1 U47590 ( .A1(n43423), .A2(n43422), .ZN(n43426) );
  NAND2HSV0 U47591 ( .A1(n43424), .A2(n56558), .ZN(n43425) );
  XOR3HSV2 U47592 ( .A1(n43427), .A2(n43426), .A3(n43425), .Z(n43428) );
  XNOR2HSV1 U47593 ( .A1(n43429), .A2(n43428), .ZN(n43431) );
  CLKNAND2HSV1 U47594 ( .A1(n55826), .A2(n43829), .ZN(n43430) );
  XOR3HSV2 U47595 ( .A1(n43432), .A2(n43431), .A3(n43430), .Z(n43433) );
  XOR2HSV0 U47596 ( .A1(n43434), .A2(n43433), .Z(n43435) );
  XOR2HSV0 U47597 ( .A1(n43436), .A2(n43435), .Z(n43439) );
  CLKNAND2HSV0 U47598 ( .A1(n46313), .A2(n43437), .ZN(n43438) );
  XOR2HSV0 U47599 ( .A1(n43439), .A2(n43438), .Z(n43441) );
  NAND2HSV0 U47600 ( .A1(n56127), .A2(n56335), .ZN(n43440) );
  XNOR2HSV1 U47601 ( .A1(n43441), .A2(n43440), .ZN(n43442) );
  XNOR2HSV1 U47602 ( .A1(n43443), .A2(n43442), .ZN(n43444) );
  XNOR2HSV1 U47603 ( .A1(n43445), .A2(n43444), .ZN(n43446) );
  XNOR2HSV1 U47604 ( .A1(n43447), .A2(n43446), .ZN(n43451) );
  NOR2HSV1 U47605 ( .A1(n43448), .A2(n37275), .ZN(n43450) );
  CLKNAND2HSV1 U47606 ( .A1(n56136), .A2(n42770), .ZN(n43449) );
  XOR3HSV2 U47607 ( .A1(n43451), .A2(n43450), .A3(n43449), .Z(n43456) );
  NOR2HSV2 U47608 ( .A1(n43577), .A2(n42827), .ZN(n43455) );
  NAND2HSV0 U47609 ( .A1(n43453), .A2(n43452), .ZN(n43454) );
  XOR3HSV2 U47610 ( .A1(n43456), .A2(n43455), .A3(n43454), .Z(n43460) );
  NOR2HSV2 U47611 ( .A1(n47430), .A2(n43457), .ZN(n43459) );
  CLKNAND2HSV1 U47612 ( .A1(n43850), .A2(n46441), .ZN(n43458) );
  XOR3HSV2 U47613 ( .A1(n43460), .A2(n43459), .A3(n43458), .Z(n43462) );
  CLKNAND2HSV1 U47614 ( .A1(n43621), .A2(n45633), .ZN(n43461) );
  NAND3HSV4 U47615 ( .A1(n43473), .A2(n43471), .A3(n43472), .ZN(n43474) );
  NAND2HSV4 U47616 ( .A1(n43475), .A2(n43474), .ZN(n43600) );
  INHSV4 U47617 ( .I(n43600), .ZN(n43612) );
  INHSV2 U47618 ( .I(n43871), .ZN(n43478) );
  NOR2HSV4 U47619 ( .A1(n43479), .A2(n43478), .ZN(n43480) );
  NAND3HSV3 U47620 ( .A1(n43609), .A2(n43600), .A3(n43482), .ZN(n43740) );
  INHSV4 U47621 ( .I(n43742), .ZN(n43738) );
  NAND3HSV2 U47622 ( .A1(n43739), .A2(n43740), .A3(n43484), .ZN(n43485) );
  AND2HSV2 U47623 ( .A1(n43139), .A2(n44669), .Z(n43489) );
  NAND2HSV0 U47624 ( .A1(n43493), .A2(n43489), .ZN(n43492) );
  CLKNAND2HSV1 U47625 ( .A1(n43490), .A2(n43139), .ZN(n43491) );
  BUFHSV4 U47626 ( .I(n43493), .Z(n56265) );
  NAND2HSV2 U47627 ( .A1(n45583), .A2(n45633), .ZN(n43590) );
  NAND2HSV2 U47628 ( .A1(n43754), .A2(n43855), .ZN(n43586) );
  NAND2HSV2 U47629 ( .A1(n59821), .A2(n55701), .ZN(n43582) );
  CLKNAND2HSV1 U47630 ( .A1(n43755), .A2(\pe3/got [18]), .ZN(n43573) );
  NAND2HSV0 U47631 ( .A1(n59625), .A2(n56335), .ZN(n43571) );
  CLKNAND2HSV0 U47632 ( .A1(n43495), .A2(n49252), .ZN(n43569) );
  NAND2HSV0 U47633 ( .A1(n55707), .A2(n43829), .ZN(n43563) );
  CLKNAND2HSV1 U47634 ( .A1(n46314), .A2(n43496), .ZN(n43561) );
  BUFHSV2 U47635 ( .I(n37017), .Z(n45950) );
  NAND2HSV0 U47636 ( .A1(n45950), .A2(n56620), .ZN(n43515) );
  CLKNAND2HSV1 U47637 ( .A1(\pe3/aot [14]), .A2(n48520), .ZN(n43498) );
  CLKNAND2HSV0 U47638 ( .A1(\pe3/aot [15]), .A2(n42530), .ZN(n43497) );
  XOR2HSV0 U47639 ( .A1(n43498), .A2(n43497), .Z(n43503) );
  NAND2HSV0 U47640 ( .A1(n56864), .A2(n43499), .ZN(n43501) );
  INHSV2 U47641 ( .I(n56778), .ZN(n56771) );
  NAND2HSV0 U47642 ( .A1(n56771), .A2(n45955), .ZN(n43500) );
  XOR2HSV0 U47643 ( .A1(n43501), .A2(n43500), .Z(n43502) );
  XOR2HSV0 U47644 ( .A1(n43503), .A2(n43502), .Z(n43511) );
  NAND2HSV0 U47645 ( .A1(n46456), .A2(n43775), .ZN(n43505) );
  NAND2HSV0 U47646 ( .A1(n56349), .A2(n49439), .ZN(n43504) );
  XOR2HSV0 U47647 ( .A1(n43505), .A2(n43504), .Z(n43509) );
  CLKNAND2HSV0 U47648 ( .A1(n55988), .A2(n56644), .ZN(n43507) );
  NAND2HSV0 U47649 ( .A1(n56182), .A2(\pe3/bq[18] ), .ZN(n43506) );
  XOR2HSV0 U47650 ( .A1(n43507), .A2(n43506), .Z(n43508) );
  XOR2HSV0 U47651 ( .A1(n43509), .A2(n43508), .Z(n43510) );
  XOR2HSV0 U47652 ( .A1(n43511), .A2(n43510), .Z(n43513) );
  CLKNAND2HSV1 U47653 ( .A1(n37131), .A2(n56855), .ZN(n43512) );
  XNOR2HSV1 U47654 ( .A1(n43513), .A2(n43512), .ZN(n43514) );
  XNOR2HSV1 U47655 ( .A1(n43515), .A2(n43514), .ZN(n43559) );
  NAND2HSV0 U47656 ( .A1(n43516), .A2(n59644), .ZN(n43556) );
  CLKNHSV0 U47657 ( .I(n46613), .ZN(n46612) );
  CLKNAND2HSV0 U47658 ( .A1(n46612), .A2(\pe3/pvq [26]), .ZN(n43517) );
  XNOR2HSV1 U47659 ( .A1(n43517), .A2(\pe3/phq [26]), .ZN(n43518) );
  NAND2HSV0 U47660 ( .A1(\pe3/aot [8]), .A2(n48538), .ZN(n48537) );
  XNOR2HSV1 U47661 ( .A1(n43518), .A2(n48537), .ZN(n43536) );
  NAND2HSV0 U47662 ( .A1(n55750), .A2(\pe3/bq[11] ), .ZN(n43520) );
  CLKNAND2HSV1 U47663 ( .A1(n56204), .A2(\pe3/bq[19] ), .ZN(n43519) );
  XOR2HSV0 U47664 ( .A1(n43520), .A2(n43519), .Z(n43524) );
  NAND2HSV0 U47665 ( .A1(n46463), .A2(n56627), .ZN(n43522) );
  CLKNHSV0 U47666 ( .I(n55755), .ZN(n55616) );
  NAND2HSV0 U47667 ( .A1(\pe3/aot [22]), .A2(n55616), .ZN(n43521) );
  XOR2HSV0 U47668 ( .A1(n43522), .A2(n43521), .Z(n43523) );
  XOR2HSV0 U47669 ( .A1(n43524), .A2(n43523), .Z(n43535) );
  CLKNAND2HSV0 U47670 ( .A1(n48496), .A2(n56785), .ZN(n46480) );
  NAND2HSV0 U47671 ( .A1(n56464), .A2(n42971), .ZN(n46367) );
  XOR2HSV0 U47672 ( .A1(n46480), .A2(n46367), .Z(n43534) );
  NAND2HSV0 U47673 ( .A1(n45676), .A2(n43780), .ZN(n43526) );
  CLKNHSV0 U47674 ( .I(n55714), .ZN(n55858) );
  CLKNAND2HSV1 U47675 ( .A1(n55858), .A2(n48499), .ZN(n43525) );
  XOR2HSV0 U47676 ( .A1(n43526), .A2(n43525), .Z(n43532) );
  CLKNHSV1 U47677 ( .I(n43527), .ZN(n59344) );
  NAND2HSV0 U47678 ( .A1(n59344), .A2(n43772), .ZN(n43530) );
  NAND2HSV0 U47679 ( .A1(n43528), .A2(n45639), .ZN(n43529) );
  XOR2HSV0 U47680 ( .A1(n43530), .A2(n43529), .Z(n43531) );
  XOR2HSV0 U47681 ( .A1(n43532), .A2(n43531), .Z(n43533) );
  XOR4HSV1 U47682 ( .A1(n43536), .A2(n43535), .A3(n43534), .A4(n43533), .Z(
        n43554) );
  NAND2HSV0 U47683 ( .A1(n46332), .A2(n43809), .ZN(n43538) );
  NAND2HSV0 U47684 ( .A1(n45645), .A2(\pe3/bq[23] ), .ZN(n43537) );
  XOR2HSV0 U47685 ( .A1(n43538), .A2(n43537), .Z(n43543) );
  CLKNAND2HSV0 U47686 ( .A1(n59623), .A2(n43539), .ZN(n43541) );
  CLKNAND2HSV0 U47687 ( .A1(n45952), .A2(\pe3/bq[26] ), .ZN(n43540) );
  XOR2HSV0 U47688 ( .A1(n43541), .A2(n43540), .Z(n43542) );
  XOR2HSV0 U47689 ( .A1(n43543), .A2(n43542), .Z(n43552) );
  NAND2HSV0 U47690 ( .A1(\pe3/aot [23]), .A2(n43544), .ZN(n43546) );
  NAND2HSV0 U47691 ( .A1(n56423), .A2(n45663), .ZN(n43545) );
  XOR2HSV0 U47692 ( .A1(n43546), .A2(n43545), .Z(n43550) );
  NAND2HSV0 U47693 ( .A1(n43547), .A2(n56827), .ZN(n45557) );
  NAND2HSV0 U47694 ( .A1(n59960), .A2(n43793), .ZN(n43548) );
  XOR2HSV0 U47695 ( .A1(n45557), .A2(n43548), .Z(n43549) );
  XOR2HSV0 U47696 ( .A1(n43550), .A2(n43549), .Z(n43551) );
  XOR2HSV0 U47697 ( .A1(n43552), .A2(n43551), .Z(n43553) );
  XNOR2HSV1 U47698 ( .A1(n43554), .A2(n43553), .ZN(n43555) );
  XNOR2HSV1 U47699 ( .A1(n43556), .A2(n43555), .ZN(n43558) );
  CLKNAND2HSV0 U47700 ( .A1(n37316), .A2(n56342), .ZN(n43557) );
  XOR3HSV2 U47701 ( .A1(n43559), .A2(n43558), .A3(n43557), .Z(n43560) );
  XOR2HSV0 U47702 ( .A1(n43561), .A2(n43560), .Z(n43562) );
  XOR2HSV0 U47703 ( .A1(n43563), .A2(n43562), .Z(n43565) );
  CLKNAND2HSV1 U47704 ( .A1(n46313), .A2(n56493), .ZN(n43564) );
  XOR2HSV0 U47705 ( .A1(n43565), .A2(n43564), .Z(n43567) );
  NAND2HSV0 U47706 ( .A1(n56127), .A2(n48584), .ZN(n43566) );
  XNOR2HSV1 U47707 ( .A1(n43567), .A2(n43566), .ZN(n43568) );
  XNOR2HSV1 U47708 ( .A1(n43569), .A2(n43568), .ZN(n43570) );
  XNOR2HSV1 U47709 ( .A1(n43571), .A2(n43570), .ZN(n43572) );
  XNOR2HSV1 U47710 ( .A1(n43573), .A2(n43572), .ZN(n43576) );
  NOR2HSV2 U47711 ( .A1(n45728), .A2(n49250), .ZN(n43575) );
  CLKNAND2HSV1 U47712 ( .A1(n56136), .A2(n45581), .ZN(n43574) );
  XOR3HSV2 U47713 ( .A1(n43576), .A2(n43575), .A3(n43574), .Z(n43580) );
  NOR2HSV1 U47714 ( .A1(n43577), .A2(n37275), .ZN(n43579) );
  NAND2HSV2 U47715 ( .A1(n45732), .A2(n42770), .ZN(n43578) );
  XOR3HSV2 U47716 ( .A1(n43580), .A2(n43579), .A3(n43578), .Z(n43581) );
  XNOR2HSV1 U47717 ( .A1(n43582), .A2(n43581), .ZN(n43584) );
  CLKNAND2HSV1 U47718 ( .A1(n43850), .A2(\pe3/got [23]), .ZN(n43583) );
  XOR2HSV0 U47719 ( .A1(n43584), .A2(n43583), .Z(n43585) );
  XNOR2HSV1 U47720 ( .A1(n43586), .A2(n43585), .ZN(n43588) );
  CLKNAND2HSV0 U47721 ( .A1(n45582), .A2(n45947), .ZN(n43587) );
  XNOR2HSV1 U47722 ( .A1(n43588), .A2(n43587), .ZN(n43589) );
  NAND2HSV4 U47723 ( .A1(n43595), .A2(n43594), .ZN(n55705) );
  NAND2HSV4 U47724 ( .A1(n43597), .A2(n43897), .ZN(n43906) );
  NOR2HSV2 U47725 ( .A1(n43598), .A2(n47428), .ZN(n43602) );
  OAI21HSV0 U47726 ( .A1(n43478), .A2(n45625), .B(n45612), .ZN(n43599) );
  INHSV2 U47727 ( .I(n43599), .ZN(n43603) );
  CLKNAND2HSV2 U47728 ( .A1(n43610), .A2(n43602), .ZN(n43606) );
  CLKNAND2HSV3 U47729 ( .A1(n43609), .A2(n43603), .ZN(n43611) );
  AOI31HSV2 U47730 ( .A1(n43611), .A2(n45779), .A3(n43612), .B(n45509), .ZN(
        n43605) );
  NAND2HSV2 U47731 ( .A1(n43606), .A2(n43605), .ZN(n43607) );
  INHSV2 U47732 ( .I(n43607), .ZN(n55612) );
  INHSV2 U47733 ( .I(n55612), .ZN(n56063) );
  INHSV2 U47734 ( .I(n45503), .ZN(n44667) );
  NOR2HSV0 U47735 ( .A1(n45509), .A2(n44664), .ZN(n45511) );
  NOR2HSV2 U47736 ( .A1(n45511), .A2(n43613), .ZN(n43616) );
  NOR2HSV0 U47737 ( .A1(n43750), .A2(n43866), .ZN(n43618) );
  INHSV1 U47738 ( .I(n43618), .ZN(n43615) );
  CLKNHSV0 U47739 ( .I(n43616), .ZN(n43617) );
  NOR2HSV0 U47740 ( .A1(n43617), .A2(n43867), .ZN(n43620) );
  NOR2HSV2 U47741 ( .A1(n43618), .A2(n59964), .ZN(n43619) );
  NAND2HSV2 U47742 ( .A1(n46312), .A2(\pe3/got [26]), .ZN(n43721) );
  CLKNAND2HSV1 U47743 ( .A1(n45583), .A2(n45634), .ZN(n43719) );
  BUFHSV2 U47744 ( .I(n43621), .Z(n53228) );
  CLKNAND2HSV1 U47745 ( .A1(n53228), .A2(n48483), .ZN(n43715) );
  INHSV2 U47746 ( .I(n47430), .ZN(n45636) );
  CLKNAND2HSV1 U47747 ( .A1(n45636), .A2(n55821), .ZN(n43711) );
  INHSV2 U47748 ( .I(n45576), .ZN(n56065) );
  NAND2HSV0 U47749 ( .A1(n43755), .A2(n56065), .ZN(n43702) );
  BUFHSV2 U47750 ( .I(n43622), .Z(n49255) );
  CLKNAND2HSV1 U47751 ( .A1(n49255), .A2(n45518), .ZN(n43700) );
  BUFHSV2 U47752 ( .I(n37151), .Z(n55706) );
  NAND2HSV0 U47753 ( .A1(n55706), .A2(n56493), .ZN(n43698) );
  NAND2HSV0 U47754 ( .A1(n45949), .A2(n56247), .ZN(n43692) );
  CLKNAND2HSV1 U47755 ( .A1(n46314), .A2(n59644), .ZN(n43690) );
  NAND2HSV0 U47756 ( .A1(n45950), .A2(n56771), .ZN(n43641) );
  NAND2HSV0 U47757 ( .A1(n55873), .A2(n46614), .ZN(n43625) );
  CLKNHSV0 U47758 ( .I(n56859), .ZN(n56734) );
  NAND2HSV0 U47759 ( .A1(n56734), .A2(n37051), .ZN(n43624) );
  XOR2HSV0 U47760 ( .A1(n43625), .A2(n43624), .Z(n43629) );
  NAND2HSV0 U47761 ( .A1(n59623), .A2(\pe3/bq[26] ), .ZN(n43627) );
  NAND2HSV0 U47762 ( .A1(n56188), .A2(\pe3/bq[23] ), .ZN(n43626) );
  XOR2HSV0 U47763 ( .A1(n43627), .A2(n43626), .Z(n43628) );
  XOR2HSV0 U47764 ( .A1(n43629), .A2(n43628), .Z(n43637) );
  NAND2HSV0 U47765 ( .A1(n56423), .A2(n55867), .ZN(n43631) );
  NAND2HSV0 U47766 ( .A1(n45676), .A2(n55976), .ZN(n43630) );
  XOR2HSV0 U47767 ( .A1(n43631), .A2(n43630), .Z(n43635) );
  NAND2HSV0 U47768 ( .A1(n45973), .A2(n48538), .ZN(n43633) );
  NAND2HSV0 U47769 ( .A1(n45645), .A2(n56218), .ZN(n43632) );
  XOR2HSV0 U47770 ( .A1(n43633), .A2(n43632), .Z(n43634) );
  XOR2HSV0 U47771 ( .A1(n43635), .A2(n43634), .Z(n43636) );
  XOR2HSV0 U47772 ( .A1(n43637), .A2(n43636), .Z(n43639) );
  NAND2HSV0 U47773 ( .A1(n59648), .A2(n56560), .ZN(n43638) );
  XNOR2HSV1 U47774 ( .A1(n43639), .A2(n43638), .ZN(n43640) );
  XNOR2HSV1 U47775 ( .A1(n43641), .A2(n43640), .ZN(n43688) );
  NAND2HSV0 U47776 ( .A1(n59671), .A2(n56855), .ZN(n43685) );
  NAND2HSV0 U47777 ( .A1(\pe3/aot [20]), .A2(n55616), .ZN(n43643) );
  NAND2HSV0 U47778 ( .A1(\pe3/aot [18]), .A2(\pe3/bq[19] ), .ZN(n43642) );
  XOR2HSV0 U47779 ( .A1(n43643), .A2(n43642), .Z(n43647) );
  NAND2HSV0 U47780 ( .A1(n42743), .A2(\pe3/bq[11] ), .ZN(n43645) );
  NAND2HSV0 U47781 ( .A1(n45952), .A2(n55872), .ZN(n43644) );
  XOR2HSV0 U47782 ( .A1(n43645), .A2(n43644), .Z(n43646) );
  XOR2HSV0 U47783 ( .A1(n43647), .A2(n43646), .Z(n43656) );
  NAND2HSV0 U47784 ( .A1(n46332), .A2(n45534), .ZN(n43649) );
  NAND2HSV0 U47785 ( .A1(n55858), .A2(n43775), .ZN(n43648) );
  XOR2HSV0 U47786 ( .A1(n43649), .A2(n43648), .Z(n43654) );
  NAND2HSV0 U47787 ( .A1(n43650), .A2(n45639), .ZN(n43652) );
  CLKNHSV0 U47788 ( .I(n46138), .ZN(n45696) );
  CLKNAND2HSV0 U47789 ( .A1(n42940), .A2(n45696), .ZN(n43651) );
  XOR2HSV0 U47790 ( .A1(n43652), .A2(n43651), .Z(n43653) );
  XOR2HSV0 U47791 ( .A1(n43654), .A2(n43653), .Z(n43655) );
  XOR2HSV0 U47792 ( .A1(n43656), .A2(n43655), .Z(n43668) );
  NAND2HSV0 U47793 ( .A1(n48500), .A2(\pe3/bq[8] ), .ZN(n43658) );
  NAND2HSV0 U47794 ( .A1(n45640), .A2(n53232), .ZN(n43657) );
  XOR2HSV0 U47795 ( .A1(n43658), .A2(n43657), .Z(n43662) );
  NAND2HSV0 U47796 ( .A1(n36809), .A2(\pe3/bq[10] ), .ZN(n43660) );
  NAND2HSV0 U47797 ( .A1(n42818), .A2(n48499), .ZN(n43659) );
  XOR2HSV0 U47798 ( .A1(n43660), .A2(n43659), .Z(n43661) );
  XOR2HSV0 U47799 ( .A1(n43662), .A2(n43661), .Z(n43666) );
  NAND2HSV0 U47800 ( .A1(n46127), .A2(\pe3/pvq [28]), .ZN(n43663) );
  XNOR2HSV1 U47801 ( .A1(n43663), .A2(\pe3/phq [28]), .ZN(n43664) );
  NAND2HSV0 U47802 ( .A1(n59627), .A2(n45663), .ZN(n48521) );
  XNOR2HSV1 U47803 ( .A1(n43664), .A2(n48521), .ZN(n43665) );
  XNOR2HSV1 U47804 ( .A1(n43666), .A2(n43665), .ZN(n43667) );
  XNOR2HSV1 U47805 ( .A1(n43668), .A2(n43667), .ZN(n43683) );
  NAND2HSV0 U47806 ( .A1(\pe3/aot [8]), .A2(n43793), .ZN(n43670) );
  BUFHSV2 U47807 ( .I(n56651), .Z(n45951) );
  NAND2HSV0 U47808 ( .A1(n45951), .A2(n43772), .ZN(n43669) );
  XOR2HSV0 U47809 ( .A1(n43670), .A2(n43669), .Z(n43674) );
  NAND2HSV0 U47810 ( .A1(n59344), .A2(n42971), .ZN(n43672) );
  CLKNHSV0 U47811 ( .I(n56914), .ZN(n56189) );
  NAND2HSV0 U47812 ( .A1(n45572), .A2(n56189), .ZN(n43671) );
  XOR2HSV0 U47813 ( .A1(n43672), .A2(n43671), .Z(n43673) );
  XOR2HSV0 U47814 ( .A1(n43674), .A2(n43673), .Z(n43681) );
  NOR2HSV0 U47815 ( .A1(n45567), .A2(n46615), .ZN(n43676) );
  NAND2HSV0 U47816 ( .A1(n59960), .A2(n43780), .ZN(n43675) );
  XOR2HSV0 U47817 ( .A1(n43676), .A2(n43675), .Z(n43679) );
  INHSV2 U47818 ( .I(n49258), .ZN(n56835) );
  NAND2HSV0 U47819 ( .A1(n43265), .A2(n56835), .ZN(n48515) );
  NAND2HSV0 U47820 ( .A1(n56464), .A2(\pe3/bq[18] ), .ZN(n43677) );
  XOR2HSV0 U47821 ( .A1(n48515), .A2(n43677), .Z(n43678) );
  XOR2HSV0 U47822 ( .A1(n43679), .A2(n43678), .Z(n43680) );
  XOR2HSV0 U47823 ( .A1(n43681), .A2(n43680), .Z(n43682) );
  XNOR2HSV1 U47824 ( .A1(n43683), .A2(n43682), .ZN(n43684) );
  XNOR2HSV1 U47825 ( .A1(n43685), .A2(n43684), .ZN(n43687) );
  CLKNAND2HSV1 U47826 ( .A1(n55826), .A2(n59645), .ZN(n43686) );
  XOR3HSV2 U47827 ( .A1(n43688), .A2(n43687), .A3(n43686), .Z(n43689) );
  XOR2HSV0 U47828 ( .A1(n43690), .A2(n43689), .Z(n43691) );
  XOR2HSV0 U47829 ( .A1(n43692), .A2(n43691), .Z(n43694) );
  NAND2HSV0 U47830 ( .A1(n46313), .A2(n43756), .ZN(n43693) );
  XOR2HSV0 U47831 ( .A1(n43694), .A2(n43693), .Z(n43696) );
  NAND2HSV0 U47832 ( .A1(n56127), .A2(n56421), .ZN(n43695) );
  XNOR2HSV1 U47833 ( .A1(n43696), .A2(n43695), .ZN(n43697) );
  XNOR2HSV1 U47834 ( .A1(n43698), .A2(n43697), .ZN(n43699) );
  XNOR2HSV1 U47835 ( .A1(n43700), .A2(n43699), .ZN(n43701) );
  XNOR2HSV1 U47836 ( .A1(n43702), .A2(n43701), .ZN(n43705) );
  NOR2HSV1 U47837 ( .A1(n43840), .A2(n44693), .ZN(n43704) );
  BUFHSV2 U47838 ( .I(n49251), .Z(n46533) );
  NOR2HSV0 U47839 ( .A1(n46519), .A2(n46533), .ZN(n43703) );
  XOR3HSV2 U47840 ( .A1(n43705), .A2(n43704), .A3(n43703), .Z(n43709) );
  BUFHSV2 U47841 ( .I(n43706), .Z(n59362) );
  INHSV2 U47842 ( .I(n59362), .ZN(n43844) );
  NOR2HSV2 U47843 ( .A1(n43844), .A2(n49250), .ZN(n43708) );
  NAND2HSV0 U47844 ( .A1(n45732), .A2(n45581), .ZN(n43707) );
  XOR3HSV2 U47845 ( .A1(n43709), .A2(n43708), .A3(n43707), .Z(n43710) );
  NAND2HSV0 U47846 ( .A1(n43850), .A2(n55945), .ZN(n43712) );
  XOR2HSV0 U47847 ( .A1(n43713), .A2(n43712), .Z(n43714) );
  XNOR2HSV1 U47848 ( .A1(n43715), .A2(n43714), .ZN(n43717) );
  NAND2HSV0 U47849 ( .A1(n45582), .A2(n59617), .ZN(n43716) );
  XNOR2HSV1 U47850 ( .A1(n43717), .A2(n43716), .ZN(n43718) );
  XNOR2HSV1 U47851 ( .A1(n43719), .A2(n43718), .ZN(n43720) );
  XNOR2HSV1 U47852 ( .A1(n43721), .A2(n43720), .ZN(n43724) );
  CLKNHSV1 U47853 ( .I(n43724), .ZN(n43722) );
  AOI21HSV2 U47854 ( .A1(n43234), .A2(n49253), .B(n43722), .ZN(n43723) );
  CLKNAND2HSV1 U47855 ( .A1(n43725), .A2(n25761), .ZN(n43737) );
  AND2HSV2 U47856 ( .A1(n43750), .A2(n55940), .Z(n43726) );
  NAND2HSV2 U47857 ( .A1(n43726), .A2(n43614), .ZN(n43733) );
  NOR2HSV1 U47858 ( .A1(pov3[24]), .A2(n43733), .ZN(n43727) );
  INHSV2 U47859 ( .I(n43727), .ZN(n43731) );
  NAND4HSV4 U47860 ( .A1(n43731), .A2(n43729), .A3(n43730), .A4(n29657), .ZN(
        n43736) );
  INHSV2 U47861 ( .I(n43733), .ZN(n43734) );
  NAND3HSV4 U47862 ( .A1(n43737), .A2(n43736), .A3(n43735), .ZN(n43747) );
  INHSV2 U47863 ( .I(n45596), .ZN(n45598) );
  OAI21HSV2 U47864 ( .A1(n45599), .A2(n45598), .B(n43745), .ZN(n43746) );
  XNOR2HSV4 U47865 ( .A1(n43747), .A2(n43746), .ZN(n43749) );
  CLKNAND2HSV3 U47866 ( .A1(n43749), .A2(n43748), .ZN(n45763) );
  NOR2HSV0 U47867 ( .A1(n44679), .A2(n43132), .ZN(n45760) );
  INAND2HSV2 U47868 ( .A1(n46092), .B1(n45760), .ZN(n43915) );
  OR2HSV1 U47869 ( .A1(n45511), .A2(n43752), .Z(n43862) );
  INHSV2 U47870 ( .I(n43862), .ZN(n43753) );
  NAND2HSV2 U47871 ( .A1(n46312), .A2(n37107), .ZN(n43861) );
  INHSV2 U47872 ( .I(n43494), .ZN(n56685) );
  NAND2HSV2 U47873 ( .A1(n56685), .A2(\pe3/got [26]), .ZN(n43859) );
  CLKNAND2HSV0 U47874 ( .A1(n43754), .A2(n55701), .ZN(n43854) );
  CLKNAND2HSV1 U47875 ( .A1(n45636), .A2(n48483), .ZN(n43849) );
  NAND2HSV0 U47876 ( .A1(n43755), .A2(n56335), .ZN(n43839) );
  NAND2HSV0 U47877 ( .A1(n59625), .A2(n49252), .ZN(n43837) );
  CLKNAND2HSV1 U47878 ( .A1(n55706), .A2(n45518), .ZN(n43835) );
  NAND2HSV0 U47879 ( .A1(n45949), .A2(n43756), .ZN(n43828) );
  NAND2HSV0 U47880 ( .A1(n46314), .A2(n59967), .ZN(n43826) );
  NAND2HSV0 U47881 ( .A1(n59608), .A2(\pe3/bq[7] ), .ZN(n43759) );
  NAND2HSV0 U47882 ( .A1(n43650), .A2(n56454), .ZN(n43758) );
  XOR2HSV0 U47883 ( .A1(n43759), .A2(n43758), .Z(n43763) );
  NAND2HSV0 U47884 ( .A1(\pe3/aot [14]), .A2(n55872), .ZN(n43761) );
  BUFHSV2 U47885 ( .I(\pe3/aot [6]), .Z(n56795) );
  NAND2HSV0 U47886 ( .A1(n56795), .A2(n46614), .ZN(n43760) );
  XOR2HSV0 U47887 ( .A1(n43761), .A2(n43760), .Z(n43762) );
  XOR2HSV0 U47888 ( .A1(n43763), .A2(n43762), .Z(n43771) );
  NAND2HSV0 U47889 ( .A1(n55750), .A2(n56627), .ZN(n43765) );
  NAND2HSV0 U47890 ( .A1(n46456), .A2(\pe3/bq[11] ), .ZN(n43764) );
  XOR2HSV0 U47891 ( .A1(n43765), .A2(n43764), .Z(n43769) );
  NAND2HSV0 U47892 ( .A1(n46332), .A2(n48499), .ZN(n43767) );
  NAND2HSV0 U47893 ( .A1(n55858), .A2(n45534), .ZN(n43766) );
  XOR2HSV0 U47894 ( .A1(n43767), .A2(n43766), .Z(n43768) );
  XOR2HSV0 U47895 ( .A1(n43769), .A2(n43768), .Z(n43770) );
  XOR2HSV0 U47896 ( .A1(n43771), .A2(n43770), .Z(n43790) );
  NAND2HSV0 U47897 ( .A1(\pe3/aot [8]), .A2(n45663), .ZN(n43774) );
  NAND2HSV0 U47898 ( .A1(n45645), .A2(n43772), .ZN(n43773) );
  XOR2HSV0 U47899 ( .A1(n43774), .A2(n43773), .Z(n43779) );
  NAND2HSV0 U47900 ( .A1(n59627), .A2(n48538), .ZN(n43777) );
  NAND2HSV0 U47901 ( .A1(n55988), .A2(n43775), .ZN(n43776) );
  XOR2HSV0 U47902 ( .A1(n43777), .A2(n43776), .Z(n43778) );
  XOR2HSV0 U47903 ( .A1(n43779), .A2(n43778), .Z(n43788) );
  NOR2HSV0 U47904 ( .A1(n45567), .A2(n46138), .ZN(n43782) );
  NAND2HSV0 U47905 ( .A1(n59623), .A2(n43780), .ZN(n43781) );
  XOR2HSV0 U47906 ( .A1(n43782), .A2(n43781), .Z(n43786) );
  NAND2HSV0 U47907 ( .A1(n56204), .A2(\pe3/bq[18] ), .ZN(n43784) );
  NAND2HSV0 U47908 ( .A1(\pe3/aot [15]), .A2(\pe3/bq[23] ), .ZN(n43783) );
  XOR2HSV0 U47909 ( .A1(n43784), .A2(n43783), .Z(n43785) );
  XOR2HSV0 U47910 ( .A1(n43786), .A2(n43785), .Z(n43787) );
  XOR2HSV0 U47911 ( .A1(n43788), .A2(n43787), .Z(n43789) );
  XOR2HSV0 U47912 ( .A1(n43790), .A2(n43789), .Z(n43792) );
  NAND2HSV0 U47913 ( .A1(n45950), .A2(n56855), .ZN(n43791) );
  XOR2HSV0 U47914 ( .A1(n43792), .A2(n43791), .Z(n43824) );
  BUFHSV2 U47915 ( .I(n59671), .Z(n48511) );
  CLKNAND2HSV1 U47916 ( .A1(n48511), .A2(n59645), .ZN(n43821) );
  NAND2HSV0 U47917 ( .A1(n59960), .A2(n43539), .ZN(n43795) );
  NAND2HSV0 U47918 ( .A1(n56423), .A2(n43793), .ZN(n43794) );
  XOR2HSV0 U47919 ( .A1(n43795), .A2(n43794), .Z(n43799) );
  NAND2HSV0 U47920 ( .A1(n56349), .A2(n42971), .ZN(n43797) );
  NAND2HSV0 U47921 ( .A1(n56464), .A2(\pe3/bq[19] ), .ZN(n43796) );
  XOR2HSV0 U47922 ( .A1(n43797), .A2(n43796), .Z(n43798) );
  XOR2HSV0 U47923 ( .A1(n43799), .A2(n43798), .Z(n43819) );
  NAND2HSV0 U47924 ( .A1(n45676), .A2(\pe3/bq[26] ), .ZN(n43801) );
  NAND2HSV0 U47925 ( .A1(n45952), .A2(n55976), .ZN(n43800) );
  XOR2HSV0 U47926 ( .A1(n43801), .A2(n43800), .Z(n43804) );
  NAND2HSV0 U47927 ( .A1(n48020), .A2(\pe3/pvq [27]), .ZN(n43802) );
  XNOR2HSV1 U47928 ( .A1(n43802), .A2(\pe3/phq [27]), .ZN(n43803) );
  XNOR2HSV1 U47929 ( .A1(n43804), .A2(n43803), .ZN(n43808) );
  NAND2HSV0 U47930 ( .A1(n48500), .A2(n56785), .ZN(n43806) );
  NAND2HSV0 U47931 ( .A1(n59344), .A2(n56218), .ZN(n43805) );
  XOR2HSV0 U47932 ( .A1(n43806), .A2(n43805), .Z(n43807) );
  XNOR2HSV1 U47933 ( .A1(n43808), .A2(n43807), .ZN(n43818) );
  NOR2HSV0 U47934 ( .A1(n42539), .A2(n55755), .ZN(n43811) );
  NAND2HSV0 U47935 ( .A1(n42818), .A2(n43809), .ZN(n43810) );
  XOR2HSV0 U47936 ( .A1(n43811), .A2(n43810), .Z(n43815) );
  NAND2HSV0 U47937 ( .A1(n45962), .A2(n56835), .ZN(n43813) );
  NAND2HSV0 U47938 ( .A1(\pe3/got [6]), .A2(n37051), .ZN(n43812) );
  XOR2HSV0 U47939 ( .A1(n43813), .A2(n43812), .Z(n43814) );
  XOR2HSV0 U47940 ( .A1(n43815), .A2(n43814), .Z(n43817) );
  NAND2HSV0 U47941 ( .A1(n59648), .A2(n56771), .ZN(n43816) );
  XOR4HSV1 U47942 ( .A1(n43819), .A2(n43818), .A3(n43817), .A4(n43816), .Z(
        n43820) );
  XNOR2HSV1 U47943 ( .A1(n43821), .A2(n43820), .ZN(n43823) );
  CLKNAND2HSV1 U47944 ( .A1(n52727), .A2(n59644), .ZN(n43822) );
  XOR3HSV2 U47945 ( .A1(n43824), .A2(n43823), .A3(n43822), .Z(n43825) );
  XOR2HSV0 U47946 ( .A1(n43826), .A2(n43825), .Z(n43827) );
  XOR2HSV0 U47947 ( .A1(n43828), .A2(n43827), .Z(n43831) );
  NAND2HSV0 U47948 ( .A1(n46313), .A2(n43829), .ZN(n43830) );
  XOR2HSV0 U47949 ( .A1(n43831), .A2(n43830), .Z(n43833) );
  NAND2HSV0 U47950 ( .A1(n55895), .A2(n56493), .ZN(n43832) );
  XNOR2HSV1 U47951 ( .A1(n43833), .A2(n43832), .ZN(n43834) );
  XNOR2HSV1 U47952 ( .A1(n43835), .A2(n43834), .ZN(n43836) );
  XNOR2HSV1 U47953 ( .A1(n43837), .A2(n43836), .ZN(n43838) );
  XNOR2HSV1 U47954 ( .A1(n43839), .A2(n43838), .ZN(n43843) );
  NOR2HSV2 U47955 ( .A1(n43840), .A2(n46533), .ZN(n43842) );
  NAND2HSV0 U47956 ( .A1(n46043), .A2(n59965), .ZN(n43841) );
  XOR3HSV2 U47957 ( .A1(n43843), .A2(n43842), .A3(n43841), .Z(n43847) );
  NOR2HSV2 U47958 ( .A1(n43844), .A2(n45635), .ZN(n43846) );
  NAND2HSV0 U47959 ( .A1(n45732), .A2(n55945), .ZN(n43845) );
  XOR3HSV2 U47960 ( .A1(n43847), .A2(n43846), .A3(n43845), .Z(n43848) );
  XNOR2HSV1 U47961 ( .A1(n43849), .A2(n43848), .ZN(n43852) );
  NAND2HSV0 U47962 ( .A1(n43850), .A2(n42770), .ZN(n43851) );
  XOR2HSV0 U47963 ( .A1(n43852), .A2(n43851), .Z(n43853) );
  XNOR2HSV1 U47964 ( .A1(n43854), .A2(n43853), .ZN(n43857) );
  CLKNAND2HSV1 U47965 ( .A1(n56662), .A2(n43855), .ZN(n43856) );
  XNOR2HSV1 U47966 ( .A1(n43857), .A2(n43856), .ZN(n43858) );
  XNOR2HSV1 U47967 ( .A1(n43859), .A2(n43858), .ZN(n43860) );
  NOR2HSV2 U47968 ( .A1(n43863), .A2(n43862), .ZN(n43864) );
  CLKBUFHSV4 U47969 ( .I(n43869), .Z(n48486) );
  NAND2HSV2 U47970 ( .A1(n48486), .A2(n37041), .ZN(n43875) );
  CLKNHSV1 U47971 ( .I(n43875), .ZN(n43865) );
  NOR2HSV2 U47972 ( .A1(n43868), .A2(n43867), .ZN(n43877) );
  CLKNAND2HSV0 U47973 ( .A1(n43870), .A2(n59575), .ZN(n43874) );
  OR2HSV1 U47974 ( .A1(n43871), .A2(n43371), .Z(n43872) );
  OAI21HSV2 U47975 ( .A1(n43874), .A2(n43873), .B(n43872), .ZN(n43876) );
  CLKNAND2HSV2 U47976 ( .A1(n43887), .A2(n43884), .ZN(n43883) );
  OAI21HSV2 U47977 ( .A1(n59515), .A2(n45598), .B(n43881), .ZN(n43882) );
  NAND3HSV4 U47978 ( .A1(n43888), .A2(n44328), .A3(n43887), .ZN(n44675) );
  NAND2HSV4 U47979 ( .A1(n44675), .A2(n44676), .ZN(n44665) );
  INHSV3 U47980 ( .I(n44665), .ZN(n48895) );
  INHSV2 U47981 ( .I(n48895), .ZN(n43910) );
  BUFHSV2 U47982 ( .I(n43906), .Z(n51011) );
  INHSV1 U47983 ( .I(n43906), .ZN(n43892) );
  NOR2HSV2 U47984 ( .A1(n43892), .A2(n43484), .ZN(n43893) );
  OAI21HSV2 U47985 ( .A1(n56175), .A2(n43899), .B(n43897), .ZN(n43901) );
  OAI21HSV2 U47986 ( .A1(n43899), .A2(n43898), .B(n44664), .ZN(n43900) );
  NOR2HSV2 U47987 ( .A1(n43901), .A2(n43900), .ZN(n43902) );
  OA21HSV2 U47988 ( .A1(\pe3/ti_7t [26]), .A2(n45625), .B(n45624), .Z(n45504)
         );
  INHSV2 U47989 ( .I(n45504), .ZN(n43904) );
  NOR2HSV4 U47990 ( .A1(n26396), .A2(n43904), .ZN(n44680) );
  CLKNAND2HSV1 U47991 ( .A1(n43906), .A2(n43905), .ZN(n43907) );
  INHSV2 U47992 ( .I(n43907), .ZN(n43908) );
  INHSV6 U47993 ( .I(n43913), .ZN(n44678) );
  NAND2HSV0 U47994 ( .A1(n47428), .A2(\pe3/ti_7t [28]), .ZN(n46085) );
  CLKNHSV2 U47995 ( .I(n46085), .ZN(n45756) );
  CLKNAND2HSV2 U47996 ( .A1(n43917), .A2(n59979), .ZN(n43922) );
  NOR2HSV4 U47997 ( .A1(n44150), .A2(n44831), .ZN(n43918) );
  AOI22HSV4 U47998 ( .A1(n43920), .A2(n43919), .B1(n39113), .B2(n43918), .ZN(
        n43921) );
  CLKNAND2HSV0 U47999 ( .A1(n38324), .A2(n51801), .ZN(n44018) );
  CLKNAND2HSV1 U48000 ( .A1(n59773), .A2(n43924), .ZN(n44016) );
  CLKNAND2HSV0 U48001 ( .A1(n45288), .A2(n43925), .ZN(n44013) );
  NAND2HSV2 U48002 ( .A1(n44713), .A2(\pe2/got [21]), .ZN(n44011) );
  NAND2HSV0 U48003 ( .A1(n51889), .A2(n52419), .ZN(n44009) );
  CLKNAND2HSV0 U48004 ( .A1(n50929), .A2(n44712), .ZN(n44006) );
  CLKNAND2HSV1 U48005 ( .A1(n44185), .A2(n43926), .ZN(n43998) );
  NAND2HSV0 U48006 ( .A1(n45150), .A2(n43927), .ZN(n43996) );
  NAND2HSV0 U48007 ( .A1(n43928), .A2(n52172), .ZN(n43992) );
  NAND2HSV0 U48008 ( .A1(n44046), .A2(n44044), .ZN(n43930) );
  NOR2HSV0 U48009 ( .A1(n52420), .A2(n44045), .ZN(n43929) );
  XNOR2HSV1 U48010 ( .A1(n43930), .A2(n43929), .ZN(n43990) );
  XOR2HSV0 U48011 ( .A1(n43932), .A2(n43931), .Z(n43937) );
  INHSV2 U48012 ( .I(n43933), .ZN(n59977) );
  CLKNAND2HSV1 U48013 ( .A1(n59977), .A2(n39020), .ZN(n43935) );
  NAND2HSV0 U48014 ( .A1(n39019), .A2(\pe2/bq[29] ), .ZN(n43934) );
  XOR2HSV0 U48015 ( .A1(n43935), .A2(n43934), .Z(n43936) );
  XOR2HSV0 U48016 ( .A1(n43937), .A2(n43936), .Z(n43953) );
  NOR2HSV0 U48017 ( .A1(n44871), .A2(n48064), .ZN(n43939) );
  NAND2HSV0 U48018 ( .A1(n53019), .A2(n36480), .ZN(n43938) );
  XOR2HSV0 U48019 ( .A1(n43939), .A2(n43938), .Z(n43943) );
  CLKNAND2HSV0 U48020 ( .A1(n45034), .A2(n39032), .ZN(n43941) );
  NAND2HSV0 U48021 ( .A1(n45024), .A2(\pe2/bq[24] ), .ZN(n43940) );
  XNOR2HSV1 U48022 ( .A1(n43941), .A2(n43940), .ZN(n43942) );
  XNOR2HSV1 U48023 ( .A1(n43943), .A2(n43942), .ZN(n43949) );
  NAND2HSV0 U48024 ( .A1(n48078), .A2(\pe2/pvq [25]), .ZN(n43944) );
  XOR2HSV0 U48025 ( .A1(n43944), .A2(\pe2/phq [25]), .Z(n43947) );
  NOR2HSV0 U48026 ( .A1(n52103), .A2(n51567), .ZN(n52225) );
  CLKNHSV0 U48027 ( .I(n52103), .ZN(n59358) );
  AOI22HSV0 U48028 ( .A1(n44750), .A2(n51825), .B1(n38054), .B2(n59358), .ZN(
        n43945) );
  AOI21HSV0 U48029 ( .A1(n44206), .A2(n52225), .B(n43945), .ZN(n43946) );
  XOR2HSV0 U48030 ( .A1(n43947), .A2(n43946), .Z(n43948) );
  XNOR2HSV1 U48031 ( .A1(n43949), .A2(n43948), .ZN(n43952) );
  BUFHSV2 U48032 ( .I(n44835), .Z(n51800) );
  CLKNHSV0 U48033 ( .I(n51800), .ZN(n44714) );
  NAND2HSV0 U48034 ( .A1(n43950), .A2(n44714), .ZN(n43951) );
  XOR3HSV2 U48035 ( .A1(n43953), .A2(n43952), .A3(n43951), .Z(n43988) );
  NAND2HSV0 U48036 ( .A1(n52294), .A2(\pe2/bq[21] ), .ZN(n43955) );
  BUFHSV2 U48037 ( .I(\pe2/bq[12] ), .Z(n51733) );
  NAND2HSV0 U48038 ( .A1(n44081), .A2(n51733), .ZN(n43954) );
  XOR2HSV0 U48039 ( .A1(n43955), .A2(n43954), .Z(n43960) );
  NAND2HSV0 U48040 ( .A1(n38048), .A2(n43956), .ZN(n43958) );
  NAND2HSV0 U48041 ( .A1(n59972), .A2(n52984), .ZN(n43957) );
  XOR2HSV0 U48042 ( .A1(n43958), .A2(n43957), .Z(n43959) );
  XOR2HSV0 U48043 ( .A1(n43960), .A2(n43959), .Z(n43969) );
  NAND2HSV0 U48044 ( .A1(n39029), .A2(n43961), .ZN(n43963) );
  CLKNAND2HSV0 U48045 ( .A1(n39052), .A2(n44197), .ZN(n43962) );
  XOR2HSV0 U48046 ( .A1(n43963), .A2(n43962), .Z(n43967) );
  NAND2HSV0 U48047 ( .A1(n50930), .A2(n44074), .ZN(n43965) );
  INHSV2 U48048 ( .I(n47511), .ZN(n52193) );
  NAND2HSV0 U48049 ( .A1(n59968), .A2(n52193), .ZN(n43964) );
  XOR2HSV0 U48050 ( .A1(n43965), .A2(n43964), .Z(n43966) );
  XOR2HSV0 U48051 ( .A1(n43967), .A2(n43966), .Z(n43968) );
  XOR2HSV0 U48052 ( .A1(n43969), .A2(n43968), .Z(n43986) );
  NAND2HSV0 U48053 ( .A1(\pe2/aot [14]), .A2(n38064), .ZN(n43971) );
  NAND2HSV0 U48054 ( .A1(n59588), .A2(n51900), .ZN(n43970) );
  XOR2HSV0 U48055 ( .A1(n43971), .A2(n43970), .Z(n43976) );
  INHSV1 U48056 ( .I(n49628), .ZN(n44231) );
  NAND2HSV0 U48057 ( .A1(n45295), .A2(n44231), .ZN(n43974) );
  INHSV2 U48058 ( .I(n47518), .ZN(n52457) );
  NAND2HSV0 U48059 ( .A1(n52457), .A2(n43972), .ZN(n43973) );
  XOR2HSV0 U48060 ( .A1(n43974), .A2(n43973), .Z(n43975) );
  XOR2HSV0 U48061 ( .A1(n43976), .A2(n43975), .Z(n43984) );
  NOR2HSV0 U48062 ( .A1(n47503), .A2(n44854), .ZN(n43978) );
  NAND2HSV0 U48063 ( .A1(n52289), .A2(n44090), .ZN(n43977) );
  XOR2HSV0 U48064 ( .A1(n43978), .A2(n43977), .Z(n43982) );
  CLKNAND2HSV0 U48065 ( .A1(\pe2/aot [17]), .A2(n52179), .ZN(n43980) );
  INHSV2 U48066 ( .I(\pe2/got [8]), .ZN(n44188) );
  NAND2HSV0 U48067 ( .A1(n59371), .A2(n45303), .ZN(n43979) );
  XOR2HSV0 U48068 ( .A1(n43980), .A2(n43979), .Z(n43981) );
  XOR2HSV0 U48069 ( .A1(n43982), .A2(n43981), .Z(n43983) );
  XOR2HSV0 U48070 ( .A1(n43984), .A2(n43983), .Z(n43985) );
  XOR2HSV0 U48071 ( .A1(n43986), .A2(n43985), .Z(n43987) );
  XNOR2HSV1 U48072 ( .A1(n43988), .A2(n43987), .ZN(n43989) );
  XNOR2HSV1 U48073 ( .A1(n43990), .A2(n43989), .ZN(n43991) );
  XNOR2HSV1 U48074 ( .A1(n43992), .A2(n43991), .ZN(n43994) );
  CLKNHSV0 U48075 ( .I(n51607), .ZN(n44186) );
  NAND2HSV0 U48076 ( .A1(n44254), .A2(n44186), .ZN(n43993) );
  XNOR2HSV1 U48077 ( .A1(n43994), .A2(n43993), .ZN(n43995) );
  XNOR2HSV1 U48078 ( .A1(n43996), .A2(n43995), .ZN(n43997) );
  XNOR2HSV1 U48079 ( .A1(n43998), .A2(n43997), .ZN(n44001) );
  BUFHSV2 U48080 ( .I(n45055), .Z(n44261) );
  CLKNAND2HSV1 U48081 ( .A1(n44261), .A2(n51796), .ZN(n44000) );
  XOR2HSV0 U48082 ( .A1(n44001), .A2(n44000), .Z(n44004) );
  INHSV2 U48083 ( .I(n51795), .ZN(n47571) );
  NAND2HSV0 U48084 ( .A1(n44120), .A2(n47571), .ZN(n44003) );
  XNOR2HSV1 U48085 ( .A1(n44004), .A2(n44003), .ZN(n44005) );
  XNOR2HSV1 U48086 ( .A1(n44006), .A2(n44005), .ZN(n44008) );
  BUFHSV2 U48087 ( .I(n51610), .Z(n45063) );
  NAND2HSV2 U48088 ( .A1(n45063), .A2(n52042), .ZN(n44007) );
  XOR3HSV2 U48089 ( .A1(n44009), .A2(n44008), .A3(n44007), .Z(n44010) );
  XNOR2HSV1 U48090 ( .A1(n44011), .A2(n44010), .ZN(n44012) );
  XNOR2HSV1 U48091 ( .A1(n44013), .A2(n44012), .ZN(n44015) );
  CLKNAND2HSV0 U48092 ( .A1(n52251), .A2(n52416), .ZN(n44014) );
  XOR3HSV2 U48093 ( .A1(n44016), .A2(n44015), .A3(n44014), .Z(n44017) );
  XNOR2HSV1 U48094 ( .A1(n44018), .A2(n44017), .ZN(n44019) );
  XNOR2HSV1 U48095 ( .A1(n44020), .A2(n44019), .ZN(n44021) );
  NAND2HSV0 U48096 ( .A1(n44022), .A2(n44145), .ZN(n44023) );
  XNOR2HSV4 U48097 ( .A1(n44024), .A2(n44023), .ZN(n44038) );
  CLKNHSV0 U48098 ( .I(n44032), .ZN(n44026) );
  NAND2HSV0 U48099 ( .A1(n44031), .A2(n38108), .ZN(n44025) );
  OAI21HSV2 U48100 ( .A1(n44026), .A2(n44025), .B(n36277), .ZN(n44029) );
  NOR2HSV2 U48101 ( .A1(n44309), .A2(n44027), .ZN(n44028) );
  AOI21HSV0 U48102 ( .A1(n44031), .A2(n44032), .B(n44030), .ZN(n44033) );
  INAND2HSV2 U48103 ( .A1(n44034), .B1(n44033), .ZN(n44035) );
  CLKNAND2HSV2 U48104 ( .A1(n45083), .A2(n59980), .ZN(n44037) );
  XNOR2HSV4 U48105 ( .A1(n44039), .A2(n44040), .ZN(n44178) );
  NAND2HSV4 U48106 ( .A1(n44178), .A2(n44309), .ZN(n44168) );
  NOR2HSV2 U48107 ( .A1(n36473), .A2(\pe2/ti_7t [25]), .ZN(n44967) );
  NOR2HSV2 U48108 ( .A1(n44967), .A2(n44307), .ZN(n44169) );
  BUFHSV2 U48109 ( .I(n44169), .Z(n44177) );
  NAND3HSV2 U48110 ( .A1(n44303), .A2(n45089), .A3(n44169), .ZN(n45106) );
  NAND2HSV2 U48111 ( .A1(n51687), .A2(n38723), .ZN(n44142) );
  NAND2HSV0 U48112 ( .A1(n44711), .A2(n45795), .ZN(n44138) );
  NAND2HSV0 U48113 ( .A1(n52416), .A2(n52173), .ZN(n44136) );
  CLKNAND2HSV0 U48114 ( .A1(n59773), .A2(n49591), .ZN(n44134) );
  BUFHSV2 U48115 ( .I(n45288), .Z(n59634) );
  CLKNAND2HSV1 U48116 ( .A1(n59634), .A2(n52167), .ZN(n44131) );
  INHSV2 U48117 ( .I(n44327), .ZN(n52042) );
  CLKNAND2HSV0 U48118 ( .A1(n44713), .A2(n52042), .ZN(n44129) );
  NAND2HSV0 U48119 ( .A1(n44712), .A2(n52419), .ZN(n44127) );
  BUFHSV4 U48120 ( .I(n38780), .Z(n52931) );
  CLKNAND2HSV1 U48121 ( .A1(n52931), .A2(n47571), .ZN(n44124) );
  CLKNAND2HSV0 U48122 ( .A1(n44185), .A2(n48084), .ZN(n44117) );
  CLKNAND2HSV1 U48123 ( .A1(n52934), .A2(n44186), .ZN(n44115) );
  NAND2HSV0 U48124 ( .A1(n44715), .A2(n44044), .ZN(n44111) );
  NAND2HSV0 U48125 ( .A1(n44046), .A2(\pe2/got [10]), .ZN(n44048) );
  NOR2HSV0 U48126 ( .A1(n44971), .A2(n51800), .ZN(n44047) );
  XNOR2HSV1 U48127 ( .A1(n44048), .A2(n44047), .ZN(n44109) );
  NOR2HSV0 U48128 ( .A1(n52200), .A2(n44699), .ZN(n53021) );
  NAND2HSV0 U48129 ( .A1(n44976), .A2(n53223), .ZN(n44209) );
  NAND2HSV0 U48130 ( .A1(n52974), .A2(n44231), .ZN(n44050) );
  XOR2HSV0 U48131 ( .A1(n44209), .A2(n44050), .Z(n44051) );
  XOR3HSV2 U48132 ( .A1(n53021), .A2(n44052), .A3(n44051), .Z(n44071) );
  NAND2HSV2 U48133 ( .A1(n38291), .A2(n59371), .ZN(n44070) );
  CLKNAND2HSV0 U48134 ( .A1(n44750), .A2(\pe2/bq[7] ), .ZN(n44055) );
  NAND2HSV0 U48135 ( .A1(n45034), .A2(n38064), .ZN(n44054) );
  XOR2HSV0 U48136 ( .A1(n44055), .A2(n44054), .Z(n44059) );
  NAND2HSV0 U48137 ( .A1(n39029), .A2(n52988), .ZN(n44057) );
  NAND2HSV0 U48138 ( .A1(n39019), .A2(n38565), .ZN(n44056) );
  XOR2HSV0 U48139 ( .A1(n44057), .A2(n44056), .Z(n44058) );
  XOR2HSV0 U48140 ( .A1(n44059), .A2(n44058), .Z(n44068) );
  NOR2HSV0 U48141 ( .A1(n50947), .A2(n52429), .ZN(n44061) );
  NAND2HSV0 U48142 ( .A1(n59972), .A2(n52337), .ZN(n44060) );
  XOR2HSV0 U48143 ( .A1(n44061), .A2(n44060), .Z(n44066) );
  NAND2HSV0 U48144 ( .A1(n44062), .A2(\pe2/bq[21] ), .ZN(n44064) );
  NAND2HSV0 U48145 ( .A1(\pe2/aot [12]), .A2(n52973), .ZN(n44063) );
  XOR2HSV0 U48146 ( .A1(n44064), .A2(n44063), .Z(n44065) );
  XOR2HSV0 U48147 ( .A1(n44066), .A2(n44065), .Z(n44067) );
  XOR2HSV0 U48148 ( .A1(n44068), .A2(n44067), .Z(n44069) );
  XOR3HSV2 U48149 ( .A1(n44071), .A2(n44070), .A3(n44069), .Z(n44107) );
  NAND2HSV0 U48150 ( .A1(n45024), .A2(n52179), .ZN(n44073) );
  NAND2HSV0 U48151 ( .A1(n44745), .A2(n52950), .ZN(n44072) );
  XOR2HSV0 U48152 ( .A1(n44073), .A2(n44072), .Z(n44078) );
  NAND2HSV0 U48153 ( .A1(\pe2/aot [22]), .A2(n44074), .ZN(n44076) );
  NAND2HSV0 U48154 ( .A1(\pe2/aot [19]), .A2(n44197), .ZN(n44075) );
  XOR2HSV0 U48155 ( .A1(n44076), .A2(n44075), .Z(n44077) );
  XOR2HSV0 U48156 ( .A1(n44078), .A2(n44077), .Z(n44087) );
  NAND2HSV0 U48157 ( .A1(\pe2/aot [17]), .A2(n52299), .ZN(n44080) );
  NAND2HSV0 U48158 ( .A1(n59585), .A2(n52984), .ZN(n44079) );
  XOR2HSV0 U48159 ( .A1(n44080), .A2(n44079), .Z(n44085) );
  CLKNAND2HSV0 U48160 ( .A1(\pe2/aot [25]), .A2(\pe2/bq[14] ), .ZN(n44083) );
  NAND2HSV0 U48161 ( .A1(n44081), .A2(n52073), .ZN(n44082) );
  XOR2HSV0 U48162 ( .A1(n44083), .A2(n44082), .Z(n44084) );
  XOR2HSV0 U48163 ( .A1(n44085), .A2(n44084), .Z(n44086) );
  XOR2HSV0 U48164 ( .A1(n44087), .A2(n44086), .Z(n44105) );
  CLKNAND2HSV0 U48165 ( .A1(n52289), .A2(n52481), .ZN(n44089) );
  NAND2HSV0 U48166 ( .A1(n59977), .A2(\pe2/bq[29] ), .ZN(n44088) );
  XOR2HSV0 U48167 ( .A1(n44089), .A2(n44088), .Z(n44094) );
  CLKNAND2HSV1 U48168 ( .A1(n59633), .A2(n53015), .ZN(n44092) );
  NAND2HSV0 U48169 ( .A1(n52485), .A2(n44090), .ZN(n44091) );
  XOR2HSV0 U48170 ( .A1(n44092), .A2(n44091), .Z(n44093) );
  XOR2HSV0 U48171 ( .A1(n44094), .A2(n44093), .Z(n44103) );
  NOR2HSV0 U48172 ( .A1(n47503), .A2(n38687), .ZN(n44097) );
  BUFHSV2 U48173 ( .I(\pe2/bq[12] ), .Z(n52438) );
  CLKNAND2HSV1 U48174 ( .A1(n45295), .A2(n52438), .ZN(n44096) );
  XOR2HSV0 U48175 ( .A1(n44097), .A2(n44096), .Z(n44101) );
  NAND2HSV0 U48176 ( .A1(n36480), .A2(n52457), .ZN(n44099) );
  INHSV2 U48177 ( .I(n50928), .ZN(n52125) );
  NAND2HSV0 U48178 ( .A1(n52125), .A2(n45303), .ZN(n44098) );
  XOR2HSV0 U48179 ( .A1(n44099), .A2(n44098), .Z(n44100) );
  XOR2HSV0 U48180 ( .A1(n44101), .A2(n44100), .Z(n44102) );
  XOR2HSV0 U48181 ( .A1(n44103), .A2(n44102), .Z(n44104) );
  XOR2HSV0 U48182 ( .A1(n44105), .A2(n44104), .Z(n44106) );
  XNOR2HSV1 U48183 ( .A1(n44107), .A2(n44106), .ZN(n44108) );
  XNOR2HSV1 U48184 ( .A1(n44109), .A2(n44108), .ZN(n44110) );
  XNOR2HSV1 U48185 ( .A1(n44111), .A2(n44110), .ZN(n44113) );
  NAND2HSV0 U48186 ( .A1(n44254), .A2(n52172), .ZN(n44112) );
  XNOR2HSV1 U48187 ( .A1(n44113), .A2(n44112), .ZN(n44114) );
  XNOR2HSV1 U48188 ( .A1(n44115), .A2(n44114), .ZN(n44116) );
  XNOR2HSV1 U48189 ( .A1(n44117), .A2(n44116), .ZN(n44119) );
  CLKNAND2HSV0 U48190 ( .A1(n44261), .A2(n51964), .ZN(n44118) );
  XOR2HSV0 U48191 ( .A1(n44119), .A2(n44118), .Z(n44122) );
  NAND2HSV0 U48192 ( .A1(n44120), .A2(\pe2/got [16]), .ZN(n44121) );
  XNOR2HSV1 U48193 ( .A1(n44122), .A2(n44121), .ZN(n44123) );
  XNOR2HSV1 U48194 ( .A1(n44124), .A2(n44123), .ZN(n44126) );
  CLKNAND2HSV1 U48195 ( .A1(n45063), .A2(n52533), .ZN(n44125) );
  XOR3HSV2 U48196 ( .A1(n44127), .A2(n44126), .A3(n44125), .Z(n44128) );
  XNOR2HSV1 U48197 ( .A1(n44129), .A2(n44128), .ZN(n44130) );
  XNOR2HSV1 U48198 ( .A1(n44131), .A2(n44130), .ZN(n44133) );
  NAND2HSV0 U48199 ( .A1(n59505), .A2(n45249), .ZN(n44132) );
  XOR3HSV2 U48200 ( .A1(n44134), .A2(n44133), .A3(n44132), .Z(n44135) );
  XNOR2HSV1 U48201 ( .A1(n44136), .A2(n44135), .ZN(n44137) );
  XNOR2HSV1 U48202 ( .A1(n44138), .A2(n44137), .ZN(n44140) );
  CLKNAND2HSV1 U48203 ( .A1(n52534), .A2(n38778), .ZN(n44139) );
  CLKNHSV0 U48204 ( .I(n60002), .ZN(n44833) );
  NOR2HSV2 U48205 ( .A1(n44833), .A2(n44143), .ZN(n44144) );
  AND2HSV2 U48206 ( .A1(n45083), .A2(n44145), .Z(n44146) );
  XNOR2HSV4 U48207 ( .A1(n44147), .A2(n44146), .ZN(n44154) );
  NAND3HSV4 U48208 ( .A1(n44148), .A2(n43917), .A3(n44149), .ZN(n44152) );
  INHSV2 U48209 ( .I(n59980), .ZN(n52411) );
  AOI31HSV2 U48210 ( .A1(n26883), .A2(n44150), .A3(n44149), .B(n52411), .ZN(
        n44151) );
  XNOR2HSV4 U48211 ( .A1(n44154), .A2(n44153), .ZN(n44164) );
  INHSV4 U48212 ( .I(n44164), .ZN(n44162) );
  AND2HSV2 U48213 ( .A1(n45409), .A2(n38890), .Z(n45407) );
  NAND3HSV2 U48214 ( .A1(n44155), .A2(n29769), .A3(n45407), .ZN(n44163) );
  CLKNAND2HSV1 U48215 ( .A1(n44158), .A2(n44157), .ZN(n44160) );
  CLKNAND2HSV1 U48216 ( .A1(n44298), .A2(n36414), .ZN(n44159) );
  INOR2HSV4 U48217 ( .A1(n44163), .B1(n44165), .ZN(n44161) );
  CLKNHSV2 U48218 ( .I(\pe2/ti_7t [26]), .ZN(n44167) );
  OR2HSV1 U48219 ( .A1(n44309), .A2(n44167), .Z(n45108) );
  NAND2HSV2 U48220 ( .A1(n44169), .A2(n44309), .ZN(n44170) );
  CLKNHSV0 U48221 ( .I(n44303), .ZN(n44171) );
  NAND2HSV2 U48222 ( .A1(n45089), .A2(n44171), .ZN(n45112) );
  INHSV2 U48223 ( .I(n45112), .ZN(n44172) );
  CLKBUFHSV4 U48224 ( .I(n47554), .Z(n47939) );
  INHSV2 U48225 ( .I(n47939), .ZN(n59929) );
  BUFHSV4 U48226 ( .I(n54729), .Z(n59736) );
  NAND3HSV4 U48227 ( .A1(n44176), .A2(n44175), .A3(n44174), .ZN(n44182) );
  NAND2HSV4 U48228 ( .A1(n44182), .A2(n38873), .ZN(n44306) );
  NAND2HSV4 U48229 ( .A1(n44183), .A2(n44300), .ZN(n44832) );
  NAND2HSV2 U48230 ( .A1(n44832), .A2(n45388), .ZN(n44293) );
  CLKBUFHSV4 U48231 ( .I(n51687), .Z(n51485) );
  CLKNAND2HSV2 U48232 ( .A1(n51687), .A2(n38512), .ZN(n44287) );
  CLKNAND2HSV0 U48233 ( .A1(n45249), .A2(n25824), .ZN(n44280) );
  NAND2HSV2 U48234 ( .A1(n59634), .A2(n38390), .ZN(n44275) );
  CLKNAND2HSV1 U48235 ( .A1(n44713), .A2(n39075), .ZN(n44273) );
  NAND2HSV0 U48236 ( .A1(n47571), .A2(n52929), .ZN(n44271) );
  BUFHSV4 U48237 ( .I(n50929), .Z(n52287) );
  NAND2HSV2 U48238 ( .A1(n52287), .A2(n51796), .ZN(n44268) );
  NAND2HSV2 U48239 ( .A1(n52932), .A2(n44186), .ZN(n44260) );
  NAND2HSV2 U48240 ( .A1(n52053), .A2(n52172), .ZN(n44258) );
  NAND2HSV0 U48241 ( .A1(n44715), .A2(\pe2/got [10]), .ZN(n44253) );
  BUFHSV2 U48242 ( .I(n44187), .Z(n59684) );
  CLKNAND2HSV1 U48243 ( .A1(n59684), .A2(n44714), .ZN(n44190) );
  NOR2HSV0 U48244 ( .A1(n44971), .A2(n44188), .ZN(n44189) );
  XOR2HSV0 U48245 ( .A1(n44190), .A2(n44189), .Z(n44251) );
  CLKNHSV0 U48246 ( .I(n50928), .ZN(n59757) );
  CLKNAND2HSV1 U48247 ( .A1(n38291), .A2(n59757), .ZN(n44249) );
  CLKNAND2HSV0 U48248 ( .A1(n45295), .A2(n51900), .ZN(n44192) );
  NAND2HSV0 U48249 ( .A1(n59768), .A2(\pe2/bq[29] ), .ZN(n44191) );
  XOR2HSV0 U48250 ( .A1(n44192), .A2(n44191), .Z(n44196) );
  CLKNAND2HSV0 U48251 ( .A1(n53009), .A2(n38565), .ZN(n44194) );
  CLKNAND2HSV0 U48252 ( .A1(n52457), .A2(n39020), .ZN(n44193) );
  XOR2HSV0 U48253 ( .A1(n44194), .A2(n44193), .Z(n44195) );
  XOR2HSV0 U48254 ( .A1(n44196), .A2(n44195), .Z(n44204) );
  CLKNHSV0 U48255 ( .I(n52103), .ZN(n52955) );
  CLKNAND2HSV1 U48256 ( .A1(n52955), .A2(n44197), .ZN(n44199) );
  NAND2HSV0 U48257 ( .A1(n39029), .A2(n44074), .ZN(n44198) );
  XOR2HSV0 U48258 ( .A1(n44199), .A2(n44198), .Z(n44202) );
  NAND2HSV0 U48259 ( .A1(n38576), .A2(\pe2/pvq [27]), .ZN(n44200) );
  XOR2HSV0 U48260 ( .A1(n44200), .A2(\pe2/phq [27]), .Z(n44201) );
  XOR2HSV0 U48261 ( .A1(n44202), .A2(n44201), .Z(n44203) );
  XOR2HSV0 U48262 ( .A1(n44204), .A2(n44203), .Z(n44216) );
  NOR2HSV0 U48263 ( .A1(n52226), .A2(n44718), .ZN(n51972) );
  INHSV2 U48264 ( .I(n44718), .ZN(n52866) );
  AOI22HSV0 U48265 ( .A1(n44750), .A2(n52866), .B1(n38054), .B2(n59973), .ZN(
        n44205) );
  AOI21HSV0 U48266 ( .A1(n44206), .A2(n51972), .B(n44205), .ZN(n44211) );
  NAND2HSV0 U48267 ( .A1(n44207), .A2(\pe2/bq[7] ), .ZN(n44767) );
  NAND2HSV0 U48268 ( .A1(n38061), .A2(\pe2/bq[7] ), .ZN(n44890) );
  OAI21HSV0 U48269 ( .A1(n51567), .A2(n38404), .B(n44890), .ZN(n44208) );
  OAI21HSV1 U48270 ( .A1(n44767), .A2(n44209), .B(n44208), .ZN(n44210) );
  XOR2HSV0 U48271 ( .A1(n44211), .A2(n44210), .Z(n44214) );
  NAND2HSV2 U48272 ( .A1(n52995), .A2(n51997), .ZN(n45182) );
  NAND2HSV0 U48273 ( .A1(\pe2/aot [17]), .A2(\pe2/bq[21] ), .ZN(n51968) );
  XOR2HSV0 U48274 ( .A1(n45182), .A2(n51968), .Z(n44213) );
  XNOR2HSV1 U48275 ( .A1(n44214), .A2(n44213), .ZN(n44215) );
  XNOR2HSV1 U48276 ( .A1(n44216), .A2(n44215), .ZN(n44248) );
  NAND2HSV0 U48277 ( .A1(n44745), .A2(n45015), .ZN(n44218) );
  NAND2HSV0 U48278 ( .A1(\pe2/aot [23]), .A2(n52337), .ZN(n44217) );
  XOR2HSV0 U48279 ( .A1(n44218), .A2(n44217), .Z(n44222) );
  NAND2HSV0 U48280 ( .A1(n59972), .A2(\pe2/bq[14] ), .ZN(n44220) );
  CLKNAND2HSV0 U48281 ( .A1(n52294), .A2(n38792), .ZN(n44219) );
  XOR2HSV0 U48282 ( .A1(n44220), .A2(n44219), .Z(n44221) );
  XOR2HSV0 U48283 ( .A1(n44222), .A2(n44221), .Z(n44230) );
  NAND2HSV0 U48284 ( .A1(\pe2/aot [22]), .A2(n38803), .ZN(n44224) );
  CLKNAND2HSV0 U48285 ( .A1(\pe2/aot [6]), .A2(n53015), .ZN(n44223) );
  XOR2HSV0 U48286 ( .A1(n44224), .A2(n44223), .Z(n44228) );
  NAND2HSV0 U48287 ( .A1(n52485), .A2(n52193), .ZN(n44226) );
  NAND2HSV0 U48288 ( .A1(\pe2/aot [12]), .A2(n38064), .ZN(n44225) );
  XOR2HSV0 U48289 ( .A1(n44226), .A2(n44225), .Z(n44227) );
  XOR2HSV0 U48290 ( .A1(n44228), .A2(n44227), .Z(n44229) );
  XOR2HSV0 U48291 ( .A1(n44230), .A2(n44229), .Z(n44246) );
  BUFHSV2 U48292 ( .I(\pe2/bq[12] ), .Z(n53006) );
  CLKNAND2HSV1 U48293 ( .A1(n52974), .A2(n53006), .ZN(n44233) );
  NAND2HSV0 U48294 ( .A1(\pe2/aot [25]), .A2(n44231), .ZN(n44232) );
  XOR2HSV0 U48295 ( .A1(n44233), .A2(n44232), .Z(n44237) );
  NAND2HSV0 U48296 ( .A1(n45034), .A2(n44987), .ZN(n44235) );
  CLKNHSV0 U48297 ( .I(n52018), .ZN(n53041) );
  CLKNAND2HSV0 U48298 ( .A1(n53041), .A2(n45008), .ZN(n44234) );
  XOR2HSV0 U48299 ( .A1(n44235), .A2(n44234), .Z(n44236) );
  XOR2HSV0 U48300 ( .A1(n44237), .A2(n44236), .Z(n44244) );
  NAND2HSV0 U48301 ( .A1(n59633), .A2(n36607), .ZN(n52443) );
  XOR2HSV0 U48302 ( .A1(n44238), .A2(n52443), .Z(n44242) );
  CLKNAND2HSV0 U48303 ( .A1(n39019), .A2(n52973), .ZN(n44240) );
  NAND2HSV0 U48304 ( .A1(n59974), .A2(n52300), .ZN(n44239) );
  XOR2HSV0 U48305 ( .A1(n44240), .A2(n44239), .Z(n44241) );
  XOR2HSV0 U48306 ( .A1(n44242), .A2(n44241), .Z(n44243) );
  XOR2HSV0 U48307 ( .A1(n44244), .A2(n44243), .Z(n44245) );
  XOR2HSV0 U48308 ( .A1(n44246), .A2(n44245), .Z(n44247) );
  XOR3HSV2 U48309 ( .A1(n44249), .A2(n44248), .A3(n44247), .Z(n44250) );
  XNOR2HSV1 U48310 ( .A1(n44251), .A2(n44250), .ZN(n44252) );
  XNOR2HSV1 U48311 ( .A1(n44253), .A2(n44252), .ZN(n44256) );
  NAND2HSV0 U48312 ( .A1(n44254), .A2(n52374), .ZN(n44255) );
  XNOR2HSV1 U48313 ( .A1(n44256), .A2(n44255), .ZN(n44257) );
  XNOR2HSV1 U48314 ( .A1(n44258), .A2(n44257), .ZN(n44259) );
  XNOR2HSV1 U48315 ( .A1(n44260), .A2(n44259), .ZN(n44263) );
  CLKNAND2HSV1 U48316 ( .A1(n44261), .A2(n48084), .ZN(n44262) );
  XOR2HSV0 U48317 ( .A1(n44263), .A2(n44262), .Z(n44266) );
  CLKNHSV1 U48318 ( .I(n44264), .ZN(n53050) );
  INHSV2 U48319 ( .I(n47573), .ZN(n51964) );
  CLKNAND2HSV1 U48320 ( .A1(n53050), .A2(n51964), .ZN(n44265) );
  XNOR2HSV1 U48321 ( .A1(n44266), .A2(n44265), .ZN(n44267) );
  XNOR2HSV1 U48322 ( .A1(n44268), .A2(n44267), .ZN(n44270) );
  CLKNAND2HSV1 U48323 ( .A1(n45063), .A2(n44712), .ZN(n44269) );
  XOR3HSV2 U48324 ( .A1(n44271), .A2(n44270), .A3(n44269), .Z(n44272) );
  XNOR2HSV1 U48325 ( .A1(n44273), .A2(n44272), .ZN(n44274) );
  NOR2HSV2 U48326 ( .A1(n45071), .A2(n45248), .ZN(n44276) );
  XNOR2HSV1 U48327 ( .A1(n44280), .A2(n44279), .ZN(n44281) );
  XNOR2HSV1 U48328 ( .A1(n44282), .A2(n44281), .ZN(n44285) );
  INHSV4 U48329 ( .I(n44283), .ZN(n59361) );
  NAND2HSV2 U48330 ( .A1(n59361), .A2(n44711), .ZN(n44284) );
  XNOR2HSV4 U48331 ( .A1(n44287), .A2(n44286), .ZN(n44289) );
  XOR2HSV2 U48332 ( .A1(n44289), .A2(n44288), .Z(n44291) );
  NAND2HSV2 U48333 ( .A1(n45083), .A2(n38327), .ZN(n44290) );
  XNOR2HSV4 U48334 ( .A1(n44291), .A2(n44290), .ZN(n44292) );
  XNOR2HSV4 U48335 ( .A1(n44293), .A2(n44292), .ZN(n44305) );
  CLKBUFHSV2 U48336 ( .I(n52827), .Z(n44299) );
  CLKNHSV0 U48337 ( .I(n44295), .ZN(n44301) );
  AOI31HSV2 U48338 ( .A1(n44301), .A2(n44300), .A3(n44296), .B(n36519), .ZN(
        n44297) );
  CLKNHSV0 U48339 ( .I(n29769), .ZN(n44302) );
  CLKNAND2HSV1 U48340 ( .A1(\pe2/ti_7t [25]), .A2(n38195), .ZN(n44304) );
  AOI21HSV4 U48341 ( .A1(n44323), .A2(n44030), .B(n44314), .ZN(n44953) );
  CLKAND2HSV1 U48342 ( .A1(n44313), .A2(n44322), .Z(n44308) );
  NAND3HSV4 U48343 ( .A1(n44954), .A2(n29680), .A3(n44955), .ZN(n44708) );
  AND2HSV2 U48344 ( .A1(n44313), .A2(n44309), .Z(n44310) );
  CLKNAND2HSV2 U48345 ( .A1(n44311), .A2(n44310), .ZN(n44320) );
  NOR2HSV4 U48346 ( .A1(n26799), .A2(n36563), .ZN(n44318) );
  INHSV2 U48347 ( .I(n44960), .ZN(n44317) );
  AOI21HSV2 U48348 ( .A1(n60028), .A2(n44318), .B(n44317), .ZN(n44319) );
  CLKNAND2HSV3 U48349 ( .A1(n44319), .A2(n44320), .ZN(n44707) );
  NOR2HSV2 U48350 ( .A1(n44323), .A2(n45114), .ZN(n44959) );
  NOR2HSV2 U48351 ( .A1(n44323), .A2(n44322), .ZN(n44324) );
  NOR2HSV4 U48352 ( .A1(n44324), .A2(n44821), .ZN(n44956) );
  NAND3HSV4 U48353 ( .A1(n44962), .A2(n44325), .A3(n44956), .ZN(n44706) );
  INHSV4 U48354 ( .I(n44326), .ZN(n59927) );
  INHSV2 U48355 ( .I(n44327), .ZN(n59685) );
  INHSV2 U48356 ( .I(n44328), .ZN(n50717) );
  INHSV1 U48357 ( .I(n50717), .ZN(n59527) );
  CLKNHSV0 U48358 ( .I(n55612), .ZN(n59359) );
  CLKNHSV0 U48359 ( .I(n44329), .ZN(n59516) );
  CLKNAND2HSV1 U48360 ( .A1(n53656), .A2(n53655), .ZN(n59521) );
  CLKNHSV0 U48361 ( .I(n48484), .ZN(n59930) );
  INHSV2 U48362 ( .I(n44330), .ZN(n58448) );
  CLKBUFHSV2 U48363 ( .I(n58448), .Z(n59918) );
  CLKNHSV0 U48364 ( .I(n54037), .ZN(n59422) );
  BUFHSV2 U48365 ( .I(n47842), .Z(n59672) );
  BUFHSV2 U48366 ( .I(n45818), .Z(n59894) );
  BUFHSV2 U48367 ( .I(n44331), .Z(n44834) );
  INHSV2 U48368 ( .I(n44834), .ZN(n59506) );
  CLKNHSV0 U48369 ( .I(n56936), .ZN(n59807) );
  CLKNHSV0 U48370 ( .I(n56778), .ZN(n59647) );
  BUFHSV2 U48371 ( .I(n37177), .Z(n59797) );
  NAND2HSV0 U48372 ( .A1(n59797), .A2(n52726), .ZN(n44334) );
  XNOR2HSV0 U48373 ( .A1(n44334), .A2(n44333), .ZN(n60029) );
  MUX2HSV1 U48374 ( .I0(bo3[30]), .I1(n45663), .S(n46127), .Z(n59760) );
  MUX2HSV1 U48375 ( .I0(bo3[4]), .I1(\pe3/bq[4] ), .S(n46128), .Z(n59561) );
  INHSV2 U48376 ( .I(\pe5/bq[1] ), .ZN(n45421) );
  MUX2HSV1 U48377 ( .I0(bo5[1]), .I1(n52581), .S(n48039), .Z(n59865) );
  MUX2HSV1 U48378 ( .I0(bo5[24]), .I1(n30891), .S(n48077), .Z(n59842) );
  MUX2HSV1 U48379 ( .I0(bo1[19]), .I1(n42092), .S(n48053), .Z(n59702) );
  MUX2HSV1 U48380 ( .I0(bo1[27]), .I1(\pe1/bq[27] ), .S(n48053), .Z(n59694) );
  MUX2HSV1 U48381 ( .I0(bo1[30]), .I1(n53411), .S(n48054), .Z(n59691) );
  BUFHSV2 U48382 ( .I(\pe6/ctrq ), .Z(n48036) );
  MUX2HSV1 U48383 ( .I0(bo6[16]), .I1(n49844), .S(n48043), .Z(n59898) );
  MUX2HSV1 U48384 ( .I0(bo6[14]), .I1(n58668), .S(n59902), .Z(n59538) );
  MUX2HSV1 U48385 ( .I0(bo6[24]), .I1(n44453), .S(n48025), .Z(n59874) );
  MUX2HSV1 U48386 ( .I0(bo6[10]), .I1(n44336), .S(n59201), .Z(n59906) );
  MUX2HSV1 U48387 ( .I0(bo1[12]), .I1(n42373), .S(n48061), .Z(n59709) );
  MUX2HSV1 U48388 ( .I0(bo1[9]), .I1(\pe1/bq[9] ), .S(n48061), .Z(n59710) );
  CLKNHSV0 U48389 ( .I(n50518), .ZN(n59881) );
  CLKNHSV1 U48390 ( .I(n44338), .ZN(n59857) );
  NOR2HSV1 U48391 ( .A1(n44339), .A2(n46549), .ZN(n44340) );
  CLKNHSV0 U48392 ( .I(n46575), .ZN(n44343) );
  CLKNAND2HSV1 U48393 ( .A1(n44343), .A2(n44342), .ZN(n44347) );
  AND2HSV2 U48394 ( .A1(n44344), .A2(n32053), .Z(n44345) );
  NAND3HSV2 U48395 ( .A1(n44347), .A2(n44346), .A3(n44345), .ZN(n44348) );
  AND2HSV2 U48396 ( .A1(n44378), .A2(n46163), .Z(n44350) );
  NOR2HSV2 U48397 ( .A1(n44354), .A2(n44353), .ZN(n44356) );
  CLKNAND2HSV1 U48398 ( .A1(n44356), .A2(n44355), .ZN(n44361) );
  XNOR2HSV4 U48399 ( .A1(n44367), .A2(n44366), .ZN(n44381) );
  NAND2HSV2 U48400 ( .A1(n44368), .A2(n44381), .ZN(n44374) );
  INHSV6 U48401 ( .I(n44381), .ZN(n45787) );
  OR2HSV1 U48402 ( .A1(n44369), .A2(n52705), .Z(n44370) );
  NOR2HSV2 U48403 ( .A1(n47932), .A2(n44370), .ZN(n44371) );
  CLKNAND2HSV3 U48404 ( .A1(n45787), .A2(n44371), .ZN(n44373) );
  CLKNAND2HSV0 U48405 ( .A1(\pe6/ti_7t [28]), .A2(n46584), .ZN(n45784) );
  OR2HSV1 U48406 ( .A1(n45784), .A2(n44372), .Z(n44382) );
  NAND3HSV4 U48407 ( .A1(n44373), .A2(n44374), .A3(n44382), .ZN(n44388) );
  INAND2HSV2 U48408 ( .A1(n44376), .B1(n44375), .ZN(n44377) );
  CLKAND2HSV2 U48409 ( .A1(n47932), .A2(n44378), .Z(n45788) );
  NOR2HSV2 U48410 ( .A1(n47932), .A2(n44380), .ZN(n45786) );
  NOR2HSV2 U48411 ( .A1(n44381), .A2(n32457), .ZN(n44384) );
  CLKNHSV0 U48412 ( .I(n44382), .ZN(n44383) );
  AOI21HSV2 U48413 ( .A1(n45786), .A2(n44384), .B(n44383), .ZN(n44385) );
  AOI22HSV4 U48414 ( .A1(n44388), .A2(n44387), .B1(n44386), .B2(n44385), .ZN(
        n44518) );
  CLKNAND2HSV1 U48415 ( .A1(n44389), .A2(n59022), .ZN(n44517) );
  NAND2HSV2 U48416 ( .A1(n58480), .A2(n49665), .ZN(n44513) );
  CLKNAND2HSV1 U48417 ( .A1(n46769), .A2(n31717), .ZN(n44506) );
  NAND2HSV0 U48418 ( .A1(n44390), .A2(n58714), .ZN(n44502) );
  NAND2HSV2 U48419 ( .A1(n58663), .A2(\pe6/got [21]), .ZN(n44500) );
  NAND2HSV2 U48420 ( .A1(n58664), .A2(n59176), .ZN(n44498) );
  INHSV2 U48421 ( .I(n53103), .ZN(n59178) );
  NAND2HSV0 U48422 ( .A1(n49667), .A2(n59178), .ZN(n44491) );
  BUFHSV2 U48423 ( .I(n44391), .Z(n59379) );
  NAND2HSV2 U48424 ( .A1(n59379), .A2(n46171), .ZN(n44489) );
  BUFHSV2 U48425 ( .I(n44392), .Z(n58813) );
  NAND2HSV0 U48426 ( .A1(n58813), .A2(\pe6/got [15]), .ZN(n44487) );
  NAND2HSV0 U48427 ( .A1(n49743), .A2(n35991), .ZN(n44485) );
  NAND2HSV0 U48428 ( .A1(n49829), .A2(n58711), .ZN(n44483) );
  NAND2HSV0 U48429 ( .A1(n58939), .A2(n59180), .ZN(n44481) );
  NAND2HSV2 U48430 ( .A1(n36107), .A2(n44393), .ZN(n44475) );
  BUFHSV2 U48431 ( .I(\pe6/got [9]), .Z(n58477) );
  NAND2HSV0 U48432 ( .A1(n59183), .A2(n58477), .ZN(n44473) );
  BUFHSV2 U48433 ( .I(n58399), .Z(n58398) );
  NAND2HSV0 U48434 ( .A1(n36108), .A2(n58398), .ZN(n44395) );
  NAND2HSV0 U48435 ( .A1(n59038), .A2(n58400), .ZN(n44394) );
  XOR2HSV0 U48436 ( .A1(n44395), .A2(n44394), .Z(n44467) );
  CLKNAND2HSV1 U48437 ( .A1(n59224), .A2(n58842), .ZN(n49026) );
  NAND2HSV0 U48438 ( .A1(n59224), .A2(n46217), .ZN(n50828) );
  OAI21HSV0 U48439 ( .A1(n44396), .A2(n35837), .B(n50828), .ZN(n44398) );
  OAI21HSV2 U48440 ( .A1(n44399), .A2(n49026), .B(n44398), .ZN(n44400) );
  NAND2HSV0 U48441 ( .A1(n46210), .A2(n58749), .ZN(n58853) );
  XNOR2HSV1 U48442 ( .A1(n44400), .A2(n58853), .ZN(n44402) );
  NAND2HSV0 U48443 ( .A1(n48051), .A2(\pe6/aot [23]), .ZN(n58974) );
  CLKNAND2HSV1 U48444 ( .A1(n36150), .A2(\pe6/aot [17]), .ZN(n46838) );
  XOR2HSV0 U48445 ( .A1(n58974), .A2(n46838), .Z(n44401) );
  XNOR2HSV1 U48446 ( .A1(n44402), .A2(n44401), .ZN(n44410) );
  CLKNAND2HSV1 U48447 ( .A1(n59202), .A2(n53115), .ZN(n49331) );
  CLKNAND2HSV1 U48448 ( .A1(n46626), .A2(\pe6/pvq [30]), .ZN(n44404) );
  XOR2HSV0 U48449 ( .A1(n49331), .A2(n44404), .Z(n44408) );
  NAND2HSV0 U48450 ( .A1(n58965), .A2(n58857), .ZN(n44406) );
  CLKNHSV0 U48451 ( .I(n46663), .ZN(n58824) );
  CLKNAND2HSV0 U48452 ( .A1(n44336), .A2(n58824), .ZN(n44405) );
  XOR2HSV0 U48453 ( .A1(n44406), .A2(n44405), .Z(n44407) );
  XOR2HSV0 U48454 ( .A1(n44408), .A2(n44407), .Z(n44409) );
  XOR2HSV0 U48455 ( .A1(n44410), .A2(n44409), .Z(n44465) );
  NAND2HSV0 U48456 ( .A1(n32252), .A2(n46197), .ZN(n44413) );
  NAND2HSV0 U48457 ( .A1(n46658), .A2(n58459), .ZN(n44412) );
  XOR2HSV0 U48458 ( .A1(n44413), .A2(n44412), .Z(n44417) );
  CLKNAND2HSV0 U48459 ( .A1(n32999), .A2(n46792), .ZN(n44415) );
  NAND2HSV0 U48460 ( .A1(n46672), .A2(n58378), .ZN(n44414) );
  XOR2HSV0 U48461 ( .A1(n44415), .A2(n44414), .Z(n44416) );
  XOR2HSV0 U48462 ( .A1(n44417), .A2(n44416), .Z(n44425) );
  INHSV2 U48463 ( .I(n49681), .ZN(n58734) );
  NAND2HSV0 U48464 ( .A1(n46627), .A2(n58734), .ZN(n44419) );
  NAND2HSV0 U48465 ( .A1(n58619), .A2(n32981), .ZN(n44418) );
  XOR2HSV0 U48466 ( .A1(n44419), .A2(n44418), .Z(n44423) );
  INHSV2 U48467 ( .I(n46146), .ZN(n58356) );
  CLKNHSV0 U48468 ( .I(n32714), .ZN(n59040) );
  NAND2HSV0 U48469 ( .A1(n58356), .A2(n59040), .ZN(n44421) );
  NAND2HSV0 U48470 ( .A1(n49862), .A2(n58943), .ZN(n44420) );
  XOR2HSV0 U48471 ( .A1(n44421), .A2(n44420), .Z(n44422) );
  XOR2HSV0 U48472 ( .A1(n44423), .A2(n44422), .Z(n44424) );
  XOR2HSV0 U48473 ( .A1(n44425), .A2(n44424), .Z(n44428) );
  NAND2HSV0 U48474 ( .A1(n44426), .A2(n46173), .ZN(n44427) );
  XNOR2HSV1 U48475 ( .A1(n44428), .A2(n44427), .ZN(n44464) );
  INHSV2 U48476 ( .I(n49327), .ZN(n58339) );
  NAND2HSV0 U48477 ( .A1(n58339), .A2(n46230), .ZN(n44430) );
  NAND2HSV0 U48478 ( .A1(n58618), .A2(n31829), .ZN(n44429) );
  XOR2HSV0 U48479 ( .A1(n44430), .A2(n44429), .Z(n44434) );
  NAND2HSV0 U48480 ( .A1(n49844), .A2(\pe6/aot [19]), .ZN(n44432) );
  NAND2HSV0 U48481 ( .A1(n58668), .A2(\pe6/aot [21]), .ZN(n44431) );
  XOR2HSV0 U48482 ( .A1(n44432), .A2(n44431), .Z(n44433) );
  XOR2HSV0 U48483 ( .A1(n44434), .A2(n44433), .Z(n44445) );
  NAND2HSV0 U48484 ( .A1(n44435), .A2(\pe6/aot [13]), .ZN(n44438) );
  NAND2HSV0 U48485 ( .A1(\pe6/bq[9] ), .A2(n32876), .ZN(n44437) );
  XOR2HSV0 U48486 ( .A1(n44438), .A2(n44437), .Z(n44443) );
  NAND2HSV0 U48487 ( .A1(\pe6/bq[15] ), .A2(n44439), .ZN(n44441) );
  NAND2HSV0 U48488 ( .A1(n59206), .A2(n58488), .ZN(n44440) );
  XOR2HSV0 U48489 ( .A1(n44441), .A2(n44440), .Z(n44442) );
  XOR2HSV0 U48490 ( .A1(n44443), .A2(n44442), .Z(n44444) );
  XOR2HSV0 U48491 ( .A1(n44445), .A2(n44444), .Z(n44462) );
  NOR2HSV0 U48492 ( .A1(n46853), .A2(n32373), .ZN(n44448) );
  NAND2HSV0 U48493 ( .A1(\pe6/bq[4] ), .A2(n44446), .ZN(n44447) );
  XOR2HSV0 U48494 ( .A1(n44448), .A2(n44447), .Z(n44452) );
  NAND2HSV0 U48495 ( .A1(n32982), .A2(n59088), .ZN(n44450) );
  NAND2HSV0 U48496 ( .A1(n59247), .A2(n59266), .ZN(n44449) );
  XOR2HSV0 U48497 ( .A1(n44450), .A2(n44449), .Z(n44451) );
  XOR2HSV0 U48498 ( .A1(n44452), .A2(n44451), .Z(n44460) );
  NOR2HSV0 U48499 ( .A1(n48041), .A2(n35816), .ZN(n44455) );
  NAND2HSV0 U48500 ( .A1(n44453), .A2(\pe6/aot [11]), .ZN(n44454) );
  XOR2HSV0 U48501 ( .A1(n44455), .A2(n44454), .Z(n44458) );
  NAND2HSV0 U48502 ( .A1(n46176), .A2(n48891), .ZN(n44456) );
  XOR2HSV0 U48503 ( .A1(n44456), .A2(\pe6/phq [30]), .Z(n44457) );
  XOR2HSV0 U48504 ( .A1(n44458), .A2(n44457), .Z(n44459) );
  XOR2HSV0 U48505 ( .A1(n44460), .A2(n44459), .Z(n44461) );
  XOR2HSV0 U48506 ( .A1(n44462), .A2(n44461), .Z(n44463) );
  XOR3HSV2 U48507 ( .A1(n44465), .A2(n44464), .A3(n44463), .Z(n44466) );
  XNOR2HSV1 U48508 ( .A1(n44467), .A2(n44466), .ZN(n44469) );
  NAND2HSV0 U48509 ( .A1(n59670), .A2(n58814), .ZN(n44468) );
  XNOR2HSV1 U48510 ( .A1(n44469), .A2(n44468), .ZN(n44471) );
  NAND2HSV0 U48511 ( .A1(n32293), .A2(n58526), .ZN(n44470) );
  XNOR2HSV1 U48512 ( .A1(n44471), .A2(n44470), .ZN(n44472) );
  XNOR2HSV1 U48513 ( .A1(n44473), .A2(n44472), .ZN(n44474) );
  XNOR2HSV1 U48514 ( .A1(n44475), .A2(n44474), .ZN(n44479) );
  BUFHSV2 U48515 ( .I(n44476), .Z(n59917) );
  NAND2HSV2 U48516 ( .A1(n58886), .A2(n44477), .ZN(n44478) );
  XNOR2HSV1 U48517 ( .A1(n44479), .A2(n44478), .ZN(n44480) );
  XOR2HSV0 U48518 ( .A1(n44481), .A2(n44480), .Z(n44482) );
  XNOR2HSV1 U48519 ( .A1(n44483), .A2(n44482), .ZN(n44484) );
  XOR2HSV0 U48520 ( .A1(n44485), .A2(n44484), .Z(n44486) );
  XOR2HSV0 U48521 ( .A1(n44487), .A2(n44486), .Z(n44488) );
  XNOR2HSV1 U48522 ( .A1(n44489), .A2(n44488), .ZN(n44490) );
  XOR2HSV0 U48523 ( .A1(n44491), .A2(n44490), .Z(n44493) );
  NAND2HSV0 U48524 ( .A1(n59144), .A2(n36104), .ZN(n44492) );
  XOR2HSV0 U48525 ( .A1(n44493), .A2(n44492), .Z(n44496) );
  NAND2HSV0 U48526 ( .A1(n59676), .A2(n58807), .ZN(n44495) );
  XOR2HSV0 U48527 ( .A1(n44496), .A2(n44495), .Z(n44497) );
  XOR2HSV0 U48528 ( .A1(n44498), .A2(n44497), .Z(n44499) );
  XNOR2HSV1 U48529 ( .A1(n44500), .A2(n44499), .ZN(n44501) );
  XNOR2HSV1 U48530 ( .A1(n44502), .A2(n44501), .ZN(n44504) );
  NAND2HSV2 U48531 ( .A1(n58601), .A2(n58808), .ZN(n44503) );
  XNOR2HSV1 U48532 ( .A1(n44504), .A2(n44503), .ZN(n44505) );
  XNOR2HSV1 U48533 ( .A1(n44506), .A2(n44505), .ZN(n44511) );
  INAND2HSV2 U48534 ( .A1(n44507), .B1(n59918), .ZN(n44510) );
  BUFHSV2 U48535 ( .I(n44508), .Z(n49078) );
  NAND2HSV2 U48536 ( .A1(n49078), .A2(n32354), .ZN(n44509) );
  XOR3HSV2 U48537 ( .A1(n44511), .A2(n44510), .A3(n44509), .Z(n44512) );
  XNOR2HSV1 U48538 ( .A1(n44513), .A2(n44512), .ZN(n44516) );
  INHSV2 U48539 ( .I(n44514), .ZN(n49400) );
  XNOR2HSV4 U48540 ( .A1(n44518), .A2(n29655), .ZN(n46167) );
  NOR2HSV4 U48541 ( .A1(n46302), .A2(n46546), .ZN(n46630) );
  CLKNAND2HSV1 U48542 ( .A1(n48001), .A2(\pe6/ti_7t [30]), .ZN(n49737) );
  INHSV4 U48543 ( .I(n49737), .ZN(n49178) );
  NOR2HSV4 U48544 ( .A1(n46630), .A2(n49178), .ZN(n58348) );
  NAND2HSV2 U48545 ( .A1(n40162), .A2(\pe5/ti_7t [31]), .ZN(n47052) );
  NAND2HSV2 U48546 ( .A1(n47141), .A2(n47052), .ZN(n59421) );
  INHSV2 U48547 ( .I(n44522), .ZN(n44523) );
  CLKNAND2HSV1 U48548 ( .A1(n44524), .A2(n51114), .ZN(n44525) );
  INHSV4 U48549 ( .I(n53503), .ZN(n55490) );
  INAND2HSV2 U48550 ( .A1(n48451), .B1(n53512), .ZN(n44643) );
  NAND2HSV0 U48551 ( .A1(n55229), .A2(\pe1/got [25]), .ZN(n44638) );
  BUFHSV2 U48552 ( .I(n59391), .Z(n53521) );
  NAND2HSV2 U48553 ( .A1(n53521), .A2(\pe1/got [23]), .ZN(n44634) );
  NOR2HSV2 U48554 ( .A1(n53391), .A2(n42209), .ZN(n44632) );
  BUFHSV2 U48555 ( .I(n55091), .Z(n53522) );
  NAND2HSV2 U48556 ( .A1(n53522), .A2(\pe1/got [21]), .ZN(n44630) );
  CLKNAND2HSV1 U48557 ( .A1(n53392), .A2(n44530), .ZN(n44628) );
  NOR2HSV2 U48558 ( .A1(n54454), .A2(n41928), .ZN(n44626) );
  NAND2HSV0 U48559 ( .A1(n59518), .A2(n54135), .ZN(n44624) );
  NAND2HSV0 U48560 ( .A1(n53913), .A2(\pe1/got [16]), .ZN(n44621) );
  CLKNAND2HSV1 U48561 ( .A1(n54041), .A2(n48339), .ZN(n44619) );
  NOR2HSV1 U48562 ( .A1(n41802), .A2(n54957), .ZN(n44615) );
  NAND2HSV0 U48563 ( .A1(n41332), .A2(\pe1/got [11]), .ZN(n44611) );
  NAND2HSV2 U48564 ( .A1(n53524), .A2(n55339), .ZN(n44604) );
  CLKNAND2HSV1 U48565 ( .A1(n53979), .A2(n53523), .ZN(n44602) );
  NAND2HSV2 U48566 ( .A1(n53795), .A2(n59750), .ZN(n44601) );
  NAND2HSV0 U48567 ( .A1(n44533), .A2(\pe1/bq[23] ), .ZN(n44535) );
  NAND2HSV0 U48568 ( .A1(\pe1/aot [22]), .A2(n54179), .ZN(n44534) );
  XOR2HSV0 U48569 ( .A1(n44535), .A2(n44534), .Z(n44539) );
  CLKNAND2HSV0 U48570 ( .A1(\pe1/aot [14]), .A2(\pe1/bq[21] ), .ZN(n44536) );
  XOR2HSV0 U48571 ( .A1(n44537), .A2(n44536), .Z(n44538) );
  XOR2HSV0 U48572 ( .A1(n44539), .A2(n44538), .Z(n44565) );
  CLKNAND2HSV0 U48573 ( .A1(n59675), .A2(n53863), .ZN(n44545) );
  NAND2HSV0 U48574 ( .A1(n59990), .A2(n55379), .ZN(n54642) );
  NOR2HSV0 U48575 ( .A1(n44540), .A2(n54642), .ZN(n44543) );
  AOI22HSV0 U48576 ( .A1(n41743), .A2(n55352), .B1(n54465), .B2(n44541), .ZN(
        n44542) );
  NOR2HSV2 U48577 ( .A1(n44543), .A2(n44542), .ZN(n44544) );
  XNOR2HSV1 U48578 ( .A1(n44545), .A2(n44544), .ZN(n44547) );
  NAND2HSV0 U48579 ( .A1(n26833), .A2(\pe1/got [5]), .ZN(n44546) );
  XOR2HSV0 U48580 ( .A1(n44547), .A2(n44546), .Z(n44564) );
  CLKNAND2HSV0 U48581 ( .A1(n41768), .A2(n48380), .ZN(n44549) );
  NAND2HSV0 U48582 ( .A1(n54307), .A2(\pe1/bq[11] ), .ZN(n44548) );
  XOR2HSV0 U48583 ( .A1(n44549), .A2(n44548), .Z(n44553) );
  CLKNAND2HSV1 U48584 ( .A1(n54500), .A2(n54995), .ZN(n44551) );
  NAND2HSV0 U48585 ( .A1(n48396), .A2(\pe1/bq[18] ), .ZN(n44550) );
  XOR2HSV0 U48586 ( .A1(n44551), .A2(n44550), .Z(n44552) );
  XOR2HSV0 U48587 ( .A1(n44553), .A2(n44552), .Z(n44562) );
  NAND2HSV0 U48588 ( .A1(n59992), .A2(n40733), .ZN(n44555) );
  NAND2HSV0 U48589 ( .A1(n54188), .A2(n41644), .ZN(n44554) );
  XOR2HSV0 U48590 ( .A1(n44555), .A2(n44554), .Z(n44560) );
  NAND2HSV0 U48591 ( .A1(n44556), .A2(n54836), .ZN(n44558) );
  NAND2HSV0 U48592 ( .A1(n53717), .A2(n53718), .ZN(n44557) );
  XOR2HSV0 U48593 ( .A1(n44558), .A2(n44557), .Z(n44559) );
  XOR2HSV0 U48594 ( .A1(n44560), .A2(n44559), .Z(n44561) );
  XOR2HSV0 U48595 ( .A1(n44562), .A2(n44561), .Z(n44563) );
  XOR3HSV2 U48596 ( .A1(n44565), .A2(n44564), .A3(n44563), .Z(n44599) );
  NAND2HSV0 U48597 ( .A1(n53673), .A2(\pe1/bq[4] ), .ZN(n44568) );
  CLKNHSV0 U48598 ( .I(n54399), .ZN(n54668) );
  NAND2HSV0 U48599 ( .A1(n44566), .A2(n54668), .ZN(n44567) );
  XOR2HSV0 U48600 ( .A1(n44568), .A2(n44567), .Z(n44573) );
  NAND2HSV0 U48601 ( .A1(\pe1/aot [16]), .A2(n42092), .ZN(n44571) );
  NAND2HSV0 U48602 ( .A1(n44569), .A2(n55231), .ZN(n44570) );
  XOR2HSV0 U48603 ( .A1(n44571), .A2(n44570), .Z(n44572) );
  XOR2HSV0 U48604 ( .A1(n44573), .A2(n44572), .Z(n44581) );
  NAND2HSV0 U48605 ( .A1(n54293), .A2(\pe1/bq[9] ), .ZN(n44575) );
  INHSV2 U48606 ( .I(n55515), .ZN(n59389) );
  NAND2HSV0 U48607 ( .A1(n59389), .A2(n40890), .ZN(n44574) );
  XOR2HSV0 U48608 ( .A1(n44575), .A2(n44574), .Z(n44579) );
  NAND2HSV0 U48609 ( .A1(n40683), .A2(n55394), .ZN(n44577) );
  NAND2HSV0 U48610 ( .A1(n54303), .A2(n53411), .ZN(n44576) );
  XOR2HSV0 U48611 ( .A1(n44577), .A2(n44576), .Z(n44578) );
  XOR2HSV0 U48612 ( .A1(n44579), .A2(n44578), .Z(n44580) );
  XOR2HSV0 U48613 ( .A1(n44581), .A2(n44580), .Z(n44597) );
  CLKNAND2HSV0 U48614 ( .A1(n42132), .A2(n54565), .ZN(n44583) );
  NAND2HSV0 U48615 ( .A1(n59985), .A2(n54289), .ZN(n44582) );
  XOR2HSV0 U48616 ( .A1(n44583), .A2(n44582), .Z(n44587) );
  NAND2HSV0 U48617 ( .A1(\pe1/aot [7]), .A2(n53805), .ZN(n44585) );
  NAND2HSV0 U48618 ( .A1(n59619), .A2(n48055), .ZN(n44584) );
  XOR2HSV0 U48619 ( .A1(n44585), .A2(n44584), .Z(n44586) );
  XOR2HSV0 U48620 ( .A1(n44587), .A2(n44586), .Z(n44595) );
  NAND2HSV0 U48621 ( .A1(n53936), .A2(n53578), .ZN(n44589) );
  NAND2HSV0 U48622 ( .A1(n54904), .A2(n40494), .ZN(n44588) );
  XOR2HSV0 U48623 ( .A1(n44589), .A2(n44588), .Z(n44593) );
  NOR2HSV0 U48624 ( .A1(n46142), .A2(n53691), .ZN(n44591) );
  BUFHSV2 U48625 ( .I(\pe1/bq[8] ), .Z(n53798) );
  NAND2HSV0 U48626 ( .A1(\pe1/aot [27]), .A2(n53798), .ZN(n44590) );
  XOR2HSV0 U48627 ( .A1(n44591), .A2(n44590), .Z(n44592) );
  XOR2HSV0 U48628 ( .A1(n44593), .A2(n44592), .Z(n44594) );
  XOR2HSV0 U48629 ( .A1(n44595), .A2(n44594), .Z(n44596) );
  XOR2HSV0 U48630 ( .A1(n44597), .A2(n44596), .Z(n44598) );
  XNOR2HSV1 U48631 ( .A1(n44599), .A2(n44598), .ZN(n44600) );
  XOR3HSV2 U48632 ( .A1(n44602), .A2(n44601), .A3(n44600), .Z(n44603) );
  XNOR2HSV1 U48633 ( .A1(n44604), .A2(n44603), .ZN(n44607) );
  NAND2HSV0 U48634 ( .A1(n40917), .A2(n44605), .ZN(n44606) );
  XOR2HSV0 U48635 ( .A1(n44607), .A2(n44606), .Z(n44609) );
  NAND2HSV0 U48636 ( .A1(n59919), .A2(n53473), .ZN(n44608) );
  XOR2HSV0 U48637 ( .A1(n44609), .A2(n44608), .Z(n44610) );
  XNOR2HSV1 U48638 ( .A1(n44611), .A2(n44610), .ZN(n44613) );
  NAND2HSV0 U48639 ( .A1(n29763), .A2(n55337), .ZN(n44612) );
  XOR2HSV0 U48640 ( .A1(n44613), .A2(n44612), .Z(n44614) );
  XNOR2HSV1 U48641 ( .A1(n44615), .A2(n44614), .ZN(n44617) );
  NAND2HSV0 U48642 ( .A1(n54115), .A2(\pe1/got [14]), .ZN(n44616) );
  XOR2HSV0 U48643 ( .A1(n44617), .A2(n44616), .Z(n44618) );
  XNOR2HSV1 U48644 ( .A1(n44619), .A2(n44618), .ZN(n44620) );
  XNOR2HSV1 U48645 ( .A1(n44621), .A2(n44620), .ZN(n44623) );
  NOR2HSV0 U48646 ( .A1(n41312), .A2(n54248), .ZN(n44622) );
  XOR3HSV2 U48647 ( .A1(n44624), .A2(n44623), .A3(n44622), .Z(n44625) );
  XNOR2HSV1 U48648 ( .A1(n44626), .A2(n44625), .ZN(n44627) );
  XNOR2HSV1 U48649 ( .A1(n44628), .A2(n44627), .ZN(n44629) );
  XNOR2HSV1 U48650 ( .A1(n44630), .A2(n44629), .ZN(n44631) );
  XNOR2HSV1 U48651 ( .A1(n44632), .A2(n44631), .ZN(n44633) );
  XNOR2HSV1 U48652 ( .A1(n44634), .A2(n44633), .ZN(n44636) );
  CLKNAND2HSV1 U48653 ( .A1(n53768), .A2(n53520), .ZN(n44635) );
  XOR2HSV0 U48654 ( .A1(n44636), .A2(n44635), .Z(n44637) );
  XOR2HSV0 U48655 ( .A1(n44638), .A2(n44637), .Z(n44641) );
  CLKNAND2HSV1 U48656 ( .A1(n48336), .A2(n41689), .ZN(n44640) );
  NOR2HSV2 U48657 ( .A1(n55144), .A2(n44337), .ZN(n44639) );
  XOR3HSV2 U48658 ( .A1(n44641), .A2(n44640), .A3(n44639), .Z(n44642) );
  CLKNAND2HSV1 U48659 ( .A1(n44643), .A2(n44644), .ZN(n44648) );
  CLKNHSV1 U48660 ( .I(n44643), .ZN(n44646) );
  CLKNHSV0 U48661 ( .I(n45781), .ZN(n48332) );
  INHSV2 U48662 ( .I(n44652), .ZN(n44655) );
  INOR2HSV1 U48663 ( .A1(n41418), .B1(n41701), .ZN(n44653) );
  CLKNAND2HSV1 U48664 ( .A1(n48314), .A2(n44653), .ZN(n44654) );
  INHSV3 U48665 ( .I(n44656), .ZN(n44659) );
  INHSV2 U48666 ( .I(n44657), .ZN(n44658) );
  CLKNAND2HSV3 U48667 ( .A1(n44659), .A2(n44658), .ZN(n44660) );
  NAND2HSV2 U48668 ( .A1(n25448), .A2(\pe1/ti_7t [30]), .ZN(n53511) );
  CLKBUFHSV4 U48669 ( .I(n54553), .Z(n59428) );
  INHSV2 U48670 ( .I(n55019), .ZN(n59750) );
  CLKNHSV2 U48671 ( .I(\pe1/got [1]), .ZN(n53978) );
  INHSV2 U48672 ( .I(n53978), .ZN(n59755) );
  INHSV2 U48673 ( .I(n44674), .ZN(n44670) );
  CLKNAND2HSV1 U48674 ( .A1(n42815), .A2(n44680), .ZN(n44682) );
  XNOR2HSV4 U48675 ( .A1(n44684), .A2(n44683), .ZN(n45617) );
  NAND3HSV3 U48676 ( .A1(n45617), .A2(n44687), .A3(n44686), .ZN(n44688) );
  INHSV2 U48677 ( .I(n50199), .ZN(n47920) );
  INHSV2 U48678 ( .I(n44832), .ZN(n51121) );
  BUFHSV2 U48679 ( .I(n56265), .Z(n59920) );
  BUFHSV2 U48680 ( .I(n44695), .Z(n59378) );
  BUFHSV2 U48681 ( .I(n44696), .Z(n59725) );
  BUFHSV2 U48682 ( .I(n52367), .Z(n59766) );
  MUX2HSV1 U48683 ( .I0(bo3[27]), .I1(n44698), .S(n46612), .Z(n59765) );
  MUX2HSV1 U48684 ( .I0(bo2[30]), .I1(n36475), .S(n53014), .Z(n59724) );
  BUFHSV2 U48685 ( .I(n48036), .Z(n53214) );
  MUX2HSV1 U48686 ( .I0(bo6[22]), .I1(n44700), .S(n48046), .Z(n59884) );
  BUFHSV2 U48687 ( .I(\pe5/bq[4] ), .Z(n51336) );
  MUX2HSV1 U48688 ( .I0(bo5[4]), .I1(n51336), .S(n48034), .Z(n59543) );
  BUFHSV2 U48689 ( .I(n48039), .Z(n48045) );
  MUX2HSV1 U48690 ( .I0(bo5[27]), .I1(n48787), .S(n48045), .Z(n59841) );
  BUFHSV2 U48691 ( .I(n46623), .Z(n48065) );
  MUX2HSV1 U48692 ( .I0(bo2[19]), .I1(n43961), .S(n48065), .Z(n59563) );
  INHSV2 U48693 ( .I(n55524), .ZN(n59373) );
  MUX2HSV1 U48694 ( .I0(bo1[23]), .I1(\pe1/bq[23] ), .S(n48061), .Z(n59698) );
  MUX2HSV1 U48695 ( .I0(bo6[17]), .I1(n32982), .S(n44701), .Z(n59890) );
  MUX2HSV1 U48696 ( .I0(bo6[18]), .I1(n36150), .S(n48025), .Z(n59885) );
  CLKNHSV0 U48697 ( .I(n45451), .ZN(n59941) );
  MUX2HSV1 U48698 ( .I0(bo6[19]), .I1(n50829), .S(n44701), .Z(n59889) );
  MUX2HSV1 U48699 ( .I0(bo6[23]), .I1(n44702), .S(n48025), .Z(n59887) );
  MUX2HSV1 U48700 ( .I0(bo1[15]), .I1(\pe1/bq[15] ), .S(n48061), .Z(n59706) );
  MUX2HSV1 U48701 ( .I0(bo1[17]), .I1(n42098), .S(n48076), .Z(n59703) );
  INHSV2 U48702 ( .I(n53032), .ZN(n59351) );
  MUX2HSV1 U48703 ( .I0(bo1[21]), .I1(\pe1/bq[21] ), .S(n48054), .Z(n59699) );
  CLKNHSV0 U48704 ( .I(n44704), .ZN(n59940) );
  CLKNHSV0 U48705 ( .I(n44705), .ZN(n59737) );
  CLKNHSV0 U48706 ( .I(n36623), .ZN(n44710) );
  INAND2HSV2 U48707 ( .A1(n44710), .B1(n52920), .ZN(n44816) );
  NOR2HSV0 U48708 ( .A1(n44833), .A2(n52285), .ZN(n44814) );
  NAND2HSV2 U48709 ( .A1(n59775), .A2(n44711), .ZN(n44811) );
  BUFHSV2 U48710 ( .I(n52924), .Z(n44970) );
  INHSV2 U48711 ( .I(n38275), .ZN(n53077) );
  NAND2HSV2 U48712 ( .A1(n44970), .A2(n53077), .ZN(n44806) );
  NAND2HSV0 U48713 ( .A1(n49591), .A2(n51801), .ZN(n44804) );
  CLKNAND2HSV1 U48714 ( .A1(n59634), .A2(n59982), .ZN(n44799) );
  CLKNAND2HSV0 U48715 ( .A1(n44713), .A2(n44712), .ZN(n44797) );
  NAND2HSV0 U48716 ( .A1(n51796), .A2(n52929), .ZN(n44795) );
  CLKNAND2HSV0 U48717 ( .A1(n52287), .A2(n45289), .ZN(n44792) );
  CLKNAND2HSV0 U48718 ( .A1(n52932), .A2(n52172), .ZN(n44786) );
  CLKNAND2HSV0 U48719 ( .A1(n52934), .A2(n52374), .ZN(n44784) );
  NAND2HSV0 U48720 ( .A1(n44715), .A2(n44714), .ZN(n44779) );
  CLKNAND2HSV0 U48721 ( .A1(n59684), .A2(\pe2/got [8]), .ZN(n44717) );
  NOR2HSV0 U48722 ( .A1(n44971), .A2(n50928), .ZN(n44716) );
  XNOR2HSV1 U48723 ( .A1(n44717), .A2(n44716), .ZN(n44777) );
  NAND2HSV0 U48724 ( .A1(n44976), .A2(\pe2/bq[6] ), .ZN(n44720) );
  NAND2HSV0 U48725 ( .A1(\pe2/aot [19]), .A2(n52988), .ZN(n44719) );
  XOR2HSV0 U48726 ( .A1(n44720), .A2(n44719), .Z(n44724) );
  NAND2HSV0 U48727 ( .A1(\pe2/aot [12]), .A2(n44987), .ZN(n44722) );
  CLKNAND2HSV0 U48728 ( .A1(\pe2/aot [15]), .A2(n45033), .ZN(n44721) );
  XOR2HSV0 U48729 ( .A1(n44722), .A2(n44721), .Z(n44723) );
  XOR2HSV0 U48730 ( .A1(n44724), .A2(n44723), .Z(n44742) );
  CLKNHSV0 U48731 ( .I(n49628), .ZN(n47598) );
  CLKNAND2HSV1 U48732 ( .A1(n38479), .A2(n47598), .ZN(n44726) );
  NAND2HSV0 U48733 ( .A1(n53015), .A2(\pe2/aot [5]), .ZN(n44725) );
  XOR2HSV0 U48734 ( .A1(n44726), .A2(n44725), .Z(n44728) );
  XNOR2HSV1 U48735 ( .A1(n44728), .A2(n44727), .ZN(n44732) );
  NOR2HSV0 U48736 ( .A1(n47575), .A2(n51567), .ZN(n45191) );
  NOR2HSV0 U48737 ( .A1(n47524), .A2(n49518), .ZN(n52097) );
  XOR2HSV0 U48738 ( .A1(n44730), .A2(n52097), .Z(n44731) );
  XNOR2HSV1 U48739 ( .A1(n44732), .A2(n44731), .ZN(n44741) );
  NOR2HSV0 U48740 ( .A1(n47574), .A2(n47580), .ZN(n44734) );
  NAND2HSV0 U48741 ( .A1(n39052), .A2(\pe2/bq[17] ), .ZN(n44733) );
  XOR2HSV0 U48742 ( .A1(n44734), .A2(n44733), .Z(n44738) );
  NAND2HSV0 U48743 ( .A1(\pe2/aot [17]), .A2(n52965), .ZN(n44736) );
  CLKNAND2HSV0 U48744 ( .A1(n52955), .A2(n43961), .ZN(n44735) );
  XOR2HSV0 U48745 ( .A1(n44736), .A2(n44735), .Z(n44737) );
  XOR2HSV0 U48746 ( .A1(n44738), .A2(n44737), .Z(n44740) );
  CLKNAND2HSV0 U48747 ( .A1(n36409), .A2(n53041), .ZN(n44739) );
  XOR4HSV1 U48748 ( .A1(n44742), .A2(n44741), .A3(n44740), .A4(n44739), .Z(
        n44775) );
  NAND2HSV0 U48749 ( .A1(n45024), .A2(\pe2/bq[21] ), .ZN(n44744) );
  CLKNHSV0 U48750 ( .I(n50908), .ZN(n53038) );
  NAND2HSV0 U48751 ( .A1(n53038), .A2(n45008), .ZN(n44743) );
  XOR2HSV0 U48752 ( .A1(n44744), .A2(n44743), .Z(n44749) );
  NAND2HSV0 U48753 ( .A1(n51636), .A2(n36607), .ZN(n44747) );
  NAND2HSV0 U48754 ( .A1(n44745), .A2(n52300), .ZN(n44746) );
  XOR2HSV0 U48755 ( .A1(n44747), .A2(n44746), .Z(n44748) );
  XOR2HSV0 U48756 ( .A1(n44749), .A2(n44748), .Z(n44758) );
  NAND2HSV0 U48757 ( .A1(n52974), .A2(n52073), .ZN(n44752) );
  CLKNHSV0 U48758 ( .I(n51131), .ZN(n52994) );
  NAND2HSV0 U48759 ( .A1(n44750), .A2(n52994), .ZN(n44751) );
  XOR2HSV0 U48760 ( .A1(n44752), .A2(n44751), .Z(n44756) );
  NAND2HSV0 U48761 ( .A1(n45034), .A2(n45015), .ZN(n44754) );
  CLKNHSV0 U48762 ( .I(n47511), .ZN(n52322) );
  NAND2HSV0 U48763 ( .A1(n44081), .A2(n52322), .ZN(n44753) );
  XOR2HSV0 U48764 ( .A1(n44754), .A2(n44753), .Z(n44755) );
  XOR2HSV0 U48765 ( .A1(n44756), .A2(n44755), .Z(n44757) );
  XOR2HSV0 U48766 ( .A1(n44758), .A2(n44757), .Z(n44773) );
  NAND2HSV0 U48767 ( .A1(n52457), .A2(n44759), .ZN(n44761) );
  NAND2HSV0 U48768 ( .A1(n59633), .A2(n36475), .ZN(n44760) );
  XOR2HSV0 U48769 ( .A1(n44761), .A2(n44760), .Z(n44765) );
  NAND2HSV0 U48770 ( .A1(n53009), .A2(n52973), .ZN(n44763) );
  NAND2HSV0 U48771 ( .A1(n59768), .A2(n38565), .ZN(n44762) );
  XOR2HSV0 U48772 ( .A1(n44763), .A2(n44762), .Z(n44764) );
  XOR2HSV0 U48773 ( .A1(n44765), .A2(n44764), .Z(n44771) );
  NOR2HSV0 U48774 ( .A1(n44871), .A2(n48066), .ZN(n52217) );
  NAND2HSV0 U48775 ( .A1(\pe2/aot [25]), .A2(n53006), .ZN(n52293) );
  XOR2HSV0 U48776 ( .A1(n52217), .A2(n52293), .Z(n44769) );
  NAND2HSV0 U48777 ( .A1(n45295), .A2(n52448), .ZN(n44766) );
  XOR2HSV0 U48778 ( .A1(n44767), .A2(n44766), .Z(n44768) );
  XOR2HSV0 U48779 ( .A1(n44769), .A2(n44768), .Z(n44770) );
  XOR2HSV0 U48780 ( .A1(n44771), .A2(n44770), .Z(n44772) );
  XOR2HSV0 U48781 ( .A1(n44773), .A2(n44772), .Z(n44774) );
  XNOR2HSV1 U48782 ( .A1(n44775), .A2(n44774), .ZN(n44776) );
  XNOR2HSV1 U48783 ( .A1(n44777), .A2(n44776), .ZN(n44778) );
  XNOR2HSV1 U48784 ( .A1(n44779), .A2(n44778), .ZN(n44782) );
  NAND2HSV0 U48785 ( .A1(n59679), .A2(\pe2/got [10]), .ZN(n44781) );
  XNOR2HSV1 U48786 ( .A1(n44782), .A2(n44781), .ZN(n44783) );
  XNOR2HSV1 U48787 ( .A1(n44784), .A2(n44783), .ZN(n44785) );
  XNOR2HSV1 U48788 ( .A1(n44786), .A2(n44785), .ZN(n44788) );
  CLKNHSV0 U48789 ( .I(n51607), .ZN(n45058) );
  NAND2HSV0 U48790 ( .A1(n45055), .A2(n45058), .ZN(n44787) );
  XOR2HSV0 U48791 ( .A1(n44788), .A2(n44787), .Z(n44790) );
  INHSV2 U48792 ( .I(n47498), .ZN(n51608) );
  CLKNAND2HSV0 U48793 ( .A1(n53050), .A2(n51608), .ZN(n44789) );
  XNOR2HSV1 U48794 ( .A1(n44790), .A2(n44789), .ZN(n44791) );
  XNOR2HSV1 U48795 ( .A1(n44792), .A2(n44791), .ZN(n44794) );
  CLKNAND2HSV0 U48796 ( .A1(n45063), .A2(n38782), .ZN(n44793) );
  XOR3HSV2 U48797 ( .A1(n44795), .A2(n44794), .A3(n44793), .Z(n44796) );
  XNOR2HSV1 U48798 ( .A1(n44797), .A2(n44796), .ZN(n44798) );
  XNOR2HSV1 U48799 ( .A1(n44799), .A2(n44798), .ZN(n44801) );
  NAND2HSV0 U48800 ( .A1(n52251), .A2(n52167), .ZN(n44800) );
  XOR3HSV2 U48801 ( .A1(n44802), .A2(n44801), .A3(n44800), .Z(n44803) );
  XNOR2HSV1 U48802 ( .A1(n44804), .A2(n44803), .ZN(n44805) );
  XNOR2HSV1 U48803 ( .A1(n44806), .A2(n44805), .ZN(n44809) );
  NAND2HSV0 U48804 ( .A1(n44807), .A2(n52416), .ZN(n44808) );
  XNOR2HSV1 U48805 ( .A1(n44809), .A2(n44808), .ZN(n44810) );
  CLKNAND2HSV0 U48806 ( .A1(n59774), .A2(n44944), .ZN(n44812) );
  XOR3HSV2 U48807 ( .A1(n44814), .A2(n44813), .A3(n44812), .Z(n44815) );
  NAND2HSV2 U48808 ( .A1(n44817), .A2(n59635), .ZN(n44818) );
  XNOR2HSV4 U48809 ( .A1(n44819), .A2(n44818), .ZN(n45119) );
  XNOR2HSV4 U48810 ( .A1(n45119), .A2(n44820), .ZN(n44826) );
  INAND2HSV2 U48811 ( .A1(n44827), .B1(n44826), .ZN(n45273) );
  CLKAND2HSV4 U48812 ( .A1(n45274), .A2(n29633), .Z(n44830) );
  CLKNAND2HSV1 U48813 ( .A1(n44829), .A2(n44828), .ZN(n45275) );
  NAND2HSV2 U48814 ( .A1(\pe2/ti_7t [28]), .A2(n38454), .ZN(n45277) );
  INHSV2 U48815 ( .I(n52285), .ZN(n53086) );
  NAND2HSV2 U48816 ( .A1(n52920), .A2(n53086), .ZN(n44942) );
  NOR2HSV1 U48817 ( .A1(n47500), .A2(n38205), .ZN(n44940) );
  CLKNAND2HSV0 U48818 ( .A1(n51687), .A2(n53077), .ZN(n44937) );
  INHSV2 U48819 ( .I(n44834), .ZN(n52814) );
  NAND2HSV2 U48820 ( .A1(n38390), .A2(n52814), .ZN(n44932) );
  CLKNAND2HSV1 U48821 ( .A1(n52286), .A2(n52925), .ZN(n44930) );
  NAND2HSV0 U48822 ( .A1(n45288), .A2(n38782), .ZN(n44927) );
  CLKNHSV1 U48823 ( .I(n45148), .ZN(n52928) );
  CLKNAND2HSV1 U48824 ( .A1(n52928), .A2(\pe2/got [16]), .ZN(n44925) );
  NAND2HSV0 U48825 ( .A1(n51608), .A2(n52929), .ZN(n44923) );
  NAND2HSV2 U48826 ( .A1(n52287), .A2(n45058), .ZN(n44920) );
  NAND2HSV2 U48827 ( .A1(n44185), .A2(\pe2/got [10]), .ZN(n44914) );
  BUFHSV2 U48828 ( .I(n44835), .Z(n49494) );
  NAND2HSV0 U48829 ( .A1(n52053), .A2(\pe2/got [9]), .ZN(n44912) );
  CLKNAND2HSV1 U48830 ( .A1(n44046), .A2(n53041), .ZN(n44837) );
  NOR2HSV0 U48831 ( .A1(n53033), .A2(n50908), .ZN(n44836) );
  XOR2HSV0 U48832 ( .A1(n44837), .A2(n44836), .Z(n44905) );
  NAND2HSV0 U48833 ( .A1(n59768), .A2(\pe2/bq[26] ), .ZN(n44839) );
  NAND2HSV0 U48834 ( .A1(n52456), .A2(n36608), .ZN(n44838) );
  XOR2HSV0 U48835 ( .A1(n44839), .A2(n44838), .Z(n44843) );
  NOR2HSV0 U48836 ( .A1(n45165), .A2(n47608), .ZN(n44841) );
  NAND2HSV0 U48837 ( .A1(n59758), .A2(\pe2/bq[14] ), .ZN(n44840) );
  XOR2HSV0 U48838 ( .A1(n44841), .A2(n44840), .Z(n44842) );
  XOR2HSV0 U48839 ( .A1(n44843), .A2(n44842), .Z(n44851) );
  NOR2HSV0 U48840 ( .A1(n38946), .A2(n44844), .ZN(n45297) );
  NOR2HSV0 U48841 ( .A1(n52103), .A2(n48064), .ZN(n45029) );
  AOI22HSV0 U48842 ( .A1(n51639), .A2(\pe2/bq[17] ), .B1(n52988), .B2(n51759), 
        .ZN(n44845) );
  AOI21HSV1 U48843 ( .A1(n45297), .A2(n45029), .B(n44845), .ZN(n44846) );
  NAND2HSV0 U48844 ( .A1(n45034), .A2(n45033), .ZN(n52433) );
  XNOR2HSV1 U48845 ( .A1(n44846), .A2(n52433), .ZN(n44849) );
  INHSV2 U48846 ( .I(n51538), .ZN(n52867) );
  NAND2HSV0 U48847 ( .A1(n52867), .A2(n53015), .ZN(n45332) );
  NAND2HSV0 U48848 ( .A1(n59973), .A2(\pe2/bq[19] ), .ZN(n44847) );
  XOR2HSV0 U48849 ( .A1(n45332), .A2(n44847), .Z(n44848) );
  XNOR2HSV1 U48850 ( .A1(n44849), .A2(n44848), .ZN(n44850) );
  XOR2HSV0 U48851 ( .A1(n44851), .A2(n44850), .Z(n44903) );
  CLKNAND2HSV0 U48852 ( .A1(n53005), .A2(n52300), .ZN(n44853) );
  NAND2HSV0 U48853 ( .A1(n39052), .A2(n52337), .ZN(n44852) );
  XOR2HSV0 U48854 ( .A1(n44853), .A2(n44852), .Z(n44858) );
  NAND2HSV0 U48855 ( .A1(n59976), .A2(\pe2/bq[24] ), .ZN(n44856) );
  NAND2HSV0 U48856 ( .A1(n53009), .A2(n44987), .ZN(n44855) );
  XOR2HSV0 U48857 ( .A1(n44856), .A2(n44855), .Z(n44857) );
  XOR2HSV0 U48858 ( .A1(n44858), .A2(n44857), .Z(n44866) );
  NAND2HSV0 U48859 ( .A1(n59633), .A2(\pe2/bq[28] ), .ZN(n44860) );
  NAND2HSV0 U48860 ( .A1(\pe2/aot [23]), .A2(n53006), .ZN(n44859) );
  XOR2HSV0 U48861 ( .A1(n44860), .A2(n44859), .Z(n44864) );
  NAND2HSV0 U48862 ( .A1(n38393), .A2(\pe2/aot [5]), .ZN(n44862) );
  NAND2HSV0 U48863 ( .A1(n52485), .A2(\pe2/bq[6] ), .ZN(n44861) );
  XOR2HSV0 U48864 ( .A1(n44862), .A2(n44861), .Z(n44863) );
  XNOR2HSV1 U48865 ( .A1(n44864), .A2(n44863), .ZN(n44865) );
  XNOR2HSV1 U48866 ( .A1(n44866), .A2(n44865), .ZN(n44868) );
  NAND2HSV0 U48867 ( .A1(n36409), .A2(n59984), .ZN(n44867) );
  XNOR2HSV1 U48868 ( .A1(n44868), .A2(n44867), .ZN(n44902) );
  CLKNAND2HSV0 U48869 ( .A1(n38479), .A2(n51900), .ZN(n44870) );
  NAND2HSV0 U48870 ( .A1(n59969), .A2(n52994), .ZN(n44869) );
  XOR2HSV0 U48871 ( .A1(n44870), .A2(n44869), .Z(n44875) );
  CLKNAND2HSV0 U48872 ( .A1(n37801), .A2(n47598), .ZN(n44873) );
  NAND2HSV0 U48873 ( .A1(n52457), .A2(n39032), .ZN(n44872) );
  XOR2HSV0 U48874 ( .A1(n44873), .A2(n44872), .Z(n44874) );
  XOR2HSV0 U48875 ( .A1(n44875), .A2(n44874), .Z(n44883) );
  INHSV2 U48876 ( .I(n51537), .ZN(n52993) );
  NAND2HSV0 U48877 ( .A1(n52993), .A2(n52444), .ZN(n44877) );
  NAND2HSV2 U48878 ( .A1(n59351), .A2(n45303), .ZN(n44876) );
  XOR2HSV0 U48879 ( .A1(n44877), .A2(n44876), .Z(n44881) );
  NOR2HSV0 U48880 ( .A1(n47503), .A2(n47599), .ZN(n44879) );
  NAND2HSV0 U48881 ( .A1(\pe2/aot [19]), .A2(n51732), .ZN(n44878) );
  XOR2HSV0 U48882 ( .A1(n44879), .A2(n44878), .Z(n44880) );
  XOR2HSV0 U48883 ( .A1(n44881), .A2(n44880), .Z(n44882) );
  XOR2HSV0 U48884 ( .A1(n44883), .A2(n44882), .Z(n44900) );
  INHSV2 U48885 ( .I(n44884), .ZN(n59497) );
  NAND2HSV0 U48886 ( .A1(n59497), .A2(\pe2/pvq [30]), .ZN(n44885) );
  XNOR2HSV1 U48887 ( .A1(n44885), .A2(\pe2/phq [30]), .ZN(n44888) );
  NOR2HSV0 U48888 ( .A1(n44049), .A2(n51567), .ZN(n45298) );
  NOR2HSV0 U48889 ( .A1(n44095), .A2(n47511), .ZN(n45030) );
  AOI22HSV0 U48890 ( .A1(n52974), .A2(n51623), .B1(n49530), .B2(n51825), .ZN(
        n44886) );
  AOI21HSV1 U48891 ( .A1(n45298), .A2(n45030), .B(n44886), .ZN(n44887) );
  XOR2HSV0 U48892 ( .A1(n44888), .A2(n44887), .Z(n44898) );
  NOR2HSV0 U48893 ( .A1(n44889), .A2(n48621), .ZN(n45293) );
  NOR2HSV0 U48894 ( .A1(n37940), .A2(n49529), .ZN(n44891) );
  NAND2HSV0 U48895 ( .A1(n52995), .A2(n51803), .ZN(n52490) );
  OAI22HSV1 U48896 ( .A1(n45293), .A2(n44891), .B1(n44890), .B2(n52490), .ZN(
        n44896) );
  NAND2HSV0 U48897 ( .A1(n52998), .A2(\pe2/bq[3] ), .ZN(n49540) );
  NOR2HSV0 U48898 ( .A1(n45294), .A2(n49540), .ZN(n44894) );
  INHSV2 U48899 ( .I(n49515), .ZN(n52448) );
  AOI22HSV0 U48900 ( .A1(n44892), .A2(n52905), .B1(n52998), .B2(n52448), .ZN(
        n44893) );
  NOR2HSV1 U48901 ( .A1(n44894), .A2(n44893), .ZN(n44895) );
  XOR2HSV0 U48902 ( .A1(n44896), .A2(n44895), .Z(n44897) );
  XNOR2HSV1 U48903 ( .A1(n44898), .A2(n44897), .ZN(n44899) );
  XNOR2HSV1 U48904 ( .A1(n44900), .A2(n44899), .ZN(n44901) );
  XOR3HSV2 U48905 ( .A1(n44903), .A2(n44902), .A3(n44901), .Z(n44904) );
  XNOR2HSV1 U48906 ( .A1(n44905), .A2(n44904), .ZN(n44908) );
  BUFHSV2 U48907 ( .I(n44906), .Z(n59669) );
  NAND2HSV0 U48908 ( .A1(n59669), .A2(n59757), .ZN(n44907) );
  XOR2HSV0 U48909 ( .A1(n44908), .A2(n44907), .Z(n44910) );
  NAND2HSV2 U48910 ( .A1(n59679), .A2(\pe2/got [8]), .ZN(n44909) );
  XNOR2HSV1 U48911 ( .A1(n44910), .A2(n44909), .ZN(n44911) );
  XNOR2HSV1 U48912 ( .A1(n44912), .A2(n44911), .ZN(n44913) );
  XNOR2HSV1 U48913 ( .A1(n44914), .A2(n44913), .ZN(n44916) );
  NAND2HSV0 U48914 ( .A1(n45055), .A2(n52374), .ZN(n44915) );
  XOR2HSV0 U48915 ( .A1(n44916), .A2(n44915), .Z(n44918) );
  NAND2HSV0 U48916 ( .A1(n53050), .A2(n52172), .ZN(n44917) );
  XNOR2HSV1 U48917 ( .A1(n44918), .A2(n44917), .ZN(n44919) );
  XNOR2HSV1 U48918 ( .A1(n44920), .A2(n44919), .ZN(n44922) );
  BUFHSV2 U48919 ( .I(n51610), .Z(n59761) );
  BUFHSV2 U48920 ( .I(n59761), .Z(n53056) );
  NAND2HSV2 U48921 ( .A1(n53056), .A2(n45289), .ZN(n44921) );
  XOR3HSV2 U48922 ( .A1(n44923), .A2(n44922), .A3(n44921), .Z(n44924) );
  XNOR2HSV1 U48923 ( .A1(n44925), .A2(n44924), .ZN(n44926) );
  XNOR2HSV1 U48924 ( .A1(n44927), .A2(n44926), .ZN(n44929) );
  NOR2HSV0 U48925 ( .A1(n45071), .A2(n47570), .ZN(n44928) );
  XOR3HSV2 U48926 ( .A1(n44930), .A2(n44929), .A3(n44928), .Z(n44931) );
  XNOR2HSV1 U48927 ( .A1(n44932), .A2(n44931), .ZN(n44935) );
  CLKNAND2HSV1 U48928 ( .A1(n44970), .A2(n52922), .ZN(n44934) );
  CLKNAND2HSV0 U48929 ( .A1(n59361), .A2(n45287), .ZN(n44933) );
  XOR3HSV2 U48930 ( .A1(n44935), .A2(n44934), .A3(n44933), .Z(n44936) );
  XNOR2HSV1 U48931 ( .A1(n44937), .A2(n44936), .ZN(n44939) );
  NAND2HSV2 U48932 ( .A1(n59774), .A2(n44711), .ZN(n44938) );
  XOR3HSV2 U48933 ( .A1(n44940), .A2(n44939), .A3(n44938), .Z(n44941) );
  XNOR2HSV1 U48934 ( .A1(n44942), .A2(n44941), .ZN(n44946) );
  INHSV4 U48935 ( .I(n44943), .ZN(n47572) );
  NAND2HSV2 U48936 ( .A1(n47572), .A2(n44944), .ZN(n44945) );
  XNOR2HSV1 U48937 ( .A1(n44946), .A2(n44945), .ZN(n44948) );
  CLKNAND2HSV2 U48938 ( .A1(n25825), .A2(n36623), .ZN(n44947) );
  NAND2HSV2 U48939 ( .A1(n45286), .A2(n59635), .ZN(n44950) );
  XNOR2HSV4 U48940 ( .A1(n44951), .A2(n44950), .ZN(n45401) );
  NAND2HSV2 U48941 ( .A1(n44954), .A2(n44953), .ZN(n44966) );
  INHSV4 U48942 ( .I(n25825), .ZN(n47499) );
  CLKNHSV0 U48943 ( .I(n44959), .ZN(n44963) );
  AND2HSV2 U48944 ( .A1(n44960), .A2(n53094), .Z(n44961) );
  INAND2HSV2 U48945 ( .A1(n44969), .B1(n44968), .ZN(n45088) );
  NOR2HSV2 U48946 ( .A1(n47500), .A2(n39088), .ZN(n45086) );
  CLKNAND2HSV1 U48947 ( .A1(n44970), .A2(n45287), .ZN(n45078) );
  NAND2HSV1 U48948 ( .A1(n52922), .A2(n59506), .ZN(n45076) );
  CLKNAND2HSV1 U48949 ( .A1(n52286), .A2(n59982), .ZN(n45074) );
  NAND2HSV0 U48950 ( .A1(n45288), .A2(n52925), .ZN(n45070) );
  CLKNAND2HSV1 U48951 ( .A1(n52928), .A2(n38782), .ZN(n45068) );
  NAND2HSV0 U48952 ( .A1(n45289), .A2(n52419), .ZN(n45066) );
  NAND2HSV0 U48953 ( .A1(n52931), .A2(n51608), .ZN(n45062) );
  NAND2HSV0 U48954 ( .A1(n52932), .A2(n52374), .ZN(n45054) );
  NAND2HSV0 U48955 ( .A1(n52288), .A2(\pe2/got [10]), .ZN(n45052) );
  NAND2HSV0 U48956 ( .A1(n59669), .A2(\pe2/got [8]), .ZN(n45048) );
  CLKNHSV0 U48957 ( .I(n50928), .ZN(n52174) );
  CLKNAND2HSV1 U48958 ( .A1(n59684), .A2(n52174), .ZN(n44973) );
  NOR2HSV0 U48959 ( .A1(n44971), .A2(n52018), .ZN(n44972) );
  XOR2HSV0 U48960 ( .A1(n44973), .A2(n44972), .Z(n45046) );
  NAND2HSV0 U48961 ( .A1(n39052), .A2(n52984), .ZN(n44975) );
  NAND2HSV0 U48962 ( .A1(n52974), .A2(n52448), .ZN(n44974) );
  XOR2HSV0 U48963 ( .A1(n44975), .A2(n44974), .Z(n44980) );
  CLKNHSV0 U48964 ( .I(n51537), .ZN(n51486) );
  NAND2HSV0 U48965 ( .A1(n51486), .A2(n53015), .ZN(n44978) );
  NAND2HSV0 U48966 ( .A1(n44976), .A2(n52994), .ZN(n44977) );
  XOR2HSV0 U48967 ( .A1(n44978), .A2(n44977), .Z(n44979) );
  XOR2HSV0 U48968 ( .A1(n44980), .A2(n44979), .Z(n45004) );
  NAND2HSV0 U48969 ( .A1(n36409), .A2(n53038), .ZN(n45003) );
  NAND2HSV0 U48970 ( .A1(n51759), .A2(n43961), .ZN(n44982) );
  INHSV2 U48971 ( .I(n48621), .ZN(n52309) );
  NAND2HSV0 U48972 ( .A1(n44892), .A2(n52309), .ZN(n44981) );
  XOR2HSV0 U48973 ( .A1(n44982), .A2(n44981), .Z(n44986) );
  NAND2HSV0 U48974 ( .A1(n52457), .A2(n36588), .ZN(n44984) );
  NAND2HSV0 U48975 ( .A1(\pe2/aot [15]), .A2(\pe2/bq[21] ), .ZN(n44983) );
  XOR2HSV0 U48976 ( .A1(n44984), .A2(n44983), .Z(n44985) );
  XOR2HSV0 U48977 ( .A1(n44986), .A2(n44985), .Z(n45002) );
  NAND2HSV0 U48978 ( .A1(\pe2/aot [25]), .A2(n52073), .ZN(n44989) );
  NAND2HSV0 U48979 ( .A1(n39019), .A2(n44987), .ZN(n44988) );
  XOR2HSV0 U48980 ( .A1(n44989), .A2(n44988), .Z(n44993) );
  NAND2HSV0 U48981 ( .A1(n53009), .A2(\pe2/bq[26] ), .ZN(n44991) );
  NAND2HSV0 U48982 ( .A1(\pe2/aot [19]), .A2(\pe2/bq[17] ), .ZN(n44990) );
  XOR2HSV0 U48983 ( .A1(n44991), .A2(n44990), .Z(n44992) );
  XOR2HSV0 U48984 ( .A1(n44993), .A2(n44992), .Z(n45000) );
  NAND2HSV0 U48985 ( .A1(n59497), .A2(\pe2/pvq [29]), .ZN(n44994) );
  XOR2HSV0 U48986 ( .A1(n44994), .A2(\pe2/phq [29]), .Z(n44998) );
  NAND2HSV0 U48987 ( .A1(\pe2/aot [22]), .A2(\pe2/bq[8] ), .ZN(n52082) );
  OAI22HSV0 U48988 ( .A1(n37940), .A2(n51567), .B1(n44871), .B2(n47580), .ZN(
        n44995) );
  OAI21HSV0 U48989 ( .A1(n44996), .A2(n52082), .B(n44995), .ZN(n44997) );
  XOR2HSV0 U48990 ( .A1(n44998), .A2(n44997), .Z(n44999) );
  XNOR2HSV1 U48991 ( .A1(n45000), .A2(n44999), .ZN(n45001) );
  XOR4HSV1 U48992 ( .A1(n45004), .A2(n45003), .A3(n45002), .A4(n45001), .Z(
        n45044) );
  CLKNAND2HSV0 U48993 ( .A1(n38479), .A2(n53006), .ZN(n45007) );
  NAND2HSV0 U48994 ( .A1(n45005), .A2(n51832), .ZN(n45006) );
  XOR2HSV0 U48995 ( .A1(n45007), .A2(n45006), .Z(n45012) );
  NAND2HSV0 U48996 ( .A1(n59768), .A2(n52973), .ZN(n45010) );
  NAND2HSV0 U48997 ( .A1(n59984), .A2(n45008), .ZN(n45009) );
  XOR2HSV0 U48998 ( .A1(n45010), .A2(n45009), .Z(n45011) );
  XOR2HSV0 U48999 ( .A1(n45012), .A2(n45011), .Z(n45021) );
  NAND2HSV0 U49000 ( .A1(\pe2/aot [23]), .A2(n47598), .ZN(n45014) );
  NAND2HSV0 U49001 ( .A1(n52289), .A2(\pe2/bq[6] ), .ZN(n45013) );
  XOR2HSV0 U49002 ( .A1(n45014), .A2(n45013), .Z(n45019) );
  NAND2HSV0 U49003 ( .A1(n29736), .A2(n36607), .ZN(n45017) );
  NAND2HSV0 U49004 ( .A1(\pe2/aot [12]), .A2(n45015), .ZN(n45016) );
  XOR2HSV0 U49005 ( .A1(n45017), .A2(n45016), .Z(n45018) );
  XOR2HSV0 U49006 ( .A1(n45019), .A2(n45018), .Z(n45020) );
  XOR2HSV0 U49007 ( .A1(n45021), .A2(n45020), .Z(n45042) );
  NAND2HSV0 U49008 ( .A1(\pe2/aot [21]), .A2(n52337), .ZN(n45023) );
  NAND2HSV0 U49009 ( .A1(n51636), .A2(n38393), .ZN(n45022) );
  XOR2HSV0 U49010 ( .A1(n45023), .A2(n45022), .Z(n45028) );
  NAND2HSV0 U49011 ( .A1(n59633), .A2(\pe2/bq[29] ), .ZN(n45026) );
  NAND2HSV0 U49012 ( .A1(n45024), .A2(n52965), .ZN(n45025) );
  XOR2HSV0 U49013 ( .A1(n45026), .A2(n45025), .Z(n45027) );
  XOR2HSV0 U49014 ( .A1(n45028), .A2(n45027), .Z(n45040) );
  INHSV2 U49015 ( .I(n45029), .ZN(n45032) );
  CLKNHSV0 U49016 ( .I(n45030), .ZN(n45031) );
  XOR2HSV0 U49017 ( .A1(n45032), .A2(n45031), .Z(n45038) );
  CLKNAND2HSV1 U49018 ( .A1(\pe2/aot [14]), .A2(n45033), .ZN(n45036) );
  NAND2HSV0 U49019 ( .A1(n45034), .A2(n52300), .ZN(n45035) );
  XOR2HSV0 U49020 ( .A1(n45036), .A2(n45035), .Z(n45037) );
  XOR2HSV0 U49021 ( .A1(n45038), .A2(n45037), .Z(n45039) );
  XOR2HSV0 U49022 ( .A1(n45040), .A2(n45039), .Z(n45041) );
  XOR2HSV0 U49023 ( .A1(n45042), .A2(n45041), .Z(n45043) );
  XNOR2HSV1 U49024 ( .A1(n45044), .A2(n45043), .ZN(n45045) );
  XNOR2HSV1 U49025 ( .A1(n45046), .A2(n45045), .ZN(n45047) );
  XNOR2HSV1 U49026 ( .A1(n45048), .A2(n45047), .ZN(n45050) );
  NAND2HSV0 U49027 ( .A1(n59679), .A2(n52052), .ZN(n45049) );
  XNOR2HSV1 U49028 ( .A1(n45050), .A2(n45049), .ZN(n45051) );
  XNOR2HSV1 U49029 ( .A1(n45052), .A2(n45051), .ZN(n45053) );
  XNOR2HSV1 U49030 ( .A1(n45054), .A2(n45053), .ZN(n45057) );
  NAND2HSV0 U49031 ( .A1(n45055), .A2(n52172), .ZN(n45056) );
  XOR2HSV0 U49032 ( .A1(n45057), .A2(n45056), .Z(n45060) );
  NAND2HSV0 U49033 ( .A1(n53050), .A2(n45058), .ZN(n45059) );
  XNOR2HSV1 U49034 ( .A1(n45060), .A2(n45059), .ZN(n45061) );
  XNOR2HSV1 U49035 ( .A1(n45062), .A2(n45061), .ZN(n45065) );
  NAND2HSV0 U49036 ( .A1(n45063), .A2(n51796), .ZN(n45064) );
  XOR3HSV2 U49037 ( .A1(n45066), .A2(n45065), .A3(n45064), .Z(n45067) );
  XNOR2HSV1 U49038 ( .A1(n45068), .A2(n45067), .ZN(n45069) );
  XNOR2HSV1 U49039 ( .A1(n45070), .A2(n45069), .ZN(n45073) );
  NOR2HSV0 U49040 ( .A1(n45071), .A2(n44327), .ZN(n45072) );
  XOR3HSV2 U49041 ( .A1(n45074), .A2(n45073), .A3(n45072), .Z(n45075) );
  XOR2HSV0 U49042 ( .A1(n45076), .A2(n45075), .Z(n45077) );
  XNOR2HSV1 U49043 ( .A1(n45078), .A2(n45077), .ZN(n45080) );
  CLKNAND2HSV1 U49044 ( .A1(n59361), .A2(n53077), .ZN(n45079) );
  XNOR2HSV1 U49045 ( .A1(n45080), .A2(n45079), .ZN(n45081) );
  XNOR2HSV1 U49046 ( .A1(n45082), .A2(n45081), .ZN(n45085) );
  CLKNAND2HSV0 U49047 ( .A1(n59774), .A2(n53086), .ZN(n45084) );
  XOR3HSV2 U49048 ( .A1(n45086), .A2(n45085), .A3(n45084), .Z(n45087) );
  CLKNAND2HSV0 U49049 ( .A1(n45089), .A2(n52415), .ZN(n45090) );
  AOI21HSV4 U49050 ( .A1(n29696), .A2(n45092), .B(n45276), .ZN(n45095) );
  INHSV2 U49051 ( .I(n45095), .ZN(n45093) );
  NAND2HSV2 U49052 ( .A1(n45094), .A2(n45093), .ZN(n45098) );
  CLKNAND2HSV2 U49053 ( .A1(n45096), .A2(n45095), .ZN(n45097) );
  CLKNHSV2 U49054 ( .I(n45102), .ZN(n45103) );
  NOR2HSV2 U49055 ( .A1(n45104), .A2(n45103), .ZN(n45107) );
  NAND3HSV2 U49056 ( .A1(n45107), .A2(n45106), .A3(n45105), .ZN(n45110) );
  OR2HSV1 U49057 ( .A1(n45108), .A2(n45267), .Z(n45109) );
  INHSV2 U49058 ( .I(n45119), .ZN(n45111) );
  INHSV2 U49059 ( .I(n45111), .ZN(n45116) );
  NOR2HSV4 U49060 ( .A1(n45115), .A2(n45114), .ZN(n45120) );
  NOR2HSV4 U49061 ( .A1(n45116), .A2(n45120), .ZN(n45117) );
  CLKNAND2HSV3 U49062 ( .A1(n45118), .A2(n45117), .ZN(n45126) );
  OAI21HSV4 U49063 ( .A1(n45121), .A2(n45120), .B(n45116), .ZN(n45124) );
  NOR2HSV4 U49064 ( .A1(n47499), .A2(n45276), .ZN(n45123) );
  CLKNAND2HSV3 U49065 ( .A1(n45122), .A2(n45123), .ZN(n45128) );
  INHSV2 U49066 ( .I(n45123), .ZN(n45125) );
  NOR2HSV1 U49067 ( .A1(n44309), .A2(\pe2/ti_7t [29]), .ZN(n45268) );
  NOR2HSV2 U49068 ( .A1(n45268), .A2(n45130), .ZN(n45131) );
  NAND2HSV2 U49069 ( .A1(n45132), .A2(n45133), .ZN(n45137) );
  INHSV3 U49070 ( .I(n45132), .ZN(n45135) );
  NAND2HSV2 U49071 ( .A1(n52910), .A2(\pe2/got [27]), .ZN(n45257) );
  OAI21HSV2 U49072 ( .A1(n36473), .A2(\pe2/ti_7t [28]), .B(n47997), .ZN(n45263) );
  INHSV2 U49073 ( .I(n45263), .ZN(n45139) );
  NAND2HSV0 U49074 ( .A1(n45140), .A2(n45139), .ZN(n45142) );
  OR2HSV1 U49075 ( .A1(n45263), .A2(n45399), .Z(n45141) );
  INAND2HSV2 U49076 ( .A1(n45265), .B1(\pe2/ti_7t [29]), .ZN(n45144) );
  INHSV2 U49077 ( .I(n59789), .ZN(n47497) );
  INHSV3 U49078 ( .I(n47497), .ZN(n52854) );
  CLKNAND2HSV1 U49079 ( .A1(n52854), .A2(n49492), .ZN(n45256) );
  CLKNHSV2 U49080 ( .I(n45277), .ZN(n45146) );
  INHSV2 U49081 ( .I(n45147), .ZN(n51120) );
  CLKNAND2HSV1 U49082 ( .A1(n51120), .A2(n44711), .ZN(n45255) );
  CLKNAND2HSV1 U49083 ( .A1(n25835), .A2(n52416), .ZN(n45254) );
  INHSV2 U49084 ( .I(n47572), .ZN(n52170) );
  NOR2HSV1 U49085 ( .A1(n52170), .A2(n38711), .ZN(n45247) );
  CLKNAND2HSV0 U49086 ( .A1(n44968), .A2(n52042), .ZN(n45245) );
  BUFHSV2 U49087 ( .I(n47500), .Z(n52921) );
  NOR2HSV2 U49088 ( .A1(n47500), .A2(n52169), .ZN(n45243) );
  CLKNAND2HSV1 U49089 ( .A1(n52923), .A2(n59983), .ZN(n45240) );
  NAND2HSV0 U49090 ( .A1(n51801), .A2(n51958), .ZN(n45234) );
  BUFHSV2 U49091 ( .I(n59773), .Z(n52926) );
  CLKNAND2HSV0 U49092 ( .A1(n52926), .A2(n52172), .ZN(n45232) );
  CLKNHSV2 U49093 ( .I(n49656), .ZN(n49493) );
  NAND2HSV0 U49094 ( .A1(n51965), .A2(n49493), .ZN(n45229) );
  NAND2HSV0 U49095 ( .A1(n51609), .A2(\pe2/got [10]), .ZN(n45227) );
  NAND2HSV0 U49096 ( .A1(\pe2/got [8]), .A2(n52929), .ZN(n45225) );
  CLKNAND2HSV0 U49097 ( .A1(n52931), .A2(n52174), .ZN(n45222) );
  NAND2HSV0 U49098 ( .A1(n38041), .A2(n51896), .ZN(n45215) );
  NAND2HSV0 U49099 ( .A1(n45150), .A2(n52239), .ZN(n45213) );
  NAND2HSV0 U49100 ( .A1(n59669), .A2(n59767), .ZN(n45209) );
  NAND2HSV0 U49101 ( .A1(n37801), .A2(n51457), .ZN(n45152) );
  NAND2HSV0 U49102 ( .A1(n51759), .A2(n51733), .ZN(n45151) );
  XOR2HSV0 U49103 ( .A1(n45152), .A2(n45151), .Z(n45156) );
  NAND2HSV0 U49104 ( .A1(n59587), .A2(n52481), .ZN(n45154) );
  NAND2HSV0 U49105 ( .A1(n52955), .A2(n52073), .ZN(n45153) );
  XOR2HSV0 U49106 ( .A1(n45154), .A2(n45153), .Z(n45155) );
  XOR2HSV0 U49107 ( .A1(n45156), .A2(n45155), .Z(n45164) );
  NAND2HSV0 U49108 ( .A1(n52070), .A2(\pe2/bq[14] ), .ZN(n45158) );
  NAND2HSV0 U49109 ( .A1(n52056), .A2(n38542), .ZN(n45157) );
  XOR2HSV0 U49110 ( .A1(n45158), .A2(n45157), .Z(n45162) );
  NAND2HSV0 U49111 ( .A1(\pe2/aot [2]), .A2(n39032), .ZN(n45160) );
  CLKNHSV0 U49112 ( .I(n49628), .ZN(n52962) );
  NAND2HSV0 U49113 ( .A1(n51743), .A2(n52962), .ZN(n45159) );
  XOR2HSV0 U49114 ( .A1(n45160), .A2(n45159), .Z(n45161) );
  XOR2HSV0 U49115 ( .A1(n45162), .A2(n45161), .Z(n45163) );
  XOR2HSV0 U49116 ( .A1(n45164), .A2(n45163), .Z(n45181) );
  NAND2HSV0 U49117 ( .A1(n51920), .A2(n43956), .ZN(n45167) );
  NAND2HSV0 U49118 ( .A1(n52310), .A2(n51493), .ZN(n45166) );
  XOR2HSV0 U49119 ( .A1(n45167), .A2(n45166), .Z(n45171) );
  NAND2HSV0 U49120 ( .A1(n59768), .A2(n51998), .ZN(n45169) );
  NAND2HSV0 U49121 ( .A1(\pe2/aot [8]), .A2(\pe2/bq[21] ), .ZN(n45168) );
  XOR2HSV0 U49122 ( .A1(n45169), .A2(n45168), .Z(n45170) );
  XOR2HSV0 U49123 ( .A1(n45171), .A2(n45170), .Z(n45179) );
  NAND2HSV0 U49124 ( .A1(n52974), .A2(n52484), .ZN(n45173) );
  NAND2HSV0 U49125 ( .A1(n53005), .A2(\pe2/bq[17] ), .ZN(n45172) );
  XOR2HSV0 U49126 ( .A1(n45173), .A2(n45172), .Z(n45177) );
  NAND2HSV0 U49127 ( .A1(\pe2/aot [7]), .A2(n45033), .ZN(n45175) );
  NAND2HSV0 U49128 ( .A1(n39019), .A2(n52988), .ZN(n45174) );
  XOR2HSV0 U49129 ( .A1(n45175), .A2(n45174), .Z(n45176) );
  XOR2HSV0 U49130 ( .A1(n45177), .A2(n45176), .Z(n45178) );
  XOR2HSV0 U49131 ( .A1(n45179), .A2(n45178), .Z(n45180) );
  XOR2HSV0 U49132 ( .A1(n45181), .A2(n45180), .Z(n45207) );
  NOR2HSV0 U49133 ( .A1(n37940), .A2(n50920), .ZN(n52291) );
  NOR2HSV0 U49134 ( .A1(n52080), .A2(n49515), .ZN(n45183) );
  CLKNAND2HSV1 U49135 ( .A1(n52294), .A2(n52851), .ZN(n51817) );
  OAI22HSV0 U49136 ( .A1(n52291), .A2(n45183), .B1(n45182), .B2(n51817), .ZN(
        n45188) );
  NAND2HSV0 U49137 ( .A1(n52998), .A2(n51803), .ZN(n49538) );
  NAND2HSV0 U49138 ( .A1(n52456), .A2(n52179), .ZN(n45186) );
  NAND2HSV2 U49139 ( .A1(n52456), .A2(n51803), .ZN(n51124) );
  NOR2HSV0 U49140 ( .A1(n45184), .A2(n51124), .ZN(n45185) );
  AOI21HSV1 U49141 ( .A1(n49538), .A2(n45186), .B(n45185), .ZN(n45187) );
  XOR2HSV0 U49142 ( .A1(n45188), .A2(n45187), .Z(n45198) );
  NOR2HSV0 U49143 ( .A1(n51537), .A2(n44854), .ZN(n45190) );
  INHSV2 U49144 ( .I(n51537), .ZN(n52184) );
  NAND2HSV2 U49145 ( .A1(n52184), .A2(\pe2/bq[8] ), .ZN(n51540) );
  OAI22HSV0 U49146 ( .A1(n45191), .A2(n45190), .B1(n45189), .B2(n51540), .ZN(
        n45196) );
  NAND2HSV2 U49147 ( .A1(n53016), .A2(n52857), .ZN(n51967) );
  NOR2HSV0 U49148 ( .A1(n45192), .A2(n51967), .ZN(n45194) );
  AOI22HSV0 U49149 ( .A1(n50956), .A2(n52994), .B1(n52987), .B2(\pe2/aot [1]), 
        .ZN(n45193) );
  NOR2HSV2 U49150 ( .A1(n45194), .A2(n45193), .ZN(n45195) );
  XNOR2HSV1 U49151 ( .A1(n45196), .A2(n45195), .ZN(n45197) );
  XNOR2HSV1 U49152 ( .A1(n45198), .A2(n45197), .ZN(n45205) );
  NAND2HSV0 U49153 ( .A1(n59792), .A2(n52952), .ZN(n49519) );
  NAND2HSV0 U49154 ( .A1(n59977), .A2(\pe2/bq[19] ), .ZN(n52432) );
  XOR2HSV0 U49155 ( .A1(n49519), .A2(n52432), .Z(n45203) );
  NOR2HSV0 U49156 ( .A1(n47574), .A2(n44718), .ZN(n45201) );
  INHSV2 U49157 ( .I(n38822), .ZN(n52966) );
  NAND2HSV0 U49158 ( .A1(n52966), .A2(\pe2/bq[16] ), .ZN(n45200) );
  XOR2HSV0 U49159 ( .A1(n45201), .A2(n45200), .Z(n45202) );
  XOR2HSV0 U49160 ( .A1(n45203), .A2(n45202), .Z(n45204) );
  XNOR2HSV1 U49161 ( .A1(n45205), .A2(n45204), .ZN(n45206) );
  XNOR2HSV1 U49162 ( .A1(n45207), .A2(n45206), .ZN(n45208) );
  XNOR2HSV1 U49163 ( .A1(n45209), .A2(n45208), .ZN(n45211) );
  NAND2HSV0 U49164 ( .A1(n44254), .A2(n51932), .ZN(n45210) );
  XNOR2HSV1 U49165 ( .A1(n45211), .A2(n45210), .ZN(n45212) );
  XNOR2HSV1 U49166 ( .A1(n45213), .A2(n45212), .ZN(n45214) );
  XNOR2HSV1 U49167 ( .A1(n45215), .A2(n45214), .ZN(n45217) );
  INHSV2 U49168 ( .I(n50908), .ZN(n52175) );
  NAND2HSV0 U49169 ( .A1(n59766), .A2(n52175), .ZN(n45216) );
  XOR2HSV0 U49170 ( .A1(n45217), .A2(n45216), .Z(n45220) );
  NAND2HSV0 U49171 ( .A1(n44120), .A2(\pe2/got [6]), .ZN(n45219) );
  XNOR2HSV1 U49172 ( .A1(n45220), .A2(n45219), .ZN(n45221) );
  XNOR2HSV1 U49173 ( .A1(n45222), .A2(n45221), .ZN(n45224) );
  NAND2HSV0 U49174 ( .A1(n59761), .A2(n44714), .ZN(n45223) );
  XOR3HSV2 U49175 ( .A1(n45225), .A2(n45224), .A3(n45223), .Z(n45226) );
  XNOR2HSV1 U49176 ( .A1(n45227), .A2(n45226), .ZN(n45228) );
  XNOR2HSV1 U49177 ( .A1(n45229), .A2(n45228), .ZN(n45231) );
  NOR2HSV0 U49178 ( .A1(n45071), .A2(n51607), .ZN(n45230) );
  XOR3HSV2 U49179 ( .A1(n45232), .A2(n45231), .A3(n45230), .Z(n45233) );
  XOR2HSV0 U49180 ( .A1(n45234), .A2(n45233), .Z(n45238) );
  CLKNHSV0 U49181 ( .I(n45235), .ZN(n45795) );
  BUFHSV2 U49182 ( .I(n45795), .Z(n52532) );
  CLKNAND2HSV0 U49183 ( .A1(n52532), .A2(n51964), .ZN(n45237) );
  INHSV2 U49184 ( .I(n29745), .ZN(n52138) );
  CLKNAND2HSV1 U49185 ( .A1(n52138), .A2(n51796), .ZN(n45236) );
  XOR3HSV2 U49186 ( .A1(n45238), .A2(n45237), .A3(n45236), .Z(n45239) );
  XNOR2HSV1 U49187 ( .A1(n45240), .A2(n45239), .ZN(n45242) );
  BUFHSV2 U49188 ( .I(n59774), .Z(n53078) );
  INHSV2 U49189 ( .I(n47570), .ZN(n52533) );
  CLKNAND2HSV0 U49190 ( .A1(n53078), .A2(n52533), .ZN(n45241) );
  XOR3HSV2 U49191 ( .A1(n45243), .A2(n45242), .A3(n45241), .Z(n45244) );
  XOR2HSV0 U49192 ( .A1(n45245), .A2(n45244), .Z(n45246) );
  XNOR2HSV1 U49193 ( .A1(n45247), .A2(n45246), .ZN(n45252) );
  INHSV2 U49194 ( .I(n45248), .ZN(n52276) );
  CLKNAND2HSV1 U49195 ( .A1(n59927), .A2(n52276), .ZN(n45251) );
  INHSV2 U49196 ( .I(n47939), .ZN(n52399) );
  CLKNAND2HSV0 U49197 ( .A1(n52399), .A2(n45249), .ZN(n45250) );
  XOR3HSV2 U49198 ( .A1(n45252), .A2(n45251), .A3(n45250), .Z(n45253) );
  CLKNAND2HSV1 U49199 ( .A1(n45257), .A2(n45258), .ZN(n45262) );
  INHSV1 U49200 ( .I(n45257), .ZN(n45260) );
  CLKNAND2HSV1 U49201 ( .A1(n45260), .A2(n45259), .ZN(n45261) );
  AND3HSV2 U49202 ( .A1(n45275), .A2(n45274), .A3(n45273), .Z(n45279) );
  NOR2HSV1 U49203 ( .A1(n45277), .A2(n45276), .ZN(n45278) );
  AOI31HSV2 U49204 ( .A1(n53388), .A2(n45279), .A3(n38873), .B(n45278), .ZN(
        n45285) );
  INHSV2 U49205 ( .I(n53388), .ZN(n45283) );
  NAND3HSV2 U49206 ( .A1(n45283), .A2(n45282), .A3(n59980), .ZN(n45284) );
  NAND2HSV2 U49207 ( .A1(n45285), .A2(n45284), .ZN(n45393) );
  NAND2HSV2 U49208 ( .A1(n59522), .A2(n38324), .ZN(n45382) );
  NOR2HSV0 U49209 ( .A1(n47500), .A2(n38275), .ZN(n45380) );
  NAND2HSV0 U49210 ( .A1(n51485), .A2(n45287), .ZN(n45377) );
  NAND2HSV0 U49211 ( .A1(n52924), .A2(n52042), .ZN(n45373) );
  NAND2HSV0 U49212 ( .A1(n52533), .A2(n52173), .ZN(n45371) );
  CLKNAND2HSV0 U49213 ( .A1(n52286), .A2(\pe2/got [17]), .ZN(n45369) );
  NAND2HSV0 U49214 ( .A1(n45288), .A2(n51796), .ZN(n45366) );
  CLKNAND2HSV0 U49215 ( .A1(n52928), .A2(n45289), .ZN(n45364) );
  INHSV2 U49216 ( .I(n51607), .ZN(n53055) );
  NAND2HSV0 U49217 ( .A1(n53055), .A2(n51966), .ZN(n45362) );
  CLKNAND2HSV1 U49218 ( .A1(n52287), .A2(n52172), .ZN(n45359) );
  CLKNAND2HSV1 U49219 ( .A1(n44185), .A2(\pe2/got [9]), .ZN(n45353) );
  NAND2HSV0 U49220 ( .A1(n45290), .A2(\pe2/got [8]), .ZN(n45351) );
  NAND2HSV0 U49221 ( .A1(n38539), .A2(n53038), .ZN(n45292) );
  NOR2HSV0 U49222 ( .A1(n53033), .A2(n50909), .ZN(n45291) );
  XOR2HSV0 U49223 ( .A1(n45292), .A2(n45291), .Z(n45345) );
  NAND2HSV0 U49224 ( .A1(\pe2/aot [19]), .A2(n52337), .ZN(n51814) );
  NAND2HSV0 U49225 ( .A1(n52994), .A2(n52485), .ZN(n48936) );
  NOR2HSV0 U49226 ( .A1(n38404), .A2(n47893), .ZN(n52947) );
  INHSV2 U49227 ( .I(n38404), .ZN(n52289) );
  NAND2HSV0 U49228 ( .A1(n38479), .A2(\pe2/bq[2] ), .ZN(n52219) );
  NAND2HSV0 U49229 ( .A1(n45295), .A2(n51457), .ZN(n49528) );
  CLKNHSV0 U49230 ( .I(n36530), .ZN(n52973) );
  NAND2HSV0 U49231 ( .A1(n59633), .A2(n52973), .ZN(n49533) );
  NAND2HSV0 U49232 ( .A1(n59768), .A2(n44987), .ZN(n52202) );
  NAND2HSV0 U49233 ( .A1(n52457), .A2(n38064), .ZN(n52455) );
  NAND2HSV0 U49234 ( .A1(n52995), .A2(\pe2/bq[6] ), .ZN(n45296) );
  XOR2HSV0 U49235 ( .A1(n45297), .A2(n45296), .Z(n45300) );
  NAND2HSV0 U49236 ( .A1(n52070), .A2(\pe2/bq[19] ), .ZN(n51843) );
  XOR2HSV0 U49237 ( .A1(n45298), .A2(n51843), .Z(n45299) );
  XOR2HSV0 U49238 ( .A1(n45300), .A2(n45299), .Z(n45309) );
  NOR2HSV0 U49239 ( .A1(n52226), .A2(n48064), .ZN(n45302) );
  NAND2HSV0 U49240 ( .A1(n39052), .A2(\pe2/bq[14] ), .ZN(n45301) );
  XOR2HSV0 U49241 ( .A1(n45302), .A2(n45301), .Z(n45307) );
  NAND2HSV0 U49242 ( .A1(n52993), .A2(n38393), .ZN(n45305) );
  NAND2HSV2 U49243 ( .A1(\pe2/got [2]), .A2(n45303), .ZN(n45304) );
  XNOR2HSV1 U49244 ( .A1(n45305), .A2(n45304), .ZN(n45306) );
  XNOR2HSV1 U49245 ( .A1(n45307), .A2(n45306), .ZN(n45308) );
  XNOR2HSV1 U49246 ( .A1(n45309), .A2(n45308), .ZN(n45311) );
  NAND2HSV0 U49247 ( .A1(n36409), .A2(n59351), .ZN(n45310) );
  XNOR2HSV1 U49248 ( .A1(n45311), .A2(n45310), .ZN(n45342) );
  CLKNAND2HSV0 U49249 ( .A1(n52966), .A2(\pe2/bq[21] ), .ZN(n45313) );
  CLKNAND2HSV0 U49250 ( .A1(n53005), .A2(n45033), .ZN(n45312) );
  XOR2HSV0 U49251 ( .A1(n45313), .A2(n45312), .Z(n45317) );
  NAND2HSV0 U49252 ( .A1(n52955), .A2(n51732), .ZN(n45315) );
  NAND2HSV0 U49253 ( .A1(\pe2/aot [11]), .A2(n52300), .ZN(n45314) );
  XOR2HSV0 U49254 ( .A1(n45315), .A2(n45314), .Z(n45316) );
  XOR2HSV0 U49255 ( .A1(n45317), .A2(n45316), .Z(n45325) );
  NAND2HSV0 U49256 ( .A1(n52456), .A2(n52987), .ZN(n45319) );
  NAND2HSV0 U49257 ( .A1(\pe2/aot [5]), .A2(n36608), .ZN(n45318) );
  XOR2HSV0 U49258 ( .A1(n45319), .A2(n45318), .Z(n45323) );
  NAND2HSV0 U49259 ( .A1(n53009), .A2(\pe2/bq[24] ), .ZN(n45321) );
  NAND2HSV0 U49260 ( .A1(n52998), .A2(n52322), .ZN(n45320) );
  XOR2HSV0 U49261 ( .A1(n45321), .A2(n45320), .Z(n45322) );
  XOR2HSV0 U49262 ( .A1(n45323), .A2(n45322), .Z(n45324) );
  XOR2HSV0 U49263 ( .A1(n45325), .A2(n45324), .Z(n45340) );
  NOR2HSV0 U49264 ( .A1(n47574), .A2(n47508), .ZN(n45327) );
  NAND2HSV0 U49265 ( .A1(n37801), .A2(n53006), .ZN(n45326) );
  XOR2HSV0 U49266 ( .A1(n45327), .A2(n45326), .Z(n45330) );
  NAND2HSV0 U49267 ( .A1(n59497), .A2(\pe2/pvq [31]), .ZN(n45328) );
  XOR2HSV0 U49268 ( .A1(n45328), .A2(\pe2/phq [31]), .Z(n45329) );
  XOR2HSV0 U49269 ( .A1(n45330), .A2(n45329), .Z(n45338) );
  NAND2HSV0 U49270 ( .A1(\pe2/aot [2]), .A2(n52444), .ZN(n52946) );
  OAI22HSV0 U49271 ( .A1(n38418), .A2(n49618), .B1(n51538), .B2(n36237), .ZN(
        n45331) );
  OAI21HSV1 U49272 ( .A1(n45332), .A2(n52946), .B(n45331), .ZN(n45336) );
  CLKNAND2HSV0 U49273 ( .A1(n44745), .A2(n52962), .ZN(n52102) );
  OAI22HSV0 U49274 ( .A1(n47575), .A2(n49628), .B1(n45165), .B2(n47599), .ZN(
        n45333) );
  OAI21HSV0 U49275 ( .A1(n52102), .A2(n45334), .B(n45333), .ZN(n45335) );
  XOR2HSV0 U49276 ( .A1(n45336), .A2(n45335), .Z(n45337) );
  XOR2HSV0 U49277 ( .A1(n45338), .A2(n45337), .Z(n45339) );
  XNOR2HSV1 U49278 ( .A1(n45340), .A2(n45339), .ZN(n45341) );
  XOR3HSV2 U49279 ( .A1(n45343), .A2(n45342), .A3(n45341), .Z(n45344) );
  XOR2HSV0 U49280 ( .A1(n45345), .A2(n45344), .Z(n45347) );
  CLKNAND2HSV1 U49281 ( .A1(n59669), .A2(n53041), .ZN(n45346) );
  XOR2HSV0 U49282 ( .A1(n45347), .A2(n45346), .Z(n45349) );
  CLKNAND2HSV0 U49283 ( .A1(n59679), .A2(n59757), .ZN(n45348) );
  XNOR2HSV1 U49284 ( .A1(n45349), .A2(n45348), .ZN(n45350) );
  XNOR2HSV1 U49285 ( .A1(n45351), .A2(n45350), .ZN(n45352) );
  XNOR2HSV1 U49286 ( .A1(n45353), .A2(n45352), .ZN(n45355) );
  NAND2HSV0 U49287 ( .A1(n52367), .A2(\pe2/got [10]), .ZN(n45354) );
  XOR2HSV0 U49288 ( .A1(n45355), .A2(n45354), .Z(n45357) );
  NAND2HSV0 U49289 ( .A1(n53050), .A2(n52374), .ZN(n45356) );
  XNOR2HSV1 U49290 ( .A1(n45357), .A2(n45356), .ZN(n45358) );
  XNOR2HSV1 U49291 ( .A1(n45359), .A2(n45358), .ZN(n45361) );
  CLKNAND2HSV1 U49292 ( .A1(n53056), .A2(n51608), .ZN(n45360) );
  XOR3HSV2 U49293 ( .A1(n45362), .A2(n45361), .A3(n45360), .Z(n45363) );
  XNOR2HSV1 U49294 ( .A1(n45364), .A2(n45363), .ZN(n45365) );
  XNOR2HSV1 U49295 ( .A1(n45366), .A2(n45365), .ZN(n45368) );
  NAND2HSV0 U49296 ( .A1(n59505), .A2(n52925), .ZN(n45367) );
  XOR3HSV2 U49297 ( .A1(n45369), .A2(n45368), .A3(n45367), .Z(n45370) );
  XOR2HSV0 U49298 ( .A1(n45371), .A2(n45370), .Z(n45372) );
  XNOR2HSV1 U49299 ( .A1(n45373), .A2(n45372), .ZN(n45375) );
  NAND2HSV0 U49300 ( .A1(n59361), .A2(\pe2/got [21]), .ZN(n45374) );
  XNOR2HSV1 U49301 ( .A1(n45375), .A2(n45374), .ZN(n45376) );
  XNOR2HSV1 U49302 ( .A1(n45377), .A2(n45376), .ZN(n45379) );
  CLKNAND2HSV1 U49303 ( .A1(n59774), .A2(n59584), .ZN(n45378) );
  XOR3HSV2 U49304 ( .A1(n45380), .A2(n45379), .A3(n45378), .Z(n45381) );
  XOR2HSV0 U49305 ( .A1(n45382), .A2(n45381), .Z(n45384) );
  NAND2HSV2 U49306 ( .A1(n47572), .A2(n38389), .ZN(n45383) );
  XOR2HSV0 U49307 ( .A1(n45384), .A2(n45383), .Z(n45385) );
  NAND2HSV2 U49308 ( .A1(n59927), .A2(n44944), .ZN(n45386) );
  XNOR2HSV4 U49309 ( .A1(n45393), .A2(n45392), .ZN(n45395) );
  INHSV2 U49310 ( .I(n45395), .ZN(n45394) );
  CLKNAND2HSV1 U49311 ( .A1(n45396), .A2(n45395), .ZN(n45397) );
  CLKNHSV0 U49312 ( .I(n45401), .ZN(n45402) );
  NAND2HSV2 U49313 ( .A1(n45400), .A2(n45402), .ZN(n45406) );
  CLKNHSV0 U49314 ( .I(n45403), .ZN(n45404) );
  AND2HSV2 U49315 ( .A1(n38184), .A2(\pe2/ti_7t [31]), .Z(n48161) );
  INAND2HSV2 U49316 ( .A1(n45411), .B1(n53097), .ZN(n45412) );
  XNOR2HSV1 U49317 ( .A1(n45413), .A2(n45412), .ZN(\pe2/poht [4]) );
  NAND2HSV2 U49318 ( .A1(\pe5/ti_7t [30]), .A2(n39702), .ZN(n53188) );
  NAND2HSV4 U49319 ( .A1(n51230), .A2(n51229), .ZN(n59580) );
  INHSV2 U49320 ( .I(n46976), .ZN(n52670) );
  CLKNAND2HSV0 U49321 ( .A1(n52670), .A2(\pe5/got [23]), .ZN(n45498) );
  BUFHSV2 U49322 ( .I(n25864), .Z(n53291) );
  CLKNAND2HSV0 U49323 ( .A1(n53291), .A2(n51228), .ZN(n45494) );
  NOR2HSV0 U49324 ( .A1(n51361), .A2(n46583), .ZN(n45488) );
  BUFHSV2 U49325 ( .I(n45818), .Z(n52569) );
  CLKNAND2HSV0 U49326 ( .A1(n52569), .A2(n51224), .ZN(n45484) );
  NAND2HSV0 U49327 ( .A1(n51158), .A2(n51157), .ZN(n45482) );
  BUFHSV2 U49328 ( .I(n45417), .Z(n52572) );
  CLKNHSV0 U49329 ( .I(n45418), .ZN(n59513) );
  INHSV2 U49330 ( .I(n51231), .ZN(n51331) );
  NAND2HSV0 U49331 ( .A1(\pe5/aot [14]), .A2(n52610), .ZN(n45420) );
  NAND2HSV0 U49332 ( .A1(\pe5/aot [16]), .A2(n52632), .ZN(n45419) );
  XOR2HSV0 U49333 ( .A1(n45420), .A2(n45419), .Z(n45425) );
  NAND2HSV0 U49334 ( .A1(n48663), .A2(\pe5/bq[1] ), .ZN(n45423) );
  NAND2HSV0 U49335 ( .A1(\pe5/aot [13]), .A2(n51176), .ZN(n45422) );
  XOR2HSV0 U49336 ( .A1(n45423), .A2(n45422), .Z(n45424) );
  XOR2HSV0 U49337 ( .A1(n45425), .A2(n45424), .Z(n45434) );
  NAND2HSV0 U49338 ( .A1(n51313), .A2(n39487), .ZN(n45428) );
  NAND2HSV0 U49339 ( .A1(\pe5/aot [20]), .A2(n53216), .ZN(n45427) );
  XOR2HSV0 U49340 ( .A1(n45428), .A2(n45427), .Z(n45432) );
  NAND2HSV0 U49341 ( .A1(n47278), .A2(n39914), .ZN(n45430) );
  NAND2HSV0 U49342 ( .A1(n37660), .A2(n51191), .ZN(n45429) );
  XOR2HSV0 U49343 ( .A1(n45430), .A2(n45429), .Z(n45431) );
  XOR2HSV0 U49344 ( .A1(n45432), .A2(n45431), .Z(n45433) );
  XOR2HSV0 U49345 ( .A1(n45434), .A2(n45433), .Z(n45450) );
  CLKNHSV0 U49346 ( .I(n48031), .ZN(n48764) );
  NAND2HSV0 U49347 ( .A1(n48829), .A2(n48764), .ZN(n45436) );
  NAND2HSV0 U49348 ( .A1(n59944), .A2(n47305), .ZN(n45435) );
  XOR2HSV0 U49349 ( .A1(n45436), .A2(n45435), .Z(n45440) );
  NAND2HSV0 U49350 ( .A1(n39266), .A2(\pe5/bq[2] ), .ZN(n45438) );
  CLKNHSV2 U49351 ( .I(n50507), .ZN(n53299) );
  NAND2HSV0 U49352 ( .A1(n53299), .A2(n51167), .ZN(n45437) );
  XOR2HSV0 U49353 ( .A1(n45438), .A2(n45437), .Z(n45439) );
  XOR2HSV0 U49354 ( .A1(n45440), .A2(n45439), .Z(n45448) );
  NAND2HSV0 U49355 ( .A1(n52611), .A2(\pe5/bq[19] ), .ZN(n45442) );
  NAND2HSV0 U49356 ( .A1(\pe5/aot [8]), .A2(n47059), .ZN(n45441) );
  XOR2HSV0 U49357 ( .A1(n45442), .A2(n45441), .Z(n45446) );
  NOR2HSV0 U49358 ( .A1(n40043), .A2(n47207), .ZN(n45444) );
  NAND2HSV0 U49359 ( .A1(n48242), .A2(n48775), .ZN(n45443) );
  XOR2HSV0 U49360 ( .A1(n45444), .A2(n45443), .Z(n45445) );
  XNOR2HSV1 U49361 ( .A1(n45446), .A2(n45445), .ZN(n45447) );
  XNOR2HSV1 U49362 ( .A1(n45448), .A2(n45447), .ZN(n45449) );
  XNOR2HSV1 U49363 ( .A1(n45450), .A2(n45449), .ZN(n45476) );
  CLKNHSV0 U49364 ( .I(n45451), .ZN(n51188) );
  NAND2HSV0 U49365 ( .A1(n51188), .A2(n52672), .ZN(n45453) );
  BUFHSV2 U49366 ( .I(\pe5/aot [6]), .Z(n53295) );
  NAND2HSV0 U49367 ( .A1(n52682), .A2(n30341), .ZN(n45452) );
  XOR2HSV0 U49368 ( .A1(n45453), .A2(n45452), .Z(n45457) );
  NAND2HSV0 U49369 ( .A1(n48199), .A2(n39592), .ZN(n45455) );
  CLKNHSV0 U49370 ( .I(n51021), .ZN(n52630) );
  NAND2HSV0 U49371 ( .A1(n48761), .A2(n52630), .ZN(n45454) );
  XOR2HSV0 U49372 ( .A1(n45455), .A2(n45454), .Z(n45456) );
  XOR2HSV0 U49373 ( .A1(n45457), .A2(n45456), .Z(n45467) );
  NOR2HSV0 U49374 ( .A1(n50518), .A2(n48050), .ZN(n45459) );
  CLKNHSV0 U49375 ( .I(n48219), .ZN(n59879) );
  BUFHSV2 U49376 ( .I(\pe5/bq[4] ), .Z(n51177) );
  NAND2HSV0 U49377 ( .A1(n59879), .A2(n51177), .ZN(n45458) );
  XOR2HSV0 U49378 ( .A1(n45459), .A2(n45458), .Z(n45465) );
  NOR2HSV0 U49379 ( .A1(n48246), .A2(n45460), .ZN(n47233) );
  NOR2HSV0 U49380 ( .A1(n45904), .A2(n45461), .ZN(n45463) );
  CLKNAND2HSV1 U49381 ( .A1(n51182), .A2(n39445), .ZN(n51025) );
  OAI22HSV0 U49382 ( .A1(n47233), .A2(n45463), .B1(n45462), .B2(n51025), .ZN(
        n45464) );
  XNOR2HSV1 U49383 ( .A1(n45465), .A2(n45464), .ZN(n45466) );
  XNOR2HSV1 U49384 ( .A1(n45467), .A2(n45466), .ZN(n45474) );
  NOR2HSV0 U49385 ( .A1(n59869), .A2(n30287), .ZN(n47242) );
  NOR2HSV0 U49386 ( .A1(n47409), .A2(n30113), .ZN(n48677) );
  AOI22HSV0 U49387 ( .A1(n50588), .A2(\pe5/bq[25] ), .B1(\pe5/bq[27] ), .B2(
        n52600), .ZN(n45468) );
  AOI21HSV2 U49388 ( .A1(n47242), .A2(n48677), .B(n45468), .ZN(n45469) );
  NAND2HSV0 U49389 ( .A1(\pe5/aot [4]), .A2(n30222), .ZN(n48674) );
  XNOR2HSV1 U49390 ( .A1(n45469), .A2(n48674), .ZN(n45472) );
  NAND2HSV0 U49391 ( .A1(\pe5/aot [18]), .A2(n39615), .ZN(n47315) );
  INHSV2 U49392 ( .I(n51232), .ZN(n48786) );
  NAND2HSV0 U49393 ( .A1(n48786), .A2(n45470), .ZN(n47311) );
  XOR2HSV0 U49394 ( .A1(n47315), .A2(n47311), .Z(n45471) );
  XOR2HSV0 U49395 ( .A1(n45472), .A2(n45471), .Z(n45473) );
  XNOR2HSV1 U49396 ( .A1(n45474), .A2(n45473), .ZN(n45475) );
  XNOR2HSV1 U49397 ( .A1(n45476), .A2(n45475), .ZN(n45478) );
  NAND2HSV0 U49398 ( .A1(n59517), .A2(n52652), .ZN(n45479) );
  XNOR2HSV1 U49399 ( .A1(n45480), .A2(n45479), .ZN(n45481) );
  XOR2HSV0 U49400 ( .A1(n45482), .A2(n45481), .Z(n45483) );
  XNOR2HSV1 U49401 ( .A1(n45484), .A2(n45483), .ZN(n45486) );
  NAND2HSV0 U49402 ( .A1(n51211), .A2(n51156), .ZN(n45485) );
  XNOR2HSV1 U49403 ( .A1(n45486), .A2(n45485), .ZN(n45487) );
  XNOR2HSV1 U49404 ( .A1(n45488), .A2(n45487), .ZN(n45492) );
  CLKNAND2HSV0 U49405 ( .A1(n48745), .A2(n39432), .ZN(n45491) );
  BUFHSV2 U49406 ( .I(n45489), .Z(n47394) );
  INHSV2 U49407 ( .I(n47394), .ZN(n52659) );
  NOR2HSV2 U49408 ( .A1(n52659), .A2(n39119), .ZN(n45490) );
  XOR3HSV2 U49409 ( .A1(n45492), .A2(n45491), .A3(n45490), .Z(n45493) );
  XNOR2HSV1 U49410 ( .A1(n45494), .A2(n45493), .ZN(n45496) );
  NAND2HSV0 U49411 ( .A1(n51092), .A2(n48744), .ZN(n45495) );
  XNOR2HSV1 U49412 ( .A1(n45496), .A2(n45495), .ZN(n45497) );
  XNOR2HSV1 U49413 ( .A1(n45498), .A2(n45497), .ZN(n45502) );
  CLKNAND2HSV0 U49414 ( .A1(n52693), .A2(n45500), .ZN(n45501) );
  CLKNAND2HSV2 U49415 ( .A1(n47141), .A2(n47052), .ZN(n52562) );
  NOR2HSV1 U49416 ( .A1(n45503), .A2(n46090), .ZN(n45507) );
  AND2HSV2 U49417 ( .A1(n45504), .A2(n29750), .Z(n45505) );
  NAND2HSV0 U49418 ( .A1(n45509), .A2(n55940), .ZN(n45510) );
  CLKNAND2HSV1 U49419 ( .A1(n45588), .A2(n45510), .ZN(n45515) );
  CLKNHSV0 U49420 ( .I(n45511), .ZN(n45512) );
  AND3HSV2 U49421 ( .A1(n45512), .A2(n37107), .A3(n59964), .Z(n45513) );
  NAND2HSV2 U49422 ( .A1(n56175), .A2(n45513), .ZN(n45514) );
  NAND2HSV2 U49423 ( .A1(n45515), .A2(n45514), .ZN(n45590) );
  INHSV2 U49424 ( .I(n45590), .ZN(n45595) );
  INHSV2 U49425 ( .I(n43457), .ZN(n45947) );
  CLKNHSV0 U49426 ( .I(n56821), .ZN(n48487) );
  CLKNHSV0 U49427 ( .I(n36694), .ZN(n48021) );
  NAND2HSV0 U49428 ( .A1(n59627), .A2(n48021), .ZN(n45520) );
  NAND2HSV0 U49429 ( .A1(n45973), .A2(n45663), .ZN(n45519) );
  XOR2HSV0 U49430 ( .A1(n45520), .A2(n45519), .Z(n45524) );
  NAND2HSV0 U49431 ( .A1(n59646), .A2(n46614), .ZN(n45522) );
  NAND2HSV2 U49432 ( .A1(n55873), .A2(n48538), .ZN(n45521) );
  XOR2HSV0 U49433 ( .A1(n45522), .A2(n45521), .Z(n45523) );
  NAND2HSV0 U49434 ( .A1(n56423), .A2(n55960), .ZN(n45527) );
  NAND2HSV0 U49435 ( .A1(\pe3/got [4]), .A2(n37007), .ZN(n45526) );
  XOR2HSV0 U49436 ( .A1(n45527), .A2(n45526), .Z(n45531) );
  BUFHSV2 U49437 ( .I(n36755), .Z(n55827) );
  NAND2HSV2 U49438 ( .A1(n55827), .A2(n56785), .ZN(n45529) );
  NAND2HSV0 U49439 ( .A1(n46332), .A2(n45982), .ZN(n45528) );
  XOR2HSV0 U49440 ( .A1(n45529), .A2(n45528), .Z(n45530) );
  INHSV2 U49441 ( .I(n56859), .ZN(n59799) );
  NAND2HSV0 U49442 ( .A1(n42728), .A2(n55616), .ZN(n45533) );
  BUFHSV2 U49443 ( .I(\pe3/aot [11]), .Z(n56197) );
  CLKNAND2HSV1 U49444 ( .A1(n56354), .A2(n55976), .ZN(n45532) );
  XOR2HSV0 U49445 ( .A1(n45533), .A2(n45532), .Z(n45538) );
  NAND2HSV0 U49446 ( .A1(n45645), .A2(n42971), .ZN(n45536) );
  CLKNAND2HSV0 U49447 ( .A1(n42818), .A2(n45534), .ZN(n45535) );
  XOR2HSV0 U49448 ( .A1(n45536), .A2(n45535), .Z(n45537) );
  XOR2HSV0 U49449 ( .A1(n45538), .A2(n45537), .Z(n45546) );
  NAND2HSV0 U49450 ( .A1(n45676), .A2(n43052), .ZN(n45540) );
  NAND2HSV0 U49451 ( .A1(\pe3/aot [8]), .A2(n55867), .ZN(n45539) );
  XOR2HSV0 U49452 ( .A1(n45540), .A2(n45539), .Z(n45544) );
  NAND2HSV0 U49453 ( .A1(n55858), .A2(\pe3/bq[11] ), .ZN(n45542) );
  CLKNAND2HSV0 U49454 ( .A1(n48500), .A2(n45639), .ZN(n45541) );
  XOR2HSV0 U49455 ( .A1(n45542), .A2(n45541), .Z(n45543) );
  XOR2HSV0 U49456 ( .A1(n45544), .A2(n45543), .Z(n45545) );
  XOR2HSV0 U49457 ( .A1(n45546), .A2(n45545), .Z(n45563) );
  NAND2HSV0 U49458 ( .A1(n46363), .A2(\pe3/bq[19] ), .ZN(n45548) );
  NAND2HSV0 U49459 ( .A1(n45952), .A2(\pe3/bq[23] ), .ZN(n45547) );
  XOR2HSV0 U49460 ( .A1(n45548), .A2(n45547), .Z(n45552) );
  CLKNAND2HSV0 U49461 ( .A1(n56188), .A2(n43146), .ZN(n45550) );
  NAND2HSV0 U49462 ( .A1(n59960), .A2(\pe3/bq[26] ), .ZN(n45549) );
  XOR2HSV0 U49463 ( .A1(n45550), .A2(n45549), .Z(n45551) );
  XOR2HSV0 U49464 ( .A1(n45552), .A2(n45551), .Z(n45561) );
  NAND2HSV0 U49465 ( .A1(n46612), .A2(\pe3/pvq [29]), .ZN(n45553) );
  XOR2HSV0 U49466 ( .A1(n45553), .A2(\pe3/phq [29]), .Z(n45559) );
  INHSV2 U49467 ( .I(n56914), .ZN(n56867) );
  NAND2HSV0 U49468 ( .A1(n56867), .A2(n45554), .ZN(n46373) );
  OAI22HSV0 U49469 ( .A1(n45691), .A2(n56914), .B1(n45555), .B2(n49272), .ZN(
        n45556) );
  OAI21HSV0 U49470 ( .A1(n46373), .A2(n45557), .B(n45556), .ZN(n45558) );
  XOR2HSV0 U49471 ( .A1(n45559), .A2(n45558), .Z(n45560) );
  XNOR2HSV1 U49472 ( .A1(n45561), .A2(n45560), .ZN(n45562) );
  CLKNAND2HSV1 U49473 ( .A1(\pe3/aot [20]), .A2(n45696), .ZN(n45566) );
  NAND2HSV0 U49474 ( .A1(n42743), .A2(n56627), .ZN(n45565) );
  XOR2HSV0 U49475 ( .A1(n45566), .A2(n45565), .Z(n45571) );
  NAND2HSV0 U49476 ( .A1(n56349), .A2(\pe3/bq[18] ), .ZN(n45569) );
  NAND2HSV0 U49477 ( .A1(\pe3/aot [22]), .A2(n48499), .ZN(n45568) );
  XOR2HSV0 U49478 ( .A1(n45569), .A2(n45568), .Z(n45570) );
  INHSV2 U49479 ( .I(n49258), .ZN(n55876) );
  NAND2HSV2 U49480 ( .A1(n37362), .A2(n55876), .ZN(n46353) );
  CLKNHSV0 U49481 ( .I(n46615), .ZN(n46323) );
  CLKNAND2HSV1 U49482 ( .A1(n42940), .A2(n46323), .ZN(n56181) );
  XOR2HSV0 U49483 ( .A1(n46353), .A2(n56181), .Z(n45575) );
  NAND2HSV0 U49484 ( .A1(\pe3/bq[4] ), .A2(n45572), .ZN(n45692) );
  NAND2HSV0 U49485 ( .A1(n45951), .A2(n56218), .ZN(n45573) );
  XOR2HSV0 U49486 ( .A1(n45692), .A2(n45573), .Z(n45574) );
  INHSV2 U49487 ( .I(n50802), .ZN(n56494) );
  NOR2HSV2 U49488 ( .A1(n45728), .A2(n45576), .ZN(n45578) );
  CLKNHSV0 U49489 ( .I(n46519), .ZN(n49468) );
  CLKNAND2HSV1 U49490 ( .A1(n49468), .A2(n56335), .ZN(n45577) );
  NOR2HSV2 U49491 ( .A1(n56475), .A2(n46533), .ZN(n45580) );
  CLKNHSV0 U49492 ( .I(n45593), .ZN(n45589) );
  INHSV1 U49493 ( .I(n45588), .ZN(n45585) );
  NAND2HSV2 U49494 ( .A1(n45586), .A2(n45585), .ZN(n45592) );
  NOR2HSV0 U49495 ( .A1(n45941), .A2(n45932), .ZN(n45587) );
  NAND3HSV2 U49496 ( .A1(n45588), .A2(pov3[24]), .A3(n45587), .ZN(n45591) );
  AOI21HSV2 U49497 ( .A1(n45596), .A2(n43591), .B(n43371), .ZN(n45597) );
  OAI21HSV2 U49498 ( .A1(n45599), .A2(n45598), .B(n45597), .ZN(n45600) );
  XNOR2HSV4 U49499 ( .A1(n45601), .A2(n45600), .ZN(n45604) );
  INHSV2 U49500 ( .I(n45604), .ZN(n45602) );
  INHSV3 U49501 ( .I(n45623), .ZN(n45626) );
  NOR2HSV1 U49502 ( .A1(n46092), .A2(n45607), .ZN(n45608) );
  CLKNAND2HSV1 U49503 ( .A1(n45626), .A2(n45608), .ZN(n46099) );
  INHSV4 U49504 ( .I(n45623), .ZN(n45614) );
  NOR2HSV4 U49505 ( .A1(n45611), .A2(n46101), .ZN(n45928) );
  CLKNAND2HSV1 U49506 ( .A1(n46092), .A2(n45612), .ZN(n45613) );
  OAI22HSV4 U49507 ( .A1(n45626), .A2(n45618), .B1(n45617), .B2(n45616), .ZN(
        n46104) );
  NAND3HSV0 U49508 ( .A1(n45927), .A2(n46104), .A3(n43484), .ZN(n45619) );
  CLKNHSV0 U49509 ( .I(n45619), .ZN(n45620) );
  NOR2HSV4 U49510 ( .A1(n60060), .A2(n45627), .ZN(n45926) );
  NOR2HSV2 U49511 ( .A1(n45926), .A2(n45628), .ZN(n45629) );
  NAND2HSV2 U49512 ( .A1(n45630), .A2(n45629), .ZN(n45631) );
  NOR2HSV2 U49513 ( .A1(n50717), .A2(n43867), .ZN(n45750) );
  CLKNAND2HSV0 U49514 ( .A1(n56063), .A2(n45633), .ZN(n45748) );
  BUFHSV2 U49515 ( .I(n46312), .Z(n55613) );
  NAND2HSV2 U49516 ( .A1(n55613), .A2(n55701), .ZN(n45746) );
  CLKNAND2HSV0 U49517 ( .A1(n56066), .A2(n48483), .ZN(n45744) );
  NAND2HSV0 U49518 ( .A1(n45636), .A2(n49404), .ZN(n45737) );
  NAND2HSV0 U49519 ( .A1(n55948), .A2(n56493), .ZN(n45726) );
  NAND2HSV0 U49520 ( .A1(n49255), .A2(n56421), .ZN(n45724) );
  NAND2HSV0 U49521 ( .A1(n56180), .A2(n56494), .ZN(n45722) );
  NAND2HSV0 U49522 ( .A1(n46313), .A2(n59644), .ZN(n45718) );
  NAND2HSV0 U49523 ( .A1(n52738), .A2(n59645), .ZN(n45716) );
  CLKNAND2HSV0 U49524 ( .A1(n48488), .A2(n56855), .ZN(n45714) );
  INHSV2 U49525 ( .I(n56859), .ZN(n56267) );
  NAND2HSV0 U49526 ( .A1(n45950), .A2(n56267), .ZN(n45659) );
  NAND2HSV0 U49527 ( .A1(n59612), .A2(n45982), .ZN(n45638) );
  NAND2HSV0 U49528 ( .A1(\pe3/aot [8]), .A2(n55960), .ZN(n45637) );
  XOR2HSV0 U49529 ( .A1(n45638), .A2(n45637), .Z(n45644) );
  CLKNAND2HSV0 U49530 ( .A1(\pe3/aot [22]), .A2(n55975), .ZN(n45642) );
  NAND2HSV0 U49531 ( .A1(n45640), .A2(n45639), .ZN(n45641) );
  XOR2HSV0 U49532 ( .A1(n45642), .A2(n45641), .Z(n45643) );
  XOR2HSV0 U49533 ( .A1(n45644), .A2(n45643), .Z(n45655) );
  NAND2HSV0 U49534 ( .A1(n55858), .A2(\pe3/bq[10] ), .ZN(n45647) );
  NAND2HSV0 U49535 ( .A1(n45645), .A2(\pe3/bq[19] ), .ZN(n45646) );
  XOR2HSV0 U49536 ( .A1(n45647), .A2(n45646), .Z(n45653) );
  NAND2HSV0 U49537 ( .A1(n45648), .A2(n55876), .ZN(n45651) );
  NAND2HSV0 U49538 ( .A1(n59627), .A2(n37280), .ZN(n45650) );
  XOR2HSV0 U49539 ( .A1(n45651), .A2(n45650), .Z(n45652) );
  XNOR2HSV1 U49540 ( .A1(n45653), .A2(n45652), .ZN(n45654) );
  XNOR2HSV1 U49541 ( .A1(n45655), .A2(n45654), .ZN(n45657) );
  NAND2HSV0 U49542 ( .A1(n59648), .A2(n56781), .ZN(n45656) );
  XNOR2HSV1 U49543 ( .A1(n45657), .A2(n45656), .ZN(n45658) );
  XNOR2HSV1 U49544 ( .A1(n45659), .A2(n45658), .ZN(n45712) );
  CLKNAND2HSV0 U49545 ( .A1(n48511), .A2(n48487), .ZN(n45709) );
  NAND2HSV0 U49546 ( .A1(n56740), .A2(n55976), .ZN(n45661) );
  NAND2HSV0 U49547 ( .A1(n56197), .A2(n43052), .ZN(n45660) );
  XOR2HSV0 U49548 ( .A1(n45661), .A2(n45660), .Z(n45667) );
  NAND2HSV0 U49549 ( .A1(n59816), .A2(n45663), .ZN(n45665) );
  NAND2HSV0 U49550 ( .A1(n45973), .A2(n48021), .ZN(n45664) );
  XOR2HSV0 U49551 ( .A1(n45665), .A2(n45664), .Z(n45666) );
  XOR2HSV0 U49552 ( .A1(n45667), .A2(n45666), .Z(n45675) );
  NAND2HSV0 U49553 ( .A1(n45951), .A2(n42971), .ZN(n45669) );
  NAND2HSV0 U49554 ( .A1(n46363), .A2(\pe3/bq[18] ), .ZN(n45668) );
  XOR2HSV0 U49555 ( .A1(n45669), .A2(n45668), .Z(n45673) );
  NOR2HSV0 U49556 ( .A1(n42539), .A2(n49281), .ZN(n45671) );
  NAND2HSV0 U49557 ( .A1(n59622), .A2(\pe3/bq[8] ), .ZN(n45670) );
  XOR2HSV0 U49558 ( .A1(n45671), .A2(n45670), .Z(n45672) );
  XOR2HSV0 U49559 ( .A1(n45673), .A2(n45672), .Z(n45674) );
  XOR2HSV0 U49560 ( .A1(n45675), .A2(n45674), .Z(n45690) );
  NAND2HSV0 U49561 ( .A1(n37362), .A2(n56189), .ZN(n45678) );
  NAND2HSV0 U49562 ( .A1(n45676), .A2(\pe3/bq[23] ), .ZN(n45677) );
  XOR2HSV0 U49563 ( .A1(n45678), .A2(n45677), .Z(n45682) );
  NOR2HSV0 U49564 ( .A1(n37357), .A2(n46615), .ZN(n45680) );
  NAND2HSV0 U49565 ( .A1(\pe3/got [3]), .A2(n45955), .ZN(n45679) );
  XOR2HSV0 U49566 ( .A1(n45680), .A2(n45679), .Z(n45681) );
  XOR2HSV0 U49567 ( .A1(n45682), .A2(n45681), .Z(n45688) );
  NAND2HSV0 U49568 ( .A1(n56520), .A2(\pe3/bq[26] ), .ZN(n45684) );
  NAND2HSV0 U49569 ( .A1(n56188), .A2(n56106), .ZN(n45683) );
  XOR2HSV0 U49570 ( .A1(n45684), .A2(n45683), .Z(n45686) );
  CLKNHSV0 U49571 ( .I(n46613), .ZN(n48019) );
  XNOR2HSV1 U49572 ( .A1(n45686), .A2(n45685), .ZN(n45687) );
  XNOR2HSV1 U49573 ( .A1(n45688), .A2(n45687), .ZN(n45689) );
  XNOR2HSV1 U49574 ( .A1(n45690), .A2(n45689), .ZN(n45707) );
  NAND2HSV0 U49575 ( .A1(\pe3/aot [18]), .A2(n55616), .ZN(n56435) );
  NOR2HSV0 U49576 ( .A1(n45691), .A2(n50722), .ZN(n46005) );
  CLKNHSV0 U49577 ( .I(n45692), .ZN(n45694) );
  AOI22HSV0 U49578 ( .A1(n45962), .A2(\pe3/bq[3] ), .B1(n43265), .B2(
        \pe3/bq[4] ), .ZN(n45693) );
  AOI21HSV2 U49579 ( .A1(n46005), .A2(n45694), .B(n45693), .ZN(n45698) );
  BUFHSV2 U49580 ( .I(n45695), .Z(n56087) );
  CLKNAND2HSV0 U49581 ( .A1(n56087), .A2(\pe3/bq[11] ), .ZN(n55635) );
  NAND2HSV0 U49582 ( .A1(\pe3/aot [19]), .A2(n45696), .ZN(n56463) );
  XOR2HSV0 U49583 ( .A1(n55635), .A2(n56463), .Z(n45697) );
  XOR3HSV2 U49584 ( .A1(n56435), .A2(n45698), .A3(n45697), .Z(n45705) );
  NAND2HSV0 U49585 ( .A1(n53250), .A2(n46614), .ZN(n45700) );
  NAND2HSV0 U49586 ( .A1(n42743), .A2(n56785), .ZN(n45699) );
  XOR2HSV0 U49587 ( .A1(n45700), .A2(n45699), .Z(n45703) );
  NAND2HSV0 U49588 ( .A1(\pe3/aot [4]), .A2(n48538), .ZN(n46350) );
  NAND2HSV0 U49589 ( .A1(n45952), .A2(n43146), .ZN(n45701) );
  XOR2HSV0 U49590 ( .A1(n46350), .A2(n45701), .Z(n45702) );
  XOR2HSV0 U49591 ( .A1(n45703), .A2(n45702), .Z(n45704) );
  XOR2HSV0 U49592 ( .A1(n45705), .A2(n45704), .Z(n45706) );
  XNOR2HSV1 U49593 ( .A1(n45707), .A2(n45706), .ZN(n45708) );
  XNOR2HSV1 U49594 ( .A1(n45709), .A2(n45708), .ZN(n45711) );
  NAND2HSV0 U49595 ( .A1(n52727), .A2(n59647), .ZN(n45710) );
  XOR3HSV2 U49596 ( .A1(n45712), .A2(n45711), .A3(n45710), .Z(n45713) );
  XNOR2HSV1 U49597 ( .A1(n45714), .A2(n45713), .ZN(n45715) );
  XNOR2HSV1 U49598 ( .A1(n45716), .A2(n45715), .ZN(n45717) );
  XNOR2HSV1 U49599 ( .A1(n45718), .A2(n45717), .ZN(n45720) );
  NAND2HSV0 U49600 ( .A1(n55895), .A2(n59967), .ZN(n45719) );
  XNOR2HSV1 U49601 ( .A1(n45720), .A2(n45719), .ZN(n45721) );
  XNOR2HSV1 U49602 ( .A1(n45722), .A2(n45721), .ZN(n45723) );
  XNOR2HSV1 U49603 ( .A1(n45724), .A2(n45723), .ZN(n45725) );
  XNOR2HSV1 U49604 ( .A1(n45726), .A2(n45725), .ZN(n45731) );
  NOR2HSV0 U49605 ( .A1(n45728), .A2(n45727), .ZN(n45730) );
  CLKNHSV0 U49606 ( .I(n46519), .ZN(n56392) );
  CLKNAND2HSV1 U49607 ( .A1(n56392), .A2(n56065), .ZN(n45729) );
  XOR3HSV1 U49608 ( .A1(n45731), .A2(n45730), .A3(n45729), .Z(n45735) );
  NOR2HSV1 U49609 ( .A1(n56475), .A2(n44693), .ZN(n45734) );
  NAND2HSV0 U49610 ( .A1(n45732), .A2(\pe3/got [18]), .ZN(n45733) );
  XOR3HSV2 U49611 ( .A1(n45735), .A2(n45734), .A3(n45733), .Z(n45736) );
  XNOR2HSV1 U49612 ( .A1(n45737), .A2(n45736), .ZN(n45739) );
  NAND2HSV0 U49613 ( .A1(n46052), .A2(\pe3/got [19]), .ZN(n45738) );
  XNOR2HSV1 U49614 ( .A1(n45739), .A2(n45738), .ZN(n45742) );
  CLKNAND2HSV0 U49615 ( .A1(n53228), .A2(n55945), .ZN(n45741) );
  NAND2HSV0 U49616 ( .A1(n45582), .A2(n48485), .ZN(n45740) );
  XOR3HSV2 U49617 ( .A1(n45742), .A2(n45741), .A3(n45740), .Z(n45743) );
  XNOR2HSV1 U49618 ( .A1(n45744), .A2(n45743), .ZN(n45745) );
  XOR2HSV0 U49619 ( .A1(n45746), .A2(n45745), .Z(n45747) );
  XOR2HSV2 U49620 ( .A1(n45750), .A2(n45749), .Z(n45751) );
  XNOR2HSV4 U49621 ( .A1(n45752), .A2(n45751), .ZN(n45770) );
  CLKNAND2HSV1 U49622 ( .A1(n45754), .A2(n45753), .ZN(n45759) );
  CLKNAND2HSV0 U49623 ( .A1(n45756), .A2(n45755), .ZN(n45757) );
  AND2HSV2 U49624 ( .A1(n45760), .A2(n46107), .Z(n45761) );
  NAND3HSV2 U49625 ( .A1(n45763), .A2(n45762), .A3(n45761), .ZN(n45764) );
  INHSV2 U49626 ( .I(n45770), .ZN(n45768) );
  NAND2HSV2 U49627 ( .A1(n45768), .A2(n45767), .ZN(n45775) );
  CLKNAND2HSV1 U49628 ( .A1(n45770), .A2(n45769), .ZN(n45774) );
  NOR2HSV2 U49629 ( .A1(n45772), .A2(n45771), .ZN(n45773) );
  INHSV4 U49630 ( .I(n45930), .ZN(n45936) );
  XNOR2HSV4 U49631 ( .A1(n45778), .A2(n45936), .ZN(n60001) );
  NAND2HSV2 U49632 ( .A1(\pe3/ti_7t [30]), .A2(n47428), .ZN(n47429) );
  BUFHSV2 U49633 ( .I(n56260), .Z(n59823) );
  NAND2HSV2 U49634 ( .A1(n29654), .A2(n53519), .ZN(n55226) );
  CLKNHSV2 U49635 ( .I(n45784), .ZN(n45785) );
  AOI21HSV2 U49636 ( .A1(n45787), .A2(n45786), .B(n45785), .ZN(n45791) );
  INHSV2 U49637 ( .I(n45787), .ZN(n45789) );
  NAND2HSV2 U49638 ( .A1(n45789), .A2(n45788), .ZN(n45790) );
  INHSV2 U49639 ( .I(n46156), .ZN(n49401) );
  INHSV2 U49640 ( .I(n45147), .ZN(n59475) );
  CLKBUFHSV4 U49641 ( .I(n46310), .Z(n56420) );
  XNOR2HSV0 U49642 ( .A1(n45793), .A2(n45792), .ZN(n60053) );
  BUFHSV4 U49643 ( .I(n47865), .Z(n59837) );
  BUFHSV2 U49644 ( .I(n45795), .Z(n59769) );
  BUFHSV2 U49645 ( .I(n45800), .Z(n59871) );
  BUFHSV2 U49646 ( .I(n45801), .Z(n59833) );
  XOR2HSV0 U49647 ( .A1(n45803), .A2(n45802), .Z(n45805) );
  XNOR2HSV0 U49648 ( .A1(n45805), .A2(n45804), .ZN(n60049) );
  BUFHSV2 U49649 ( .I(n34595), .Z(n59681) );
  CLKNHSV0 U49650 ( .I(n50091), .ZN(n59832) );
  MUX2HSV1 U49651 ( .I0(bo3[22]), .I1(n45807), .S(n59537), .Z(n59762) );
  MUX2HSV1 U49652 ( .I0(bo3[13]), .I1(n56460), .S(n45808), .Z(n59788) );
  MUX2HSV1 U49653 ( .I0(bo3[14]), .I1(n48499), .S(n46129), .Z(n59787) );
  MUX2HSV1 U49654 ( .I0(bo3[18]), .I1(\pe3/bq[18] ), .S(n45809), .Z(n59559) );
  MUX2HSV1 U49655 ( .I0(bo3[20]), .I1(n42971), .S(n46132), .Z(n59771) );
  MUX2HSV1 U49656 ( .I0(bo5[21]), .I1(n48206), .S(n37707), .Z(n59847) );
  MUX2HSV1 U49657 ( .I0(bo4[22]), .I1(n34044), .S(n48072), .Z(n59813) );
  BUFHSV2 U49658 ( .I(n45811), .Z(n48052) );
  MUX2HSV1 U49659 ( .I0(bo2[22]), .I1(n38054), .S(n48057), .Z(n59734) );
  BUFHSV2 U49660 ( .I(n45811), .Z(n46619) );
  MUX2HSV1 U49661 ( .I0(bo2[31]), .I1(n36607), .S(n46619), .Z(n59722) );
  MUX2HSV1 U49662 ( .I0(bo2[20]), .I1(n51998), .S(n53225), .Z(n59738) );
  MUX2HSV1 U49663 ( .I0(bo6[27]), .I1(n45812), .S(n46621), .Z(n59876) );
  MUX2HSV1 U49664 ( .I0(bo6[30]), .I1(n59071), .S(n48025), .Z(n59870) );
  MUX2HSV1 U49665 ( .I0(bo3[10]), .I1(n56627), .S(n46140), .Z(n59784) );
  MUX2HSV1 U49666 ( .I0(bo6[21]), .I1(n45813), .S(n48025), .Z(n59886) );
  MUX2HSV1 U49667 ( .I0(bo1[16]), .I1(n55100), .S(n48054), .Z(n59705) );
  INHSV2 U49668 ( .I(n47139), .ZN(n53287) );
  INHSV2 U49669 ( .I(n25830), .ZN(n53288) );
  INHSV2 U49670 ( .I(n46976), .ZN(n53290) );
  CLKNAND2HSV1 U49671 ( .A1(n53291), .A2(n52658), .ZN(n45897) );
  NOR2HSV0 U49672 ( .A1(n47057), .A2(n45817), .ZN(n45892) );
  BUFHSV2 U49673 ( .I(n45818), .Z(n53294) );
  INHSV2 U49674 ( .I(n47143), .ZN(n53349) );
  NAND2HSV0 U49675 ( .A1(n53294), .A2(n53349), .ZN(n45888) );
  NAND2HSV0 U49676 ( .A1(n52570), .A2(n53289), .ZN(n45886) );
  NAND2HSV0 U49677 ( .A1(n51018), .A2(n47144), .ZN(n45882) );
  BUFHSV2 U49678 ( .I(n45819), .Z(n59878) );
  NAND2HSV0 U49679 ( .A1(n59878), .A2(n51200), .ZN(n45878) );
  NAND2HSV0 U49680 ( .A1(n45820), .A2(n52576), .ZN(n45876) );
  BUFHSV2 U49681 ( .I(n59871), .Z(n52575) );
  NAND2HSV0 U49682 ( .A1(n52575), .A2(n51302), .ZN(n45874) );
  NAND2HSV0 U49683 ( .A1(n29770), .A2(n53211), .ZN(n45872) );
  NAND2HSV0 U49684 ( .A1(n52578), .A2(\pe5/got [2]), .ZN(n45870) );
  NAND2HSV0 U49685 ( .A1(n59381), .A2(n51362), .ZN(n45868) );
  NAND2HSV0 U49686 ( .A1(n59880), .A2(n51176), .ZN(n45823) );
  INHSV2 U49687 ( .I(n48204), .ZN(n53323) );
  NAND2HSV0 U49688 ( .A1(n53323), .A2(n39472), .ZN(n45822) );
  XOR2HSV0 U49689 ( .A1(n45823), .A2(n45822), .Z(n45827) );
  CLKNHSV0 U49690 ( .I(n48822), .ZN(n52618) );
  NAND2HSV0 U49691 ( .A1(n53304), .A2(n52618), .ZN(n45825) );
  NAND2HSV0 U49692 ( .A1(\pe5/aot [10]), .A2(n53314), .ZN(n45824) );
  XOR2HSV0 U49693 ( .A1(n45825), .A2(n45824), .Z(n45826) );
  XOR2HSV0 U49694 ( .A1(n45827), .A2(n45826), .Z(n45835) );
  NAND2HSV0 U49695 ( .A1(n52584), .A2(n39471), .ZN(n45829) );
  INHSV2 U49696 ( .I(n45904), .ZN(n59895) );
  NAND2HSV0 U49697 ( .A1(n59895), .A2(n30891), .ZN(n45828) );
  XOR2HSV0 U49698 ( .A1(n45829), .A2(n45828), .Z(n45833) );
  NAND2HSV0 U49699 ( .A1(n39887), .A2(\pe5/bq[16] ), .ZN(n45831) );
  CLKNHSV0 U49700 ( .I(n50518), .ZN(n52607) );
  NAND2HSV0 U49701 ( .A1(n52607), .A2(n52672), .ZN(n45830) );
  XOR2HSV0 U49702 ( .A1(n45831), .A2(n45830), .Z(n45832) );
  XOR2HSV0 U49703 ( .A1(n45833), .A2(n45832), .Z(n45834) );
  XOR2HSV0 U49704 ( .A1(n45835), .A2(n45834), .Z(n45850) );
  CLKNHSV0 U49705 ( .I(n45451), .ZN(n52631) );
  NAND2HSV0 U49706 ( .A1(n52631), .A2(n53200), .ZN(n45837) );
  NAND2HSV0 U49707 ( .A1(n40190), .A2(n51191), .ZN(n45836) );
  XOR2HSV0 U49708 ( .A1(n45837), .A2(n45836), .Z(n45841) );
  NAND2HSV0 U49709 ( .A1(\pe5/aot [16]), .A2(n51307), .ZN(n45839) );
  NAND2HSV0 U49710 ( .A1(\pe5/aot [13]), .A2(\pe5/bq[12] ), .ZN(n45838) );
  XOR2HSV0 U49711 ( .A1(n45839), .A2(n45838), .Z(n45840) );
  XOR2HSV0 U49712 ( .A1(n45841), .A2(n45840), .Z(n45848) );
  NAND2HSV0 U49713 ( .A1(\pe5/aot [4]), .A2(n46933), .ZN(n45843) );
  NAND2HSV0 U49714 ( .A1(n51310), .A2(\pe5/bq[19] ), .ZN(n45842) );
  XOR2HSV0 U49715 ( .A1(n45843), .A2(n45842), .Z(n45846) );
  NOR2HSV0 U49716 ( .A1(n47409), .A2(n45426), .ZN(n47303) );
  NAND2HSV0 U49717 ( .A1(\pe5/aot [3]), .A2(n48237), .ZN(n46920) );
  CLKNHSV0 U49718 ( .I(n47409), .ZN(n52623) );
  CLKNHSV0 U49719 ( .I(n45844), .ZN(n47291) );
  NAND2HSV0 U49720 ( .A1(n52623), .A2(n47291), .ZN(n52627) );
  XNOR2HSV1 U49721 ( .A1(n45846), .A2(n45845), .ZN(n45847) );
  XNOR2HSV1 U49722 ( .A1(n45848), .A2(n45847), .ZN(n45849) );
  XNOR2HSV1 U49723 ( .A1(n45850), .A2(n45849), .ZN(n45866) );
  NAND2HSV0 U49724 ( .A1(n59943), .A2(n48170), .ZN(n45852) );
  NAND2HSV0 U49725 ( .A1(n59940), .A2(n52581), .ZN(n45851) );
  XOR2HSV0 U49726 ( .A1(n45852), .A2(n45851), .Z(n45856) );
  NAND2HSV0 U49727 ( .A1(n52591), .A2(n52630), .ZN(n45854) );
  BUFHSV2 U49728 ( .I(\pe5/bq[4] ), .Z(n53307) );
  NAND2HSV0 U49729 ( .A1(n48242), .A2(n53307), .ZN(n45853) );
  XOR2HSV0 U49730 ( .A1(n45854), .A2(n45853), .Z(n45855) );
  XOR2HSV0 U49731 ( .A1(n45856), .A2(n45855), .Z(n45864) );
  NOR2HSV0 U49732 ( .A1(n51232), .A2(n37564), .ZN(n47238) );
  NAND2HSV0 U49733 ( .A1(n48681), .A2(\pe5/bq[11] ), .ZN(n45857) );
  XOR2HSV0 U49734 ( .A1(n47238), .A2(n45857), .Z(n45862) );
  NOR2HSV0 U49735 ( .A1(n45858), .A2(n47207), .ZN(n45860) );
  NAND2HSV0 U49736 ( .A1(\pe5/aot [23]), .A2(\pe5/bq[2] ), .ZN(n45859) );
  XOR2HSV0 U49737 ( .A1(n45860), .A2(n45859), .Z(n45861) );
  XOR2HSV0 U49738 ( .A1(n45862), .A2(n45861), .Z(n45863) );
  XOR2HSV0 U49739 ( .A1(n45864), .A2(n45863), .Z(n45865) );
  XNOR2HSV1 U49740 ( .A1(n45866), .A2(n45865), .ZN(n45867) );
  XNOR2HSV1 U49741 ( .A1(n45868), .A2(n45867), .ZN(n45869) );
  XNOR2HSV1 U49742 ( .A1(n45870), .A2(n45869), .ZN(n45871) );
  XNOR2HSV1 U49743 ( .A1(n45872), .A2(n45871), .ZN(n45873) );
  XNOR2HSV1 U49744 ( .A1(n45874), .A2(n45873), .ZN(n45875) );
  XNOR2HSV1 U49745 ( .A1(n45876), .A2(n45875), .ZN(n45877) );
  XNOR2HSV1 U49746 ( .A1(n45878), .A2(n45877), .ZN(n45880) );
  NAND2HSV0 U49747 ( .A1(n44694), .A2(n51359), .ZN(n45879) );
  XOR2HSV0 U49748 ( .A1(n45880), .A2(n45879), .Z(n45881) );
  XNOR2HSV1 U49749 ( .A1(n45882), .A2(n45881), .ZN(n45884) );
  CLKNHSV0 U49750 ( .I(n51205), .ZN(n50617) );
  NOR2HSV0 U49751 ( .A1(n50617), .A2(n46119), .ZN(n45883) );
  XNOR2HSV1 U49752 ( .A1(n45884), .A2(n45883), .ZN(n45885) );
  XNOR2HSV1 U49753 ( .A1(n45886), .A2(n45885), .ZN(n45887) );
  XNOR2HSV1 U49754 ( .A1(n45888), .A2(n45887), .ZN(n45890) );
  NAND2HSV0 U49755 ( .A1(n52653), .A2(n48167), .ZN(n45889) );
  XNOR2HSV1 U49756 ( .A1(n45890), .A2(n45889), .ZN(n45891) );
  XNOR2HSV1 U49757 ( .A1(n45892), .A2(n45891), .ZN(n45895) );
  INHSV2 U49758 ( .I(n51217), .ZN(n53338) );
  CLKNAND2HSV0 U49759 ( .A1(n53338), .A2(n53285), .ZN(n45894) );
  NOR2HSV2 U49760 ( .A1(n51273), .A2(n48722), .ZN(n45893) );
  XOR3HSV2 U49761 ( .A1(n45895), .A2(n45894), .A3(n45893), .Z(n45896) );
  XNOR2HSV1 U49762 ( .A1(n45897), .A2(n45896), .ZN(n45899) );
  NAND2HSV0 U49763 ( .A1(n59516), .A2(n59949), .ZN(n45898) );
  NAND2HSV2 U49764 ( .A1(n51230), .A2(n51229), .ZN(n53198) );
  INHSV2 U49765 ( .I(n45902), .ZN(n47926) );
  INHSV2 U49766 ( .I(n47926), .ZN(n52669) );
  INHSV2 U49767 ( .I(n46976), .ZN(n47268) );
  NAND2HSV0 U49768 ( .A1(n59893), .A2(\pe5/got [1]), .ZN(n45920) );
  CLKNAND2HSV1 U49769 ( .A1(n59895), .A2(n48775), .ZN(n45906) );
  BUFHSV2 U49770 ( .I(\pe5/aot [6]), .Z(n51310) );
  NAND2HSV0 U49771 ( .A1(n51310), .A2(n51336), .ZN(n45905) );
  XOR2HSV0 U49772 ( .A1(n45906), .A2(n45905), .Z(n45918) );
  NAND2HSV0 U49773 ( .A1(\pe5/aot [3]), .A2(\pe5/bq[7] ), .ZN(n45908) );
  INHSV2 U49774 ( .I(n48031), .ZN(n51420) );
  NAND2HSV0 U49775 ( .A1(n51247), .A2(n51420), .ZN(n45907) );
  XOR2HSV0 U49776 ( .A1(n45908), .A2(n45907), .Z(n45909) );
  NAND2HSV2 U49777 ( .A1(n51363), .A2(n48686), .ZN(n48176) );
  XNOR2HSV1 U49778 ( .A1(n45909), .A2(n48176), .ZN(n45917) );
  NAND2HSV0 U49779 ( .A1(n50501), .A2(\pe5/bq[6] ), .ZN(n45911) );
  NAND2HSV0 U49780 ( .A1(n50511), .A2(\pe5/bq[2] ), .ZN(n45910) );
  XOR2HSV0 U49781 ( .A1(n45911), .A2(n45910), .Z(n45915) );
  NAND2HSV0 U49782 ( .A1(n53203), .A2(n50675), .ZN(n45913) );
  INHSV2 U49783 ( .I(\pe5/bq[1] ), .ZN(n51235) );
  NAND2HSV0 U49784 ( .A1(n39887), .A2(n51276), .ZN(n45912) );
  XOR2HSV0 U49785 ( .A1(n45913), .A2(n45912), .Z(n45914) );
  XOR2HSV0 U49786 ( .A1(n45915), .A2(n45914), .Z(n45916) );
  XOR3HSV2 U49787 ( .A1(n45918), .A2(n45917), .A3(n45916), .Z(n45919) );
  XNOR2HSV1 U49788 ( .A1(n45920), .A2(n45919), .ZN(n45922) );
  CLKNHSV0 U49789 ( .I(n39992), .ZN(n51399) );
  CLKNAND2HSV0 U49790 ( .A1(n51399), .A2(n51161), .ZN(n45921) );
  INHSV4 U49791 ( .I(n59535), .ZN(n45923) );
  INHSV6 U49792 ( .I(n45923), .ZN(n51404) );
  INHSV2 U49793 ( .I(n46118), .ZN(n47496) );
  NOR2HSV4 U49794 ( .A1(n46116), .A2(n46114), .ZN(n45940) );
  OAI22HSV2 U49795 ( .A1(n45935), .A2(n46114), .B1(n45934), .B2(n45933), .ZN(
        n45937) );
  AOI21HSV4 U49796 ( .A1(n55820), .A2(n45940), .B(n45939), .ZN(n46113) );
  NAND2HSV2 U49797 ( .A1(n56863), .A2(n37516), .ZN(n46070) );
  BUFHSV2 U49798 ( .I(n55612), .Z(n50718) );
  INHSV2 U49799 ( .I(n50718), .ZN(n48482) );
  NAND2HSV2 U49800 ( .A1(n48482), .A2(n45947), .ZN(n46068) );
  INAND2HSV2 U49801 ( .A1(n48484), .B1(n42508), .ZN(n46066) );
  CLKNAND2HSV0 U49802 ( .A1(n49253), .A2(n43452), .ZN(n46064) );
  NAND2HSV0 U49803 ( .A1(n46312), .A2(n48483), .ZN(n46062) );
  CLKNAND2HSV0 U49804 ( .A1(n56066), .A2(n48485), .ZN(n46060) );
  NAND2HSV2 U49805 ( .A1(n55947), .A2(n49404), .ZN(n46056) );
  CLKNHSV0 U49806 ( .I(n47430), .ZN(n56178) );
  CLKNAND2HSV1 U49807 ( .A1(n56178), .A2(n59965), .ZN(n46051) );
  NAND2HSV0 U49808 ( .A1(n55948), .A2(n56421), .ZN(n46041) );
  BUFHSV2 U49809 ( .I(n49255), .Z(n56179) );
  NAND2HSV0 U49810 ( .A1(n56179), .A2(n56494), .ZN(n46039) );
  NAND2HSV0 U49811 ( .A1(n56180), .A2(n56557), .ZN(n46037) );
  NAND2HSV0 U49812 ( .A1(n45949), .A2(n56855), .ZN(n46030) );
  NAND2HSV0 U49813 ( .A1(n46314), .A2(n59647), .ZN(n46028) );
  NAND2HSV0 U49814 ( .A1(n45950), .A2(n56684), .ZN(n45972) );
  NAND2HSV0 U49815 ( .A1(n45951), .A2(\pe3/bq[19] ), .ZN(n45954) );
  NAND2HSV0 U49816 ( .A1(n45952), .A2(n56106), .ZN(n45953) );
  XOR2HSV0 U49817 ( .A1(n45954), .A2(n45953), .Z(n45959) );
  NAND2HSV0 U49818 ( .A1(n59627), .A2(n55960), .ZN(n45957) );
  CLKNHSV0 U49819 ( .I(n56936), .ZN(n55950) );
  NAND2HSV0 U49820 ( .A1(n55950), .A2(n45955), .ZN(n45956) );
  XOR2HSV0 U49821 ( .A1(n45957), .A2(n45956), .Z(n45958) );
  XOR2HSV0 U49822 ( .A1(n45959), .A2(n45958), .Z(n45968) );
  CLKNAND2HSV1 U49823 ( .A1(n42818), .A2(\pe3/bq[11] ), .ZN(n45961) );
  NAND2HSV0 U49824 ( .A1(n56087), .A2(\pe3/bq[10] ), .ZN(n45960) );
  XOR2HSV0 U49825 ( .A1(n45961), .A2(n45960), .Z(n45966) );
  INHSV2 U49826 ( .I(n48495), .ZN(n56969) );
  NAND2HSV0 U49827 ( .A1(n45962), .A2(n56969), .ZN(n45964) );
  NAND2HSV0 U49828 ( .A1(n36809), .A2(\pe3/bq[7] ), .ZN(n45963) );
  XOR2HSV0 U49829 ( .A1(n45964), .A2(n45963), .Z(n45965) );
  XOR2HSV0 U49830 ( .A1(n45966), .A2(n45965), .Z(n45967) );
  XOR2HSV0 U49831 ( .A1(n45968), .A2(n45967), .Z(n45970) );
  NAND2HSV0 U49832 ( .A1(n59648), .A2(n56735), .ZN(n45969) );
  XNOR2HSV1 U49833 ( .A1(n45970), .A2(n45969), .ZN(n45971) );
  XNOR2HSV1 U49834 ( .A1(n45972), .A2(n45971), .ZN(n46026) );
  INHSV2 U49835 ( .I(n56914), .ZN(n56428) );
  NAND2HSV0 U49836 ( .A1(n48500), .A2(n56428), .ZN(n45975) );
  NAND2HSV0 U49837 ( .A1(n45973), .A2(n43539), .ZN(n45974) );
  XOR2HSV0 U49838 ( .A1(n45975), .A2(n45974), .Z(n45979) );
  NAND2HSV0 U49839 ( .A1(\pe3/aot [3]), .A2(n48538), .ZN(n45977) );
  NAND2HSV0 U49840 ( .A1(\pe3/aot [5]), .A2(n48021), .ZN(n45976) );
  XOR2HSV0 U49841 ( .A1(n45977), .A2(n45976), .Z(n45978) );
  XOR2HSV0 U49842 ( .A1(n45979), .A2(n45978), .Z(n45988) );
  NAND2HSV0 U49843 ( .A1(n37362), .A2(\pe3/bq[4] ), .ZN(n45981) );
  NAND2HSV0 U49844 ( .A1(n59960), .A2(n55872), .ZN(n45980) );
  XOR2HSV0 U49845 ( .A1(n45981), .A2(n45980), .Z(n45986) );
  NAND2HSV0 U49846 ( .A1(\pe3/aot [4]), .A2(n48522), .ZN(n45984) );
  NAND2HSV0 U49847 ( .A1(\pe3/aot [22]), .A2(n45982), .ZN(n45983) );
  XOR2HSV0 U49848 ( .A1(n45984), .A2(n45983), .Z(n45985) );
  XOR2HSV0 U49849 ( .A1(n45986), .A2(n45985), .Z(n45987) );
  XOR2HSV0 U49850 ( .A1(n45988), .A2(n45987), .Z(n46004) );
  BUFHSV2 U49851 ( .I(\pe3/bq[18] ), .Z(n55727) );
  NAND2HSV2 U49852 ( .A1(\pe3/aot [16]), .A2(n55727), .ZN(n45990) );
  NAND2HSV0 U49853 ( .A1(n42728), .A2(n46323), .ZN(n45989) );
  XOR2HSV0 U49854 ( .A1(n45990), .A2(n45989), .Z(n45994) );
  NAND2HSV0 U49855 ( .A1(n56188), .A2(n42971), .ZN(n45992) );
  NAND2HSV0 U49856 ( .A1(n56972), .A2(n46614), .ZN(n45991) );
  XOR2HSV0 U49857 ( .A1(n45992), .A2(n45991), .Z(n45993) );
  XOR2HSV0 U49858 ( .A1(n45994), .A2(n45993), .Z(n46002) );
  NOR2HSV0 U49859 ( .A1(n42539), .A2(n49423), .ZN(n45996) );
  NAND2HSV0 U49860 ( .A1(\pe3/aot [20]), .A2(n48499), .ZN(n45995) );
  XOR2HSV0 U49861 ( .A1(n45996), .A2(n45995), .Z(n46000) );
  NAND2HSV0 U49862 ( .A1(n56197), .A2(\pe3/bq[23] ), .ZN(n45998) );
  CLKNHSV0 U49863 ( .I(n53229), .ZN(n56370) );
  NAND2HSV0 U49864 ( .A1(n56370), .A2(n43146), .ZN(n45997) );
  XOR2HSV0 U49865 ( .A1(n45998), .A2(n45997), .Z(n45999) );
  XOR2HSV0 U49866 ( .A1(n46000), .A2(n45999), .Z(n46001) );
  XOR2HSV0 U49867 ( .A1(n46002), .A2(n46001), .Z(n46003) );
  XOR2HSV0 U49868 ( .A1(n46004), .A2(n46003), .Z(n46021) );
  CLKNHSV1 U49869 ( .I(n46005), .ZN(n46006) );
  NAND2HSV0 U49870 ( .A1(n55876), .A2(n55750), .ZN(n46483) );
  XOR2HSV0 U49871 ( .A1(n46006), .A2(n46483), .Z(n46019) );
  NAND2HSV0 U49872 ( .A1(n48020), .A2(\pe3/pvq [31]), .ZN(n46007) );
  XOR2HSV0 U49873 ( .A1(n46007), .A2(\pe3/phq [31]), .Z(n46010) );
  OAI22HSV0 U49874 ( .A1(n56295), .A2(n46138), .B1(n43527), .B2(n55755), .ZN(
        n46008) );
  OAI21HSV0 U49875 ( .A1(n56435), .A2(n46364), .B(n46008), .ZN(n46009) );
  XNOR2HSV1 U49876 ( .A1(n46010), .A2(n46009), .ZN(n46018) );
  NAND2HSV0 U49877 ( .A1(n42743), .A2(n56454), .ZN(n46012) );
  NAND2HSV0 U49878 ( .A1(n59808), .A2(n56071), .ZN(n46011) );
  XOR2HSV0 U49879 ( .A1(n46012), .A2(n46011), .Z(n46016) );
  NAND2HSV0 U49880 ( .A1(\pe3/aot [8]), .A2(\pe3/bq[26] ), .ZN(n46013) );
  XOR2HSV0 U49881 ( .A1(n46014), .A2(n46013), .Z(n46015) );
  XOR2HSV0 U49882 ( .A1(n46016), .A2(n46015), .Z(n46017) );
  XOR3HSV2 U49883 ( .A1(n46019), .A2(n46018), .A3(n46017), .Z(n46020) );
  XNOR2HSV1 U49884 ( .A1(n46021), .A2(n46020), .ZN(n46023) );
  NAND2HSV0 U49885 ( .A1(n48511), .A2(n59799), .ZN(n46022) );
  XNOR2HSV1 U49886 ( .A1(n46023), .A2(n46022), .ZN(n46025) );
  NAND2HSV0 U49887 ( .A1(n55826), .A2(n48487), .ZN(n46024) );
  XOR3HSV2 U49888 ( .A1(n46026), .A2(n46025), .A3(n46024), .Z(n46027) );
  XOR2HSV0 U49889 ( .A1(n46028), .A2(n46027), .Z(n46029) );
  XOR2HSV0 U49890 ( .A1(n46030), .A2(n46029), .Z(n46033) );
  BUFHSV2 U49891 ( .I(n42767), .Z(n56070) );
  NAND2HSV0 U49892 ( .A1(n56070), .A2(n59645), .ZN(n46032) );
  XNOR2HSV1 U49893 ( .A1(n46033), .A2(n46032), .ZN(n46035) );
  NAND2HSV0 U49894 ( .A1(n56127), .A2(n59644), .ZN(n46034) );
  XNOR2HSV1 U49895 ( .A1(n46035), .A2(n46034), .ZN(n46036) );
  XNOR2HSV1 U49896 ( .A1(n46037), .A2(n46036), .ZN(n46038) );
  XNOR2HSV1 U49897 ( .A1(n46039), .A2(n46038), .ZN(n46040) );
  XNOR2HSV1 U49898 ( .A1(n46041), .A2(n46040), .ZN(n46046) );
  NOR2HSV1 U49899 ( .A1(n56391), .A2(n46042), .ZN(n46045) );
  NAND2HSV0 U49900 ( .A1(n46043), .A2(n48584), .ZN(n46044) );
  XOR3HSV2 U49901 ( .A1(n46046), .A2(n46045), .A3(n46044), .Z(n46049) );
  CLKNHSV0 U49902 ( .I(n59362), .ZN(n48583) );
  NOR2HSV2 U49903 ( .A1(n48583), .A2(n45576), .ZN(n46048) );
  NAND2HSV0 U49904 ( .A1(n59810), .A2(n56335), .ZN(n46047) );
  XOR3HSV2 U49905 ( .A1(n46049), .A2(n46048), .A3(n46047), .Z(n46050) );
  XNOR2HSV1 U49906 ( .A1(n46051), .A2(n46050), .ZN(n46054) );
  NAND2HSV0 U49907 ( .A1(n46052), .A2(\pe3/got [18]), .ZN(n46053) );
  XOR2HSV0 U49908 ( .A1(n46054), .A2(n46053), .Z(n46055) );
  XNOR2HSV1 U49909 ( .A1(n46056), .A2(n46055), .ZN(n46058) );
  CLKNHSV1 U49910 ( .I(n55917), .ZN(n56662) );
  CLKNAND2HSV1 U49911 ( .A1(n56662), .A2(n56171), .ZN(n46057) );
  XNOR2HSV1 U49912 ( .A1(n46058), .A2(n46057), .ZN(n46059) );
  XNOR2HSV1 U49913 ( .A1(n46060), .A2(n46059), .ZN(n46061) );
  XNOR2HSV1 U49914 ( .A1(n46062), .A2(n46061), .ZN(n46063) );
  XNOR2HSV1 U49915 ( .A1(n46064), .A2(n46063), .ZN(n46065) );
  XNOR2HSV1 U49916 ( .A1(n46066), .A2(n46065), .ZN(n46067) );
  XNOR2HSV1 U49917 ( .A1(n46068), .A2(n46067), .ZN(n46069) );
  CLKNAND2HSV1 U49918 ( .A1(n46073), .A2(n46074), .ZN(n46078) );
  NAND3HSV2 U49919 ( .A1(n46078), .A2(n46077), .A3(n46076), .ZN(n46079) );
  INHSV2 U49920 ( .I(n46083), .ZN(n46088) );
  NOR2HSV0 U49921 ( .A1(n46085), .A2(n46084), .ZN(n46086) );
  OR2HSV1 U49922 ( .A1(n46091), .A2(n46090), .Z(n46093) );
  NOR2HSV1 U49923 ( .A1(n46093), .A2(n46092), .ZN(n46094) );
  CLKNAND2HSV2 U49924 ( .A1(n46099), .A2(n46107), .ZN(n46100) );
  CLKNAND2HSV1 U49925 ( .A1(n46108), .A2(n46107), .ZN(n46109) );
  CLKAND2HSV2 U49926 ( .A1(n46559), .A2(\pe3/ti_7t [31]), .Z(n46112) );
  AOI21HSV4 U49927 ( .A1(n46113), .A2(n25888), .B(n46112), .ZN(n46117) );
  OR2HSV1 U49928 ( .A1(n46114), .A2(n36967), .Z(n46115) );
  INHSV4 U49929 ( .I(n46308), .ZN(n56854) );
  INHSV2 U49930 ( .I(n50799), .ZN(n59967) );
  BUFHSV2 U49931 ( .I(n51687), .Z(n59775) );
  BUFHSV2 U49932 ( .I(n49726), .Z(n59915) );
  BUFHSV2 U49933 ( .I(n46170), .Z(n59177) );
  MUX2HSV1 U49934 ( .I0(bo3[5]), .I1(n56937), .S(n46124), .Z(n59793) );
  MUX2HSV1 U49935 ( .I0(bo3[23]), .I1(n56213), .S(n46127), .Z(n59558) );
  MUX2HSV1 U49936 ( .I0(bo3[26]), .I1(\pe3/bq[26] ), .S(n46128), .Z(n59555) );
  MUX2HSV1 U49937 ( .I0(bo3[31]), .I1(n48538), .S(n46129), .Z(n59554) );
  MUX2HSV1 U49938 ( .I0(bo3[25]), .I1(n56071), .S(n46130), .Z(n59556) );
  MUX2HSV1 U49939 ( .I0(bo3[19]), .I1(\pe3/bq[19] ), .S(n46132), .Z(n59770) );
  MUX2HSV1 U49940 ( .I0(bo2[23]), .I1(n52300), .S(n48079), .Z(n59562) );
  MUX2HSV1 U49941 ( .I0(bo4[31]), .I1(n33423), .S(n48072), .Z(n59800) );
  MUX2HSV1 U49942 ( .I0(bo3[21]), .I1(n56218), .S(n46140), .Z(n59772) );
  MUX2HSV1 U49943 ( .I0(bo5[19]), .I1(n39454), .S(n30925), .Z(n59850) );
  MUX2HSV1 U49944 ( .I0(bo6[28]), .I1(n46135), .S(n46621), .Z(n59873) );
  MUX2HSV1 U49945 ( .I0(bo5[6]), .I1(n50526), .S(n48049), .Z(n59863) );
  MUX2HSV1 U49946 ( .I0(bo6[20]), .I1(n46137), .S(n48025), .Z(n59888) );
  MUX2HSV1 U49947 ( .I0(bo3[16]), .I1(n43544), .S(n46140), .Z(n59780) );
  MUX2HSV1 U49948 ( .I0(bo3[9]), .I1(n53232), .S(n46139), .Z(n59786) );
  MUX2HSV1 U49949 ( .I0(bo3[8]), .I1(n55970), .S(n46140), .Z(n59785) );
  MUX2HSV1 U49950 ( .I0(bo3[2]), .I1(n56892), .S(n46141), .Z(n59795) );
  INHSV2 U49951 ( .I(n54472), .ZN(n59495) );
  NAND2HSV2 U49952 ( .A1(n46151), .A2(n46152), .ZN(n46145) );
  BUFHSV2 U49953 ( .I(n49317), .Z(n46823) );
  BUFHSV2 U49954 ( .I(\pe6/got [2]), .Z(n58724) );
  BUFHSV2 U49955 ( .I(n58724), .Z(n58816) );
  BUFHSV2 U49956 ( .I(n49078), .Z(n58805) );
  CLKNAND2HSV1 U49957 ( .A1(n58805), .A2(n58403), .ZN(n46149) );
  INHSV2 U49958 ( .I(n46146), .ZN(n58452) );
  INHSV1 U49959 ( .I(n49327), .ZN(n58496) );
  INHSV2 U49960 ( .I(n46147), .ZN(n58405) );
  INHSV2 U49961 ( .I(n48041), .ZN(n58460) );
  CLKNHSV0 U49962 ( .I(n58483), .ZN(n58449) );
  BUFHSV2 U49963 ( .I(n58479), .Z(n58401) );
  INHSV2 U49964 ( .I(n46302), .ZN(n46150) );
  AND2HSV2 U49965 ( .A1(n46155), .A2(n46154), .Z(n46153) );
  CLKNAND2HSV0 U49966 ( .A1(n46153), .A2(n46156), .ZN(n46158) );
  CLKNAND2HSV2 U49967 ( .A1(n58369), .A2(n46154), .ZN(n46157) );
  NAND2HSV2 U49968 ( .A1(n46156), .A2(n46155), .ZN(n46552) );
  NAND2HSV2 U49969 ( .A1(n46584), .A2(\pe6/ti_7t [31]), .ZN(n46303) );
  INOR2HSV0 U49970 ( .A1(n46303), .B1(n46159), .ZN(n46160) );
  NAND2HSV2 U49971 ( .A1(n46299), .A2(n46160), .ZN(n46161) );
  CLKNAND2HSV1 U49972 ( .A1(n46552), .A2(n51438), .ZN(n46168) );
  NOR2HSV2 U49973 ( .A1(n46168), .A2(n46553), .ZN(n46164) );
  NOR2HSV2 U49974 ( .A1(n46164), .A2(n46546), .ZN(n46166) );
  NOR2HSV1 U49975 ( .A1(n46552), .A2(n25463), .ZN(n46169) );
  INHSV2 U49976 ( .I(n46303), .ZN(n46305) );
  AOI21HSV4 U49977 ( .A1(n46166), .A2(n46165), .B(n46305), .ZN(n58435) );
  NAND2HSV2 U49978 ( .A1(n46819), .A2(n46299), .ZN(n58439) );
  CLKNHSV0 U49979 ( .I(n46169), .ZN(n46296) );
  NAND2HSV2 U49980 ( .A1(n59166), .A2(n46822), .ZN(n46294) );
  INHSV2 U49981 ( .I(n46823), .ZN(n58402) );
  NAND2HSV2 U49982 ( .A1(n58402), .A2(n49665), .ZN(n46292) );
  NAND2HSV2 U49983 ( .A1(n58611), .A2(n32242), .ZN(n46288) );
  NAND2HSV0 U49984 ( .A1(n46769), .A2(n58808), .ZN(n46282) );
  BUFHSV2 U49985 ( .I(n46170), .Z(n58662) );
  NAND2HSV2 U49986 ( .A1(n58662), .A2(n59328), .ZN(n46278) );
  CLKNAND2HSV0 U49987 ( .A1(n58663), .A2(n59176), .ZN(n46276) );
  CLKNAND2HSV0 U49988 ( .A1(n58664), .A2(n58807), .ZN(n46274) );
  NAND2HSV2 U49989 ( .A1(n59032), .A2(n46171), .ZN(n46267) );
  NAND2HSV0 U49990 ( .A1(n46172), .A2(\pe6/got [15]), .ZN(n46265) );
  NAND2HSV0 U49991 ( .A1(n58813), .A2(n58713), .ZN(n46263) );
  NAND2HSV0 U49992 ( .A1(n49743), .A2(n58711), .ZN(n46261) );
  NAND2HSV0 U49993 ( .A1(n49829), .A2(n59180), .ZN(n46259) );
  INHSV2 U49994 ( .I(n53110), .ZN(n58572) );
  NAND2HSV0 U49995 ( .A1(n26109), .A2(n58572), .ZN(n46257) );
  NAND2HSV0 U49996 ( .A1(n36107), .A2(n58477), .ZN(n46253) );
  NAND2HSV0 U49997 ( .A1(n59183), .A2(n58526), .ZN(n46251) );
  BUFHSV2 U49998 ( .I(n58400), .Z(n58384) );
  NAND2HSV0 U49999 ( .A1(n36108), .A2(n58384), .ZN(n46175) );
  NAND2HSV0 U50000 ( .A1(n59038), .A2(n46173), .ZN(n46174) );
  XOR2HSV0 U50001 ( .A1(n46175), .A2(n46174), .Z(n46245) );
  NAND2HSV0 U50002 ( .A1(n59202), .A2(\pe6/aot [11]), .ZN(n46654) );
  NAND2HSV0 U50003 ( .A1(n59247), .A2(n58378), .ZN(n59109) );
  XOR2HSV0 U50004 ( .A1(n46654), .A2(n59109), .Z(n46189) );
  BUFHSV2 U50005 ( .I(\pe6/got [2]), .Z(n58331) );
  NAND2HSV0 U50006 ( .A1(n46176), .A2(n58331), .ZN(n46177) );
  XOR2HSV0 U50007 ( .A1(n46177), .A2(\pe6/phq [31]), .Z(n46181) );
  CLKNAND2HSV1 U50008 ( .A1(\pe6/bq[4] ), .A2(n58459), .ZN(n58395) );
  OAI22HSV0 U50009 ( .A1(n32484), .A2(n58530), .B1(n46642), .B2(n32193), .ZN(
        n46178) );
  OAI21HSV0 U50010 ( .A1(n46179), .A2(n58395), .B(n46178), .ZN(n46180) );
  XNOR2HSV1 U50011 ( .A1(n46181), .A2(n46180), .ZN(n46188) );
  NAND2HSV0 U50012 ( .A1(n44701), .A2(\pe6/pvq [31]), .ZN(n46182) );
  XOR2HSV0 U50013 ( .A1(n49026), .A2(n46182), .Z(n46186) );
  NAND2HSV0 U50014 ( .A1(n32999), .A2(n59266), .ZN(n46184) );
  NAND2HSV0 U50015 ( .A1(n59084), .A2(n58824), .ZN(n46183) );
  XOR2HSV0 U50016 ( .A1(n46184), .A2(n46183), .Z(n46185) );
  XOR2HSV0 U50017 ( .A1(n46186), .A2(n46185), .Z(n46187) );
  XOR3HSV2 U50018 ( .A1(n46189), .A2(n46188), .A3(n46187), .Z(n46243) );
  INAND2HSV2 U50019 ( .A1(n32723), .B1(n58339), .ZN(n46191) );
  NAND2HSV0 U50020 ( .A1(n58991), .A2(n58618), .ZN(n46190) );
  XOR2HSV0 U50021 ( .A1(n46191), .A2(n46190), .Z(n46196) );
  NAND2HSV0 U50022 ( .A1(n48051), .A2(n33004), .ZN(n46194) );
  NAND2HSV0 U50023 ( .A1(n59217), .A2(n58449), .ZN(n46193) );
  XOR2HSV0 U50024 ( .A1(n46194), .A2(n46193), .Z(n46195) );
  XOR2HSV0 U50025 ( .A1(n46196), .A2(n46195), .Z(n46205) );
  NAND2HSV0 U50026 ( .A1(n44435), .A2(n53115), .ZN(n46199) );
  NAND2HSV0 U50027 ( .A1(n59206), .A2(n46197), .ZN(n46198) );
  XOR2HSV0 U50028 ( .A1(n46199), .A2(n46198), .Z(n46203) );
  NAND2HSV0 U50029 ( .A1(n33005), .A2(n58943), .ZN(n46201) );
  NAND2HSV0 U50030 ( .A1(n36143), .A2(\pe6/aot [21]), .ZN(n46200) );
  XOR2HSV0 U50031 ( .A1(n46201), .A2(n46200), .Z(n46202) );
  XOR2HSV0 U50032 ( .A1(n46203), .A2(n46202), .Z(n46204) );
  XOR2HSV0 U50033 ( .A1(n46205), .A2(n46204), .Z(n46207) );
  NAND2HSV0 U50034 ( .A1(n31454), .A2(n48891), .ZN(n46206) );
  XNOR2HSV1 U50035 ( .A1(n46207), .A2(n46206), .ZN(n46242) );
  INHSV2 U50036 ( .I(n49681), .ZN(n58404) );
  NAND2HSV0 U50037 ( .A1(n46658), .A2(n58404), .ZN(n46209) );
  NAND2HSV0 U50038 ( .A1(n35751), .A2(\pe6/aot [19]), .ZN(n46208) );
  XOR2HSV0 U50039 ( .A1(n46209), .A2(n46208), .Z(n46214) );
  NAND2HSV0 U50040 ( .A1(n46210), .A2(\pe6/aot [23]), .ZN(n46212) );
  CLKNHSV0 U50041 ( .I(n35607), .ZN(n59264) );
  NAND2HSV0 U50042 ( .A1(n58668), .A2(n59264), .ZN(n46211) );
  XOR2HSV0 U50043 ( .A1(n46212), .A2(n46211), .Z(n46213) );
  XOR2HSV0 U50044 ( .A1(n46214), .A2(n46213), .Z(n46223) );
  NAND2HSV0 U50045 ( .A1(n58619), .A2(n59272), .ZN(n46216) );
  NAND2HSV0 U50046 ( .A1(n49844), .A2(n59088), .ZN(n46215) );
  XOR2HSV0 U50047 ( .A1(n46216), .A2(n46215), .Z(n46221) );
  NAND2HSV0 U50048 ( .A1(n49862), .A2(\pe6/aot [13]), .ZN(n46219) );
  NAND2HSV0 U50049 ( .A1(\pe6/bq[18] ), .A2(n46217), .ZN(n46218) );
  XOR2HSV0 U50050 ( .A1(n46219), .A2(n46218), .Z(n46220) );
  XOR2HSV0 U50051 ( .A1(n46221), .A2(n46220), .Z(n46222) );
  XOR2HSV0 U50052 ( .A1(n46223), .A2(n46222), .Z(n46240) );
  NAND2HSV0 U50053 ( .A1(n58965), .A2(n46792), .ZN(n46225) );
  NAND2HSV0 U50054 ( .A1(n58675), .A2(n32588), .ZN(n46224) );
  XOR2HSV0 U50055 ( .A1(n46225), .A2(n46224), .Z(n46229) );
  NAND2HSV0 U50056 ( .A1(\pe6/bq[10] ), .A2(n58749), .ZN(n46227) );
  NAND2HSV0 U50057 ( .A1(n59050), .A2(n58488), .ZN(n46226) );
  XOR2HSV0 U50058 ( .A1(n46227), .A2(n46226), .Z(n46228) );
  XOR2HSV0 U50059 ( .A1(n46229), .A2(n46228), .Z(n46238) );
  NAND2HSV0 U50060 ( .A1(n46627), .A2(\pe6/aot [2]), .ZN(n46232) );
  NAND2HSV0 U50061 ( .A1(n58360), .A2(n46230), .ZN(n46231) );
  XOR2HSV0 U50062 ( .A1(n46232), .A2(n46231), .Z(n46236) );
  NAND2HSV0 U50063 ( .A1(n58356), .A2(n31829), .ZN(n46234) );
  CLKNAND2HSV0 U50064 ( .A1(n32982), .A2(\pe6/aot [17]), .ZN(n46233) );
  XOR2HSV0 U50065 ( .A1(n46234), .A2(n46233), .Z(n46235) );
  XOR2HSV0 U50066 ( .A1(n46236), .A2(n46235), .Z(n46237) );
  XOR2HSV0 U50067 ( .A1(n46238), .A2(n46237), .Z(n46239) );
  XOR2HSV0 U50068 ( .A1(n46240), .A2(n46239), .Z(n46241) );
  XOR3HSV2 U50069 ( .A1(n46243), .A2(n46242), .A3(n46241), .Z(n46244) );
  XNOR2HSV1 U50070 ( .A1(n46245), .A2(n46244), .ZN(n46247) );
  NAND2HSV0 U50071 ( .A1(n59121), .A2(n58398), .ZN(n46246) );
  XNOR2HSV1 U50072 ( .A1(n46247), .A2(n46246), .ZN(n46249) );
  NAND2HSV0 U50073 ( .A1(n25218), .A2(n58814), .ZN(n46248) );
  XNOR2HSV1 U50074 ( .A1(n46249), .A2(n46248), .ZN(n46250) );
  XNOR2HSV1 U50075 ( .A1(n46251), .A2(n46250), .ZN(n46252) );
  XNOR2HSV1 U50076 ( .A1(n46253), .A2(n46252), .ZN(n46255) );
  CLKNAND2HSV1 U50077 ( .A1(n58886), .A2(n44393), .ZN(n46254) );
  XNOR2HSV1 U50078 ( .A1(n46255), .A2(n46254), .ZN(n46256) );
  XOR2HSV0 U50079 ( .A1(n46257), .A2(n46256), .Z(n46258) );
  XNOR2HSV1 U50080 ( .A1(n46259), .A2(n46258), .ZN(n46260) );
  XOR2HSV0 U50081 ( .A1(n46261), .A2(n46260), .Z(n46262) );
  XOR2HSV0 U50082 ( .A1(n46263), .A2(n46262), .Z(n46264) );
  XNOR2HSV1 U50083 ( .A1(n46265), .A2(n46264), .ZN(n46266) );
  XOR2HSV0 U50084 ( .A1(n46267), .A2(n46266), .Z(n46269) );
  NAND2HSV0 U50085 ( .A1(n59144), .A2(n59178), .ZN(n46268) );
  XOR2HSV0 U50086 ( .A1(n46269), .A2(n46268), .Z(n46272) );
  NAND2HSV0 U50087 ( .A1(n59676), .A2(n58715), .ZN(n46271) );
  XOR2HSV0 U50088 ( .A1(n46272), .A2(n46271), .Z(n46273) );
  XNOR2HSV1 U50089 ( .A1(n46274), .A2(n46273), .ZN(n46275) );
  XNOR2HSV1 U50090 ( .A1(n46276), .A2(n46275), .ZN(n46277) );
  XNOR2HSV1 U50091 ( .A1(n46278), .A2(n46277), .ZN(n46280) );
  CLKNAND2HSV0 U50092 ( .A1(n58601), .A2(n58714), .ZN(n46279) );
  XNOR2HSV1 U50093 ( .A1(n46280), .A2(n46279), .ZN(n46281) );
  XNOR2HSV1 U50094 ( .A1(n46282), .A2(n46281), .ZN(n46286) );
  INAND2HSV2 U50095 ( .A1(n32631), .B1(n59918), .ZN(n46285) );
  CLKNAND2HSV1 U50096 ( .A1(n49078), .A2(n46283), .ZN(n46284) );
  XOR3HSV2 U50097 ( .A1(n46286), .A2(n46285), .A3(n46284), .Z(n46287) );
  XNOR2HSV1 U50098 ( .A1(n46288), .A2(n46287), .ZN(n46291) );
  XOR3HSV2 U50099 ( .A1(n46292), .A2(n46291), .A3(n46290), .Z(n46293) );
  XNOR2HSV4 U50100 ( .A1(n46294), .A2(n46293), .ZN(n46551) );
  NOR2HSV2 U50101 ( .A1(n46551), .A2(n36050), .ZN(n46295) );
  OAI21HSV2 U50102 ( .A1(n46553), .A2(n46296), .B(n46295), .ZN(n46297) );
  NOR2HSV4 U50103 ( .A1(n46819), .A2(n46300), .ZN(n58441) );
  NOR2HSV4 U50104 ( .A1(n46306), .A2(n58441), .ZN(n48890) );
  NOR2HSV4 U50105 ( .A1(n46301), .A2(n48890), .ZN(n49173) );
  INHSV2 U50106 ( .I(n49173), .ZN(n46817) );
  NOR2HSV4 U50107 ( .A1(n49177), .A2(n46304), .ZN(n58442) );
  NOR2HSV2 U50108 ( .A1(n46551), .A2(n46305), .ZN(n58434) );
  NOR2HSV2 U50109 ( .A1(n58442), .A2(n58434), .ZN(n46307) );
  NOR2HSV4 U50110 ( .A1(n46306), .A2(n58441), .ZN(n49402) );
  INHSV4 U50111 ( .I(n46308), .ZN(n50752) );
  CLKNAND2HSV1 U50112 ( .A1(n56676), .A2(n52726), .ZN(n46440) );
  INHSV3 U50113 ( .I(n50716), .ZN(n56780) );
  CLKNAND2HSV0 U50114 ( .A1(n56780), .A2(n46309), .ZN(n46437) );
  CLKNAND2HSV0 U50115 ( .A1(n48481), .A2(n36958), .ZN(n46435) );
  CLKNAND2HSV0 U50116 ( .A1(n48482), .A2(n59384), .ZN(n46431) );
  INAND2HSV2 U50117 ( .A1(n48484), .B1(n59617), .ZN(n46429) );
  CLKNAND2HSV0 U50118 ( .A1(n49253), .A2(n42673), .ZN(n46427) );
  BUFHSV2 U50119 ( .I(n46312), .Z(n56737) );
  NAND2HSV0 U50120 ( .A1(n56737), .A2(n48485), .ZN(n46425) );
  NAND2HSV0 U50121 ( .A1(n56066), .A2(n55945), .ZN(n46423) );
  NAND2HSV0 U50122 ( .A1(n53228), .A2(\pe3/got [19]), .ZN(n46419) );
  NAND2HSV0 U50123 ( .A1(n56178), .A2(\pe3/got [18]), .ZN(n46414) );
  CLKNAND2HSV0 U50124 ( .A1(n43755), .A2(n56494), .ZN(n46405) );
  INHSV2 U50125 ( .I(n50799), .ZN(n56247) );
  NAND2HSV0 U50126 ( .A1(n56179), .A2(n56247), .ZN(n46403) );
  NAND2HSV0 U50127 ( .A1(n56180), .A2(n59644), .ZN(n46401) );
  NAND2HSV0 U50128 ( .A1(n46313), .A2(n56855), .ZN(n46397) );
  CLKNHSV0 U50129 ( .I(n56778), .ZN(n56241) );
  NAND2HSV0 U50130 ( .A1(n55707), .A2(n56241), .ZN(n46395) );
  NAND2HSV0 U50131 ( .A1(n48488), .A2(n48487), .ZN(n46393) );
  NAND2HSV0 U50132 ( .A1(\pe3/aot [8]), .A2(n55976), .ZN(n46316) );
  NAND2HSV0 U50133 ( .A1(n56197), .A2(n43146), .ZN(n46315) );
  XOR2HSV0 U50134 ( .A1(n46316), .A2(n46315), .Z(n46320) );
  INHSV2 U50135 ( .I(n56567), .ZN(n56373) );
  NAND2HSV0 U50136 ( .A1(n56373), .A2(n55872), .ZN(n46318) );
  NAND2HSV0 U50137 ( .A1(n56864), .A2(\pe3/bq[26] ), .ZN(n46317) );
  XOR2HSV0 U50138 ( .A1(n46318), .A2(n46317), .Z(n46319) );
  XOR2HSV0 U50139 ( .A1(n46320), .A2(n46319), .Z(n46329) );
  NAND2HSV0 U50140 ( .A1(n56740), .A2(n56213), .ZN(n46322) );
  NAND2HSV0 U50141 ( .A1(n55864), .A2(n55727), .ZN(n46321) );
  XOR2HSV0 U50142 ( .A1(n46322), .A2(n46321), .Z(n46327) );
  NAND2HSV0 U50143 ( .A1(n56349), .A2(n46323), .ZN(n46325) );
  NAND2HSV0 U50144 ( .A1(n55873), .A2(n37280), .ZN(n46324) );
  XOR2HSV0 U50145 ( .A1(n46325), .A2(n46324), .Z(n46326) );
  XOR2HSV0 U50146 ( .A1(n46327), .A2(n46326), .Z(n46328) );
  XOR2HSV0 U50147 ( .A1(n46329), .A2(n46328), .Z(n46331) );
  NAND2HSV0 U50148 ( .A1(n59648), .A2(n55950), .ZN(n46330) );
  XNOR2HSV1 U50149 ( .A1(n46331), .A2(n46330), .ZN(n46389) );
  NAND2HSV0 U50150 ( .A1(\pe3/aot [14]), .A2(\pe3/bq[19] ), .ZN(n46334) );
  NAND2HSV0 U50151 ( .A1(n46332), .A2(n56785), .ZN(n46333) );
  XOR2HSV0 U50152 ( .A1(n46334), .A2(n46333), .Z(n46338) );
  NAND2HSV0 U50153 ( .A1(n42818), .A2(n56187), .ZN(n46336) );
  NAND2HSV0 U50154 ( .A1(n56508), .A2(n55616), .ZN(n46335) );
  XOR2HSV0 U50155 ( .A1(n46336), .A2(n46335), .Z(n46337) );
  XOR2HSV0 U50156 ( .A1(n46338), .A2(n46337), .Z(n46346) );
  NAND2HSV0 U50157 ( .A1(\pe3/aot [22]), .A2(\pe3/bq[11] ), .ZN(n46340) );
  NAND2HSV0 U50158 ( .A1(n48500), .A2(\pe3/bq[4] ), .ZN(n46339) );
  XOR2HSV0 U50159 ( .A1(n46340), .A2(n46339), .Z(n46344) );
  NOR2HSV0 U50160 ( .A1(n55714), .A2(n49272), .ZN(n46342) );
  NAND2HSV0 U50161 ( .A1(n42743), .A2(n45639), .ZN(n46341) );
  XOR2HSV0 U50162 ( .A1(n46342), .A2(n46341), .Z(n46343) );
  XOR2HSV0 U50163 ( .A1(n46344), .A2(n46343), .Z(n46345) );
  XOR2HSV0 U50164 ( .A1(n46346), .A2(n46345), .Z(n46362) );
  NAND2HSV0 U50165 ( .A1(n56106), .A2(n56970), .ZN(n47434) );
  NAND2HSV0 U50166 ( .A1(\pe3/pq ), .A2(n48020), .ZN(n46349) );
  CLKNHSV0 U50167 ( .I(\pe3/bq[12] ), .ZN(n48545) );
  NAND2HSV0 U50168 ( .A1(n56182), .A2(n56688), .ZN(n46348) );
  XOR2HSV0 U50169 ( .A1(n46349), .A2(n46348), .Z(n46359) );
  NAND2HSV0 U50170 ( .A1(n59961), .A2(n48527), .ZN(n46473) );
  NOR2HSV0 U50171 ( .A1(n46350), .A2(n46473), .ZN(n46352) );
  AOI22HSV0 U50172 ( .A1(n56074), .A2(n48527), .B1(n48538), .B2(n56972), .ZN(
        n46351) );
  NOR2HSV2 U50173 ( .A1(n46352), .A2(n46351), .ZN(n46357) );
  NAND2HSV0 U50174 ( .A1(n55827), .A2(\pe3/bq[3] ), .ZN(n55725) );
  NOR2HSV0 U50175 ( .A1(n46353), .A2(n55725), .ZN(n46355) );
  AOI22HSV0 U50176 ( .A1(n48496), .A2(\pe3/bq[3] ), .B1(n56272), .B2(n36755), 
        .ZN(n46354) );
  NOR2HSV1 U50177 ( .A1(n46355), .A2(n46354), .ZN(n46356) );
  XOR2HSV0 U50178 ( .A1(n46357), .A2(n46356), .Z(n46358) );
  XOR3HSV2 U50179 ( .A1(n46360), .A2(n46359), .A3(n46358), .Z(n46361) );
  XNOR2HSV1 U50180 ( .A1(n46362), .A2(n46361), .ZN(n46385) );
  NAND2HSV0 U50181 ( .A1(n46363), .A2(n56824), .ZN(n56514) );
  OAI21HSV0 U50182 ( .A1(n59606), .A2(n49275), .B(n46364), .ZN(n46365) );
  OAI21HSV0 U50183 ( .A1(n46366), .A2(n56514), .B(n46365), .ZN(n46371) );
  NAND2HSV0 U50184 ( .A1(n53249), .A2(\pe3/bq[14] ), .ZN(n49419) );
  NOR2HSV0 U50185 ( .A1(n46367), .A2(n49419), .ZN(n46369) );
  AOI22HSV0 U50186 ( .A1(n56464), .A2(n56379), .B1(n42971), .B2(n53249), .ZN(
        n46368) );
  NOR2HSV2 U50187 ( .A1(n46369), .A2(n46368), .ZN(n46370) );
  XNOR2HSV1 U50188 ( .A1(n46371), .A2(n46370), .ZN(n46375) );
  NAND2HSV0 U50189 ( .A1(\pe3/aot [6]), .A2(n55960), .ZN(n46372) );
  XOR2HSV0 U50190 ( .A1(n46373), .A2(n46372), .Z(n46374) );
  XNOR2HSV1 U50191 ( .A1(n46375), .A2(n46374), .ZN(n46383) );
  CLKNHSV2 U50192 ( .I(\pe3/got [1]), .ZN(n47431) );
  NAND2HSV0 U50193 ( .A1(n56975), .A2(n45955), .ZN(n46377) );
  CLKNHSV0 U50194 ( .I(n48495), .ZN(n55828) );
  NAND2HSV0 U50195 ( .A1(n43547), .A2(n55828), .ZN(n46376) );
  XOR2HSV0 U50196 ( .A1(n46377), .A2(n46376), .Z(n46381) );
  NAND2HSV0 U50197 ( .A1(n56204), .A2(n55975), .ZN(n46379) );
  NAND2HSV0 U50198 ( .A1(\pe3/aot [3]), .A2(n48522), .ZN(n46378) );
  XOR2HSV0 U50199 ( .A1(n46379), .A2(n46378), .Z(n46380) );
  XOR2HSV0 U50200 ( .A1(n46381), .A2(n46380), .Z(n46382) );
  XOR2HSV0 U50201 ( .A1(n46383), .A2(n46382), .Z(n46384) );
  XNOR2HSV1 U50202 ( .A1(n46385), .A2(n46384), .ZN(n46388) );
  NAND2HSV0 U50203 ( .A1(n59797), .A2(n59356), .ZN(n46387) );
  NAND2HSV0 U50204 ( .A1(n48511), .A2(n56781), .ZN(n46386) );
  XOR4HSV1 U50205 ( .A1(n46389), .A2(n46388), .A3(n46387), .A4(n46386), .Z(
        n46391) );
  NAND2HSV0 U50206 ( .A1(n52727), .A2(n59799), .ZN(n46390) );
  XNOR2HSV1 U50207 ( .A1(n46391), .A2(n46390), .ZN(n46392) );
  XNOR2HSV1 U50208 ( .A1(n46393), .A2(n46392), .ZN(n46394) );
  XNOR2HSV1 U50209 ( .A1(n46395), .A2(n46394), .ZN(n46396) );
  XNOR2HSV1 U50210 ( .A1(n46397), .A2(n46396), .ZN(n46399) );
  NAND2HSV0 U50211 ( .A1(n55895), .A2(n56177), .ZN(n46398) );
  XNOR2HSV1 U50212 ( .A1(n46399), .A2(n46398), .ZN(n46400) );
  XNOR2HSV1 U50213 ( .A1(n46401), .A2(n46400), .ZN(n46402) );
  XNOR2HSV1 U50214 ( .A1(n46403), .A2(n46402), .ZN(n46404) );
  XNOR2HSV1 U50215 ( .A1(n46405), .A2(n46404), .ZN(n46409) );
  NOR2HSV0 U50216 ( .A1(n56391), .A2(n46406), .ZN(n46408) );
  NAND2HSV0 U50217 ( .A1(n49468), .A2(n56493), .ZN(n46407) );
  XOR3HSV1 U50218 ( .A1(n46409), .A2(n46408), .A3(n46407), .Z(n46412) );
  NOR2HSV1 U50219 ( .A1(n48583), .A2(n45727), .ZN(n46411) );
  BUFHSV2 U50220 ( .I(n59810), .Z(n56396) );
  NAND2HSV0 U50221 ( .A1(n56396), .A2(n56065), .ZN(n46410) );
  XOR3HSV2 U50222 ( .A1(n46412), .A2(n46411), .A3(n46410), .Z(n46413) );
  XNOR2HSV1 U50223 ( .A1(n46414), .A2(n46413), .ZN(n46417) );
  BUFHSV2 U50224 ( .I(n46415), .Z(n59811) );
  NAND2HSV0 U50225 ( .A1(n55912), .A2(n56335), .ZN(n46416) );
  XNOR2HSV1 U50226 ( .A1(n46417), .A2(n46416), .ZN(n46418) );
  XNOR2HSV1 U50227 ( .A1(n46419), .A2(n46418), .ZN(n46421) );
  NOR2HSV0 U50228 ( .A1(n55917), .A2(n45635), .ZN(n46420) );
  XNOR2HSV1 U50229 ( .A1(n46421), .A2(n46420), .ZN(n46422) );
  XNOR2HSV1 U50230 ( .A1(n46423), .A2(n46422), .ZN(n46424) );
  XOR2HSV0 U50231 ( .A1(n46425), .A2(n46424), .Z(n46426) );
  XNOR2HSV1 U50232 ( .A1(n46427), .A2(n46426), .ZN(n46428) );
  XNOR2HSV1 U50233 ( .A1(n46429), .A2(n46428), .ZN(n46430) );
  XNOR2HSV1 U50234 ( .A1(n46431), .A2(n46430), .ZN(n46432) );
  XNOR2HSV1 U50235 ( .A1(n46433), .A2(n46432), .ZN(n46434) );
  XNOR2HSV1 U50236 ( .A1(n46435), .A2(n46434), .ZN(n46436) );
  XNOR2HSV1 U50237 ( .A1(n46440), .A2(n46439), .ZN(po3) );
  INAND2HSV2 U50238 ( .A1(n48484), .B1(n48485), .ZN(n46543) );
  CLKNAND2HSV0 U50239 ( .A1(n49253), .A2(n43262), .ZN(n46541) );
  NAND2HSV0 U50240 ( .A1(n55613), .A2(n42996), .ZN(n46539) );
  NAND2HSV0 U50241 ( .A1(n56562), .A2(\pe3/got [19]), .ZN(n46537) );
  NAND2HSV0 U50242 ( .A1(n43754), .A2(n56064), .ZN(n46531) );
  NAND2HSV0 U50243 ( .A1(n55824), .A2(n56065), .ZN(n46527) );
  CLKNAND2HSV0 U50244 ( .A1(n56067), .A2(n56558), .ZN(n46518) );
  NAND2HSV0 U50245 ( .A1(n49255), .A2(n56177), .ZN(n46516) );
  BUFHSV2 U50246 ( .I(n47991), .Z(n55949) );
  NAND2HSV0 U50247 ( .A1(n55949), .A2(n56855), .ZN(n46514) );
  NAND2HSV0 U50248 ( .A1(n56070), .A2(n48487), .ZN(n46510) );
  NAND2HSV0 U50249 ( .A1(n56267), .A2(n55825), .ZN(n46508) );
  INHSV1 U50250 ( .I(n56904), .ZN(n56068) );
  NAND2HSV0 U50251 ( .A1(n48488), .A2(n56068), .ZN(n46506) );
  NAND2HSV0 U50252 ( .A1(n59797), .A2(n56975), .ZN(n46502) );
  NAND2HSV0 U50253 ( .A1(n48511), .A2(n59807), .ZN(n46501) );
  NAND2HSV0 U50254 ( .A1(n42950), .A2(n55975), .ZN(n46443) );
  NAND2HSV0 U50255 ( .A1(n56113), .A2(\pe3/bq[14] ), .ZN(n46442) );
  XOR2HSV0 U50256 ( .A1(n46443), .A2(n46442), .Z(n46447) );
  CLKNHSV0 U50257 ( .I(n46138), .ZN(n56640) );
  NAND2HSV0 U50258 ( .A1(n55864), .A2(n56640), .ZN(n46445) );
  NAND2HSV0 U50259 ( .A1(n56439), .A2(\pe3/bq[26] ), .ZN(n46444) );
  XOR2HSV0 U50260 ( .A1(n46445), .A2(n46444), .Z(n46446) );
  XOR2HSV0 U50261 ( .A1(n46447), .A2(n46446), .Z(n46455) );
  NAND2HSV0 U50262 ( .A1(\pe3/aot [6]), .A2(n48520), .ZN(n46449) );
  NAND2HSV0 U50263 ( .A1(\pe3/aot [23]), .A2(n55970), .ZN(n46448) );
  XOR2HSV0 U50264 ( .A1(n46449), .A2(n46448), .Z(n46453) );
  NAND2HSV0 U50265 ( .A1(n56087), .A2(\pe3/bq[7] ), .ZN(n46451) );
  NAND2HSV0 U50266 ( .A1(n53249), .A2(n55727), .ZN(n46450) );
  XOR2HSV0 U50267 ( .A1(n46451), .A2(n46450), .Z(n46452) );
  XOR2HSV0 U50268 ( .A1(n46453), .A2(n46452), .Z(n46454) );
  XOR2HSV0 U50269 ( .A1(n46455), .A2(n46454), .Z(n46472) );
  CLKNHSV0 U50270 ( .I(n46615), .ZN(n56094) );
  NAND2HSV0 U50271 ( .A1(n43030), .A2(n56094), .ZN(n46458) );
  NAND2HSV0 U50272 ( .A1(n46456), .A2(\pe3/bq[4] ), .ZN(n46457) );
  XOR2HSV0 U50273 ( .A1(n46458), .A2(n46457), .Z(n46462) );
  NAND2HSV0 U50274 ( .A1(n56188), .A2(n55616), .ZN(n46460) );
  NAND2HSV0 U50275 ( .A1(n56370), .A2(\pe3/bq[19] ), .ZN(n46459) );
  XOR2HSV0 U50276 ( .A1(n46460), .A2(n46459), .Z(n46461) );
  XOR2HSV0 U50277 ( .A1(n46462), .A2(n46461), .Z(n46470) );
  NAND2HSV0 U50278 ( .A1(n59511), .A2(n48522), .ZN(n46465) );
  NAND2HSV0 U50279 ( .A1(n46463), .A2(n55828), .ZN(n46464) );
  XOR2HSV0 U50280 ( .A1(n46465), .A2(n46464), .Z(n46468) );
  NAND2HSV0 U50281 ( .A1(n42743), .A2(n56428), .ZN(n49414) );
  NAND2HSV0 U50282 ( .A1(n56197), .A2(\pe3/bq[20] ), .ZN(n46466) );
  XOR2HSV0 U50283 ( .A1(n49414), .A2(n46466), .Z(n46467) );
  XOR2HSV0 U50284 ( .A1(n46468), .A2(n46467), .Z(n46469) );
  XOR2HSV0 U50285 ( .A1(n46470), .A2(n46469), .Z(n46471) );
  XOR2HSV0 U50286 ( .A1(n46472), .A2(n46471), .Z(n46499) );
  NAND2HSV0 U50287 ( .A1(\pe3/aot [19]), .A2(n56507), .ZN(n47448) );
  XOR2HSV0 U50288 ( .A1(n46473), .A2(n47448), .Z(n46497) );
  NAND2HSV0 U50289 ( .A1(\pe3/aot [3]), .A2(n42634), .ZN(n46475) );
  NAND2HSV0 U50290 ( .A1(n56788), .A2(n55960), .ZN(n46474) );
  XOR2HSV0 U50291 ( .A1(n46475), .A2(n46474), .Z(n46479) );
  NAND2HSV0 U50292 ( .A1(\pe3/aot [8]), .A2(n56213), .ZN(n46477) );
  NAND2HSV0 U50293 ( .A1(n56373), .A2(n45807), .ZN(n46476) );
  XOR2HSV0 U50294 ( .A1(n46477), .A2(n46476), .Z(n46478) );
  XNOR2HSV1 U50295 ( .A1(n46479), .A2(n46478), .ZN(n46496) );
  NOR2HSV0 U50296 ( .A1(n42643), .A2(n49275), .ZN(n46482) );
  NOR2HSV0 U50297 ( .A1(n45567), .A2(n56277), .ZN(n46481) );
  NAND2HSV0 U50298 ( .A1(\pe3/aot [22]), .A2(n56824), .ZN(n49413) );
  OAI22HSV0 U50299 ( .A1(n46482), .A2(n46481), .B1(n46480), .B2(n49413), .ZN(
        n46487) );
  NAND2HSV0 U50300 ( .A1(n55858), .A2(\pe3/bq[3] ), .ZN(n56000) );
  NOR2HSV0 U50301 ( .A1(n46483), .A2(n56000), .ZN(n46485) );
  AOI22HSV0 U50302 ( .A1(n59809), .A2(n56529), .B1(n48530), .B2(n56272), .ZN(
        n46484) );
  NOR2HSV2 U50303 ( .A1(n46485), .A2(n46484), .ZN(n46486) );
  XNOR2HSV1 U50304 ( .A1(n46487), .A2(n46486), .ZN(n46495) );
  NAND2HSV0 U50305 ( .A1(n42940), .A2(n56627), .ZN(n46489) );
  NAND2HSV0 U50306 ( .A1(n56204), .A2(\pe3/bq[11] ), .ZN(n46488) );
  XOR2HSV0 U50307 ( .A1(n46489), .A2(n46488), .Z(n46493) );
  NAND2HSV0 U50308 ( .A1(n59627), .A2(n55872), .ZN(n46491) );
  NAND2HSV0 U50309 ( .A1(n56740), .A2(n56106), .ZN(n46490) );
  XOR2HSV0 U50310 ( .A1(n46491), .A2(n46490), .Z(n46492) );
  XOR2HSV0 U50311 ( .A1(n46493), .A2(n46492), .Z(n46494) );
  XOR4HSV1 U50312 ( .A1(n46497), .A2(n46496), .A3(n46495), .A4(n46494), .Z(
        n46498) );
  XNOR2HSV1 U50313 ( .A1(n46499), .A2(n46498), .ZN(n46500) );
  XOR3HSV2 U50314 ( .A1(n46502), .A2(n46501), .A3(n46500), .Z(n46504) );
  NAND2HSV0 U50315 ( .A1(n55826), .A2(n56069), .ZN(n46503) );
  XNOR2HSV1 U50316 ( .A1(n46504), .A2(n46503), .ZN(n46505) );
  XNOR2HSV1 U50317 ( .A1(n46506), .A2(n46505), .ZN(n46507) );
  XNOR2HSV1 U50318 ( .A1(n46508), .A2(n46507), .ZN(n46509) );
  XNOR2HSV1 U50319 ( .A1(n46510), .A2(n46509), .ZN(n46512) );
  NAND2HSV0 U50320 ( .A1(n55895), .A2(n56241), .ZN(n46511) );
  XNOR2HSV1 U50321 ( .A1(n46512), .A2(n46511), .ZN(n46513) );
  XNOR2HSV1 U50322 ( .A1(n46514), .A2(n46513), .ZN(n46515) );
  XNOR2HSV1 U50323 ( .A1(n46516), .A2(n46515), .ZN(n46517) );
  XNOR2HSV1 U50324 ( .A1(n46518), .A2(n46517), .ZN(n46522) );
  NOR2HSV0 U50325 ( .A1(n43840), .A2(n50799), .ZN(n46521) );
  CLKNHSV0 U50326 ( .I(n46519), .ZN(n56422) );
  NAND2HSV0 U50327 ( .A1(n56422), .A2(n56176), .ZN(n46520) );
  XOR3HSV1 U50328 ( .A1(n46522), .A2(n46521), .A3(n46520), .Z(n46525) );
  NOR2HSV1 U50329 ( .A1(n48583), .A2(n46406), .ZN(n46524) );
  NAND2HSV0 U50330 ( .A1(n56396), .A2(n56493), .ZN(n46523) );
  XOR3HSV2 U50331 ( .A1(n46525), .A2(n46524), .A3(n46523), .Z(n46526) );
  XNOR2HSV1 U50332 ( .A1(n46527), .A2(n46526), .ZN(n46529) );
  CLKNAND2HSV0 U50333 ( .A1(n55912), .A2(n48584), .ZN(n46528) );
  XNOR2HSV1 U50334 ( .A1(n46529), .A2(n46528), .ZN(n46530) );
  XNOR2HSV1 U50335 ( .A1(n46531), .A2(n46530), .ZN(n46535) );
  BUFHSV2 U50336 ( .I(n46532), .Z(n56406) );
  NOR2HSV0 U50337 ( .A1(n56406), .A2(n46533), .ZN(n46534) );
  XNOR2HSV1 U50338 ( .A1(n46535), .A2(n46534), .ZN(n46536) );
  XNOR2HSV1 U50339 ( .A1(n46537), .A2(n46536), .ZN(n46538) );
  XOR2HSV0 U50340 ( .A1(n46539), .A2(n46538), .Z(n46540) );
  XNOR2HSV1 U50341 ( .A1(n46541), .A2(n46540), .ZN(n46542) );
  XNOR2HSV1 U50342 ( .A1(n46543), .A2(n46542), .ZN(n46544) );
  NAND2HSV2 U50343 ( .A1(n49177), .A2(n46546), .ZN(n46547) );
  INHSV2 U50344 ( .I(n46547), .ZN(n46548) );
  BUFHSV2 U50345 ( .I(\pe2/bq[2] ), .Z(n51493) );
  NOR2HSV0 U50346 ( .A1(n49737), .A2(n46549), .ZN(n46550) );
  XNOR2HSV1 U50347 ( .A1(n46551), .A2(n46550), .ZN(n46555) );
  XOR2HSV0 U50348 ( .A1(n46553), .A2(n46552), .Z(n46554) );
  XOR2HSV0 U50349 ( .A1(n46555), .A2(n46554), .Z(n46556) );
  NOR2HSV2 U50350 ( .A1(n46556), .A2(n52701), .ZN(n46557) );
  XOR2HSV0 U50351 ( .A1(n46557), .A2(poh6[31]), .Z(po[32]) );
  CLKBUFHSV0 U50352 ( .I(n25888), .Z(n46562) );
  INHSV4 U50353 ( .I(n50111), .ZN(n50318) );
  CLKNAND2HSV1 U50354 ( .A1(n59026), .A2(n46567), .ZN(n46571) );
  XOR2HSV0 U50355 ( .A1(n46569), .A2(n46568), .Z(n46570) );
  XNOR2HSV1 U50356 ( .A1(n46571), .A2(n46570), .ZN(n46572) );
  NOR2HSV2 U50357 ( .A1(n46572), .A2(n33089), .ZN(n46573) );
  CLKNAND2HSV0 U50358 ( .A1(n58402), .A2(n46574), .ZN(n46576) );
  CLKXOR2HSV1 U50359 ( .A1(n46576), .A2(n26462), .Z(n46577) );
  XNOR2HSV1 U50360 ( .A1(n46578), .A2(n46577), .ZN(n46579) );
  CLKNAND2HSV1 U50361 ( .A1(n46579), .A2(n48001), .ZN(n46580) );
  XNOR2HSV1 U50362 ( .A1(n46580), .A2(poh6[27]), .ZN(po[28]) );
  INHSV2 U50363 ( .I(n55144), .ZN(n59751) );
  BUFHSV3 U50364 ( .I(n49921), .Z(n58193) );
  BUFHSV2 U50365 ( .I(n50301), .Z(n50094) );
  NAND2HSV0 U50366 ( .A1(n46585), .A2(n46584), .ZN(n46586) );
  XNOR2HSV1 U50367 ( .A1(n46586), .A2(poh6[24]), .ZN(po[25]) );
  BUFHSV2 U50368 ( .I(n46825), .Z(n59680) );
  CLKNHSV0 U50369 ( .I(n43131), .ZN(n59500) );
  BUFHSV2 U50370 ( .I(n46592), .Z(n59916) );
  CLKNHSV0 U50371 ( .I(n46595), .ZN(n46598) );
  NAND3HSV0 U50372 ( .A1(n46598), .A2(n46597), .A3(n46596), .ZN(n46600) );
  XNOR2HSV0 U50373 ( .A1(n46600), .A2(n46599), .ZN(pov4[15]) );
  BUFHSV2 U50374 ( .I(n46601), .Z(n59835) );
  NAND2HSV0 U50375 ( .A1(n46603), .A2(n46602), .ZN(n46605) );
  INAND2HSV0 U50376 ( .A1(n46605), .B1(n46604), .ZN(n46606) );
  XNOR2HSV0 U50377 ( .A1(n46606), .A2(n52757), .ZN(n60027) );
  NAND2HSV0 U50378 ( .A1(n59681), .A2(n47772), .ZN(n46608) );
  XNOR2HSV0 U50379 ( .A1(n46608), .A2(n46607), .ZN(n60079) );
  CLKNHSV0 U50380 ( .I(rst), .ZN(n48477) );
  CLKNHSV0 U50381 ( .I(n48477), .ZN(n59434) );
  BUFHSV2 U50382 ( .I(n46611), .Z(n59524) );
  MUX2HSV2 U50383 ( .I0(bo3[6]), .I1(n56272), .S(n46612), .Z(n59791) );
  MUX2HSV2 U50384 ( .I0(bo3[32]), .I1(n46614), .S(n48020), .Z(n59688) );
  MUX2HSV2 U50385 ( .I0(bo3[15]), .I1(n56641), .S(n53221), .Z(n59779) );
  MUX2HSV1 U50386 ( .I0(bo3[17]), .I1(n56519), .S(n46616), .Z(n59776) );
  MUX2HSV1 U50387 ( .I0(bo4[30]), .I1(n46617), .S(n48058), .Z(n59804) );
  MUX2HSV2 U50388 ( .I0(bo2[26]), .I1(\pe2/bq[26] ), .S(n46619), .Z(n59728) );
  MUX2HSV2 U50389 ( .I0(bo6[29]), .I1(n35768), .S(n46621), .Z(n59872) );
  MUX2HSV1 U50390 ( .I0(bo5[22]), .I1(n47291), .S(n46628), .Z(n59849) );
  MUX2HSV1 U50391 ( .I0(bo1[26]), .I1(n41644), .S(n48081), .Z(n59695) );
  BUFHSV2 U50392 ( .I(n48039), .Z(n48027) );
  MUX2HSV1 U50393 ( .I0(bo5[25]), .I1(n46622), .S(n48027), .Z(n59843) );
  INHSV2 U50394 ( .I(n55504), .ZN(n59730) );
  BUFHSV2 U50395 ( .I(n48062), .Z(n48033) );
  MUX2HSV1 U50396 ( .I0(bo2[32]), .I1(n38303), .S(n48033), .Z(n59721) );
  INHSV2 U50397 ( .I(\pe4/aot [3]), .ZN(n57776) );
  MUX2HSV1 U50398 ( .I0(bo6[25]), .I1(n46624), .S(n48048), .Z(n59877) );
  BUFHSV2 U50399 ( .I(n48043), .Z(n46626) );
  MUX2HSV1 U50400 ( .I0(bo6[31]), .I1(n46625), .S(n46626), .Z(n59868) );
  MUX2HSV2 U50401 ( .I0(bo6[32]), .I1(n46627), .S(n46626), .Z(n59867) );
  CLKNHSV0 U50402 ( .I(n29892), .ZN(n48804) );
  MUX2HSV1 U50403 ( .I0(bo5[30]), .I1(n48804), .S(n46628), .Z(n59568) );
  NOR2HSV4 U50404 ( .A1(n46630), .A2(n49178), .ZN(n59338) );
  NAND2HSV2 U50405 ( .A1(n59167), .A2(n59168), .ZN(n46764) );
  CLKNAND2HSV0 U50406 ( .A1(n58809), .A2(n32815), .ZN(n46756) );
  BUFHSV2 U50407 ( .I(n46824), .Z(n59028) );
  CLKNAND2HSV0 U50408 ( .A1(n59028), .A2(n32970), .ZN(n46749) );
  NAND2HSV0 U50409 ( .A1(n58448), .A2(n59175), .ZN(n46745) );
  NAND2HSV0 U50410 ( .A1(n59680), .A2(n59328), .ZN(n46743) );
  NAND2HSV0 U50411 ( .A1(n59177), .A2(n49096), .ZN(n46739) );
  NAND2HSV0 U50412 ( .A1(n53112), .A2(n53101), .ZN(n46737) );
  NAND2HSV0 U50413 ( .A1(n58938), .A2(n49174), .ZN(n46735) );
  BUFHSV2 U50414 ( .I(n46631), .Z(n59179) );
  INHSV2 U50415 ( .I(n49666), .ZN(n58937) );
  NAND2HSV0 U50416 ( .A1(n59179), .A2(n58937), .ZN(n46733) );
  NAND2HSV0 U50417 ( .A1(n46632), .A2(n58810), .ZN(n46729) );
  NAND2HSV0 U50418 ( .A1(n59379), .A2(\pe6/got [13]), .ZN(n46727) );
  INHSV2 U50419 ( .I(n53110), .ZN(n59181) );
  NAND2HSV0 U50420 ( .A1(n59036), .A2(n59181), .ZN(n46723) );
  NAND2HSV0 U50421 ( .A1(n49829), .A2(\pe6/got [10]), .ZN(n46721) );
  NAND2HSV0 U50422 ( .A1(n49319), .A2(n46633), .ZN(n46719) );
  NAND2HSV0 U50423 ( .A1(n59678), .A2(n58814), .ZN(n46715) );
  BUFHSV2 U50424 ( .I(\pe6/got [6]), .Z(n58723) );
  NAND2HSV0 U50425 ( .A1(n59597), .A2(n58723), .ZN(n46713) );
  NAND2HSV0 U50426 ( .A1(n36108), .A2(\pe6/got [3]), .ZN(n46635) );
  BUFHSV2 U50427 ( .I(\pe6/got [2]), .Z(n59039) );
  NAND2HSV0 U50428 ( .A1(n59038), .A2(n59039), .ZN(n46634) );
  XNOR2HSV1 U50429 ( .A1(n46635), .A2(n46634), .ZN(n46707) );
  NAND2HSV0 U50430 ( .A1(n31454), .A2(n59235), .ZN(n46705) );
  NAND2HSV0 U50431 ( .A1(n59265), .A2(n58378), .ZN(n49191) );
  NOR2HSV0 U50432 ( .A1(n46636), .A2(n49191), .ZN(n46639) );
  CLKNHSV0 U50433 ( .I(n46853), .ZN(n59089) );
  AOI22HSV0 U50434 ( .A1(n45812), .A2(n58378), .B1(\pe6/aot [19]), .B2(n59089), 
        .ZN(n46638) );
  NOR2HSV1 U50435 ( .A1(n46639), .A2(n46638), .ZN(n46653) );
  NAND2HSV0 U50436 ( .A1(\pe6/bq[8] ), .A2(n59074), .ZN(n46641) );
  NAND2HSV0 U50437 ( .A1(n50829), .A2(\pe6/aot [13]), .ZN(n46640) );
  XOR2HSV0 U50438 ( .A1(n46641), .A2(n46640), .Z(n46652) );
  NAND2HSV2 U50439 ( .A1(n49106), .A2(n58404), .ZN(n58382) );
  NAND2HSV0 U50440 ( .A1(n59062), .A2(n46643), .ZN(n58988) );
  OAI21HSV0 U50441 ( .A1(n49681), .A2(n46620), .B(n58988), .ZN(n46644) );
  OAI21HSV0 U50442 ( .A1(n58382), .A2(n46645), .B(n46644), .ZN(n46650) );
  NAND2HSV0 U50443 ( .A1(n58833), .A2(n46217), .ZN(n58986) );
  NAND2HSV0 U50444 ( .A1(n59251), .A2(n58459), .ZN(n46648) );
  CLKNAND2HSV0 U50445 ( .A1(n49844), .A2(\pe6/aot [4]), .ZN(n49112) );
  NOR2HSV0 U50446 ( .A1(n46646), .A2(n49112), .ZN(n46647) );
  AOI21HSV0 U50447 ( .A1(n58986), .A2(n46648), .B(n46647), .ZN(n46649) );
  XNOR2HSV1 U50448 ( .A1(n46650), .A2(n46649), .ZN(n46651) );
  XOR3HSV2 U50449 ( .A1(n46653), .A2(n46652), .A3(n46651), .Z(n46669) );
  CLKNHSV0 U50450 ( .I(n46654), .ZN(n46656) );
  NOR2HSV0 U50451 ( .A1(n59205), .A2(n59193), .ZN(n49685) );
  AOI22HSV0 U50452 ( .A1(n59054), .A2(n58999), .B1(n32172), .B2(\pe6/aot [11]), 
        .ZN(n46655) );
  AOI21HSV2 U50453 ( .A1(n46656), .A2(n49685), .B(n46655), .ZN(n46660) );
  NAND2HSV0 U50454 ( .A1(n44435), .A2(\pe6/aot [1]), .ZN(n49841) );
  XNOR2HSV1 U50455 ( .A1(n46660), .A2(n46659), .ZN(n46667) );
  NAND2HSV0 U50456 ( .A1(n58731), .A2(n49760), .ZN(n49852) );
  NOR2HSV0 U50457 ( .A1(n48041), .A2(n46663), .ZN(n46664) );
  XNOR2HSV1 U50458 ( .A1(n46665), .A2(n46664), .ZN(n46666) );
  XNOR2HSV1 U50459 ( .A1(n46667), .A2(n46666), .ZN(n46668) );
  XNOR2HSV1 U50460 ( .A1(n46669), .A2(n46668), .ZN(n46704) );
  NAND2HSV0 U50461 ( .A1(n58976), .A2(n58856), .ZN(n46671) );
  NAND2HSV0 U50462 ( .A1(\pe6/bq[11] ), .A2(\pe6/aot [21]), .ZN(n46670) );
  XOR2HSV0 U50463 ( .A1(n46671), .A2(n46670), .Z(n46676) );
  NAND2HSV0 U50464 ( .A1(n46672), .A2(n58464), .ZN(n46674) );
  NAND2HSV0 U50465 ( .A1(n58962), .A2(n49831), .ZN(n46673) );
  XOR2HSV0 U50466 ( .A1(n46674), .A2(n46673), .Z(n46675) );
  XOR2HSV0 U50467 ( .A1(n46676), .A2(n46675), .Z(n46685) );
  CLKNHSV0 U50468 ( .I(n49327), .ZN(n59066) );
  NAND2HSV0 U50469 ( .A1(n59066), .A2(n46677), .ZN(n46679) );
  NAND2HSV0 U50470 ( .A1(n59084), .A2(\pe6/aot [23]), .ZN(n46678) );
  XOR2HSV0 U50471 ( .A1(n46679), .A2(n46678), .Z(n46683) );
  NAND2HSV0 U50472 ( .A1(n36150), .A2(n49208), .ZN(n46681) );
  NAND2HSV0 U50473 ( .A1(n59098), .A2(n58631), .ZN(n46680) );
  XOR2HSV0 U50474 ( .A1(n46681), .A2(n46680), .Z(n46682) );
  XOR2HSV0 U50475 ( .A1(n46683), .A2(n46682), .Z(n46684) );
  XOR2HSV0 U50476 ( .A1(n46685), .A2(n46684), .Z(n46702) );
  NAND2HSV0 U50477 ( .A1(n59206), .A2(n46792), .ZN(n46687) );
  CLKNHSV0 U50478 ( .I(n46147), .ZN(n58975) );
  NAND2HSV0 U50479 ( .A1(n58975), .A2(n59272), .ZN(n46686) );
  XOR2HSV0 U50480 ( .A1(n46687), .A2(n46686), .Z(n46692) );
  NAND2HSV0 U50481 ( .A1(n59045), .A2(\pe6/aot [17]), .ZN(n46690) );
  NAND2HSV0 U50482 ( .A1(\pe6/bq[17] ), .A2(\pe6/aot [15]), .ZN(n46689) );
  XOR2HSV0 U50483 ( .A1(n46690), .A2(n46689), .Z(n46691) );
  XOR2HSV0 U50484 ( .A1(n46692), .A2(n46691), .Z(n46700) );
  NAND2HSV0 U50485 ( .A1(n59217), .A2(n59266), .ZN(n46694) );
  NAND2HSV0 U50486 ( .A1(n59050), .A2(n58857), .ZN(n46693) );
  XOR2HSV0 U50487 ( .A1(n46694), .A2(n46693), .Z(n46698) );
  NOR2HSV0 U50488 ( .A1(n48887), .A2(n32086), .ZN(n46696) );
  NAND2HSV0 U50489 ( .A1(n59041), .A2(n59040), .ZN(n46695) );
  XOR2HSV0 U50490 ( .A1(n46696), .A2(n46695), .Z(n46697) );
  XOR2HSV0 U50491 ( .A1(n46698), .A2(n46697), .Z(n46699) );
  XOR2HSV0 U50492 ( .A1(n46700), .A2(n46699), .Z(n46701) );
  XOR2HSV0 U50493 ( .A1(n46702), .A2(n46701), .Z(n46703) );
  XOR3HSV2 U50494 ( .A1(n46705), .A2(n46704), .A3(n46703), .Z(n46706) );
  XNOR2HSV1 U50495 ( .A1(n46707), .A2(n46706), .ZN(n46709) );
  NAND2HSV0 U50496 ( .A1(n58940), .A2(\pe6/got [4]), .ZN(n46708) );
  XNOR2HSV1 U50497 ( .A1(n46709), .A2(n46708), .ZN(n46711) );
  BUFHSV2 U50498 ( .I(\pe6/got [5]), .Z(n59292) );
  NAND2HSV0 U50499 ( .A1(n59295), .A2(n59292), .ZN(n46710) );
  XNOR2HSV1 U50500 ( .A1(n46711), .A2(n46710), .ZN(n46712) );
  XNOR2HSV1 U50501 ( .A1(n46713), .A2(n46712), .ZN(n46714) );
  XNOR2HSV1 U50502 ( .A1(n46715), .A2(n46714), .ZN(n46717) );
  NAND2HSV0 U50503 ( .A1(n59917), .A2(n59182), .ZN(n46716) );
  XNOR2HSV1 U50504 ( .A1(n46717), .A2(n46716), .ZN(n46718) );
  XNOR2HSV1 U50505 ( .A1(n46719), .A2(n46718), .ZN(n46720) );
  XNOR2HSV1 U50506 ( .A1(n46721), .A2(n46720), .ZN(n46722) );
  XNOR2HSV1 U50507 ( .A1(n46723), .A2(n46722), .ZN(n46724) );
  XNOR2HSV1 U50508 ( .A1(n46725), .A2(n46724), .ZN(n46726) );
  XNOR2HSV1 U50509 ( .A1(n46727), .A2(n46726), .ZN(n46728) );
  XNOR2HSV1 U50510 ( .A1(n46729), .A2(n46728), .ZN(n46731) );
  BUFHSV2 U50511 ( .I(n35898), .Z(n59144) );
  NAND2HSV0 U50512 ( .A1(n59144), .A2(\pe6/got [15]), .ZN(n46730) );
  XNOR2HSV1 U50513 ( .A1(n46731), .A2(n46730), .ZN(n46732) );
  XOR2HSV0 U50514 ( .A1(n46733), .A2(n46732), .Z(n46734) );
  XOR2HSV0 U50515 ( .A1(n46735), .A2(n46734), .Z(n46736) );
  XNOR2HSV1 U50516 ( .A1(n46737), .A2(n46736), .ZN(n46738) );
  XNOR2HSV1 U50517 ( .A1(n46739), .A2(n46738), .ZN(n46741) );
  NAND2HSV0 U50518 ( .A1(n59915), .A2(n46818), .ZN(n46740) );
  XNOR2HSV1 U50519 ( .A1(n46741), .A2(n46740), .ZN(n46742) );
  XNOR2HSV1 U50520 ( .A1(n46743), .A2(n46742), .ZN(n46744) );
  XOR2HSV0 U50521 ( .A1(n46745), .A2(n46744), .Z(n46747) );
  NAND2HSV0 U50522 ( .A1(n58805), .A2(n49002), .ZN(n46746) );
  XOR2HSV0 U50523 ( .A1(n46747), .A2(n46746), .Z(n46748) );
  XNOR2HSV1 U50524 ( .A1(n46749), .A2(n46748), .ZN(n46752) );
  NOR2HSV0 U50525 ( .A1(n46823), .A2(n46750), .ZN(n46751) );
  XNOR2HSV1 U50526 ( .A1(n46752), .A2(n46751), .ZN(n46754) );
  NAND2HSV0 U50527 ( .A1(n53172), .A2(n59025), .ZN(n46753) );
  XNOR2HSV1 U50528 ( .A1(n46754), .A2(n46753), .ZN(n46755) );
  XNOR2HSV1 U50529 ( .A1(n46756), .A2(n46755), .ZN(n46757) );
  AO21HSV1 U50530 ( .A1(n59514), .A2(n59022), .B(n46757), .Z(n46759) );
  NAND3HSV1 U50531 ( .A1(n46757), .A2(n59514), .A3(n59171), .ZN(n46758) );
  NAND2HSV2 U50532 ( .A1(n46759), .A2(n46758), .ZN(n46762) );
  BUFHSV2 U50533 ( .I(n59570), .Z(n58712) );
  CLKNAND2HSV0 U50534 ( .A1(n46760), .A2(n58712), .ZN(n46761) );
  XOR2HSV0 U50535 ( .A1(n46762), .A2(n46761), .Z(n46763) );
  XNOR2HSV1 U50536 ( .A1(n46764), .A2(n46763), .ZN(n46768) );
  XOR2HSV0 U50537 ( .A1(n46768), .A2(n46767), .Z(\pe6/poht [1]) );
  INHSV2 U50538 ( .I(n49316), .ZN(n59169) );
  BUFHSV4 U50539 ( .I(n46822), .Z(n58657) );
  BUFHSV2 U50540 ( .I(n58448), .Z(n58660) );
  CLKNAND2HSV1 U50541 ( .A1(n58660), .A2(n58562), .ZN(n46813) );
  BUFHSV2 U50542 ( .I(\pe6/got [6]), .Z(n58659) );
  BUFHSV2 U50543 ( .I(n58659), .Z(n58513) );
  CLKNAND2HSV0 U50544 ( .A1(n58936), .A2(n58513), .ZN(n46811) );
  NAND2HSV0 U50545 ( .A1(n58662), .A2(n58479), .ZN(n46807) );
  NAND2HSV0 U50546 ( .A1(n58663), .A2(n58527), .ZN(n46805) );
  NAND2HSV0 U50547 ( .A1(n58664), .A2(n58724), .ZN(n46803) );
  BUFHSV2 U50548 ( .I(n50805), .Z(n49099) );
  CLKNAND2HSV1 U50549 ( .A1(n53114), .A2(n58403), .ZN(n46801) );
  NAND2HSV0 U50550 ( .A1(n59240), .A2(\pe6/aot [5]), .ZN(n46771) );
  INHSV2 U50551 ( .I(n58537), .ZN(n58495) );
  NAND2HSV0 U50552 ( .A1(n59246), .A2(n58495), .ZN(n46770) );
  XOR2HSV0 U50553 ( .A1(n46771), .A2(n46770), .Z(n46775) );
  NAND2HSV0 U50554 ( .A1(n35750), .A2(n53134), .ZN(n46773) );
  NAND2HSV0 U50555 ( .A1(n49205), .A2(n49208), .ZN(n46772) );
  XOR2HSV0 U50556 ( .A1(n46773), .A2(n46772), .Z(n46774) );
  XOR2HSV0 U50557 ( .A1(n46775), .A2(n46774), .Z(n46782) );
  CLKNAND2HSV0 U50558 ( .A1(n58405), .A2(\pe6/aot [11]), .ZN(n46777) );
  CLKNAND2HSV0 U50559 ( .A1(n58731), .A2(n32972), .ZN(n46776) );
  XOR2HSV0 U50560 ( .A1(n46777), .A2(n46776), .Z(n46780) );
  CLKNAND2HSV1 U50561 ( .A1(n58668), .A2(n59252), .ZN(n49330) );
  CLKNAND2HSV0 U50562 ( .A1(n58360), .A2(n58842), .ZN(n46778) );
  XOR2HSV0 U50563 ( .A1(n49330), .A2(n46778), .Z(n46779) );
  XOR2HSV0 U50564 ( .A1(n46780), .A2(n46779), .Z(n46781) );
  XOR2HSV0 U50565 ( .A1(n46782), .A2(n46781), .Z(n46799) );
  NAND2HSV0 U50566 ( .A1(n49106), .A2(\pe6/aot [13]), .ZN(n46784) );
  NAND2HSV0 U50567 ( .A1(n49844), .A2(\pe6/aot [1]), .ZN(n46783) );
  XOR2HSV0 U50568 ( .A1(n46784), .A2(n46783), .Z(n46788) );
  NOR2HSV0 U50569 ( .A1(n50847), .A2(n58483), .ZN(n46786) );
  BUFHSV2 U50570 ( .I(\pe6/aot [2]), .Z(n59260) );
  NAND2HSV0 U50571 ( .A1(n58682), .A2(n59260), .ZN(n46785) );
  XOR2HSV0 U50572 ( .A1(n46786), .A2(n46785), .Z(n46787) );
  XNOR2HSV1 U50573 ( .A1(n46788), .A2(n46787), .ZN(n46797) );
  NOR2HSV0 U50574 ( .A1(n46853), .A2(n58530), .ZN(n46791) );
  CLKNAND2HSV0 U50575 ( .A1(n58990), .A2(n35732), .ZN(n46790) );
  XOR2HSV0 U50576 ( .A1(n46791), .A2(n46790), .Z(n46795) );
  NOR2HSV0 U50577 ( .A1(n49680), .A2(n58463), .ZN(n49102) );
  NOR2HSV0 U50578 ( .A1(n48041), .A2(n58392), .ZN(n58598) );
  CLKNHSV0 U50579 ( .I(n48041), .ZN(n59075) );
  AOI22HSV0 U50580 ( .A1(n58962), .A2(n46792), .B1(\pe6/aot [10]), .B2(n59075), 
        .ZN(n46793) );
  AOI21HSV0 U50581 ( .A1(n49102), .A2(n58598), .B(n46793), .ZN(n46794) );
  XNOR2HSV1 U50582 ( .A1(n46795), .A2(n46794), .ZN(n46796) );
  XNOR2HSV1 U50583 ( .A1(n46797), .A2(n46796), .ZN(n46798) );
  XNOR2HSV1 U50584 ( .A1(n46799), .A2(n46798), .ZN(n46800) );
  XNOR2HSV1 U50585 ( .A1(n46801), .A2(n46800), .ZN(n46802) );
  XNOR2HSV1 U50586 ( .A1(n46803), .A2(n46802), .ZN(n46804) );
  XNOR2HSV1 U50587 ( .A1(n46805), .A2(n46804), .ZN(n46806) );
  XNOR2HSV1 U50588 ( .A1(n46807), .A2(n46806), .ZN(n46809) );
  BUFHSV2 U50589 ( .I(\pe6/got [5]), .Z(n58661) );
  CLKNAND2HSV0 U50590 ( .A1(n58702), .A2(n58478), .ZN(n46808) );
  XNOR2HSV1 U50591 ( .A1(n46809), .A2(n46808), .ZN(n46810) );
  XNOR2HSV1 U50592 ( .A1(n46811), .A2(n46810), .ZN(n46812) );
  XNOR2HSV1 U50593 ( .A1(n46813), .A2(n46812), .ZN(n46815) );
  BUFHSV2 U50594 ( .I(n49078), .Z(n59161) );
  CLKNAND2HSV0 U50595 ( .A1(n59161), .A2(n59182), .ZN(n46814) );
  XOR2HSV0 U50596 ( .A1(n46815), .A2(n46814), .Z(n46816) );
  CLKNHSV2 U50597 ( .I(n46819), .ZN(n46820) );
  INHSV2 U50598 ( .I(n46820), .ZN(n49738) );
  CLKNAND2HSV2 U50599 ( .A1(n49738), .A2(n49737), .ZN(n53106) );
  NOR2HSV1 U50600 ( .A1(n49178), .A2(n52710), .ZN(n53104) );
  NOR2HSV1 U50601 ( .A1(n53104), .A2(n32696), .ZN(n46821) );
  NAND2HSV2 U50602 ( .A1(n53106), .A2(n46821), .ZN(n46899) );
  BUFHSV4 U50603 ( .I(n49181), .Z(n53107) );
  NAND2HSV2 U50604 ( .A1(n53107), .A2(n59178), .ZN(n46895) );
  INHSV2 U50605 ( .I(n58447), .ZN(n58385) );
  CLKNAND2HSV1 U50606 ( .A1(n58385), .A2(n59031), .ZN(n46893) );
  CLKNAND2HSV0 U50607 ( .A1(n53109), .A2(n49741), .ZN(n46891) );
  CLKNAND2HSV1 U50608 ( .A1(n58717), .A2(n58811), .ZN(n46888) );
  CLKNAND2HSV0 U50609 ( .A1(n59918), .A2(n49742), .ZN(n46884) );
  NAND2HSV0 U50610 ( .A1(n58936), .A2(\pe6/got [10]), .ZN(n46882) );
  BUFHSV2 U50611 ( .I(n58662), .Z(n53111) );
  CLKNAND2HSV0 U50612 ( .A1(n53111), .A2(n59182), .ZN(n46878) );
  BUFHSV2 U50613 ( .I(n53112), .Z(n59030) );
  CLKNAND2HSV1 U50614 ( .A1(n59030), .A2(n58709), .ZN(n46876) );
  NAND2HSV0 U50615 ( .A1(n53113), .A2(n58513), .ZN(n46874) );
  NAND2HSV0 U50616 ( .A1(n53114), .A2(n58478), .ZN(n46872) );
  NAND2HSV0 U50617 ( .A1(n49667), .A2(\pe6/got [3]), .ZN(n46868) );
  BUFHSV2 U50618 ( .I(n59039), .Z(n59231) );
  NAND2HSV0 U50619 ( .A1(n59379), .A2(n59231), .ZN(n46866) );
  NAND2HSV0 U50620 ( .A1(n58813), .A2(n59235), .ZN(n46864) );
  NOR2HSV0 U50621 ( .A1(n46147), .A2(n44396), .ZN(n49101) );
  NAND2HSV0 U50622 ( .A1(n32606), .A2(\pe6/aot [1]), .ZN(n46826) );
  XOR2HSV0 U50623 ( .A1(n49101), .A2(n46826), .Z(n46830) );
  NOR2HSV0 U50624 ( .A1(n46688), .A2(n58530), .ZN(n46828) );
  NAND2HSV0 U50625 ( .A1(n58962), .A2(\pe6/aot [11]), .ZN(n46827) );
  XOR2HSV0 U50626 ( .A1(n46828), .A2(n46827), .Z(n46829) );
  XOR2HSV0 U50627 ( .A1(n46830), .A2(n46829), .Z(n46862) );
  CLKNAND2HSV0 U50628 ( .A1(n58668), .A2(\pe6/aot [7]), .ZN(n46832) );
  NAND2HSV0 U50629 ( .A1(n48044), .A2(n53115), .ZN(n46831) );
  XOR2HSV0 U50630 ( .A1(n46832), .A2(n46831), .Z(n46836) );
  NOR2HSV0 U50631 ( .A1(n58984), .A2(n58359), .ZN(n46834) );
  NAND2HSV0 U50632 ( .A1(n35751), .A2(n53134), .ZN(n46833) );
  XOR2HSV0 U50633 ( .A1(n46834), .A2(n46833), .Z(n46835) );
  XNOR2HSV1 U50634 ( .A1(n46836), .A2(n46835), .ZN(n46843) );
  NAND2HSV0 U50635 ( .A1(n49106), .A2(\pe6/aot [17]), .ZN(n58852) );
  OAI21HSV0 U50636 ( .A1(n49681), .A2(n59105), .B(n58852), .ZN(n46837) );
  OAI21HSV0 U50637 ( .A1(n58382), .A2(n46838), .B(n46837), .ZN(n46841) );
  NOR2HSV0 U50638 ( .A1(n48041), .A2(n46789), .ZN(n49835) );
  NOR2HSV0 U50639 ( .A1(n46146), .A2(n32858), .ZN(n53129) );
  AOI22HSV1 U50640 ( .A1(n59075), .A2(n49208), .B1(n59189), .B2(\pe6/bq[5] ), 
        .ZN(n46839) );
  AOI21HSV1 U50641 ( .A1(n49835), .A2(n53129), .B(n46839), .ZN(n46840) );
  XOR2HSV0 U50642 ( .A1(n46841), .A2(n46840), .Z(n46842) );
  XNOR2HSV1 U50643 ( .A1(n46843), .A2(n46842), .ZN(n46861) );
  NAND2HSV0 U50644 ( .A1(n59051), .A2(\pe6/aot [2]), .ZN(n46845) );
  NAND2HSV0 U50645 ( .A1(n58976), .A2(n58495), .ZN(n46844) );
  XOR2HSV0 U50646 ( .A1(n46845), .A2(n46844), .Z(n46849) );
  NAND2HSV0 U50647 ( .A1(n58360), .A2(\pe6/aot [19]), .ZN(n46847) );
  CLKNHSV0 U50648 ( .I(n48887), .ZN(n59277) );
  NAND2HSV0 U50649 ( .A1(n59277), .A2(n59264), .ZN(n46846) );
  XOR2HSV0 U50650 ( .A1(n46847), .A2(n46846), .Z(n46848) );
  XOR2HSV0 U50651 ( .A1(n46849), .A2(n46848), .Z(n46859) );
  NAND2HSV0 U50652 ( .A1(n35750), .A2(\pe6/aot [10]), .ZN(n46852) );
  NAND2HSV0 U50653 ( .A1(\pe6/bq[8] ), .A2(\pe6/aot [13]), .ZN(n46851) );
  XOR2HSV0 U50654 ( .A1(n46852), .A2(n46851), .Z(n46857) );
  NOR2HSV0 U50655 ( .A1(n49327), .A2(n32245), .ZN(n46855) );
  NAND2HSV0 U50656 ( .A1(n59265), .A2(\pe6/aot [8]), .ZN(n46854) );
  XOR2HSV0 U50657 ( .A1(n46855), .A2(n46854), .Z(n46856) );
  XOR2HSV0 U50658 ( .A1(n46857), .A2(n46856), .Z(n46858) );
  XOR2HSV0 U50659 ( .A1(n46859), .A2(n46858), .Z(n46860) );
  XOR3HSV2 U50660 ( .A1(n46862), .A2(n46861), .A3(n46860), .Z(n46863) );
  XNOR2HSV1 U50661 ( .A1(n46864), .A2(n46863), .ZN(n46865) );
  XNOR2HSV1 U50662 ( .A1(n46866), .A2(n46865), .ZN(n46867) );
  XNOR2HSV1 U50663 ( .A1(n46868), .A2(n46867), .ZN(n46870) );
  NAND2HSV0 U50664 ( .A1(n58901), .A2(n58479), .ZN(n46869) );
  XNOR2HSV1 U50665 ( .A1(n46870), .A2(n46869), .ZN(n46871) );
  XNOR2HSV1 U50666 ( .A1(n46872), .A2(n46871), .ZN(n46873) );
  XNOR2HSV1 U50667 ( .A1(n46874), .A2(n46873), .ZN(n46875) );
  XNOR2HSV1 U50668 ( .A1(n46876), .A2(n46875), .ZN(n46877) );
  XNOR2HSV1 U50669 ( .A1(n46878), .A2(n46877), .ZN(n46880) );
  CLKNAND2HSV1 U50670 ( .A1(n49726), .A2(\pe6/got [9]), .ZN(n46879) );
  XNOR2HSV1 U50671 ( .A1(n46880), .A2(n46879), .ZN(n46881) );
  XNOR2HSV1 U50672 ( .A1(n46882), .A2(n46881), .ZN(n46883) );
  XNOR2HSV1 U50673 ( .A1(n46884), .A2(n46883), .ZN(n46886) );
  NAND2HSV0 U50674 ( .A1(n58805), .A2(\pe6/got [12]), .ZN(n46885) );
  XOR2HSV0 U50675 ( .A1(n46886), .A2(n46885), .Z(n46887) );
  XNOR2HSV1 U50676 ( .A1(n46888), .A2(n46887), .ZN(n46890) );
  XOR3HSV2 U50677 ( .A1(n46891), .A2(n46890), .A3(n46889), .Z(n46892) );
  XNOR2HSV1 U50678 ( .A1(n46893), .A2(n46892), .ZN(n46894) );
  XOR2HSV0 U50679 ( .A1(n46895), .A2(n46894), .Z(n46897) );
  CLKNAND2HSV0 U50680 ( .A1(n58712), .A2(n58715), .ZN(n46896) );
  XOR2HSV0 U50681 ( .A1(n46897), .A2(n46896), .Z(n46898) );
  XNOR2HSV1 U50682 ( .A1(n46899), .A2(n46898), .ZN(n46900) );
  XNOR2HSV1 U50683 ( .A1(n46901), .A2(n46900), .ZN(\pe6/poht [12]) );
  CLKNAND2HSV1 U50684 ( .A1(n51016), .A2(n53285), .ZN(n46971) );
  BUFHSV2 U50685 ( .I(n59883), .Z(n46977) );
  NOR2HSV2 U50686 ( .A1(n53293), .A2(n47143), .ZN(n46965) );
  CLKNAND2HSV0 U50687 ( .A1(n53294), .A2(n59891), .ZN(n46959) );
  CLKNAND2HSV0 U50688 ( .A1(n48747), .A2(n50698), .ZN(n46957) );
  NAND2HSV0 U50689 ( .A1(n51018), .A2(n51200), .ZN(n46953) );
  NAND2HSV0 U50690 ( .A1(n59878), .A2(n51302), .ZN(n46949) );
  NAND2HSV0 U50691 ( .A1(n59392), .A2(n53211), .ZN(n46947) );
  NAND2HSV0 U50692 ( .A1(n52575), .A2(n53197), .ZN(n46945) );
  NAND2HSV0 U50693 ( .A1(n25854), .A2(n51362), .ZN(n46943) );
  NAND2HSV0 U50694 ( .A1(n50588), .A2(n52618), .ZN(n46903) );
  INHSV2 U50695 ( .I(n48031), .ZN(n53200) );
  NAND2HSV0 U50696 ( .A1(n52591), .A2(n53200), .ZN(n46902) );
  XOR2HSV0 U50697 ( .A1(n46903), .A2(n46902), .Z(n46907) );
  NAND2HSV2 U50698 ( .A1(\pe5/aot [13]), .A2(\pe5/bq[10] ), .ZN(n46905) );
  NAND2HSV0 U50699 ( .A1(\pe5/aot [16]), .A2(\pe5/bq[7] ), .ZN(n46904) );
  XOR2HSV0 U50700 ( .A1(n46905), .A2(n46904), .Z(n46906) );
  XOR2HSV0 U50701 ( .A1(n46907), .A2(n46906), .Z(n46915) );
  NAND2HSV0 U50702 ( .A1(n53299), .A2(\pe5/bq[11] ), .ZN(n46909) );
  NAND2HSV0 U50703 ( .A1(n59941), .A2(n53199), .ZN(n46908) );
  XOR2HSV0 U50704 ( .A1(n46909), .A2(n46908), .Z(n46913) );
  NOR2HSV0 U50705 ( .A1(n48246), .A2(n48186), .ZN(n46911) );
  NAND2HSV0 U50706 ( .A1(n59881), .A2(n50526), .ZN(n46910) );
  XOR2HSV0 U50707 ( .A1(n46911), .A2(n46910), .Z(n46912) );
  XOR2HSV0 U50708 ( .A1(n46913), .A2(n46912), .Z(n46914) );
  XOR2HSV0 U50709 ( .A1(n46915), .A2(n46914), .Z(n46925) );
  NOR2HSV0 U50710 ( .A1(n48823), .A2(n47162), .ZN(n51174) );
  NOR2HSV0 U50711 ( .A1(n59641), .A2(n46916), .ZN(n51028) );
  AOI22HSV0 U50712 ( .A1(n48681), .A2(n51307), .B1(n50653), .B2(n50675), .ZN(
        n46917) );
  AOI21HSV1 U50713 ( .A1(n51174), .A2(n51028), .B(n46917), .ZN(n46923) );
  NAND2HSV0 U50714 ( .A1(n59638), .A2(\pe5/bq[2] ), .ZN(n46919) );
  NAND2HSV0 U50715 ( .A1(n53296), .A2(n50500), .ZN(n46918) );
  XOR2HSV0 U50716 ( .A1(n46919), .A2(n46918), .Z(n46922) );
  CLKNAND2HSV1 U50717 ( .A1(n51182), .A2(n47291), .ZN(n48809) );
  XOR2HSV0 U50718 ( .A1(n48809), .A2(n46920), .Z(n46921) );
  XOR3HSV2 U50719 ( .A1(n46923), .A2(n46922), .A3(n46921), .Z(n46924) );
  XNOR2HSV1 U50720 ( .A1(n46925), .A2(n46924), .ZN(n46941) );
  NAND2HSV0 U50721 ( .A1(\pe5/aot [4]), .A2(n39454), .ZN(n46927) );
  NAND2HSV0 U50722 ( .A1(n40190), .A2(n53307), .ZN(n46926) );
  XOR2HSV0 U50723 ( .A1(n46927), .A2(n46926), .Z(n46931) );
  NAND2HSV0 U50724 ( .A1(\pe5/aot [18]), .A2(n52671), .ZN(n46929) );
  NAND2HSV0 U50725 ( .A1(\pe5/aot [7]), .A2(n48181), .ZN(n46928) );
  XOR2HSV0 U50726 ( .A1(n46929), .A2(n46928), .Z(n46930) );
  XOR2HSV0 U50727 ( .A1(n46931), .A2(n46930), .Z(n46939) );
  CLKNAND2HSV0 U50728 ( .A1(n53295), .A2(n51176), .ZN(n48679) );
  XOR2HSV0 U50729 ( .A1(n46932), .A2(n48679), .Z(n46937) );
  NAND2HSV0 U50730 ( .A1(\pe5/aot [10]), .A2(n39471), .ZN(n46935) );
  NAND2HSV0 U50731 ( .A1(n53203), .A2(n46933), .ZN(n46934) );
  XOR2HSV0 U50732 ( .A1(n46935), .A2(n46934), .Z(n46936) );
  XOR2HSV0 U50733 ( .A1(n46937), .A2(n46936), .Z(n46938) );
  XOR2HSV0 U50734 ( .A1(n46939), .A2(n46938), .Z(n46940) );
  XNOR2HSV1 U50735 ( .A1(n46941), .A2(n46940), .ZN(n46942) );
  XNOR2HSV1 U50736 ( .A1(n46943), .A2(n46942), .ZN(n46944) );
  XNOR2HSV1 U50737 ( .A1(n46945), .A2(n46944), .ZN(n46946) );
  XNOR2HSV1 U50738 ( .A1(n46947), .A2(n46946), .ZN(n46948) );
  XNOR2HSV1 U50739 ( .A1(n46949), .A2(n46948), .ZN(n46951) );
  NAND2HSV0 U50740 ( .A1(n44694), .A2(n52576), .ZN(n46950) );
  XOR2HSV0 U50741 ( .A1(n46951), .A2(n46950), .Z(n46952) );
  XNOR2HSV1 U50742 ( .A1(n46953), .A2(n46952), .ZN(n46955) );
  NAND2HSV0 U50743 ( .A1(n51205), .A2(n51359), .ZN(n46954) );
  XNOR2HSV1 U50744 ( .A1(n46955), .A2(n46954), .ZN(n46956) );
  XNOR2HSV1 U50745 ( .A1(n46957), .A2(n46956), .ZN(n46958) );
  XNOR2HSV1 U50746 ( .A1(n46959), .A2(n46958), .ZN(n46963) );
  INHSV4 U50747 ( .I(n46961), .ZN(n50424) );
  CLKNAND2HSV0 U50748 ( .A1(n51211), .A2(n50424), .ZN(n46962) );
  XNOR2HSV1 U50749 ( .A1(n46963), .A2(n46962), .ZN(n46964) );
  XNOR2HSV1 U50750 ( .A1(n46965), .A2(n46964), .ZN(n46969) );
  CLKNAND2HSV1 U50751 ( .A1(n53338), .A2(\pe5/got [12]), .ZN(n46968) );
  NOR2HSV2 U50752 ( .A1(n52659), .A2(n45817), .ZN(n46967) );
  XOR3HSV2 U50753 ( .A1(n46969), .A2(n46968), .A3(n46967), .Z(n46970) );
  XNOR2HSV1 U50754 ( .A1(n46971), .A2(n46970), .ZN(n46973) );
  CLKNHSV0 U50755 ( .I(n39554), .ZN(n51092) );
  CLKNAND2HSV0 U50756 ( .A1(n51092), .A2(n50643), .ZN(n46972) );
  INHSV2 U50757 ( .I(n53188), .ZN(n53190) );
  INHSV4 U50758 ( .I(n53358), .ZN(n50421) );
  INHSV4 U50759 ( .I(n50421), .ZN(n51013) );
  CLKNAND2HSV1 U50760 ( .A1(n53188), .A2(n39241), .ZN(n53359) );
  CLKNAND2HSV0 U50761 ( .A1(n53359), .A2(n51103), .ZN(n46975) );
  NOR2HSV2 U50762 ( .A1(n51013), .A2(n46975), .ZN(n47051) );
  NAND2HSV2 U50763 ( .A1(n52563), .A2(n59949), .ZN(n47047) );
  INHSV2 U50764 ( .I(n47199), .ZN(n51014) );
  CLKNAND2HSV1 U50765 ( .A1(n52835), .A2(n52658), .ZN(n47045) );
  INHSV2 U50766 ( .I(n46976), .ZN(n52565) );
  CLKNAND2HSV1 U50767 ( .A1(n52565), .A2(n52652), .ZN(n47040) );
  CLKNAND2HSV1 U50768 ( .A1(n51016), .A2(\pe5/got [12]), .ZN(n47036) );
  NOR2HSV1 U50769 ( .A1(n53293), .A2(n46119), .ZN(n47031) );
  CLKNHSV0 U50770 ( .I(n46978), .ZN(n51017) );
  CLKNAND2HSV1 U50771 ( .A1(n53294), .A2(n51017), .ZN(n47027) );
  NAND2HSV0 U50772 ( .A1(n59882), .A2(n51200), .ZN(n47025) );
  CLKNAND2HSV0 U50773 ( .A1(n51018), .A2(\pe5/got [4]), .ZN(n47021) );
  BUFHSV2 U50774 ( .I(n59878), .Z(n51019) );
  CLKNAND2HSV0 U50775 ( .A1(n51019), .A2(n53197), .ZN(n47017) );
  NAND2HSV0 U50776 ( .A1(n59392), .A2(n51362), .ZN(n47015) );
  NOR2HSV0 U50777 ( .A1(n48246), .A2(n50428), .ZN(n52622) );
  NAND2HSV0 U50778 ( .A1(n51363), .A2(n48181), .ZN(n50499) );
  XOR2HSV0 U50779 ( .A1(n52622), .A2(n50499), .Z(n46982) );
  NOR2HSV0 U50780 ( .A1(n59869), .A2(n48822), .ZN(n46980) );
  NAND2HSV0 U50781 ( .A1(\pe5/aot [13]), .A2(n50675), .ZN(n46979) );
  XOR2HSV0 U50782 ( .A1(n46980), .A2(n46979), .Z(n46981) );
  XOR2HSV0 U50783 ( .A1(n46982), .A2(n46981), .Z(n47013) );
  NAND2HSV0 U50784 ( .A1(n59943), .A2(n50526), .ZN(n46984) );
  NAND2HSV0 U50785 ( .A1(\pe5/aot [18]), .A2(n51281), .ZN(n46983) );
  XOR2HSV0 U50786 ( .A1(n46984), .A2(n46983), .Z(n46988) );
  NAND2HSV0 U50787 ( .A1(n48199), .A2(\pe5/bq[2] ), .ZN(n46986) );
  NAND2HSV0 U50788 ( .A1(n52607), .A2(n53307), .ZN(n46985) );
  XOR2HSV0 U50789 ( .A1(n46986), .A2(n46985), .Z(n46987) );
  XOR2HSV0 U50790 ( .A1(n46988), .A2(n46987), .Z(n46996) );
  NAND2HSV0 U50791 ( .A1(n53299), .A2(n50533), .ZN(n46990) );
  NAND2HSV0 U50792 ( .A1(\pe5/aot [14]), .A2(\pe5/bq[7] ), .ZN(n46989) );
  XOR2HSV0 U50793 ( .A1(n46990), .A2(n46989), .Z(n46994) );
  CLKNAND2HSV0 U50794 ( .A1(n59866), .A2(\pe5/bq[11] ), .ZN(n51163) );
  NAND2HSV0 U50795 ( .A1(n51313), .A2(\pe5/bq[19] ), .ZN(n47324) );
  NOR2HSV0 U50796 ( .A1(n51163), .A2(n47324), .ZN(n46992) );
  AOI22HSV0 U50797 ( .A1(n51313), .A2(n39592), .B1(\pe5/bq[19] ), .B2(n51419), 
        .ZN(n46991) );
  NOR2HSV2 U50798 ( .A1(n46992), .A2(n46991), .ZN(n46993) );
  XNOR2HSV1 U50799 ( .A1(n46994), .A2(n46993), .ZN(n46995) );
  XNOR2HSV1 U50800 ( .A1(n46996), .A2(n46995), .ZN(n47012) );
  NAND2HSV0 U50801 ( .A1(n53304), .A2(\pe5/bq[14] ), .ZN(n46998) );
  NAND2HSV0 U50802 ( .A1(\pe5/aot [4]), .A2(n51176), .ZN(n46997) );
  XOR2HSV0 U50803 ( .A1(n46998), .A2(n46997), .Z(n47002) );
  INHSV2 U50804 ( .I(n48204), .ZN(n59897) );
  NAND2HSV0 U50805 ( .A1(n59897), .A2(n53216), .ZN(n47000) );
  NAND2HSV0 U50806 ( .A1(\pe5/aot [16]), .A2(n50504), .ZN(n46999) );
  XOR2HSV0 U50807 ( .A1(n47000), .A2(n46999), .Z(n47001) );
  XOR2HSV0 U50808 ( .A1(n47002), .A2(n47001), .Z(n47010) );
  NAND2HSV0 U50809 ( .A1(n53296), .A2(\pe5/bq[13] ), .ZN(n47004) );
  NAND2HSV0 U50810 ( .A1(n53295), .A2(n53314), .ZN(n47003) );
  XOR2HSV0 U50811 ( .A1(n47004), .A2(n47003), .Z(n47008) );
  NOR2HSV0 U50812 ( .A1(n45904), .A2(n45426), .ZN(n47006) );
  NAND2HSV0 U50813 ( .A1(n52591), .A2(n51276), .ZN(n47005) );
  XOR2HSV0 U50814 ( .A1(n47006), .A2(n47005), .Z(n47007) );
  XOR2HSV0 U50815 ( .A1(n47008), .A2(n47007), .Z(n47009) );
  XOR2HSV0 U50816 ( .A1(n47010), .A2(n47009), .Z(n47011) );
  XOR3HSV2 U50817 ( .A1(n47013), .A2(n47012), .A3(n47011), .Z(n47014) );
  XNOR2HSV1 U50818 ( .A1(n47015), .A2(n47014), .ZN(n47016) );
  XNOR2HSV1 U50819 ( .A1(n47017), .A2(n47016), .ZN(n47019) );
  NAND2HSV0 U50820 ( .A1(n44694), .A2(n53211), .ZN(n47018) );
  XOR2HSV0 U50821 ( .A1(n47019), .A2(n47018), .Z(n47020) );
  XNOR2HSV1 U50822 ( .A1(n47021), .A2(n47020), .ZN(n47023) );
  NOR2HSV0 U50823 ( .A1(n50617), .A2(n53292), .ZN(n47022) );
  XNOR2HSV1 U50824 ( .A1(n47023), .A2(n47022), .ZN(n47024) );
  XNOR2HSV1 U50825 ( .A1(n47025), .A2(n47024), .ZN(n47026) );
  XNOR2HSV1 U50826 ( .A1(n47027), .A2(n47026), .ZN(n47029) );
  NAND2HSV0 U50827 ( .A1(n52653), .A2(n50698), .ZN(n47028) );
  XNOR2HSV1 U50828 ( .A1(n47029), .A2(n47028), .ZN(n47030) );
  XNOR2HSV1 U50829 ( .A1(n47031), .A2(n47030), .ZN(n47034) );
  CLKNAND2HSV0 U50830 ( .A1(n48745), .A2(n50424), .ZN(n47033) );
  NOR2HSV1 U50831 ( .A1(n51273), .A2(n47143), .ZN(n47032) );
  XOR3HSV2 U50832 ( .A1(n47034), .A2(n47033), .A3(n47032), .Z(n47035) );
  XNOR2HSV1 U50833 ( .A1(n47036), .A2(n47035), .ZN(n47038) );
  INHSV2 U50834 ( .I(n45817), .ZN(n53286) );
  NAND2HSV0 U50835 ( .A1(n51092), .A2(n53286), .ZN(n47037) );
  XOR2HSV0 U50836 ( .A1(n47038), .A2(n47037), .Z(n47039) );
  XNOR2HSV1 U50837 ( .A1(n47040), .A2(n47039), .ZN(n47043) );
  BUFHSV2 U50838 ( .I(n47041), .Z(n51227) );
  CLKBUFHSV4 U50839 ( .I(n51227), .Z(n51335) );
  CLKNAND2HSV1 U50840 ( .A1(n51335), .A2(n50643), .ZN(n47042) );
  XNOR2HSV1 U50841 ( .A1(n47043), .A2(n47042), .ZN(n47044) );
  XNOR2HSV1 U50842 ( .A1(n47045), .A2(n47044), .ZN(n47046) );
  NAND2HSV2 U50843 ( .A1(n29775), .A2(n50495), .ZN(n47048) );
  XOR2HSV2 U50844 ( .A1(n47051), .A2(n47050), .Z(n47055) );
  INHSV2 U50845 ( .I(n47052), .ZN(n47389) );
  INHSV2 U50846 ( .I(n47389), .ZN(n47195) );
  CLKNAND2HSV0 U50847 ( .A1(n47387), .A2(n47052), .ZN(n53361) );
  AND2HSV2 U50848 ( .A1(n53361), .A2(n45816), .Z(n47053) );
  CLKNAND2HSV1 U50849 ( .A1(n53363), .A2(n47053), .ZN(n47054) );
  XNOR2HSV1 U50850 ( .A1(n47055), .A2(n47054), .ZN(\pe5/poht [12]) );
  CLKNAND2HSV1 U50851 ( .A1(n53291), .A2(n51156), .ZN(n47136) );
  NOR2HSV0 U50852 ( .A1(n47057), .A2(n31199), .ZN(n47131) );
  NAND2HSV0 U50853 ( .A1(n52570), .A2(n53349), .ZN(n47126) );
  NAND2HSV0 U50854 ( .A1(n51018), .A2(n59891), .ZN(n47122) );
  CLKNAND2HSV1 U50855 ( .A1(n51019), .A2(n52573), .ZN(n47118) );
  NAND2HSV0 U50856 ( .A1(n45820), .A2(n51200), .ZN(n47116) );
  CLKNAND2HSV0 U50857 ( .A1(n52575), .A2(n52576), .ZN(n47114) );
  NAND2HSV0 U50858 ( .A1(n39745), .A2(n52577), .ZN(n47112) );
  INHSV2 U50859 ( .I(n51231), .ZN(n52579) );
  NAND2HSV0 U50860 ( .A1(n52578), .A2(n52579), .ZN(n47110) );
  NAND2HSV0 U50861 ( .A1(n59381), .A2(n51161), .ZN(n47108) );
  NAND2HSV0 U50862 ( .A1(n47338), .A2(n51362), .ZN(n47106) );
  NAND2HSV0 U50863 ( .A1(n59940), .A2(\pe5/bq[2] ), .ZN(n47061) );
  NAND2HSV0 U50864 ( .A1(\pe5/aot [4]), .A2(n47059), .ZN(n47060) );
  XOR2HSV0 U50865 ( .A1(n47061), .A2(n47060), .Z(n47065) );
  NAND2HSV0 U50866 ( .A1(n59866), .A2(n30891), .ZN(n47063) );
  NAND2HSV0 U50867 ( .A1(n59881), .A2(n51307), .ZN(n47062) );
  XOR2HSV0 U50868 ( .A1(n47063), .A2(n47062), .Z(n47064) );
  XOR2HSV0 U50869 ( .A1(n47065), .A2(n47064), .Z(n47073) );
  NAND2HSV0 U50870 ( .A1(n48681), .A2(n52619), .ZN(n47067) );
  NAND2HSV0 U50871 ( .A1(n53323), .A2(n39914), .ZN(n47066) );
  XOR2HSV0 U50872 ( .A1(n47067), .A2(n47066), .Z(n47071) );
  NAND2HSV0 U50873 ( .A1(n47278), .A2(\pe5/bq[11] ), .ZN(n47069) );
  NAND2HSV0 U50874 ( .A1(n52600), .A2(n30607), .ZN(n47068) );
  XOR2HSV0 U50875 ( .A1(n47069), .A2(n47068), .Z(n47070) );
  XOR2HSV0 U50876 ( .A1(n47071), .A2(n47070), .Z(n47072) );
  XOR2HSV0 U50877 ( .A1(n47073), .A2(n47072), .Z(n47089) );
  CLKNAND2HSV0 U50878 ( .A1(n37700), .A2(n52630), .ZN(n47075) );
  NAND2HSV0 U50879 ( .A1(n48761), .A2(n52581), .ZN(n47074) );
  XOR2HSV0 U50880 ( .A1(n47075), .A2(n47074), .Z(n47079) );
  NAND2HSV0 U50881 ( .A1(\pe5/aot [23]), .A2(n53200), .ZN(n47077) );
  NAND2HSV0 U50882 ( .A1(n59880), .A2(n52618), .ZN(n47076) );
  XOR2HSV0 U50883 ( .A1(n47077), .A2(n47076), .Z(n47078) );
  XOR2HSV0 U50884 ( .A1(n47079), .A2(n47078), .Z(n47087) );
  NAND2HSV0 U50885 ( .A1(\pe5/aot [18]), .A2(\pe5/bq[8] ), .ZN(n47081) );
  NAND2HSV0 U50886 ( .A1(n52591), .A2(n50526), .ZN(n47080) );
  XOR2HSV0 U50887 ( .A1(n47081), .A2(n47080), .Z(n47085) );
  NAND2HSV0 U50888 ( .A1(n53295), .A2(n48237), .ZN(n47083) );
  NAND2HSV0 U50889 ( .A1(n59942), .A2(\pe5/bq[7] ), .ZN(n47082) );
  XOR2HSV0 U50890 ( .A1(n47083), .A2(n47082), .Z(n47084) );
  XOR2HSV0 U50891 ( .A1(n47085), .A2(n47084), .Z(n47086) );
  XOR2HSV0 U50892 ( .A1(n47087), .A2(n47086), .Z(n47088) );
  XOR2HSV0 U50893 ( .A1(n47089), .A2(n47088), .Z(n47104) );
  NOR2HSV0 U50894 ( .A1(n47230), .A2(n46134), .ZN(n47232) );
  NAND2HSV0 U50895 ( .A1(n50588), .A2(n46933), .ZN(n47090) );
  XOR2HSV0 U50896 ( .A1(n47232), .A2(n47090), .Z(n47102) );
  NAND2HSV0 U50897 ( .A1(n52584), .A2(n52632), .ZN(n47092) );
  CLKNAND2HSV0 U50898 ( .A1(n52631), .A2(n51177), .ZN(n47091) );
  XOR2HSV0 U50899 ( .A1(n47092), .A2(n47091), .Z(n47093) );
  NAND2HSV0 U50900 ( .A1(n39887), .A2(n52595), .ZN(n51040) );
  XNOR2HSV1 U50901 ( .A1(n47093), .A2(n51040), .ZN(n47101) );
  NAND2HSV0 U50902 ( .A1(\pe5/aot [13]), .A2(n50668), .ZN(n47095) );
  NAND2HSV0 U50903 ( .A1(n51313), .A2(n52610), .ZN(n47094) );
  XOR2HSV0 U50904 ( .A1(n47095), .A2(n47094), .Z(n47099) );
  NOR2HSV0 U50905 ( .A1(n45904), .A2(n30287), .ZN(n47097) );
  NAND2HSV0 U50906 ( .A1(\pe5/aot [16]), .A2(\pe5/bq[10] ), .ZN(n47096) );
  XOR2HSV0 U50907 ( .A1(n47097), .A2(n47096), .Z(n47098) );
  XOR2HSV0 U50908 ( .A1(n47099), .A2(n47098), .Z(n47100) );
  XOR3HSV2 U50909 ( .A1(n47102), .A2(n47101), .A3(n47100), .Z(n47103) );
  XNOR2HSV1 U50910 ( .A1(n47104), .A2(n47103), .ZN(n47105) );
  XNOR2HSV1 U50911 ( .A1(n47106), .A2(n47105), .ZN(n47107) );
  XNOR2HSV1 U50912 ( .A1(n47108), .A2(n47107), .ZN(n47109) );
  XNOR2HSV1 U50913 ( .A1(n47110), .A2(n47109), .ZN(n47111) );
  XNOR2HSV1 U50914 ( .A1(n47112), .A2(n47111), .ZN(n47113) );
  XNOR2HSV1 U50915 ( .A1(n47114), .A2(n47113), .ZN(n47115) );
  XNOR2HSV1 U50916 ( .A1(n47116), .A2(n47115), .ZN(n47117) );
  XNOR2HSV1 U50917 ( .A1(n47118), .A2(n47117), .ZN(n47120) );
  NAND2HSV0 U50918 ( .A1(n44694), .A2(n47144), .ZN(n47119) );
  XOR2HSV0 U50919 ( .A1(n47120), .A2(n47119), .Z(n47121) );
  XNOR2HSV1 U50920 ( .A1(n47122), .A2(n47121), .ZN(n47124) );
  NAND2HSV0 U50921 ( .A1(n51205), .A2(n50424), .ZN(n47123) );
  XNOR2HSV1 U50922 ( .A1(n47124), .A2(n47123), .ZN(n47125) );
  XNOR2HSV1 U50923 ( .A1(n47126), .A2(n47125), .ZN(n47129) );
  CLKNAND2HSV1 U50924 ( .A1(n53294), .A2(n48167), .ZN(n47128) );
  NAND2HSV0 U50925 ( .A1(n52653), .A2(n53286), .ZN(n47127) );
  XOR3HSV2 U50926 ( .A1(n47129), .A2(n47128), .A3(n47127), .Z(n47130) );
  XNOR2HSV1 U50927 ( .A1(n47131), .A2(n47130), .ZN(n47134) );
  CLKNAND2HSV0 U50928 ( .A1(n53338), .A2(n50643), .ZN(n47133) );
  NOR2HSV1 U50929 ( .A1(n51273), .A2(n30888), .ZN(n47132) );
  XOR3HSV2 U50930 ( .A1(n47134), .A2(n47133), .A3(n47132), .Z(n47135) );
  XNOR2HSV1 U50931 ( .A1(n47136), .A2(n47135), .ZN(n47138) );
  NAND2HSV0 U50932 ( .A1(n59516), .A2(n52566), .ZN(n47137) );
  NAND2HSV4 U50933 ( .A1(n47141), .A2(n47195), .ZN(n48886) );
  NAND2HSV0 U50934 ( .A1(n53359), .A2(n59367), .ZN(n47142) );
  NOR2HSV2 U50935 ( .A1(n51013), .A2(n47142), .ZN(n47194) );
  INHSV2 U50936 ( .I(n47139), .ZN(n52563) );
  NAND2HSV2 U50937 ( .A1(n52563), .A2(n53349), .ZN(n47191) );
  CLKNAND2HSV1 U50938 ( .A1(n51272), .A2(n53289), .ZN(n47189) );
  CLKNAND2HSV1 U50939 ( .A1(n47268), .A2(n47144), .ZN(n47186) );
  NAND2HSV0 U50940 ( .A1(n59893), .A2(n51200), .ZN(n47183) );
  NOR2HSV1 U50941 ( .A1(n51273), .A2(n53292), .ZN(n47181) );
  NAND2HSV0 U50942 ( .A1(n59903), .A2(n51418), .ZN(n47179) );
  NOR2HSV1 U50943 ( .A1(n53293), .A2(n51231), .ZN(n47177) );
  NAND2HSV0 U50944 ( .A1(n59894), .A2(n51362), .ZN(n47173) );
  NAND2HSV0 U50945 ( .A1(\pe5/aot [14]), .A2(n53199), .ZN(n47147) );
  NAND2HSV0 U50946 ( .A1(n52675), .A2(\pe5/bq[7] ), .ZN(n47146) );
  XOR2HSV0 U50947 ( .A1(n47147), .A2(n47146), .Z(n47151) );
  NAND2HSV0 U50948 ( .A1(n51247), .A2(n52672), .ZN(n47149) );
  NAND2HSV0 U50949 ( .A1(n59896), .A2(n51281), .ZN(n47148) );
  XOR2HSV0 U50950 ( .A1(n47149), .A2(n47148), .Z(n47150) );
  XOR2HSV0 U50951 ( .A1(n47151), .A2(n47150), .Z(n47159) );
  NAND2HSV0 U50952 ( .A1(\pe5/aot [13]), .A2(\pe5/bq[2] ), .ZN(n47153) );
  NAND2HSV0 U50953 ( .A1(n51313), .A2(n52671), .ZN(n47152) );
  XOR2HSV0 U50954 ( .A1(n47153), .A2(n47152), .Z(n47157) );
  NAND2HSV0 U50955 ( .A1(\pe5/aot [9]), .A2(n50526), .ZN(n47155) );
  NAND2HSV0 U50956 ( .A1(n51339), .A2(n52632), .ZN(n47154) );
  XOR2HSV0 U50957 ( .A1(n47155), .A2(n47154), .Z(n47156) );
  XOR2HSV0 U50958 ( .A1(n47157), .A2(n47156), .Z(n47158) );
  XOR2HSV0 U50959 ( .A1(n47159), .A2(n47158), .Z(n47171) );
  NAND2HSV0 U50960 ( .A1(n50588), .A2(n53216), .ZN(n47161) );
  CLKNAND2HSV0 U50961 ( .A1(\pe5/aot [3]), .A2(n31045), .ZN(n47160) );
  XOR2HSV0 U50962 ( .A1(n47161), .A2(n47160), .Z(n47166) );
  NAND2HSV0 U50963 ( .A1(\pe5/aot [4]), .A2(\pe5/bq[11] ), .ZN(n47164) );
  NAND2HSV0 U50964 ( .A1(n51310), .A2(\pe5/bq[9] ), .ZN(n47163) );
  XOR2HSV0 U50965 ( .A1(n47164), .A2(n47163), .Z(n47165) );
  XNOR2HSV1 U50966 ( .A1(n47166), .A2(n47165), .ZN(n47169) );
  CLKNAND2HSV1 U50967 ( .A1(n48786), .A2(n50668), .ZN(n48196) );
  NAND2HSV0 U50968 ( .A1(n53323), .A2(n51370), .ZN(n47167) );
  XOR2HSV0 U50969 ( .A1(n48196), .A2(n47167), .Z(n47168) );
  XNOR2HSV1 U50970 ( .A1(n47169), .A2(n47168), .ZN(n47170) );
  XNOR2HSV1 U50971 ( .A1(n47171), .A2(n47170), .ZN(n47172) );
  XNOR2HSV1 U50972 ( .A1(n47173), .A2(n47172), .ZN(n47175) );
  NAND2HSV0 U50973 ( .A1(n52653), .A2(\pe5/got [2]), .ZN(n47174) );
  XNOR2HSV1 U50974 ( .A1(n47175), .A2(n47174), .ZN(n47176) );
  XNOR2HSV1 U50975 ( .A1(n47177), .A2(n47176), .ZN(n47178) );
  XNOR2HSV1 U50976 ( .A1(n47179), .A2(n47178), .ZN(n47180) );
  XOR2HSV0 U50977 ( .A1(n47181), .A2(n47180), .Z(n47182) );
  XNOR2HSV1 U50978 ( .A1(n47183), .A2(n47182), .ZN(n47185) );
  NAND2HSV0 U50979 ( .A1(n51399), .A2(n59905), .ZN(n47184) );
  CLKNAND2HSV0 U50980 ( .A1(n51404), .A2(n51358), .ZN(n47187) );
  NAND2HSV2 U50981 ( .A1(n29778), .A2(n48167), .ZN(n47192) );
  CLKXOR2HSV2 U50982 ( .A1(n47194), .A2(n47193), .Z(n47198) );
  NAND2HSV4 U50983 ( .A1(n47196), .A2(n47195), .ZN(n51109) );
  BUFHSV2 U50984 ( .I(n53361), .Z(n51108) );
  NAND3HSV2 U50985 ( .A1(n51109), .A2(n40186), .A3(n51108), .ZN(n47197) );
  XNOR2HSV1 U50986 ( .A1(n47198), .A2(n47197), .ZN(\pe5/poht [18]) );
  CLKNAND2HSV0 U50987 ( .A1(n48165), .A2(n39432), .ZN(n47264) );
  NOR2HSV0 U50988 ( .A1(n51361), .A2(n30888), .ZN(n47259) );
  CLKNAND2HSV0 U50989 ( .A1(n52569), .A2(n52652), .ZN(n47255) );
  NAND2HSV0 U50990 ( .A1(n52570), .A2(n52568), .ZN(n47253) );
  NAND2HSV0 U50991 ( .A1(n52572), .A2(n51305), .ZN(n47249) );
  NAND2HSV0 U50992 ( .A1(n59878), .A2(n59891), .ZN(n47245) );
  NAND2HSV0 U50993 ( .A1(n50501), .A2(\pe5/bq[24] ), .ZN(n47202) );
  NAND2HSV0 U50994 ( .A1(n52682), .A2(n47291), .ZN(n47201) );
  XOR2HSV0 U50995 ( .A1(n47202), .A2(n47201), .Z(n47206) );
  NAND2HSV0 U50996 ( .A1(n59879), .A2(\pe5/bq[2] ), .ZN(n47204) );
  NAND2HSV0 U50997 ( .A1(n48199), .A2(n48775), .ZN(n47203) );
  XOR2HSV0 U50998 ( .A1(n47204), .A2(n47203), .Z(n47205) );
  XOR2HSV0 U50999 ( .A1(n47206), .A2(n47205), .Z(n47215) );
  NAND2HSV0 U51000 ( .A1(n48829), .A2(n52581), .ZN(n47209) );
  NAND2HSV0 U51001 ( .A1(n51187), .A2(\pe5/bq[7] ), .ZN(n47208) );
  XOR2HSV0 U51002 ( .A1(n47209), .A2(n47208), .Z(n47213) );
  NAND2HSV0 U51003 ( .A1(n48681), .A2(n52632), .ZN(n47211) );
  NAND2HSV0 U51004 ( .A1(\pe5/aot [18]), .A2(n48778), .ZN(n47210) );
  XOR2HSV0 U51005 ( .A1(n47211), .A2(n47210), .Z(n47212) );
  XOR2HSV0 U51006 ( .A1(n47213), .A2(n47212), .Z(n47214) );
  NAND2HSV0 U51007 ( .A1(n37660), .A2(n51177), .ZN(n47217) );
  NAND2HSV0 U51008 ( .A1(\pe5/aot [20]), .A2(\pe5/bq[8] ), .ZN(n47216) );
  XOR2HSV0 U51009 ( .A1(n47217), .A2(n47216), .Z(n47221) );
  NAND2HSV0 U51010 ( .A1(n48761), .A2(n53200), .ZN(n47219) );
  NAND2HSV0 U51011 ( .A1(n52584), .A2(n52610), .ZN(n47218) );
  XOR2HSV0 U51012 ( .A1(n47219), .A2(n47218), .Z(n47220) );
  XOR2HSV0 U51013 ( .A1(n47221), .A2(n47220), .Z(n47229) );
  NAND2HSV0 U51014 ( .A1(n52611), .A2(n51176), .ZN(n47223) );
  NAND2HSV0 U51015 ( .A1(n51188), .A2(n51191), .ZN(n47222) );
  XOR2HSV0 U51016 ( .A1(n47223), .A2(n47222), .Z(n47227) );
  NAND2HSV0 U51017 ( .A1(n47278), .A2(n50668), .ZN(n47224) );
  XOR2HSV0 U51018 ( .A1(n47225), .A2(n47224), .Z(n47226) );
  XOR2HSV0 U51019 ( .A1(n47227), .A2(n47226), .Z(n47228) );
  AOI22HSV0 U51020 ( .A1(\pe5/aot [9]), .A2(n39454), .B1(n48206), .B2(n59944), 
        .ZN(n47231) );
  AOI21HSV1 U51021 ( .A1(n47233), .A2(n47232), .B(n47231), .ZN(n47235) );
  NAND2HSV0 U51022 ( .A1(n59895), .A2(n47234), .ZN(n47310) );
  NAND2HSV0 U51023 ( .A1(n50511), .A2(n39487), .ZN(n47237) );
  NAND2HSV0 U51024 ( .A1(n51313), .A2(n51167), .ZN(n47236) );
  XOR2HSV0 U51025 ( .A1(n47237), .A2(n47236), .Z(n47240) );
  NOR2HSV0 U51026 ( .A1(n47409), .A2(n39772), .ZN(n48675) );
  INHSV2 U51027 ( .I(n51232), .ZN(n59866) );
  NAND2HSV0 U51028 ( .A1(n52607), .A2(\pe5/bq[11] ), .ZN(n47314) );
  NAND2HSV0 U51029 ( .A1(\pe5/aot [16]), .A2(n52619), .ZN(n50510) );
  XOR2HSV0 U51030 ( .A1(n47242), .A2(n47241), .Z(n47243) );
  XNOR2HSV1 U51031 ( .A1(n47245), .A2(n47244), .ZN(n47247) );
  NAND2HSV0 U51032 ( .A1(n44694), .A2(n52571), .ZN(n47246) );
  XOR2HSV0 U51033 ( .A1(n47247), .A2(n47246), .Z(n47248) );
  XNOR2HSV1 U51034 ( .A1(n47249), .A2(n47248), .ZN(n47251) );
  NAND2HSV0 U51035 ( .A1(n51205), .A2(n48167), .ZN(n47250) );
  XNOR2HSV1 U51036 ( .A1(n47251), .A2(n47250), .ZN(n47252) );
  XNOR2HSV1 U51037 ( .A1(n47253), .A2(n47252), .ZN(n47254) );
  XNOR2HSV1 U51038 ( .A1(n47255), .A2(n47254), .ZN(n47257) );
  NAND2HSV0 U51039 ( .A1(n51211), .A2(n51157), .ZN(n47256) );
  XNOR2HSV1 U51040 ( .A1(n47257), .A2(n47256), .ZN(n47258) );
  XNOR2HSV1 U51041 ( .A1(n47259), .A2(n47258), .ZN(n47262) );
  CLKNAND2HSV0 U51042 ( .A1(n48745), .A2(n51156), .ZN(n47261) );
  NOR2HSV2 U51043 ( .A1(n52659), .A2(n46583), .ZN(n47260) );
  XOR3HSV2 U51044 ( .A1(n47262), .A2(n47261), .A3(n47260), .Z(n47263) );
  XNOR2HSV1 U51045 ( .A1(n47264), .A2(n47263), .ZN(n47266) );
  NAND2HSV0 U51046 ( .A1(n53344), .A2(n45816), .ZN(n47265) );
  NAND2HSV2 U51047 ( .A1(n51155), .A2(\pe5/got [25]), .ZN(n47381) );
  CLKNAND2HSV1 U51048 ( .A1(n52835), .A2(n37654), .ZN(n47379) );
  CLKNAND2HSV1 U51049 ( .A1(n47268), .A2(n47267), .ZN(n47375) );
  CLKNAND2HSV0 U51050 ( .A1(n48165), .A2(n45816), .ZN(n47371) );
  NOR2HSV0 U51051 ( .A1(n51361), .A2(n50422), .ZN(n47366) );
  CLKNAND2HSV0 U51052 ( .A1(n52569), .A2(n51157), .ZN(n47362) );
  NAND2HSV0 U51053 ( .A1(n51158), .A2(n52652), .ZN(n47360) );
  NAND2HSV0 U51054 ( .A1(n52572), .A2(n48167), .ZN(n47356) );
  NAND2HSV0 U51055 ( .A1(n59878), .A2(n50424), .ZN(n47352) );
  NAND2HSV0 U51056 ( .A1(n52574), .A2(n52641), .ZN(n47350) );
  CLKNAND2HSV0 U51057 ( .A1(n52575), .A2(n50698), .ZN(n47348) );
  NAND2HSV0 U51058 ( .A1(n25854), .A2(n51159), .ZN(n47346) );
  NAND2HSV2 U51059 ( .A1(n51162), .A2(n51200), .ZN(n47344) );
  NAND2HSV0 U51060 ( .A1(n52580), .A2(n51334), .ZN(n47342) );
  NAND2HSV0 U51061 ( .A1(n39654), .A2(n51331), .ZN(n47337) );
  NAND2HSV0 U51062 ( .A1(n59936), .A2(n51161), .ZN(n47335) );
  NAND2HSV0 U51063 ( .A1(n48169), .A2(n51362), .ZN(n47333) );
  NAND2HSV0 U51064 ( .A1(n52600), .A2(n30542), .ZN(n47271) );
  NAND2HSV0 U51065 ( .A1(n48681), .A2(n39914), .ZN(n47270) );
  XOR2HSV0 U51066 ( .A1(n47271), .A2(n47270), .Z(n47275) );
  NAND2HSV0 U51067 ( .A1(n39266), .A2(\pe5/bq[1] ), .ZN(n47273) );
  NAND2HSV0 U51068 ( .A1(n51188), .A2(\pe5/bq[7] ), .ZN(n47272) );
  XOR2HSV0 U51069 ( .A1(n47273), .A2(n47272), .Z(n47274) );
  XOR2HSV0 U51070 ( .A1(n47275), .A2(n47274), .Z(n47284) );
  NAND2HSV0 U51071 ( .A1(\pe5/aot [20]), .A2(n48775), .ZN(n47277) );
  NAND2HSV0 U51072 ( .A1(n48199), .A2(n48778), .ZN(n47276) );
  XOR2HSV0 U51073 ( .A1(n47277), .A2(n47276), .Z(n47282) );
  NAND2HSV0 U51074 ( .A1(n47278), .A2(n52632), .ZN(n47280) );
  NAND2HSV0 U51075 ( .A1(n59640), .A2(n50668), .ZN(n47279) );
  XOR2HSV0 U51076 ( .A1(n47280), .A2(n47279), .Z(n47281) );
  XOR2HSV0 U51077 ( .A1(n47282), .A2(n47281), .Z(n47283) );
  XOR2HSV0 U51078 ( .A1(n47284), .A2(n47283), .Z(n47301) );
  NAND2HSV0 U51079 ( .A1(n52611), .A2(n51167), .ZN(n47286) );
  NAND2HSV0 U51080 ( .A1(n37660), .A2(n52630), .ZN(n47285) );
  XOR2HSV0 U51081 ( .A1(n47286), .A2(n47285), .Z(n47290) );
  NAND2HSV0 U51082 ( .A1(n53299), .A2(n52595), .ZN(n47288) );
  NAND2HSV0 U51083 ( .A1(\pe5/aot [13]), .A2(n52610), .ZN(n47287) );
  XOR2HSV0 U51084 ( .A1(n47288), .A2(n47287), .Z(n47289) );
  XOR2HSV0 U51085 ( .A1(n47290), .A2(n47289), .Z(n47299) );
  NAND2HSV0 U51086 ( .A1(\pe5/aot [7]), .A2(n47291), .ZN(n47293) );
  NAND2HSV0 U51087 ( .A1(\pe5/aot [4]), .A2(n52585), .ZN(n47292) );
  XOR2HSV0 U51088 ( .A1(n47293), .A2(n47292), .Z(n47297) );
  NAND2HSV0 U51089 ( .A1(n48761), .A2(n51177), .ZN(n47295) );
  NAND2HSV0 U51090 ( .A1(\pe5/aot [8]), .A2(n46933), .ZN(n47294) );
  XOR2HSV0 U51091 ( .A1(n47295), .A2(n47294), .Z(n47296) );
  XOR2HSV0 U51092 ( .A1(n47297), .A2(n47296), .Z(n47298) );
  XOR2HSV0 U51093 ( .A1(n47299), .A2(n47298), .Z(n47300) );
  XOR2HSV0 U51094 ( .A1(n47301), .A2(n47300), .Z(n47331) );
  NOR2HSV0 U51095 ( .A1(n48246), .A2(n30452), .ZN(n48824) );
  AOI22HSV0 U51096 ( .A1(\pe5/aot [9]), .A2(n48237), .B1(n30341), .B2(n59945), 
        .ZN(n47302) );
  AOI21HSV1 U51097 ( .A1(n47303), .A2(n48824), .B(n47302), .ZN(n47309) );
  CLKNAND2HSV1 U51098 ( .A1(n52682), .A2(n52672), .ZN(n51382) );
  NOR2HSV0 U51099 ( .A1(n47304), .A2(n51382), .ZN(n47307) );
  AOI22HSV0 U51100 ( .A1(\pe5/aot [21]), .A2(n50675), .B1(n47305), .B2(n51310), 
        .ZN(n47306) );
  NOR2HSV1 U51101 ( .A1(n47307), .A2(n47306), .ZN(n47308) );
  XOR2HSV0 U51102 ( .A1(n47309), .A2(n47308), .Z(n47321) );
  NOR2HSV0 U51103 ( .A1(n51232), .A2(n30113), .ZN(n47313) );
  NOR2HSV0 U51104 ( .A1(n45904), .A2(n30116), .ZN(n47312) );
  OAI22HSV2 U51105 ( .A1(n47313), .A2(n47312), .B1(n47311), .B2(n47310), .ZN(
        n47319) );
  NOR2HSV0 U51106 ( .A1(n47315), .A2(n47314), .ZN(n47317) );
  AOI22HSV0 U51107 ( .A1(\pe5/aot [18]), .A2(\pe5/bq[11] ), .B1(n51022), .B2(
        n52619), .ZN(n47316) );
  NOR2HSV2 U51108 ( .A1(n47317), .A2(n47316), .ZN(n47318) );
  XNOR2HSV1 U51109 ( .A1(n47319), .A2(n47318), .ZN(n47320) );
  XNOR2HSV1 U51110 ( .A1(n47321), .A2(n47320), .ZN(n47329) );
  XOR2HSV0 U51111 ( .A1(n47323), .A2(n47322), .Z(n47327) );
  XOR2HSV0 U51112 ( .A1(n47325), .A2(n47324), .Z(n47326) );
  XOR2HSV0 U51113 ( .A1(n47327), .A2(n47326), .Z(n47328) );
  XNOR2HSV1 U51114 ( .A1(n47329), .A2(n47328), .ZN(n47330) );
  XNOR2HSV1 U51115 ( .A1(n47331), .A2(n47330), .ZN(n47332) );
  XNOR2HSV1 U51116 ( .A1(n47333), .A2(n47332), .ZN(n47334) );
  XNOR2HSV1 U51117 ( .A1(n47335), .A2(n47334), .ZN(n47336) );
  XNOR2HSV1 U51118 ( .A1(n47337), .A2(n47336), .ZN(n47340) );
  NAND2HSV0 U51119 ( .A1(n47338), .A2(n52577), .ZN(n47339) );
  XOR2HSV0 U51120 ( .A1(n47340), .A2(n47339), .Z(n47341) );
  XNOR2HSV1 U51121 ( .A1(n47342), .A2(n47341), .ZN(n47343) );
  XNOR2HSV1 U51122 ( .A1(n47344), .A2(n47343), .ZN(n47345) );
  XNOR2HSV1 U51123 ( .A1(n47346), .A2(n47345), .ZN(n47347) );
  XNOR2HSV1 U51124 ( .A1(n47348), .A2(n47347), .ZN(n47349) );
  XNOR2HSV1 U51125 ( .A1(n47350), .A2(n47349), .ZN(n47351) );
  XNOR2HSV1 U51126 ( .A1(n47352), .A2(n47351), .ZN(n47354) );
  NAND2HSV0 U51127 ( .A1(n44694), .A2(n51305), .ZN(n47353) );
  XOR2HSV0 U51128 ( .A1(n47354), .A2(n47353), .Z(n47355) );
  XNOR2HSV1 U51129 ( .A1(n47356), .A2(n47355), .ZN(n47358) );
  NAND2HSV0 U51130 ( .A1(n59517), .A2(n52568), .ZN(n47357) );
  XNOR2HSV1 U51131 ( .A1(n47358), .A2(n47357), .ZN(n47359) );
  XNOR2HSV1 U51132 ( .A1(n47360), .A2(n47359), .ZN(n47361) );
  XNOR2HSV1 U51133 ( .A1(n47362), .A2(n47361), .ZN(n47364) );
  NAND2HSV0 U51134 ( .A1(n51211), .A2(n52658), .ZN(n47363) );
  XNOR2HSV1 U51135 ( .A1(n47364), .A2(n47363), .ZN(n47365) );
  XNOR2HSV1 U51136 ( .A1(n47366), .A2(n47365), .ZN(n47369) );
  CLKNAND2HSV0 U51137 ( .A1(n48745), .A2(n52566), .ZN(n47368) );
  CLKNHSV0 U51138 ( .I(n47394), .ZN(n51218) );
  NOR2HSV1 U51139 ( .A1(n51218), .A2(n30686), .ZN(n47367) );
  XOR3HSV2 U51140 ( .A1(n47369), .A2(n47368), .A3(n47367), .Z(n47370) );
  XNOR2HSV1 U51141 ( .A1(n47371), .A2(n47370), .ZN(n47373) );
  NAND2HSV0 U51142 ( .A1(n53344), .A2(n51228), .ZN(n47372) );
  XNOR2HSV1 U51143 ( .A1(n47373), .A2(n47372), .ZN(n47374) );
  XNOR2HSV1 U51144 ( .A1(n47375), .A2(n47374), .ZN(n47377) );
  CLKNAND2HSV0 U51145 ( .A1(n59535), .A2(n47200), .ZN(n47376) );
  XNOR2HSV1 U51146 ( .A1(n47377), .A2(n47376), .ZN(n47378) );
  XNOR2HSV1 U51147 ( .A1(n47379), .A2(n47378), .ZN(n47380) );
  XNOR2HSV1 U51148 ( .A1(n47381), .A2(n47380), .ZN(n47383) );
  NAND2HSV2 U51149 ( .A1(n29775), .A2(\pe5/got [26]), .ZN(n47382) );
  XNOR2HSV1 U51150 ( .A1(n47386), .A2(n47385), .ZN(\pe5/poht [4]) );
  NOR2HSV4 U51151 ( .A1(n47388), .A2(n47387), .ZN(n47390) );
  NOR2HSV4 U51152 ( .A1(n47390), .A2(n47389), .ZN(n47427) );
  NAND3HSV2 U51153 ( .A1(n47392), .A2(n47391), .A3(n37767), .ZN(n47426) );
  NAND2HSV0 U51154 ( .A1(n29771), .A2(n51362), .ZN(n47393) );
  NAND2HSV0 U51155 ( .A1(n59893), .A2(n51418), .ZN(n47424) );
  INHSV2 U51156 ( .I(n47394), .ZN(n51360) );
  NOR2HSV2 U51157 ( .A1(n51360), .A2(n51231), .ZN(n47422) );
  NAND2HSV0 U51158 ( .A1(n59903), .A2(n59357), .ZN(n47420) );
  NOR2HSV0 U51159 ( .A1(n52567), .A2(n48625), .ZN(n47418) );
  CLKNAND2HSV1 U51160 ( .A1(\pe5/aot [4]), .A2(n51307), .ZN(n47396) );
  NAND2HSV0 U51161 ( .A1(\pe5/aot [3]), .A2(n53216), .ZN(n47395) );
  XOR2HSV0 U51162 ( .A1(n47396), .A2(n47395), .Z(n47400) );
  CLKNAND2HSV1 U51163 ( .A1(n51310), .A2(\pe5/bq[7] ), .ZN(n47398) );
  NAND2HSV0 U51164 ( .A1(n52675), .A2(n52671), .ZN(n47397) );
  XOR2HSV0 U51165 ( .A1(n47398), .A2(n47397), .Z(n47399) );
  XOR2HSV0 U51166 ( .A1(n47400), .A2(n47399), .Z(n47408) );
  NAND2HSV0 U51167 ( .A1(\pe5/aot [9]), .A2(n51336), .ZN(n47402) );
  NAND2HSV0 U51168 ( .A1(n51313), .A2(n51420), .ZN(n47401) );
  XOR2HSV0 U51169 ( .A1(n47402), .A2(n47401), .Z(n47406) );
  CLKNAND2HSV0 U51170 ( .A1(n53323), .A2(\pe5/bq[2] ), .ZN(n47404) );
  NAND2HSV0 U51171 ( .A1(n51247), .A2(n50526), .ZN(n47403) );
  XOR2HSV0 U51172 ( .A1(n47404), .A2(n47403), .Z(n47405) );
  XOR2HSV0 U51173 ( .A1(n47406), .A2(n47405), .Z(n47407) );
  XOR2HSV0 U51174 ( .A1(n47408), .A2(n47407), .Z(n47416) );
  NAND2HSV0 U51175 ( .A1(n59945), .A2(n50675), .ZN(n47411) );
  NAND2HSV0 U51176 ( .A1(n48658), .A2(n53199), .ZN(n47410) );
  XOR2HSV0 U51177 ( .A1(n47411), .A2(n47410), .Z(n47414) );
  CLKNAND2HSV0 U51178 ( .A1(n51339), .A2(n39615), .ZN(n47412) );
  XOR2HSV0 U51179 ( .A1(n51163), .A2(n47412), .Z(n47413) );
  XOR2HSV0 U51180 ( .A1(n47414), .A2(n47413), .Z(n47415) );
  XNOR2HSV1 U51181 ( .A1(n47416), .A2(n47415), .ZN(n47417) );
  XOR2HSV0 U51182 ( .A1(n47418), .A2(n47417), .Z(n47419) );
  XNOR2HSV1 U51183 ( .A1(n47420), .A2(n47419), .ZN(n47421) );
  XNOR2HSV1 U51184 ( .A1(n47422), .A2(n47421), .ZN(n47423) );
  XNOR2HSV1 U51185 ( .A1(n47424), .A2(n47423), .ZN(n47425) );
  INAND2HSV2 U51186 ( .A1(n60001), .B1(n47429), .ZN(n56418) );
  NAND2HSV0 U51187 ( .A1(n47429), .A2(n47428), .ZN(n56417) );
  INHSV1 U51188 ( .I(n45727), .ZN(n56174) );
  INHSV2 U51189 ( .I(n50718), .ZN(n56621) );
  CLKNAND2HSV0 U51190 ( .A1(n56621), .A2(\pe3/got [14]), .ZN(n47495) );
  CLKNHSV0 U51191 ( .I(n53227), .ZN(n56783) );
  CLKNAND2HSV0 U51192 ( .A1(n56783), .A2(n56421), .ZN(n47493) );
  CLKNAND2HSV1 U51193 ( .A1(n56561), .A2(n56176), .ZN(n47491) );
  CLKNAND2HSV0 U51194 ( .A1(n55613), .A2(n56247), .ZN(n47489) );
  INHSV2 U51195 ( .I(n50756), .ZN(n56619) );
  CLKNAND2HSV0 U51196 ( .A1(n56562), .A2(n56619), .ZN(n47487) );
  CLKNAND2HSV1 U51197 ( .A1(n56178), .A2(n56241), .ZN(n47480) );
  INAND2HSV0 U51198 ( .A1(n47431), .B1(n59620), .ZN(n47472) );
  NAND2HSV0 U51199 ( .A1(n42940), .A2(\pe3/bq[11] ), .ZN(n48523) );
  CLKNAND2HSV1 U51200 ( .A1(n56197), .A2(n56824), .ZN(n56747) );
  NOR2HSV0 U51201 ( .A1(n48523), .A2(n56747), .ZN(n47433) );
  AOI22HSV0 U51202 ( .A1(n56182), .A2(n56971), .B1(n59623), .B2(\pe3/bq[11] ), 
        .ZN(n47432) );
  NOR2HSV2 U51203 ( .A1(n47433), .A2(n47432), .ZN(n47435) );
  XOR2HSV0 U51204 ( .A1(n47435), .A2(n47434), .Z(n47438) );
  NOR2HSV0 U51205 ( .A1(n49265), .A2(n49258), .ZN(n56274) );
  NAND2HSV0 U51206 ( .A1(n56204), .A2(n56348), .ZN(n47436) );
  XOR2HSV0 U51207 ( .A1(n56274), .A2(n47436), .Z(n47437) );
  XNOR2HSV1 U51208 ( .A1(n47438), .A2(n47437), .ZN(n47470) );
  NAND2HSV0 U51209 ( .A1(n56370), .A2(n56187), .ZN(n47440) );
  NAND2HSV0 U51210 ( .A1(n56188), .A2(n56827), .ZN(n47439) );
  XOR2HSV0 U51211 ( .A1(n47440), .A2(n47439), .Z(n47444) );
  NAND2HSV0 U51212 ( .A1(\pe3/aot [8]), .A2(n48499), .ZN(n47442) );
  NAND2HSV0 U51213 ( .A1(n56373), .A2(n45534), .ZN(n47441) );
  XOR2HSV0 U51214 ( .A1(n47442), .A2(n47441), .Z(n47443) );
  XOR2HSV0 U51215 ( .A1(n47444), .A2(n47443), .Z(n47453) );
  NOR2HSV0 U51216 ( .A1(n56382), .A2(n56277), .ZN(n47446) );
  NAND2HSV0 U51217 ( .A1(n56221), .A2(n56094), .ZN(n47445) );
  XOR2HSV0 U51218 ( .A1(n47446), .A2(n47445), .Z(n47451) );
  NOR2HSV0 U51219 ( .A1(n42835), .A2(n50722), .ZN(n56351) );
  NOR2HSV0 U51220 ( .A1(n47447), .A2(n48545), .ZN(n47449) );
  NAND2HSV2 U51221 ( .A1(\pe3/aot [10]), .A2(\pe3/bq[3] ), .ZN(n56703) );
  OAI22HSV0 U51222 ( .A1(n56351), .A2(n47449), .B1(n47448), .B2(n56703), .ZN(
        n47450) );
  XNOR2HSV1 U51223 ( .A1(n47451), .A2(n47450), .ZN(n47452) );
  XNOR2HSV1 U51224 ( .A1(n47453), .A2(n47452), .ZN(n47469) );
  NAND2HSV0 U51225 ( .A1(n55864), .A2(n56832), .ZN(n47455) );
  NAND2HSV0 U51226 ( .A1(n59344), .A2(n56189), .ZN(n47454) );
  XOR2HSV0 U51227 ( .A1(n47455), .A2(n47454), .Z(n47459) );
  BUFHSV2 U51228 ( .I(\pe3/aot [6]), .Z(n55967) );
  CLKNAND2HSV0 U51229 ( .A1(n55967), .A2(n56640), .ZN(n47457) );
  NAND2HSV0 U51230 ( .A1(n59961), .A2(n42971), .ZN(n47456) );
  XOR2HSV0 U51231 ( .A1(n47457), .A2(n47456), .Z(n47458) );
  XOR2HSV0 U51232 ( .A1(n47459), .A2(n47458), .Z(n47467) );
  CLKNAND2HSV1 U51233 ( .A1(\pe3/aot [18]), .A2(\pe3/bq[4] ), .ZN(n47461) );
  BUFHSV2 U51234 ( .I(\pe3/aot [4]), .Z(n56074) );
  NAND2HSV0 U51235 ( .A1(n56074), .A2(n55727), .ZN(n47460) );
  XOR2HSV0 U51236 ( .A1(n47461), .A2(n47460), .Z(n47465) );
  NOR2HSV0 U51237 ( .A1(n45662), .A2(n55755), .ZN(n47463) );
  CLKNAND2HSV0 U51238 ( .A1(\pe3/aot [3]), .A2(\pe3/bq[19] ), .ZN(n47462) );
  XOR2HSV0 U51239 ( .A1(n47463), .A2(n47462), .Z(n47464) );
  XOR2HSV0 U51240 ( .A1(n47465), .A2(n47464), .Z(n47466) );
  XOR2HSV0 U51241 ( .A1(n47467), .A2(n47466), .Z(n47468) );
  XOR3HSV2 U51242 ( .A1(n47470), .A2(n47469), .A3(n47468), .Z(n47471) );
  XNOR2HSV1 U51243 ( .A1(n47472), .A2(n47471), .ZN(n47475) );
  NOR2HSV0 U51244 ( .A1(n56391), .A2(n56936), .ZN(n47474) );
  CLKNHSV0 U51245 ( .I(n56906), .ZN(n56069) );
  NAND2HSV0 U51246 ( .A1(n49468), .A2(n56069), .ZN(n47473) );
  XOR3HSV1 U51247 ( .A1(n47475), .A2(n47474), .A3(n47473), .Z(n47478) );
  NOR2HSV1 U51248 ( .A1(n56475), .A2(n56904), .ZN(n47477) );
  BUFHSV2 U51249 ( .I(n59810), .Z(n56242) );
  CLKNAND2HSV0 U51250 ( .A1(n56242), .A2(n56267), .ZN(n47476) );
  XOR3HSV2 U51251 ( .A1(n47478), .A2(n47477), .A3(n47476), .Z(n47479) );
  XNOR2HSV1 U51252 ( .A1(n47480), .A2(n47479), .ZN(n47482) );
  INHSV2 U51253 ( .I(n56821), .ZN(n56683) );
  NAND2HSV0 U51254 ( .A1(n43850), .A2(n56683), .ZN(n47481) );
  XNOR2HSV1 U51255 ( .A1(n47482), .A2(n47481), .ZN(n47485) );
  CLKNAND2HSV1 U51256 ( .A1(n56624), .A2(\pe3/got [8]), .ZN(n47484) );
  NAND2HSV0 U51257 ( .A1(n56662), .A2(n56177), .ZN(n47483) );
  XOR3HSV2 U51258 ( .A1(n47485), .A2(n47484), .A3(n47483), .Z(n47486) );
  XNOR2HSV1 U51259 ( .A1(n47487), .A2(n47486), .ZN(n47488) );
  XOR2HSV0 U51260 ( .A1(n47489), .A2(n47488), .Z(n47490) );
  XNOR2HSV1 U51261 ( .A1(n47491), .A2(n47490), .ZN(n47492) );
  XNOR2HSV1 U51262 ( .A1(n47493), .A2(n47492), .ZN(n47494) );
  INHSV2 U51263 ( .I(n47496), .ZN(n56172) );
  INHSV2 U51264 ( .I(n47497), .ZN(n52902) );
  CLKNAND2HSV1 U51265 ( .A1(n52902), .A2(n45289), .ZN(n47562) );
  INHSV2 U51266 ( .I(n47498), .ZN(n51958) );
  CLKNAND2HSV1 U51267 ( .A1(n25831), .A2(n51958), .ZN(n47561) );
  CLKNAND2HSV1 U51268 ( .A1(n25835), .A2(n59375), .ZN(n47559) );
  CLKNAND2HSV1 U51269 ( .A1(n51893), .A2(n49493), .ZN(n47553) );
  NOR2HSV1 U51270 ( .A1(n52170), .A2(n44045), .ZN(n47551) );
  NAND2HSV0 U51271 ( .A1(n59522), .A2(n52052), .ZN(n47549) );
  BUFHSV2 U51272 ( .I(n47500), .Z(n52171) );
  NOR2HSV1 U51273 ( .A1(n47500), .A2(n50928), .ZN(n47547) );
  CLKNAND2HSV1 U51274 ( .A1(n51485), .A2(n59777), .ZN(n47544) );
  INHSV1 U51275 ( .I(n53032), .ZN(n51933) );
  NAND2HSV0 U51276 ( .A1(n51933), .A2(n59506), .ZN(n47538) );
  NOR2HSV1 U51277 ( .A1(n53065), .A2(n50926), .ZN(n47536) );
  NAND2HSV0 U51278 ( .A1(n59773), .A2(n52896), .ZN(n47534) );
  NAND2HSV0 U51279 ( .A1(n52867), .A2(n49619), .ZN(n47502) );
  NAND2HSV0 U51280 ( .A1(\pe2/aot [2]), .A2(n52984), .ZN(n47501) );
  XOR2HSV0 U51281 ( .A1(n47502), .A2(n47501), .Z(n47507) );
  CLKNAND2HSV0 U51282 ( .A1(\pe2/aot [15]), .A2(n52905), .ZN(n47505) );
  NAND2HSV0 U51283 ( .A1(n51759), .A2(n52851), .ZN(n47504) );
  XOR2HSV0 U51284 ( .A1(n47505), .A2(n47504), .Z(n47506) );
  XOR2HSV0 U51285 ( .A1(n47507), .A2(n47506), .Z(n47517) );
  NAND2HSV0 U51286 ( .A1(n59633), .A2(n51900), .ZN(n47510) );
  NAND2HSV0 U51287 ( .A1(n51920), .A2(n51803), .ZN(n47509) );
  XOR2HSV0 U51288 ( .A1(n47510), .A2(n47509), .Z(n47515) );
  NAND2HSV0 U51289 ( .A1(\pe2/aot [9]), .A2(n51623), .ZN(n47513) );
  NAND2HSV0 U51290 ( .A1(n51921), .A2(n51897), .ZN(n47512) );
  XOR2HSV0 U51291 ( .A1(n47513), .A2(n47512), .Z(n47514) );
  XOR2HSV0 U51292 ( .A1(n47515), .A2(n47514), .Z(n47516) );
  XOR2HSV0 U51293 ( .A1(n47517), .A2(n47516), .Z(n47532) );
  CLKNHSV0 U51294 ( .I(n49628), .ZN(n51729) );
  NAND2HSV0 U51295 ( .A1(n52951), .A2(n51729), .ZN(n51611) );
  NAND2HSV0 U51296 ( .A1(n52063), .A2(n29736), .ZN(n51563) );
  NOR2HSV0 U51297 ( .A1(n51611), .A2(n51563), .ZN(n47520) );
  AOI22HSV0 U51298 ( .A1(n52951), .A2(n52448), .B1(n51839), .B2(n29736), .ZN(
        n47519) );
  NOR2HSV2 U51299 ( .A1(n47520), .A2(n47519), .ZN(n47521) );
  NAND2HSV0 U51300 ( .A1(n51636), .A2(\pe2/bq[12] ), .ZN(n51808) );
  XOR2HSV0 U51301 ( .A1(n47521), .A2(n51808), .Z(n47523) );
  NAND2HSV0 U51302 ( .A1(n53005), .A2(\pe2/bq[6] ), .ZN(n51621) );
  NAND2HSV0 U51303 ( .A1(n51743), .A2(n51919), .ZN(n51804) );
  XOR2HSV0 U51304 ( .A1(n51621), .A2(n51804), .Z(n47522) );
  XOR2HSV0 U51305 ( .A1(n47523), .A2(n47522), .Z(n47530) );
  NAND2HSV0 U51306 ( .A1(n51547), .A2(\pe2/bq[17] ), .ZN(n52201) );
  CLKNAND2HSV1 U51307 ( .A1(n51824), .A2(\pe2/bq[14] ), .ZN(n49629) );
  XOR2HSV0 U51308 ( .A1(n52201), .A2(n49629), .Z(n47528) );
  NAND2HSV0 U51309 ( .A1(n51460), .A2(n51825), .ZN(n47526) );
  NAND2HSV0 U51310 ( .A1(n59976), .A2(n51832), .ZN(n47525) );
  XOR2HSV0 U51311 ( .A1(n47526), .A2(n47525), .Z(n47527) );
  XNOR2HSV1 U51312 ( .A1(n47528), .A2(n47527), .ZN(n47529) );
  XNOR2HSV1 U51313 ( .A1(n47530), .A2(n47529), .ZN(n47531) );
  XOR2HSV0 U51314 ( .A1(n47532), .A2(n47531), .Z(n47533) );
  XNOR2HSV1 U51315 ( .A1(n47534), .A2(n47533), .ZN(n47535) );
  XNOR2HSV1 U51316 ( .A1(n47536), .A2(n47535), .ZN(n47537) );
  XNOR2HSV1 U51317 ( .A1(n47538), .A2(n47537), .ZN(n47542) );
  BUFHSV2 U51318 ( .I(n52532), .Z(n51861) );
  NAND2HSV2 U51319 ( .A1(n51861), .A2(n51896), .ZN(n47541) );
  CLKNHSV0 U51320 ( .I(n29746), .ZN(n51862) );
  CLKNAND2HSV1 U51321 ( .A1(n51862), .A2(n59778), .ZN(n47540) );
  XOR3HSV2 U51322 ( .A1(n47542), .A2(n47541), .A3(n47540), .Z(n47543) );
  XNOR2HSV1 U51323 ( .A1(n47544), .A2(n47543), .ZN(n47546) );
  BUFHSV2 U51324 ( .I(n59774), .Z(n51868) );
  CLKNAND2HSV1 U51325 ( .A1(n51868), .A2(\pe2/got [8]), .ZN(n47545) );
  XOR3HSV2 U51326 ( .A1(n47547), .A2(n47546), .A3(n47545), .Z(n47548) );
  XOR2HSV0 U51327 ( .A1(n47549), .A2(n47548), .Z(n47550) );
  XNOR2HSV1 U51328 ( .A1(n47551), .A2(n47550), .ZN(n47552) );
  XNOR2HSV1 U51329 ( .A1(n47553), .A2(n47552), .ZN(n47557) );
  INHSV2 U51330 ( .I(n47939), .ZN(n51878) );
  CLKNAND2HSV1 U51331 ( .A1(n51878), .A2(\pe2/got [12]), .ZN(n47556) );
  XNOR2HSV1 U51332 ( .A1(n47557), .A2(n47556), .ZN(n47558) );
  XOR2HSV0 U51333 ( .A1(n47559), .A2(n47558), .Z(n47560) );
  CLKNAND2HSV1 U51334 ( .A1(n47563), .A2(n47564), .ZN(n47566) );
  CLKNAND2HSV2 U51335 ( .A1(n47566), .A2(n47565), .ZN(n47569) );
  XNOR2HSV1 U51336 ( .A1(n47569), .A2(n47568), .ZN(\pe2/poht [15]) );
  INHSV2 U51337 ( .I(n47570), .ZN(n51889) );
  INHSV2 U51338 ( .I(n49606), .ZN(n51728) );
  CLKNAND2HSV1 U51339 ( .A1(n51728), .A2(n47571), .ZN(n47647) );
  CLKNHSV0 U51340 ( .I(n47572), .ZN(n52049) );
  NOR2HSV1 U51341 ( .A1(n52049), .A2(n52526), .ZN(n47645) );
  BUFHSV2 U51342 ( .I(n52920), .Z(n51799) );
  INHSV2 U51343 ( .I(n47573), .ZN(n52051) );
  CLKNAND2HSV0 U51344 ( .A1(n51799), .A2(n52051), .ZN(n47643) );
  NOR2HSV1 U51345 ( .A1(n52171), .A2(n51607), .ZN(n47641) );
  NAND2HSV0 U51346 ( .A1(n44714), .A2(n52814), .ZN(n47633) );
  NAND2HSV0 U51347 ( .A1(n52926), .A2(n52125), .ZN(n47631) );
  CLKNAND2HSV0 U51348 ( .A1(n52927), .A2(n51939), .ZN(n47628) );
  CLKNHSV0 U51349 ( .I(n52773), .ZN(n51609) );
  NAND2HSV0 U51350 ( .A1(n51609), .A2(n52175), .ZN(n47626) );
  NAND2HSV0 U51351 ( .A1(n51933), .A2(n51966), .ZN(n47624) );
  NAND2HSV0 U51352 ( .A1(n50929), .A2(n51932), .ZN(n47621) );
  NAND2HSV0 U51353 ( .A1(n44120), .A2(n59767), .ZN(n47619) );
  NAND2HSV2 U51354 ( .A1(n50930), .A2(\pe2/bq[3] ), .ZN(n52223) );
  CLKNHSV0 U51355 ( .I(n52223), .ZN(n47577) );
  NOR2HSV0 U51356 ( .A1(n47575), .A2(n50920), .ZN(n52204) );
  AOI22HSV0 U51357 ( .A1(n50930), .A2(n51614), .B1(n52104), .B2(n52484), .ZN(
        n47576) );
  AOI21HSV2 U51358 ( .A1(n47577), .A2(n52204), .B(n47576), .ZN(n47585) );
  NAND2HSV0 U51359 ( .A1(n59973), .A2(n53223), .ZN(n47579) );
  NAND2HSV0 U51360 ( .A1(\pe2/aot [12]), .A2(n51733), .ZN(n47578) );
  XOR2HSV0 U51361 ( .A1(n47579), .A2(n47578), .Z(n47584) );
  NOR2HSV0 U51362 ( .A1(n52200), .A2(n47580), .ZN(n48106) );
  NOR2HSV0 U51363 ( .A1(n52431), .A2(n48066), .ZN(n50971) );
  AOI22HSV0 U51364 ( .A1(n53019), .A2(n49619), .B1(\pe2/bq[14] ), .B2(n51460), 
        .ZN(n47581) );
  AOI21HSV1 U51365 ( .A1(n48106), .A2(n50971), .B(n47581), .ZN(n47582) );
  NAND2HSV0 U51366 ( .A1(n59974), .A2(n52481), .ZN(n51622) );
  XNOR2HSV1 U51367 ( .A1(n47582), .A2(n51622), .ZN(n47583) );
  XOR3HSV2 U51368 ( .A1(n47585), .A2(n47584), .A3(n47583), .Z(n47617) );
  NAND2HSV0 U51369 ( .A1(\pe2/aot [2]), .A2(n52299), .ZN(n47587) );
  NAND2HSV0 U51370 ( .A1(n51759), .A2(n51457), .ZN(n47586) );
  XOR2HSV0 U51371 ( .A1(n47587), .A2(n47586), .Z(n47591) );
  NAND2HSV0 U51372 ( .A1(\pe2/aot [7]), .A2(\pe2/bq[17] ), .ZN(n47589) );
  NAND2HSV0 U51373 ( .A1(n59783), .A2(n52179), .ZN(n47588) );
  XOR2HSV0 U51374 ( .A1(n47589), .A2(n47588), .Z(n47590) );
  XOR2HSV0 U51375 ( .A1(n47591), .A2(n47590), .Z(n47597) );
  NAND2HSV0 U51376 ( .A1(n51920), .A2(n52063), .ZN(n50952) );
  NAND2HSV0 U51377 ( .A1(\pe2/aot [19]), .A2(n52857), .ZN(n52081) );
  XOR2HSV0 U51378 ( .A1(n50952), .A2(n52081), .Z(n47595) );
  NAND2HSV0 U51379 ( .A1(\pe2/aot [20]), .A2(\pe2/bq[4] ), .ZN(n47593) );
  NAND2HSV0 U51380 ( .A1(n52955), .A2(\pe2/bq[6] ), .ZN(n47592) );
  XOR2HSV0 U51381 ( .A1(n47593), .A2(n47592), .Z(n47594) );
  XOR2HSV0 U51382 ( .A1(n47595), .A2(n47594), .Z(n47596) );
  XOR2HSV0 U51383 ( .A1(n47597), .A2(n47596), .Z(n47616) );
  NAND2HSV0 U51384 ( .A1(\pe2/aot [11]), .A2(n47598), .ZN(n47601) );
  INHSV2 U51385 ( .I(n51537), .ZN(n52858) );
  NAND2HSV0 U51386 ( .A1(n52858), .A2(n44197), .ZN(n47600) );
  XOR2HSV0 U51387 ( .A1(n47601), .A2(n47600), .Z(n47605) );
  NAND2HSV0 U51388 ( .A1(\pe2/aot [6]), .A2(n52988), .ZN(n47603) );
  NAND2HSV0 U51389 ( .A1(n37801), .A2(n51805), .ZN(n47602) );
  XOR2HSV0 U51390 ( .A1(n47603), .A2(n47602), .Z(n47604) );
  XOR2HSV0 U51391 ( .A1(n47605), .A2(n47604), .Z(n47614) );
  NAND2HSV0 U51392 ( .A1(n59975), .A2(n52073), .ZN(n47607) );
  NAND2HSV0 U51393 ( .A1(n52056), .A2(n43961), .ZN(n47606) );
  XOR2HSV0 U51394 ( .A1(n47607), .A2(n47606), .Z(n47612) );
  NAND2HSV0 U51395 ( .A1(n52951), .A2(\pe2/bq[16] ), .ZN(n47610) );
  NAND2HSV0 U51396 ( .A1(n52344), .A2(\pe2/bq[21] ), .ZN(n47609) );
  XOR2HSV0 U51397 ( .A1(n47610), .A2(n47609), .Z(n47611) );
  XOR2HSV0 U51398 ( .A1(n47612), .A2(n47611), .Z(n47613) );
  XOR2HSV0 U51399 ( .A1(n47614), .A2(n47613), .Z(n47615) );
  XOR3HSV2 U51400 ( .A1(n47617), .A2(n47616), .A3(n47615), .Z(n47618) );
  XNOR2HSV1 U51401 ( .A1(n47619), .A2(n47618), .ZN(n47620) );
  XNOR2HSV1 U51402 ( .A1(n47621), .A2(n47620), .ZN(n47623) );
  NAND2HSV0 U51403 ( .A1(n51610), .A2(n51896), .ZN(n47622) );
  XOR3HSV2 U51404 ( .A1(n47624), .A2(n47623), .A3(n47622), .Z(n47625) );
  XNOR2HSV1 U51405 ( .A1(n47626), .A2(n47625), .ZN(n47627) );
  XNOR2HSV1 U51406 ( .A1(n47628), .A2(n47627), .ZN(n47630) );
  NOR2HSV0 U51407 ( .A1(n53065), .A2(n44188), .ZN(n47629) );
  XOR3HSV2 U51408 ( .A1(n47631), .A2(n47630), .A3(n47629), .Z(n47632) );
  XOR2HSV0 U51409 ( .A1(n47633), .A2(n47632), .Z(n47636) );
  NAND2HSV0 U51410 ( .A1(n59769), .A2(\pe2/got [10]), .ZN(n47635) );
  CLKNHSV0 U51411 ( .I(n49656), .ZN(n52930) );
  CLKNAND2HSV0 U51412 ( .A1(n51862), .A2(n52930), .ZN(n47634) );
  XOR3HSV2 U51413 ( .A1(n47636), .A2(n47635), .A3(n47634), .Z(n47637) );
  XNOR2HSV1 U51414 ( .A1(n47638), .A2(n47637), .ZN(n47640) );
  BUFHSV2 U51415 ( .I(n59774), .Z(n51782) );
  CLKNAND2HSV0 U51416 ( .A1(n51782), .A2(n51958), .ZN(n47639) );
  XOR3HSV2 U51417 ( .A1(n47641), .A2(n47640), .A3(n47639), .Z(n47642) );
  XOR2HSV0 U51418 ( .A1(n47643), .A2(n47642), .Z(n47644) );
  XNOR2HSV1 U51419 ( .A1(n47645), .A2(n47644), .ZN(n47646) );
  CLKNAND2HSV0 U51420 ( .A1(n52399), .A2(n52050), .ZN(n47649) );
  CLKNAND2HSV1 U51421 ( .A1(n58219), .A2(n58299), .ZN(n47654) );
  CLKNAND2HSV0 U51422 ( .A1(\pe4/aot [1]), .A2(n58196), .ZN(n47651) );
  CLKNAND2HSV0 U51423 ( .A1(\pe4/aot [2]), .A2(\pe4/bq[2] ), .ZN(n47650) );
  XOR2HSV0 U51424 ( .A1(n47651), .A2(n47650), .Z(n47652) );
  NOR2HSV2 U51425 ( .A1(n58194), .A2(n58013), .ZN(n57344) );
  XNOR2HSV1 U51426 ( .A1(n47652), .A2(n57344), .ZN(n47653) );
  XOR2HSV0 U51427 ( .A1(n47654), .A2(n47653), .Z(n47792) );
  NAND2HSV0 U51428 ( .A1(n59601), .A2(n50065), .ZN(n47766) );
  NAND2HSV2 U51429 ( .A1(n57984), .A2(\pe4/got [18]), .ZN(n47759) );
  CLKNAND2HSV1 U51430 ( .A1(n49966), .A2(n47656), .ZN(n47755) );
  NAND2HSV0 U51431 ( .A1(n57324), .A2(n57424), .ZN(n47753) );
  CLKNAND2HSV0 U51432 ( .A1(n59833), .A2(n47657), .ZN(n47750) );
  NAND2HSV0 U51433 ( .A1(n34352), .A2(n58153), .ZN(n47746) );
  NAND2HSV0 U51434 ( .A1(n59667), .A2(n57177), .ZN(n47739) );
  NAND2HSV0 U51435 ( .A1(\pe4/aot [20]), .A2(n57139), .ZN(n57217) );
  NAND2HSV0 U51436 ( .A1(n47658), .A2(n58130), .ZN(n57123) );
  XOR2HSV0 U51437 ( .A1(n57217), .A2(n57123), .Z(n47674) );
  NAND2HSV0 U51438 ( .A1(n47659), .A2(\pe4/pvq [31]), .ZN(n47660) );
  XOR2HSV0 U51439 ( .A1(n47660), .A2(\pe4/phq [31]), .Z(n47665) );
  NAND2HSV0 U51440 ( .A1(n57210), .A2(n58010), .ZN(n57114) );
  NAND2HSV0 U51441 ( .A1(n57837), .A2(n57138), .ZN(n57222) );
  OAI21HSV0 U51442 ( .A1(n50351), .A2(n47661), .B(n57222), .ZN(n47662) );
  OAI21HSV0 U51443 ( .A1(n47663), .A2(n57114), .B(n47662), .ZN(n47664) );
  XNOR2HSV1 U51444 ( .A1(n47665), .A2(n47664), .ZN(n47673) );
  NAND2HSV0 U51445 ( .A1(n33867), .A2(\pe4/bq[16] ), .ZN(n47667) );
  NAND2HSV0 U51446 ( .A1(n57014), .A2(n57926), .ZN(n47666) );
  XOR2HSV0 U51447 ( .A1(n47667), .A2(n47666), .Z(n47671) );
  NAND2HSV0 U51448 ( .A1(n57510), .A2(n57684), .ZN(n47668) );
  XOR2HSV0 U51449 ( .A1(n47669), .A2(n47668), .Z(n47670) );
  XOR2HSV0 U51450 ( .A1(n47671), .A2(n47670), .Z(n47672) );
  XOR3HSV2 U51451 ( .A1(n47674), .A2(n47673), .A3(n47672), .Z(n47676) );
  CLKNHSV0 U51452 ( .I(n50091), .ZN(n57744) );
  NAND2HSV0 U51453 ( .A1(n57251), .A2(n57744), .ZN(n47675) );
  XOR2HSV0 U51454 ( .A1(n47676), .A2(n47675), .Z(n47732) );
  NAND2HSV0 U51455 ( .A1(n59501), .A2(n57677), .ZN(n47731) );
  NAND2HSV0 U51456 ( .A1(\pe4/aot [11]), .A2(\pe4/bq[23] ), .ZN(n47678) );
  NAND2HSV0 U51457 ( .A1(n57463), .A2(n34254), .ZN(n47677) );
  XOR2HSV0 U51458 ( .A1(n47678), .A2(n47677), .Z(n47683) );
  NAND2HSV0 U51459 ( .A1(n58198), .A2(n33427), .ZN(n47681) );
  NAND2HSV0 U51460 ( .A1(n59346), .A2(n47679), .ZN(n47680) );
  XOR2HSV0 U51461 ( .A1(n47681), .A2(n47680), .Z(n47682) );
  XOR2HSV0 U51462 ( .A1(n47683), .A2(n47682), .Z(n47691) );
  NAND2HSV0 U51463 ( .A1(n57504), .A2(n57691), .ZN(n47685) );
  NAND2HSV0 U51464 ( .A1(n33965), .A2(n58077), .ZN(n47684) );
  XOR2HSV0 U51465 ( .A1(n47685), .A2(n47684), .Z(n47689) );
  NAND2HSV0 U51466 ( .A1(n59523), .A2(n58196), .ZN(n47687) );
  NAND2HSV0 U51467 ( .A1(n57727), .A2(n58116), .ZN(n47686) );
  XOR2HSV0 U51468 ( .A1(n47687), .A2(n47686), .Z(n47688) );
  XOR2HSV0 U51469 ( .A1(n47689), .A2(n47688), .Z(n47690) );
  XOR2HSV0 U51470 ( .A1(n47691), .A2(n47690), .Z(n47708) );
  NAND2HSV0 U51471 ( .A1(n59953), .A2(n57929), .ZN(n47694) );
  NAND2HSV0 U51472 ( .A1(n47692), .A2(\pe4/bq[2] ), .ZN(n47693) );
  XOR2HSV0 U51473 ( .A1(n47694), .A2(n47693), .Z(n47698) );
  NAND2HSV0 U51474 ( .A1(n57460), .A2(n59668), .ZN(n47696) );
  NAND2HSV0 U51475 ( .A1(n33716), .A2(\pe4/bq[11] ), .ZN(n47695) );
  XOR2HSV0 U51476 ( .A1(n47696), .A2(n47695), .Z(n47697) );
  XOR2HSV0 U51477 ( .A1(n47698), .A2(n47697), .Z(n47706) );
  NOR2HSV0 U51478 ( .A1(n50008), .A2(n53219), .ZN(n47700) );
  NAND2HSV0 U51479 ( .A1(n57230), .A2(n34021), .ZN(n47699) );
  XOR2HSV0 U51480 ( .A1(n47700), .A2(n47699), .Z(n47704) );
  NAND2HSV0 U51481 ( .A1(\pe4/aot [2]), .A2(n57098), .ZN(n47702) );
  NAND2HSV0 U51482 ( .A1(n59954), .A2(\pe4/bq[31] ), .ZN(n47701) );
  XOR2HSV0 U51483 ( .A1(n47702), .A2(n47701), .Z(n47703) );
  XOR2HSV0 U51484 ( .A1(n47704), .A2(n47703), .Z(n47705) );
  XOR2HSV0 U51485 ( .A1(n47706), .A2(n47705), .Z(n47707) );
  XOR2HSV0 U51486 ( .A1(n47708), .A2(n47707), .Z(n47729) );
  NAND2HSV0 U51487 ( .A1(n59343), .A2(n33711), .ZN(n47711) );
  NAND2HSV0 U51488 ( .A1(n47709), .A2(n57595), .ZN(n47710) );
  XOR2HSV0 U51489 ( .A1(n47711), .A2(n47710), .Z(n47715) );
  NAND2HSV0 U51490 ( .A1(n59831), .A2(n33533), .ZN(n47713) );
  NAND2HSV0 U51491 ( .A1(n57338), .A2(n35194), .ZN(n47712) );
  XOR2HSV0 U51492 ( .A1(n47713), .A2(n47712), .Z(n47714) );
  XOR2HSV0 U51493 ( .A1(n47715), .A2(n47714), .Z(n47724) );
  NAND2HSV0 U51494 ( .A1(\pe4/aot [25]), .A2(n57135), .ZN(n47717) );
  NAND2HSV0 U51495 ( .A1(n57140), .A2(n58084), .ZN(n47716) );
  XOR2HSV0 U51496 ( .A1(n47717), .A2(n47716), .Z(n47722) );
  NAND2HSV0 U51497 ( .A1(n57234), .A2(n57089), .ZN(n47720) );
  NAND2HSV0 U51498 ( .A1(n47718), .A2(\pe4/bq[24] ), .ZN(n47719) );
  XOR2HSV0 U51499 ( .A1(n47720), .A2(n47719), .Z(n47721) );
  XOR2HSV0 U51500 ( .A1(n47722), .A2(n47721), .Z(n47723) );
  XOR2HSV0 U51501 ( .A1(n47724), .A2(n47723), .Z(n47727) );
  CLKNHSV0 U51502 ( .I(n47725), .ZN(n57584) );
  NAND2HSV0 U51503 ( .A1(n34127), .A2(n57584), .ZN(n47726) );
  XNOR2HSV1 U51504 ( .A1(n47727), .A2(n47726), .ZN(n47728) );
  XNOR2HSV1 U51505 ( .A1(n47729), .A2(n47728), .ZN(n47730) );
  XOR3HSV2 U51506 ( .A1(n47732), .A2(n47731), .A3(n47730), .Z(n47735) );
  NAND2HSV0 U51507 ( .A1(n47733), .A2(n58184), .ZN(n47734) );
  XOR2HSV0 U51508 ( .A1(n47735), .A2(n47734), .Z(n47737) );
  NAND2HSV0 U51509 ( .A1(n59662), .A2(n58036), .ZN(n47736) );
  XNOR2HSV1 U51510 ( .A1(n47737), .A2(n47736), .ZN(n47738) );
  XNOR2HSV1 U51511 ( .A1(n47739), .A2(n47738), .ZN(n47741) );
  CLKNAND2HSV0 U51512 ( .A1(n57405), .A2(n57180), .ZN(n47740) );
  XNOR2HSV1 U51513 ( .A1(n47741), .A2(n47740), .ZN(n47744) );
  NAND2HSV0 U51514 ( .A1(n47742), .A2(n59663), .ZN(n47743) );
  XOR2HSV0 U51515 ( .A1(n47744), .A2(n47743), .Z(n47745) );
  XNOR2HSV1 U51516 ( .A1(n47746), .A2(n47745), .ZN(n47748) );
  CLKNAND2HSV0 U51517 ( .A1(n57183), .A2(n58110), .ZN(n47747) );
  XNOR2HSV1 U51518 ( .A1(n47748), .A2(n47747), .ZN(n47749) );
  XNOR2HSV1 U51519 ( .A1(n47750), .A2(n47749), .ZN(n47752) );
  CLKNAND2HSV1 U51520 ( .A1(n25243), .A2(n57982), .ZN(n47751) );
  XOR3HSV2 U51521 ( .A1(n47753), .A2(n47752), .A3(n47751), .Z(n47754) );
  XNOR2HSV1 U51522 ( .A1(n47755), .A2(n47754), .ZN(n47757) );
  CLKNAND2HSV0 U51523 ( .A1(n57547), .A2(n57753), .ZN(n47756) );
  XNOR2HSV1 U51524 ( .A1(n47757), .A2(n47756), .ZN(n47758) );
  XNOR2HSV1 U51525 ( .A1(n47759), .A2(n47758), .ZN(n47761) );
  CLKNAND2HSV1 U51526 ( .A1(n49951), .A2(n57770), .ZN(n47760) );
  XNOR2HSV1 U51527 ( .A1(n47761), .A2(n47760), .ZN(n47764) );
  NAND2HSV0 U51528 ( .A1(n47835), .A2(n57567), .ZN(n47763) );
  CLKNAND2HSV0 U51529 ( .A1(n50288), .A2(n57564), .ZN(n47762) );
  XOR3HSV1 U51530 ( .A1(n47764), .A2(n47763), .A3(n47762), .Z(n47765) );
  XNOR2HSV1 U51531 ( .A1(n47766), .A2(n47765), .ZN(n47769) );
  NAND2HSV2 U51532 ( .A1(n58183), .A2(\pe4/got [24]), .ZN(n47768) );
  CLKNAND2HSV0 U51533 ( .A1(n58037), .A2(n57309), .ZN(n47767) );
  NAND2HSV0 U51534 ( .A1(n47774), .A2(n47773), .ZN(n47776) );
  INHSV2 U51535 ( .I(n47776), .ZN(n47779) );
  INHSV2 U51536 ( .I(n60077), .ZN(n47775) );
  NOR2HSV0 U51537 ( .A1(n47776), .A2(n35007), .ZN(n47782) );
  INHSV0 U51538 ( .I(n47782), .ZN(n47783) );
  CLKAND2HSV2 U51539 ( .A1(n47788), .A2(\pe4/ti_7t [31]), .Z(n47789) );
  INHSV2 U51540 ( .I(n26413), .ZN(n58254) );
  INHSV2 U51541 ( .I(\pe4/got [3]), .ZN(n58294) );
  NAND2HSV2 U51542 ( .A1(n58254), .A2(n58298), .ZN(n47790) );
  XNOR3HSV1 U51543 ( .A1(n47792), .A2(n47791), .A3(n47790), .ZN(\pe4/poht [29]) );
  INHSV2 U51544 ( .I(n50294), .ZN(n57974) );
  BUFHSV3 U51545 ( .I(n49921), .Z(n57673) );
  CLKNHSV2 U51546 ( .I(n49954), .ZN(n50189) );
  CLKNAND2HSV1 U51547 ( .A1(n57673), .A2(n50189), .ZN(n47852) );
  INHSV2 U51548 ( .I(n50064), .ZN(n58102) );
  NAND2HSV0 U51549 ( .A1(n50213), .A2(n58102), .ZN(n47840) );
  NAND2HSV0 U51550 ( .A1(n59378), .A2(n58219), .ZN(n47829) );
  CLKNAND2HSV0 U51551 ( .A1(n58087), .A2(\pe4/bq[11] ), .ZN(n47795) );
  NAND2HSV0 U51552 ( .A1(\pe4/aot [9]), .A2(\pe4/bq[10] ), .ZN(n47794) );
  XOR2HSV0 U51553 ( .A1(n47795), .A2(n47794), .Z(n47799) );
  CLKNAND2HSV1 U51554 ( .A1(n59683), .A2(n58130), .ZN(n47797) );
  NAND2HSV0 U51555 ( .A1(n59343), .A2(n58003), .ZN(n47796) );
  XOR2HSV0 U51556 ( .A1(n47797), .A2(n47796), .Z(n47798) );
  XOR2HSV0 U51557 ( .A1(n47799), .A2(n47798), .Z(n47827) );
  INHSV2 U51558 ( .I(n58013), .ZN(n57911) );
  CLKNAND2HSV0 U51559 ( .A1(n59605), .A2(n57911), .ZN(n47801) );
  CLKNHSV0 U51560 ( .I(n53217), .ZN(n58126) );
  NAND2HSV0 U51561 ( .A1(n58306), .A2(n58126), .ZN(n47800) );
  XOR2HSV0 U51562 ( .A1(n47801), .A2(n47800), .Z(n47806) );
  CLKNAND2HSV0 U51563 ( .A1(n57338), .A2(\pe4/bq[13] ), .ZN(n47804) );
  INHSV2 U51564 ( .I(n47905), .ZN(n57692) );
  NAND2HSV0 U51565 ( .A1(n57692), .A2(n57906), .ZN(n47803) );
  XOR2HSV0 U51566 ( .A1(n47804), .A2(n47803), .Z(n47805) );
  XNOR2HSV1 U51567 ( .A1(n47806), .A2(n47805), .ZN(n47808) );
  NAND2HSV0 U51568 ( .A1(\pe4/aot [17]), .A2(\pe4/bq[2] ), .ZN(n50354) );
  NAND2HSV0 U51569 ( .A1(n57234), .A2(n58301), .ZN(n49968) );
  XOR2HSV0 U51570 ( .A1(n50354), .A2(n49968), .Z(n47807) );
  XNOR2HSV1 U51571 ( .A1(n47808), .A2(n47807), .ZN(n47826) );
  NAND2HSV0 U51572 ( .A1(\pe4/aot [2]), .A2(n57926), .ZN(n47811) );
  NAND2HSV0 U51573 ( .A1(n58163), .A2(n57784), .ZN(n47810) );
  XOR2HSV0 U51574 ( .A1(n47811), .A2(n47810), .Z(n47815) );
  NAND2HSV0 U51575 ( .A1(n35347), .A2(\pe4/bq[4] ), .ZN(n47813) );
  NAND2HSV0 U51576 ( .A1(\pe4/aot [14]), .A2(n57837), .ZN(n47812) );
  XOR2HSV0 U51577 ( .A1(n47813), .A2(n47812), .Z(n47814) );
  XOR2HSV0 U51578 ( .A1(n47815), .A2(n47814), .Z(n47824) );
  CLKNAND2HSV1 U51579 ( .A1(n58198), .A2(n57986), .ZN(n47817) );
  BUFHSV2 U51580 ( .I(n47718), .Z(n57683) );
  CLKNAND2HSV0 U51581 ( .A1(n57683), .A2(n57135), .ZN(n47816) );
  XOR2HSV0 U51582 ( .A1(n47817), .A2(n47816), .Z(n47822) );
  NAND2HSV0 U51583 ( .A1(n58283), .A2(n49943), .ZN(n47820) );
  NAND2HSV0 U51584 ( .A1(n57230), .A2(n34879), .ZN(n47819) );
  XOR2HSV0 U51585 ( .A1(n47820), .A2(n47819), .Z(n47821) );
  XOR2HSV0 U51586 ( .A1(n47822), .A2(n47821), .Z(n47823) );
  XOR2HSV0 U51587 ( .A1(n47824), .A2(n47823), .Z(n47825) );
  XOR3HSV2 U51588 ( .A1(n47827), .A2(n47826), .A3(n47825), .Z(n47828) );
  XNOR2HSV1 U51589 ( .A1(n47829), .A2(n47828), .ZN(n47831) );
  NOR2HSV0 U51590 ( .A1(n57816), .A2(n58325), .ZN(n47830) );
  XNOR2HSV1 U51591 ( .A1(n47831), .A2(n47830), .ZN(n47834) );
  NAND2HSV0 U51592 ( .A1(n57550), .A2(n58298), .ZN(n47833) );
  BUFHSV2 U51593 ( .I(n58060), .Z(n57817) );
  NAND2HSV0 U51594 ( .A1(n57817), .A2(n58206), .ZN(n47832) );
  XOR3HSV2 U51595 ( .A1(n47834), .A2(n47833), .A3(n47832), .Z(n47838) );
  BUFHSV2 U51596 ( .I(n47835), .Z(n57308) );
  CLKNAND2HSV0 U51597 ( .A1(n57308), .A2(\pe4/got [6]), .ZN(n47837) );
  BUFHSV2 U51598 ( .I(n47969), .Z(n58097) );
  CLKNAND2HSV1 U51599 ( .A1(n58097), .A2(n58246), .ZN(n47836) );
  XOR3HSV2 U51600 ( .A1(n47838), .A2(n47837), .A3(n47836), .Z(n47839) );
  XNOR2HSV1 U51601 ( .A1(n47840), .A2(n47839), .ZN(n47845) );
  CLKNHSV2 U51602 ( .I(\pe4/got [9]), .ZN(n57836) );
  NAND2HSV2 U51603 ( .A1(n47841), .A2(n57818), .ZN(n47844) );
  BUFHSV2 U51604 ( .I(n47842), .Z(n58037) );
  CLKNAND2HSV0 U51605 ( .A1(n58037), .A2(\pe4/got [8]), .ZN(n47843) );
  XOR3HSV2 U51606 ( .A1(n47845), .A2(n47844), .A3(n47843), .Z(n47848) );
  CLKNAND2HSV1 U51607 ( .A1(n57889), .A2(n59663), .ZN(n47847) );
  XNOR2HSV1 U51608 ( .A1(n47848), .A2(n47847), .ZN(n47850) );
  CLKNAND2HSV0 U51609 ( .A1(n57755), .A2(\pe4/got [11]), .ZN(n47849) );
  XNOR2HSV1 U51610 ( .A1(n47850), .A2(n47849), .ZN(n47851) );
  XNOR2HSV1 U51611 ( .A1(n47852), .A2(n47851), .ZN(n47856) );
  CLKNAND2HSV0 U51612 ( .A1(n58141), .A2(n35400), .ZN(n47855) );
  NAND2HSV0 U51613 ( .A1(n57424), .A2(n50199), .ZN(n47854) );
  XOR3HSV2 U51614 ( .A1(n47856), .A2(n47855), .A3(n47854), .Z(n47858) );
  INHSV2 U51615 ( .I(n50212), .ZN(n57982) );
  CLKNAND2HSV0 U51616 ( .A1(n58207), .A2(n57982), .ZN(n47857) );
  XNOR2HSV1 U51617 ( .A1(n47858), .A2(n47857), .ZN(n47859) );
  XOR2HSV0 U51618 ( .A1(n47860), .A2(n47859), .Z(n47864) );
  NAND2HSV2 U51619 ( .A1(n58254), .A2(n57834), .ZN(n47862) );
  XNOR3HSV1 U51620 ( .A1(n47864), .A2(n47863), .A3(n47862), .ZN(\pe4/poht [14]) );
  CLKNAND2HSV1 U51621 ( .A1(n58299), .A2(n58140), .ZN(n47887) );
  BUFHSV2 U51622 ( .I(n47865), .Z(n58218) );
  NAND2HSV0 U51623 ( .A1(\pe4/aot [2]), .A2(n58116), .ZN(n47867) );
  NAND2HSV0 U51624 ( .A1(n59683), .A2(n57241), .ZN(n47866) );
  XOR2HSV0 U51625 ( .A1(n47867), .A2(n47866), .Z(n47871) );
  NAND2HSV0 U51626 ( .A1(n57993), .A2(n57595), .ZN(n47869) );
  NAND2HSV0 U51627 ( .A1(\pe4/aot [9]), .A2(n58301), .ZN(n47868) );
  XOR2HSV0 U51628 ( .A1(n47869), .A2(n47868), .Z(n47870) );
  XOR2HSV0 U51629 ( .A1(n47871), .A2(n47870), .Z(n47876) );
  INHSV2 U51630 ( .I(n57011), .ZN(n58199) );
  CLKNAND2HSV1 U51631 ( .A1(n58199), .A2(n58130), .ZN(n47873) );
  NAND2HSV0 U51632 ( .A1(n58223), .A2(n58197), .ZN(n47872) );
  XOR2HSV0 U51633 ( .A1(n47873), .A2(n47872), .Z(n47874) );
  NOR2HSV2 U51634 ( .A1(n35042), .A2(n48032), .ZN(n57840) );
  XNOR2HSV1 U51635 ( .A1(n47874), .A2(n57840), .ZN(n47875) );
  XNOR2HSV1 U51636 ( .A1(n47876), .A2(n47875), .ZN(n47883) );
  NAND2HSV0 U51637 ( .A1(n58230), .A2(\pe4/bq[11] ), .ZN(n47878) );
  BUFHSV2 U51638 ( .I(\pe4/bq[9] ), .Z(n58113) );
  CLKNAND2HSV0 U51639 ( .A1(n58283), .A2(n58113), .ZN(n47877) );
  XOR2HSV0 U51640 ( .A1(n47878), .A2(n47877), .Z(n47881) );
  CLKNAND2HSV1 U51641 ( .A1(\pe4/aot [6]), .A2(n58265), .ZN(n49985) );
  NAND2HSV0 U51642 ( .A1(n47718), .A2(\pe4/bq[2] ), .ZN(n47879) );
  XOR2HSV0 U51643 ( .A1(n49985), .A2(n47879), .Z(n47880) );
  XOR2HSV0 U51644 ( .A1(n47881), .A2(n47880), .Z(n47882) );
  NAND2HSV2 U51645 ( .A1(n47841), .A2(n58314), .ZN(n47884) );
  INHSV2 U51646 ( .I(n50298), .ZN(n58220) );
  INHSV2 U51647 ( .I(n50091), .ZN(n58258) );
  INHSV2 U51648 ( .I(n50064), .ZN(n58216) );
  XOR2HSV0 U51649 ( .A1(n47887), .A2(n47886), .Z(n47890) );
  NAND2HSV2 U51650 ( .A1(n58254), .A2(n58153), .ZN(n47888) );
  XNOR3HSV1 U51651 ( .A1(n47890), .A2(n47889), .A3(n47888), .ZN(\pe4/poht [21]) );
  INHSV2 U51652 ( .I(n50910), .ZN(n52901) );
  CLKNAND2HSV0 U51653 ( .A1(n52456), .A2(n51532), .ZN(n47892) );
  NAND2HSV0 U51654 ( .A1(n59499), .A2(n51493), .ZN(n47891) );
  XOR2HSV0 U51655 ( .A1(n47892), .A2(n47891), .Z(n47897) );
  INHSV2 U51656 ( .I(\pe2/bq[5] ), .ZN(n51842) );
  NOR2HSV2 U51657 ( .A1(n49618), .A2(n51842), .ZN(n47895) );
  INHSV2 U51658 ( .I(n47893), .ZN(n52905) );
  NAND2HSV0 U51659 ( .A1(n51486), .A2(n52905), .ZN(n47894) );
  XOR2HSV0 U51660 ( .A1(n47895), .A2(n47894), .Z(n47896) );
  XNOR2HSV1 U51661 ( .A1(n47897), .A2(n47896), .ZN(n47900) );
  CLKNAND2HSV1 U51662 ( .A1(n52867), .A2(n52309), .ZN(n51452) );
  NAND2HSV0 U51663 ( .A1(n51547), .A2(\pe2/bq[6] ), .ZN(n47898) );
  XOR2HSV0 U51664 ( .A1(n51452), .A2(n47898), .Z(n47899) );
  CLKNAND2HSV1 U51665 ( .A1(n58299), .A2(\pe4/got [8]), .ZN(n47922) );
  NOR2HSV1 U51666 ( .A1(n57011), .A2(n50114), .ZN(n57231) );
  CLKNAND2HSV1 U51667 ( .A1(\pe4/aot [1]), .A2(n58116), .ZN(n47906) );
  CLKNAND2HSV0 U51668 ( .A1(n58283), .A2(n58130), .ZN(n47908) );
  NAND2HSV0 U51669 ( .A1(\pe4/aot [2]), .A2(n57798), .ZN(n47907) );
  XOR2HSV0 U51670 ( .A1(n47908), .A2(n47907), .Z(n47912) );
  NOR2HSV1 U51671 ( .A1(n49929), .A2(n50351), .ZN(n47910) );
  NAND2HSV0 U51672 ( .A1(n47718), .A2(\pe4/bq[1] ), .ZN(n47909) );
  XOR2HSV0 U51673 ( .A1(n47910), .A2(n47909), .Z(n47911) );
  XNOR2HSV1 U51674 ( .A1(n47912), .A2(n47911), .ZN(n47919) );
  CLKNAND2HSV0 U51675 ( .A1(n58070), .A2(n58155), .ZN(n47914) );
  NAND2HSV0 U51676 ( .A1(n58198), .A2(n58156), .ZN(n47913) );
  XOR2HSV0 U51677 ( .A1(n47914), .A2(n47913), .Z(n47918) );
  NOR2HSV1 U51678 ( .A1(n57775), .A2(n57010), .ZN(n47916) );
  NAND2HSV0 U51679 ( .A1(\pe4/aot [9]), .A2(\pe4/bq[2] ), .ZN(n47915) );
  XOR2HSV0 U51680 ( .A1(n47916), .A2(n47915), .Z(n47917) );
  XNOR2HSV1 U51681 ( .A1(n47922), .A2(n47921), .ZN(n47925) );
  NOR2HSV2 U51682 ( .A1(n29774), .A2(n57836), .ZN(n47924) );
  NOR2HSV0 U51683 ( .A1(n26413), .A2(n49922), .ZN(n47923) );
  INHSV2 U51684 ( .I(n50211), .ZN(n58048) );
  CLKNAND2HSV0 U51685 ( .A1(n58048), .A2(n34843), .ZN(n47929) );
  XNOR2HSV0 U51686 ( .A1(n47929), .A2(n29739), .ZN(n47931) );
  XNOR2HSV0 U51687 ( .A1(n47931), .A2(n47930), .ZN(n60055) );
  INHSV2 U51688 ( .I(n54146), .ZN(n55512) );
  INAND2HSV2 U51689 ( .A1(n55512), .B1(n52831), .ZN(n47937) );
  XNOR2HSV0 U51690 ( .A1(n47937), .A2(n47936), .ZN(n60063) );
  INHSV1 U51691 ( .I(n47939), .ZN(n51949) );
  CLKNHSV0 U51692 ( .I(n47943), .ZN(n47945) );
  NAND2HSV2 U51693 ( .A1(n58183), .A2(n47772), .ZN(n47944) );
  XNOR2HSV1 U51694 ( .A1(n47945), .A2(n47944), .ZN(pov4[23]) );
  OAI21HSV0 U51695 ( .A1(n39669), .A2(n47948), .B(n47947), .ZN(n60007) );
  INHSV0 U51696 ( .I(n47952), .ZN(n47954) );
  XOR2HSV0 U51697 ( .A1(n47954), .A2(n47953), .Z(n47955) );
  CLKNAND2HSV1 U51698 ( .A1(n47955), .A2(n46546), .ZN(n47956) );
  XNOR2HSV1 U51699 ( .A1(n47956), .A2(poh6[20]), .ZN(po[21]) );
  NAND2HSV0 U51700 ( .A1(n59360), .A2(n53649), .ZN(n47959) );
  XOR3HSV0 U51701 ( .A1(n25858), .A2(n47959), .A3(n47958), .Z(pov1[21]) );
  NAND3HSV0 U51702 ( .A1(n47964), .A2(n47963), .A3(n47962), .ZN(n47966) );
  XNOR2HSV0 U51703 ( .A1(n47966), .A2(n47965), .ZN(n47968) );
  XNOR2HSV0 U51704 ( .A1(n47968), .A2(n47967), .ZN(pov4[20]) );
  BUFHSV2 U51705 ( .I(n47969), .Z(n59935) );
  XNOR2HSV0 U51706 ( .A1(n47974), .A2(n47973), .ZN(n47975) );
  NAND2HSV0 U51707 ( .A1(n47975), .A2(n46546), .ZN(n47976) );
  XNOR2HSV1 U51708 ( .A1(n47976), .A2(poh6[15]), .ZN(po[16]) );
  CLKBUFHSV0 U51709 ( .I(n47981), .Z(n47982) );
  CLKNHSV0 U51710 ( .I(n47983), .ZN(n47986) );
  NAND2HSV0 U51711 ( .A1(n54513), .A2(n53650), .ZN(n47985) );
  XOR3HSV0 U51712 ( .A1(n47987), .A2(n47986), .A3(n47985), .Z(pov1[12]) );
  CLKNHSV0 U51713 ( .I(n48083), .ZN(n59443) );
  BUFHSV2 U51714 ( .I(n59491), .Z(n59659) );
  BUFHSV2 U51715 ( .I(n59925), .Z(n59656) );
  CLKBUFHSV2 U51716 ( .I(n47988), .Z(n47989) );
  NAND2HSV0 U51717 ( .A1(n47991), .A2(n52726), .ZN(n47993) );
  XNOR2HSV0 U51718 ( .A1(n47993), .A2(n47992), .ZN(n60090) );
  NAND2HSV0 U51719 ( .A1(n52580), .A2(n52767), .ZN(n47995) );
  XNOR2HSV0 U51720 ( .A1(n47995), .A2(n47994), .ZN(n60071) );
  BUFHSV2 U51721 ( .I(n47999), .Z(n54456) );
  BUFHSV2 U51722 ( .I(n48007), .Z(n48008) );
  CLKNHSV0 U51723 ( .I(n59461), .ZN(n48473) );
  INHSV2 U51724 ( .I(n49967), .ZN(n59958) );
  NAND2HSV0 U51725 ( .A1(n34127), .A2(n52723), .ZN(n48016) );
  MUX2HSV2 U51726 ( .I0(bo3[1]), .I1(n56971), .S(n48019), .Z(n59796) );
  MUX2HSV2 U51727 ( .I0(bo3[11]), .I1(\pe3/bq[11] ), .S(n48019), .Z(n59781) );
  MUX2HSV2 U51728 ( .I0(bo3[29]), .I1(n48021), .S(n48020), .Z(n59763) );
  MUX2HSV2 U51729 ( .I0(bo3[28]), .I1(n42634), .S(n59537), .Z(n59764) );
  MUX2HSV2 U51730 ( .I0(bo5[23]), .I1(\pe5/bq[23] ), .S(n48077), .Z(n59846) );
  MUX2HSV2 U51731 ( .I0(bo5[20]), .I1(n39487), .S(n48045), .Z(n59848) );
  MUX2HSV2 U51732 ( .I0(bo4[3]), .I1(n58301), .S(n48073), .Z(n59828) );
  MUX2HSV2 U51733 ( .I0(bo2[7]), .I1(n52859), .S(n53222), .Z(n59746) );
  MUX2HSV2 U51734 ( .I0(bo4[19]), .I1(n57929), .S(n59486), .Z(n59817) );
  MUX2HSV2 U51735 ( .I0(bo4[20]), .I1(n57785), .S(n34770), .Z(n59815) );
  MUX2HSV2 U51736 ( .I0(bo4[16]), .I1(n49943), .S(n48072), .Z(n59819) );
  MUX2HSV2 U51737 ( .I0(bo6[11]), .I1(n46210), .S(n48025), .Z(n59904) );
  MUX2HSV2 U51738 ( .I0(bo6[13]), .I1(n59089), .S(n59902), .Z(n59901) );
  MUX2HSV2 U51739 ( .I0(bo4[18]), .I1(\pe4/bq[18] ), .S(n48072), .Z(n59818) );
  MUX2HSV2 U51740 ( .I0(bo5[17]), .I1(n48236), .S(n44335), .Z(n59853) );
  MUX2HSV2 U51741 ( .I0(bo5[18]), .I1(n52618), .S(n48077), .Z(n59855) );
  MUX2HSV2 U51742 ( .I0(bo5[26]), .I1(n52594), .S(n48027), .Z(n59844) );
  MUX2HSV2 U51743 ( .I0(bo4[8]), .I1(n58130), .S(n48073), .Z(n59824) );
  MUX2HSV2 U51744 ( .I0(bo5[8]), .I1(n52672), .S(n48077), .Z(n59859) );
  MUX2HSV2 U51745 ( .I0(bo5[9]), .I1(n48775), .S(n53215), .Z(n59858) );
  MUX2HSV2 U51746 ( .I0(bo5[15]), .I1(n53314), .S(n48039), .Z(n59856) );
  MUX2HSV1 U51747 ( .I0(bo5[12]), .I1(\pe5/bq[12] ), .S(n48029), .Z(n59860) );
  CLKNHSV1 U51748 ( .I(n48030), .ZN(n55241) );
  BUFHSV2 U51749 ( .I(\pe1/ctrq ), .Z(n48081) );
  MUX2HSV2 U51750 ( .I0(bo1[11]), .I1(n55241), .S(n48081), .Z(n59712) );
  MUX2HSV2 U51751 ( .I0(bo2[13]), .I1(n51729), .S(n48062), .Z(n59744) );
  MUX2HSV2 U51752 ( .I0(bo5[3]), .I1(n53200), .S(n48027), .Z(n59864) );
  MUX2HSV2 U51753 ( .I0(bo5[29]), .I1(n30547), .S(n53215), .Z(n59836) );
  MUX2HSV2 U51754 ( .I0(bo4[5]), .I1(n58155), .S(n53218), .Z(n59825) );
  MUX2HSV2 U51755 ( .I0(bo1[3]), .I1(n55577), .S(\pe1/ctrq ), .Z(n59720) );
  INHSV2 U51756 ( .I(n54093), .ZN(n55505) );
  MUX2HSV2 U51757 ( .I0(bo1[7]), .I1(n55505), .S(\pe1/ctrq ), .Z(n59716) );
  MUX2HSV2 U51758 ( .I0(bo1[28]), .I1(n53805), .S(n48054), .Z(n59689) );
  MUX2HSV2 U51759 ( .I0(bo1[10]), .I1(n55379), .S(n48080), .Z(n59713) );
  BUFHSV2 U51760 ( .I(n48065), .Z(n48057) );
  MUX2HSV2 U51761 ( .I0(bo2[6]), .I1(n52866), .S(n48057), .Z(n59749) );
  MUX2HSV2 U51762 ( .I0(bo2[10]), .I1(n51997), .S(n53222), .Z(n59747) );
  MUX2HSV2 U51763 ( .I0(bo2[4]), .I1(n52309), .S(n53224), .Z(n59752) );
  MUX2HSV2 U51764 ( .I0(bo2[3]), .I1(n52905), .S(n48033), .Z(n59754) );
  MUX2HSV2 U51765 ( .I0(bo2[9]), .I1(n51623), .S(n48062), .Z(n59748) );
  MUX2HSV1 U51766 ( .I0(bo5[7]), .I1(\pe5/bq[7] ), .S(n48029), .Z(n59861) );
  MUX2HSV1 U51767 ( .I0(bo5[5]), .I1(n52671), .S(n48034), .Z(n59862) );
  MUX2HSV1 U51768 ( .I0(bo6[26]), .I1(n48035), .S(n48025), .Z(n59875) );
  MUX2HSV2 U51769 ( .I0(bo6[5]), .I1(n48037), .S(n44701), .Z(n59911) );
  MUX2HSV2 U51770 ( .I0(bo2[1]), .I1(n51532), .S(n53225), .Z(n59753) );
  MUX2HSV2 U51771 ( .I0(bo6[6]), .I1(n48038), .S(n48025), .Z(n59910) );
  MUX2HSV2 U51772 ( .I0(bo6[7]), .I1(n58460), .S(n48025), .Z(n59909) );
  MUX2HSV2 U51773 ( .I0(bo5[32]), .I1(n31192), .S(n48077), .Z(n59830) );
  BUFHSV2 U51774 ( .I(n48043), .Z(n48048) );
  MUX2HSV2 U51775 ( .I0(bo6[8]), .I1(n58619), .S(n48048), .Z(n59907) );
  MUX2HSV2 U51776 ( .I0(bo6[9]), .I1(n48044), .S(n48025), .Z(n59908) );
  MUX2HSV2 U51777 ( .I0(bo5[28]), .I1(n30164), .S(n48045), .Z(n59840) );
  MUX2HSV2 U51778 ( .I0(bo6[1]), .I1(n58336), .S(n48025), .Z(n59687) );
  MUX2HSV2 U51779 ( .I0(bo6[3]), .I1(n49205), .S(n53214), .Z(n59913) );
  MUX2HSV2 U51780 ( .I0(bo6[4]), .I1(n59062), .S(n48046), .Z(n59912) );
  MUX2HSV2 U51781 ( .I0(bo6[15]), .I1(n58682), .S(n48048), .Z(n59900) );
  MUX2HSV2 U51782 ( .I0(bo5[16]), .I1(n48181), .S(n48077), .Z(n59851) );
  MUX2HSV2 U51783 ( .I0(bo5[13]), .I1(n50668), .S(n48077), .Z(n59854) );
  MUX2HSV2 U51784 ( .I0(bo6[12]), .I1(n48051), .S(n48025), .Z(n59899) );
  MUX2HSV2 U51785 ( .I0(bo2[25]), .I1(n44987), .S(n48052), .Z(n59729) );
  MUX2HSV2 U51786 ( .I0(bo4[1]), .I1(n58322), .S(n48073), .Z(n59829) );
  MUX2HSV2 U51787 ( .I0(bo2[24]), .I1(n38542), .S(n48052), .Z(n59731) );
  MUX2HSV2 U51788 ( .I0(bo1[29]), .I1(n40553), .S(n48053), .Z(n59693) );
  MUX2HSV2 U51789 ( .I0(bo1[31]), .I1(n48055), .S(n48054), .Z(n59690) );
  MUX2HSV2 U51790 ( .I0(bo4[23]), .I1(n57476), .S(n48073), .Z(n59812) );
  MUX2HSV2 U51791 ( .I0(bo2[21]), .I1(\pe2/bq[21] ), .S(n48057), .Z(n59735) );
  MUX2HSV2 U51792 ( .I0(bo4[12]), .I1(n58077), .S(n48073), .Z(n59822) );
  MUX2HSV2 U51793 ( .I0(bo1[32]), .I1(n40684), .S(n48076), .Z(n59692) );
  MUX2HSV2 U51794 ( .I0(bo4[15]), .I1(n34879), .S(n48068), .Z(n59820) );
  MUX2HSV2 U51795 ( .I0(bo4[24]), .I1(\pe4/bq[24] ), .S(n48058), .Z(n59814) );
  MUX2HSV2 U51796 ( .I0(bo2[28]), .I1(n52987), .S(n59497), .Z(n59726) );
  MUX2HSV2 U51797 ( .I0(bo1[13]), .I1(\pe1/bq[13] ), .S(n48081), .Z(n59707) );
  CLKNHSV0 U51798 ( .I(n54185), .ZN(n53949) );
  MUX2HSV2 U51799 ( .I0(bo1[24]), .I1(n53949), .S(n48080), .Z(n59696) );
  MUX2HSV2 U51800 ( .I0(bo1[20]), .I1(n42238), .S(n48061), .Z(n59701) );
  CLKNHSV0 U51801 ( .I(n54281), .ZN(n54999) );
  MUX2HSV2 U51802 ( .I0(bo1[14]), .I1(n54999), .S(n48053), .Z(n59708) );
  MUX2HSV2 U51803 ( .I0(bo1[25]), .I1(n41173), .S(n48061), .Z(n59697) );
  INHSV2 U51804 ( .I(n51537), .ZN(n59978) );
  MUX2HSV2 U51805 ( .I0(bo1[5]), .I1(n54289), .S(n48080), .Z(n59715) );
  MUX2HSV2 U51806 ( .I0(bo1[2]), .I1(n55451), .S(\pe1/ctrq ), .Z(n59719) );
  MUX2HSV2 U51807 ( .I0(bo1[1]), .I1(n55495), .S(n48053), .Z(n59718) );
  MUX2HSV2 U51808 ( .I0(bo2[11]), .I1(n51900), .S(n48052), .Z(n59745) );
  MUX2HSV2 U51809 ( .I0(bo2[16]), .I1(n51732), .S(n48067), .Z(n59741) );
  MUX2HSV2 U51810 ( .I0(bo2[18]), .I1(n52988), .S(n53224), .Z(n59739) );
  MUX2HSV2 U51811 ( .I0(bo2[15]), .I1(n49619), .S(n48033), .Z(n59743) );
  MUX2HSV2 U51812 ( .I0(bo2[14]), .I1(\pe2/bq[14] ), .S(n48067), .Z(n59742) );
  MUX2HSV1 U51813 ( .I0(bo4[28]), .I1(n48069), .S(n48068), .Z(n59806) );
  MUX2HSV2 U51814 ( .I0(bo4[29]), .I1(n33533), .S(n48072), .Z(n59805) );
  CLKNHSV0 U51815 ( .I(n48070), .ZN(n57337) );
  BUFHSV2 U51816 ( .I(n53218), .Z(n53220) );
  MUX2HSV2 U51817 ( .I0(bo4[25]), .I1(n57337), .S(n53220), .Z(n59801) );
  MUX2HSV1 U51818 ( .I0(bo4[26]), .I1(n48071), .S(n53220), .Z(n59803) );
  MUX2HSV2 U51819 ( .I0(bo4[27]), .I1(\pe4/bq[27] ), .S(n48072), .Z(n59802) );
  MUX2HSV1 U51820 ( .I0(bo4[32]), .I1(n48074), .S(n48073), .Z(n59798) );
  MUX2HSV1 U51821 ( .I0(bo3[12]), .I1(n56507), .S(n46139), .Z(n59782) );
  MUX2HSV2 U51822 ( .I0(bo1[18]), .I1(\pe1/bq[18] ), .S(n48076), .Z(n59704) );
  MUX2HSV2 U51823 ( .I0(bo5[14]), .I1(n39472), .S(n48077), .Z(n59852) );
  MUX2HSV2 U51824 ( .I0(bo1[22]), .I1(n54465), .S(n48080), .Z(n59700) );
  MUX2HSV2 U51825 ( .I0(bo2[29]), .I1(n36608), .S(n48079), .Z(n59723) );
  MUX2HSV2 U51826 ( .I0(bo2[27]), .I1(n52973), .S(n48079), .Z(n59727) );
  MUX2HSV2 U51827 ( .I0(bo1[4]), .I1(n55544), .S(n48061), .Z(n59717) );
  MUX2HSV2 U51828 ( .I0(bo1[6]), .I1(n55231), .S(n48080), .Z(n59714) );
  BUFHSV2 U51829 ( .I(\pe1/bq[8] ), .Z(n55501) );
  MUX2HSV2 U51830 ( .I0(bo1[8]), .I1(n55501), .S(n48081), .Z(n59711) );
  MUX2HSV2 U51831 ( .I0(bo2[17]), .I1(\pe2/bq[17] ), .S(n48067), .Z(n59740) );
  MUX2HSV2 U51832 ( .I0(bo4[7]), .I1(\pe4/bq[7] ), .S(n34138), .Z(n59826) );
  MUX2HSV2 U51833 ( .I0(bo4[6]), .I1(n58265), .S(n48082), .Z(n59827) );
  CLKNHSV0 U51834 ( .I(n59474), .ZN(n48472) );
  CLKNHSV0 U51835 ( .I(n48472), .ZN(n59396) );
  CLKNHSV0 U51836 ( .I(n48478), .ZN(n59397) );
  CLKNHSV0 U51837 ( .I(n59660), .ZN(n59399) );
  CLKNHSV0 U51838 ( .I(n59455), .ZN(n48475) );
  CLKNHSV0 U51839 ( .I(n59655), .ZN(n48478) );
  CLKNHSV0 U51840 ( .I(n59660), .ZN(n59400) );
  CLKNHSV0 U51841 ( .I(n48478), .ZN(n59401) );
  BUFHSV2 U51842 ( .I(n48474), .Z(n48479) );
  CLKNHSV0 U51843 ( .I(n48479), .ZN(n59402) );
  CLKNHSV0 U51844 ( .I(n48479), .ZN(n59403) );
  CLKNHSV0 U51845 ( .I(n48015), .ZN(n59404) );
  CLKNHSV0 U51846 ( .I(n48472), .ZN(n59405) );
  CLKNHSV0 U51847 ( .I(n48015), .ZN(n59406) );
  CLKNHSV0 U51848 ( .I(n59660), .ZN(n59407) );
  CLKNHSV0 U51849 ( .I(n48015), .ZN(n59408) );
  CLKNHSV0 U51850 ( .I(n48015), .ZN(n59409) );
  CLKNHSV0 U51851 ( .I(n48477), .ZN(n59410) );
  CLKNHSV0 U51852 ( .I(n48479), .ZN(n59468) );
  CLKNHSV0 U51853 ( .I(n48477), .ZN(n59411) );
  CLKNHSV0 U51854 ( .I(n48477), .ZN(n59412) );
  CLKNHSV0 U51855 ( .I(n48473), .ZN(n59413) );
  BUFHSV2 U51856 ( .I(n59452), .Z(n59924) );
  CLKNHSV0 U51857 ( .I(n59650), .ZN(n48476) );
  CLKNHSV0 U51858 ( .I(n48477), .ZN(n59433) );
  CLKNHSV0 U51859 ( .I(n48479), .ZN(n59414) );
  CLKNHSV0 U51860 ( .I(n48478), .ZN(n59415) );
  CLKNHSV0 U51861 ( .I(n48475), .ZN(n59416) );
  CLKNHSV0 U51862 ( .I(n48015), .ZN(n59450) );
  CLKNHSV0 U51863 ( .I(n48472), .ZN(n59417) );
  CLKNAND2HSV1 U51864 ( .A1(n59475), .A2(n51889), .ZN(n48159) );
  CLKNAND2HSV1 U51865 ( .A1(n25835), .A2(n52050), .ZN(n48157) );
  NAND2HSV0 U51866 ( .A1(n59790), .A2(n52051), .ZN(n48152) );
  CLKNAND2HSV1 U51867 ( .A1(n51799), .A2(n48084), .ZN(n48150) );
  NOR2HSV1 U51868 ( .A1(n44833), .A2(n47555), .ZN(n48148) );
  NAND2HSV0 U51869 ( .A1(n59506), .A2(\pe2/got [8]), .ZN(n48140) );
  CLKNAND2HSV0 U51870 ( .A1(n52926), .A2(n59777), .ZN(n48138) );
  CLKNAND2HSV0 U51871 ( .A1(n51965), .A2(n59778), .ZN(n48135) );
  CLKNAND2HSV0 U51872 ( .A1(n51609), .A2(\pe2/got [4]), .ZN(n48133) );
  NAND2HSV0 U51873 ( .A1(\pe2/got [2]), .A2(n52419), .ZN(n48131) );
  NAND2HSV0 U51874 ( .A1(n50929), .A2(n52896), .ZN(n48128) );
  NAND2HSV0 U51875 ( .A1(n59636), .A2(n52481), .ZN(n48086) );
  NAND2HSV0 U51876 ( .A1(n59633), .A2(n51732), .ZN(n48085) );
  XOR2HSV0 U51877 ( .A1(n48086), .A2(n48085), .Z(n48090) );
  NAND2HSV0 U51878 ( .A1(n51460), .A2(n51729), .ZN(n48088) );
  NAND2HSV0 U51879 ( .A1(n39052), .A2(\pe2/bq[3] ), .ZN(n48087) );
  XOR2HSV0 U51880 ( .A1(n48088), .A2(n48087), .Z(n48089) );
  XOR2HSV0 U51881 ( .A1(n48090), .A2(n48089), .Z(n48098) );
  NAND2HSV0 U51882 ( .A1(\pe2/aot [16]), .A2(n51832), .ZN(n48092) );
  NAND2HSV0 U51883 ( .A1(\pe2/aot [11]), .A2(n51733), .ZN(n48091) );
  XOR2HSV0 U51884 ( .A1(n48092), .A2(n48091), .Z(n48096) );
  NAND2HSV0 U51885 ( .A1(\pe2/aot [12]), .A2(n52073), .ZN(n48094) );
  NAND2HSV0 U51886 ( .A1(n52104), .A2(n51805), .ZN(n48093) );
  XOR2HSV0 U51887 ( .A1(n48094), .A2(n48093), .Z(n48095) );
  XOR2HSV0 U51888 ( .A1(n48096), .A2(n48095), .Z(n48097) );
  XOR2HSV0 U51889 ( .A1(n48098), .A2(n48097), .Z(n48110) );
  NOR2HSV0 U51890 ( .A1(n47503), .A2(n51567), .ZN(n48100) );
  NAND2HSV0 U51891 ( .A1(\pe2/aot [8]), .A2(n49619), .ZN(n48099) );
  XOR2HSV0 U51892 ( .A1(n48100), .A2(n48099), .Z(n48104) );
  NOR2HSV0 U51893 ( .A1(n44871), .A2(n48621), .ZN(n52214) );
  CLKNHSV0 U51894 ( .I(n52214), .ZN(n48102) );
  NAND2HSV0 U51895 ( .A1(n37801), .A2(n51614), .ZN(n52446) );
  OAI21HSV0 U51896 ( .A1(n48621), .A2(n52080), .B(n52446), .ZN(n48101) );
  OAI21HSV2 U51897 ( .A1(n48102), .A2(n51817), .B(n48101), .ZN(n48103) );
  XNOR2HSV1 U51898 ( .A1(n48104), .A2(n48103), .ZN(n48108) );
  NAND2HSV0 U51899 ( .A1(n52056), .A2(n52988), .ZN(n48105) );
  XOR2HSV0 U51900 ( .A1(n48106), .A2(n48105), .Z(n48107) );
  XNOR2HSV1 U51901 ( .A1(n48108), .A2(n48107), .ZN(n48109) );
  XNOR2HSV1 U51902 ( .A1(n48110), .A2(n48109), .ZN(n48126) );
  CLKNAND2HSV0 U51903 ( .A1(n59975), .A2(n52063), .ZN(n48112) );
  CLKNAND2HSV0 U51904 ( .A1(n52344), .A2(n44197), .ZN(n48111) );
  XOR2HSV0 U51905 ( .A1(n48112), .A2(n48111), .Z(n48116) );
  NAND2HSV0 U51906 ( .A1(n52858), .A2(n43961), .ZN(n48114) );
  NAND2HSV0 U51907 ( .A1(\pe2/aot [6]), .A2(\pe2/bq[17] ), .ZN(n48113) );
  XOR2HSV0 U51908 ( .A1(n48114), .A2(n48113), .Z(n48115) );
  XOR2HSV0 U51909 ( .A1(n48116), .A2(n48115), .Z(n48124) );
  NAND2HSV0 U51910 ( .A1(\pe2/aot [2]), .A2(\pe2/bq[21] ), .ZN(n48118) );
  NAND2HSV0 U51911 ( .A1(n59783), .A2(n52299), .ZN(n48117) );
  XOR2HSV0 U51912 ( .A1(n48118), .A2(n48117), .Z(n48122) );
  NOR2HSV0 U51913 ( .A1(n52103), .A2(n51842), .ZN(n48120) );
  NAND2HSV0 U51914 ( .A1(n51759), .A2(\pe2/bq[6] ), .ZN(n48119) );
  XOR2HSV0 U51915 ( .A1(n48120), .A2(n48119), .Z(n48121) );
  XOR2HSV0 U51916 ( .A1(n48122), .A2(n48121), .Z(n48123) );
  XOR2HSV0 U51917 ( .A1(n48124), .A2(n48123), .Z(n48125) );
  XNOR2HSV1 U51918 ( .A1(n48126), .A2(n48125), .ZN(n48127) );
  XNOR2HSV1 U51919 ( .A1(n48128), .A2(n48127), .ZN(n48130) );
  NAND2HSV0 U51920 ( .A1(n51610), .A2(n52900), .ZN(n48129) );
  XOR3HSV2 U51921 ( .A1(n48131), .A2(n48130), .A3(n48129), .Z(n48132) );
  XNOR2HSV1 U51922 ( .A1(n48133), .A2(n48132), .ZN(n48134) );
  XNOR2HSV1 U51923 ( .A1(n48135), .A2(n48134), .ZN(n48137) );
  NAND2HSV0 U51924 ( .A1(n52251), .A2(n52125), .ZN(n48136) );
  XOR3HSV2 U51925 ( .A1(n48138), .A2(n48137), .A3(n48136), .Z(n48139) );
  XNOR2HSV1 U51926 ( .A1(n48140), .A2(n48139), .ZN(n48143) );
  NAND2HSV2 U51927 ( .A1(n51861), .A2(n52052), .ZN(n48142) );
  CLKNAND2HSV1 U51928 ( .A1(n52138), .A2(\pe2/got [10]), .ZN(n48141) );
  XOR3HSV2 U51929 ( .A1(n48143), .A2(n48142), .A3(n48141), .Z(n48144) );
  XNOR2HSV1 U51930 ( .A1(n48145), .A2(n48144), .ZN(n48147) );
  CLKNAND2HSV1 U51931 ( .A1(n51782), .A2(n53055), .ZN(n48146) );
  XOR3HSV2 U51932 ( .A1(n48148), .A2(n48147), .A3(n48146), .Z(n48149) );
  XOR2HSV0 U51933 ( .A1(n48150), .A2(n48149), .Z(n48151) );
  XOR2HSV0 U51934 ( .A1(n48152), .A2(n48151), .Z(n48155) );
  NAND2HSV2 U51935 ( .A1(n51728), .A2(n51796), .ZN(n48154) );
  INHSV2 U51936 ( .I(n47939), .ZN(n51792) );
  CLKNAND2HSV0 U51937 ( .A1(n51792), .A2(n47571), .ZN(n48153) );
  XOR3HSV2 U51938 ( .A1(n48155), .A2(n48154), .A3(n48153), .Z(n48156) );
  XOR2HSV0 U51939 ( .A1(n48157), .A2(n48156), .Z(n48158) );
  XOR2HSV0 U51940 ( .A1(n48159), .A2(n48158), .Z(n48160) );
  INHSV4 U51941 ( .I(n59789), .ZN(n51727) );
  NOR2HSV4 U51942 ( .A1(n48162), .A2(n48161), .ZN(n51150) );
  CLKNAND2HSV0 U51943 ( .A1(n52558), .A2(n52276), .ZN(n48163) );
  NAND2HSV2 U51944 ( .A1(n59933), .A2(n39430), .ZN(n48308) );
  CLKNAND2HSV0 U51945 ( .A1(n51014), .A2(\pe5/got [27]), .ZN(n48306) );
  CLKNAND2HSV0 U51946 ( .A1(n52670), .A2(\pe5/got [25]), .ZN(n48302) );
  CLKNAND2HSV0 U51947 ( .A1(n51016), .A2(\pe5/got [23]), .ZN(n48298) );
  NOR2HSV0 U51948 ( .A1(n50692), .A2(n47140), .ZN(n48296) );
  NAND2HSV0 U51949 ( .A1(n48745), .A2(n51228), .ZN(n48294) );
  NOR2HSV0 U51950 ( .A1(n48166), .A2(n39119), .ZN(n48292) );
  NAND2HSV0 U51951 ( .A1(n48746), .A2(n52566), .ZN(n48288) );
  NAND2HSV0 U51952 ( .A1(n48747), .A2(n51156), .ZN(n48286) );
  NAND2HSV0 U51953 ( .A1(n51018), .A2(n51015), .ZN(n48282) );
  NAND2HSV0 U51954 ( .A1(n51160), .A2(n52568), .ZN(n48278) );
  NAND2HSV0 U51955 ( .A1(n59392), .A2(n48167), .ZN(n48276) );
  NAND2HSV0 U51956 ( .A1(n59871), .A2(n48749), .ZN(n48274) );
  NAND2HSV0 U51957 ( .A1(n39745), .A2(n50424), .ZN(n48272) );
  NAND2HSV0 U51958 ( .A1(n48624), .A2(n52641), .ZN(n48270) );
  NAND2HSV0 U51959 ( .A1(n52580), .A2(n50698), .ZN(n48268) );
  NAND2HSV0 U51960 ( .A1(n48750), .A2(\pe5/got [6]), .ZN(n48264) );
  NAND2HSV0 U51961 ( .A1(n48168), .A2(n48841), .ZN(n48262) );
  NAND2HSV0 U51962 ( .A1(n48169), .A2(n51302), .ZN(n48260) );
  NAND2HSV0 U51963 ( .A1(n48751), .A2(n51331), .ZN(n48218) );
  NAND2HSV0 U51964 ( .A1(n48171), .A2(n48170), .ZN(n48174) );
  NAND2HSV0 U51965 ( .A1(n48172), .A2(\pe5/bq[1] ), .ZN(n48173) );
  XOR2HSV0 U51966 ( .A1(n48174), .A2(n48173), .Z(n48180) );
  NOR2HSV0 U51967 ( .A1(n48175), .A2(n51021), .ZN(n48178) );
  OAI22HSV0 U51968 ( .A1(n48677), .A2(n48178), .B1(n48177), .B2(n48176), .ZN(
        n48179) );
  XNOR2HSV1 U51969 ( .A1(n48180), .A2(n48179), .ZN(n48192) );
  NAND2HSV0 U51970 ( .A1(\pe5/aot [1]), .A2(n48181), .ZN(n53322) );
  NOR2HSV0 U51971 ( .A1(n48182), .A2(n53322), .ZN(n48184) );
  CLKNHSV0 U51972 ( .I(n45904), .ZN(n48810) );
  AOI22HSV0 U51973 ( .A1(\pe5/aot [16]), .A2(n52610), .B1(n30698), .B2(n48810), 
        .ZN(n48183) );
  NOR2HSV2 U51974 ( .A1(n48184), .A2(n48183), .ZN(n48190) );
  NAND2HSV0 U51975 ( .A1(\pe5/aot [18]), .A2(\pe5/bq[2] ), .ZN(n50517) );
  NOR2HSV0 U51976 ( .A1(n48185), .A2(n50517), .ZN(n48188) );
  AOI22HSV0 U51977 ( .A1(n39472), .A2(\pe5/aot [18]), .B1(n59427), .B2(
        \pe5/bq[2] ), .ZN(n48187) );
  NOR2HSV1 U51978 ( .A1(n48188), .A2(n48187), .ZN(n48189) );
  XOR2HSV0 U51979 ( .A1(n48190), .A2(n48189), .Z(n48191) );
  XNOR2HSV1 U51980 ( .A1(n48192), .A2(n48191), .ZN(n48214) );
  CLKNAND2HSV0 U51981 ( .A1(n59944), .A2(\pe5/bq[7] ), .ZN(n51386) );
  NOR2HSV0 U51982 ( .A1(n48193), .A2(n51386), .ZN(n48195) );
  AOI22HSV0 U51983 ( .A1(n52590), .A2(\pe5/bq[7] ), .B1(\pe5/bq[25] ), .B2(
        n59944), .ZN(n48194) );
  NOR2HSV2 U51984 ( .A1(n48195), .A2(n48194), .ZN(n48203) );
  NOR2HSV0 U51985 ( .A1(n48197), .A2(n48196), .ZN(n48201) );
  AOI22HSV0 U51986 ( .A1(n48199), .A2(n39471), .B1(n48198), .B2(n59866), .ZN(
        n48200) );
  NOR2HSV1 U51987 ( .A1(n48201), .A2(n48200), .ZN(n48202) );
  XOR2HSV0 U51988 ( .A1(n48203), .A2(n48202), .Z(n48212) );
  NOR2HSV0 U51989 ( .A1(n48204), .A2(n48031), .ZN(n51383) );
  AOI22HSV0 U51990 ( .A1(n48816), .A2(n51420), .B1(n48206), .B2(n48205), .ZN(
        n48207) );
  AOI21HSV0 U51991 ( .A1(n51383), .A2(n48208), .B(n48207), .ZN(n48210) );
  NOR2HSV0 U51992 ( .A1(n59641), .A2(n48822), .ZN(n48209) );
  XNOR2HSV1 U51993 ( .A1(n48210), .A2(n48209), .ZN(n48211) );
  XNOR2HSV1 U51994 ( .A1(n48212), .A2(n48211), .ZN(n48213) );
  XNOR2HSV1 U51995 ( .A1(n48214), .A2(n48213), .ZN(n48216) );
  NAND2HSV0 U51996 ( .A1(n39278), .A2(\pe5/got [1]), .ZN(n48215) );
  XNOR2HSV1 U51997 ( .A1(n48216), .A2(n48215), .ZN(n48217) );
  XNOR2HSV1 U51998 ( .A1(n48218), .A2(n48217), .ZN(n48258) );
  NAND2HSV0 U51999 ( .A1(n51313), .A2(n47291), .ZN(n48221) );
  CLKNHSV0 U52000 ( .I(n48219), .ZN(n48796) );
  NAND2HSV0 U52001 ( .A1(n48796), .A2(n51191), .ZN(n48220) );
  XOR2HSV0 U52002 ( .A1(n48221), .A2(n48220), .Z(n48225) );
  NAND2HSV0 U52003 ( .A1(\pe5/aot [13]), .A2(\pe5/bq[19] ), .ZN(n48223) );
  NAND2HSV0 U52004 ( .A1(n52600), .A2(n48755), .ZN(n48222) );
  XOR2HSV0 U52005 ( .A1(n48223), .A2(n48222), .Z(n48224) );
  XOR2HSV0 U52006 ( .A1(n48225), .A2(n48224), .Z(n48233) );
  NAND2HSV0 U52007 ( .A1(n52591), .A2(n31045), .ZN(n48227) );
  NAND2HSV0 U52008 ( .A1(n40234), .A2(n51177), .ZN(n48226) );
  XOR2HSV0 U52009 ( .A1(n48227), .A2(n48226), .Z(n48231) );
  NAND2HSV0 U52010 ( .A1(\pe5/aot [4]), .A2(n48802), .ZN(n48229) );
  NAND2HSV0 U52011 ( .A1(n53295), .A2(n30542), .ZN(n48228) );
  XOR2HSV0 U52012 ( .A1(n48229), .A2(n48228), .Z(n48230) );
  XOR2HSV0 U52013 ( .A1(n48231), .A2(n48230), .Z(n48232) );
  XOR2HSV0 U52014 ( .A1(n48233), .A2(n48232), .Z(n48254) );
  NAND2HSV0 U52015 ( .A1(n52675), .A2(n30341), .ZN(n48235) );
  NAND2HSV0 U52016 ( .A1(n52607), .A2(n50500), .ZN(n48234) );
  XOR2HSV0 U52017 ( .A1(n48235), .A2(n48234), .Z(n48241) );
  NAND2HSV0 U52018 ( .A1(n50505), .A2(n48236), .ZN(n48239) );
  NAND2HSV0 U52019 ( .A1(n52584), .A2(n48237), .ZN(n48238) );
  XOR2HSV0 U52020 ( .A1(n48239), .A2(n48238), .Z(n48240) );
  XOR2HSV0 U52021 ( .A1(n48241), .A2(n48240), .Z(n48252) );
  NAND2HSV0 U52022 ( .A1(n48242), .A2(\pe5/bq[11] ), .ZN(n48245) );
  NAND2HSV0 U52023 ( .A1(n48243), .A2(n48760), .ZN(n48244) );
  XOR2HSV0 U52024 ( .A1(n48245), .A2(n48244), .Z(n48250) );
  NOR2HSV0 U52025 ( .A1(n48246), .A2(n37564), .ZN(n48248) );
  NAND2HSV0 U52026 ( .A1(\pe5/aot [23]), .A2(n48775), .ZN(n48247) );
  XOR2HSV0 U52027 ( .A1(n48248), .A2(n48247), .Z(n48249) );
  XOR2HSV0 U52028 ( .A1(n48250), .A2(n48249), .Z(n48251) );
  XOR2HSV0 U52029 ( .A1(n48252), .A2(n48251), .Z(n48253) );
  XOR2HSV0 U52030 ( .A1(n48254), .A2(n48253), .Z(n48256) );
  NAND2HSV0 U52031 ( .A1(n30270), .A2(n59357), .ZN(n48255) );
  XNOR2HSV1 U52032 ( .A1(n48256), .A2(n48255), .ZN(n48257) );
  XNOR2HSV1 U52033 ( .A1(n48258), .A2(n48257), .ZN(n48259) );
  XNOR2HSV1 U52034 ( .A1(n48260), .A2(n48259), .ZN(n48261) );
  XNOR2HSV1 U52035 ( .A1(n48262), .A2(n48261), .ZN(n48263) );
  XNOR2HSV1 U52036 ( .A1(n48264), .A2(n48263), .ZN(n48266) );
  NAND2HSV0 U52037 ( .A1(n48848), .A2(n51159), .ZN(n48265) );
  XOR2HSV0 U52038 ( .A1(n48266), .A2(n48265), .Z(n48267) );
  XNOR2HSV1 U52039 ( .A1(n48268), .A2(n48267), .ZN(n48269) );
  XNOR2HSV1 U52040 ( .A1(n48270), .A2(n48269), .ZN(n48271) );
  XNOR2HSV1 U52041 ( .A1(n48272), .A2(n48271), .ZN(n48273) );
  XNOR2HSV1 U52042 ( .A1(n48274), .A2(n48273), .ZN(n48275) );
  XNOR2HSV1 U52043 ( .A1(n48276), .A2(n48275), .ZN(n48277) );
  XNOR2HSV1 U52044 ( .A1(n48278), .A2(n48277), .ZN(n48280) );
  NAND2HSV0 U52045 ( .A1(n30752), .A2(\pe5/got [14]), .ZN(n48279) );
  XOR2HSV0 U52046 ( .A1(n48280), .A2(n48279), .Z(n48281) );
  XNOR2HSV1 U52047 ( .A1(n48282), .A2(n48281), .ZN(n48284) );
  NAND2HSV0 U52048 ( .A1(n51205), .A2(n51224), .ZN(n48283) );
  XNOR2HSV1 U52049 ( .A1(n48284), .A2(n48283), .ZN(n48285) );
  XNOR2HSV1 U52050 ( .A1(n48286), .A2(n48285), .ZN(n48287) );
  XNOR2HSV1 U52051 ( .A1(n48288), .A2(n48287), .ZN(n48290) );
  NAND2HSV0 U52052 ( .A1(n52653), .A2(n39432), .ZN(n48289) );
  XNOR2HSV1 U52053 ( .A1(n48290), .A2(n48289), .ZN(n48291) );
  XNOR2HSV1 U52054 ( .A1(n48292), .A2(n48291), .ZN(n48293) );
  XNOR2HSV1 U52055 ( .A1(n48294), .A2(n48293), .ZN(n48295) );
  XNOR2HSV1 U52056 ( .A1(n48296), .A2(n48295), .ZN(n48297) );
  XNOR2HSV1 U52057 ( .A1(n48298), .A2(n48297), .ZN(n48300) );
  NAND2HSV0 U52058 ( .A1(n59516), .A2(n48743), .ZN(n48299) );
  XNOR2HSV1 U52059 ( .A1(n48300), .A2(n48299), .ZN(n48301) );
  XNOR2HSV1 U52060 ( .A1(n48302), .A2(n48301), .ZN(n48304) );
  XNOR2HSV1 U52061 ( .A1(n48304), .A2(n48303), .ZN(n48305) );
  XNOR2HSV1 U52062 ( .A1(n48306), .A2(n48305), .ZN(n48307) );
  CLKNHSV0 U52063 ( .I(n48477), .ZN(n59418) );
  CLKNHSV0 U52064 ( .I(n48477), .ZN(n59419) );
  CLKNHSV0 U52065 ( .I(n48312), .ZN(n48310) );
  CLKNAND2HSV1 U52066 ( .A1(n48315), .A2(n48314), .ZN(n48318) );
  CLKNAND2HSV0 U52067 ( .A1(n48315), .A2(n48314), .ZN(n48316) );
  AOI21HSV4 U52068 ( .A1(n48319), .A2(n48318), .B(n48317), .ZN(n48323) );
  NOR2HSV2 U52069 ( .A1(n48321), .A2(n48320), .ZN(n48322) );
  AOI21HSV4 U52070 ( .A1(n53368), .A2(n48323), .B(n48322), .ZN(n48465) );
  NOR2HSV4 U52071 ( .A1(n48325), .A2(n48324), .ZN(n48327) );
  CLKNAND2HSV2 U52072 ( .A1(n48327), .A2(n48326), .ZN(n48464) );
  AO21HSV1 U52073 ( .A1(n48332), .A2(n48331), .B(n40936), .Z(n48333) );
  CLKNAND2HSV0 U52074 ( .A1(n48336), .A2(\pe1/got [25]), .ZN(n48445) );
  NAND2HSV0 U52075 ( .A1(n55229), .A2(n53520), .ZN(n48443) );
  CLKNAND2HSV1 U52076 ( .A1(n53521), .A2(n53390), .ZN(n48439) );
  NOR2HSV1 U52077 ( .A1(n53391), .A2(n48337), .ZN(n48437) );
  CLKNAND2HSV1 U52078 ( .A1(n53522), .A2(\pe1/got [20]), .ZN(n48435) );
  CLKNAND2HSV1 U52079 ( .A1(n53392), .A2(\pe1/got [19]), .ZN(n48433) );
  NOR2HSV1 U52080 ( .A1(n54040), .A2(n54248), .ZN(n48431) );
  NAND2HSV0 U52081 ( .A1(n59518), .A2(n54161), .ZN(n48429) );
  CLKNAND2HSV1 U52082 ( .A1(n54600), .A2(n54135), .ZN(n48428) );
  NAND2HSV2 U52083 ( .A1(n59725), .A2(n48339), .ZN(n48426) );
  NAND2HSV0 U52084 ( .A1(n54041), .A2(\pe1/got [14]), .ZN(n48424) );
  NAND2HSV0 U52085 ( .A1(n41332), .A2(n53473), .ZN(n48417) );
  NAND2HSV0 U52086 ( .A1(n41144), .A2(n54894), .ZN(n48411) );
  CLKNAND2HSV0 U52087 ( .A1(n53795), .A2(n53523), .ZN(n48341) );
  CLKNAND2HSV0 U52088 ( .A1(n53979), .A2(n55475), .ZN(n48340) );
  XNOR2HSV1 U52089 ( .A1(n48341), .A2(n48340), .ZN(n48409) );
  NAND2HSV0 U52090 ( .A1(n40683), .A2(n55231), .ZN(n53446) );
  XOR2HSV0 U52091 ( .A1(n48342), .A2(n53446), .Z(n48346) );
  XOR2HSV0 U52092 ( .A1(n48344), .A2(n48343), .Z(n48345) );
  XOR2HSV0 U52093 ( .A1(n48346), .A2(n48345), .Z(n48355) );
  NOR2HSV0 U52094 ( .A1(n54901), .A2(n48347), .ZN(n48349) );
  NAND2HSV0 U52095 ( .A1(n55496), .A2(n25179), .ZN(n48348) );
  XOR2HSV0 U52096 ( .A1(n48349), .A2(n48348), .Z(n48353) );
  NAND2HSV0 U52097 ( .A1(n41153), .A2(n53798), .ZN(n48351) );
  NAND2HSV0 U52098 ( .A1(n54303), .A2(n41339), .ZN(n48350) );
  XOR2HSV0 U52099 ( .A1(n48351), .A2(n48350), .Z(n48352) );
  XOR2HSV0 U52100 ( .A1(n48353), .A2(n48352), .Z(n48354) );
  XOR2HSV0 U52101 ( .A1(n48355), .A2(n48354), .Z(n48407) );
  CLKNHSV0 U52102 ( .I(n54399), .ZN(n55491) );
  NAND2HSV0 U52103 ( .A1(n53673), .A2(n55491), .ZN(n48357) );
  NAND2HSV0 U52104 ( .A1(n25226), .A2(\pe1/bq[2] ), .ZN(n48356) );
  XOR2HSV0 U52105 ( .A1(n48357), .A2(n48356), .Z(n48361) );
  NAND2HSV0 U52106 ( .A1(n59619), .A2(n25428), .ZN(n48359) );
  CLKNHSV0 U52107 ( .I(n53957), .ZN(n53538) );
  CLKNAND2HSV0 U52108 ( .A1(n53538), .A2(n54289), .ZN(n48358) );
  XOR2HSV0 U52109 ( .A1(n48359), .A2(n48358), .Z(n48360) );
  XOR2HSV0 U52110 ( .A1(n48361), .A2(n48360), .Z(n48364) );
  NAND2HSV0 U52111 ( .A1(n59675), .A2(\pe1/got [3]), .ZN(n48362) );
  NAND2HSV0 U52112 ( .A1(n55595), .A2(n40684), .ZN(n53525) );
  XNOR2HSV1 U52113 ( .A1(n48362), .A2(n53525), .ZN(n48363) );
  XNOR2HSV1 U52114 ( .A1(n48364), .A2(n48363), .ZN(n48371) );
  NAND2HSV0 U52115 ( .A1(n41248), .A2(n53863), .ZN(n48369) );
  INHSV2 U52116 ( .I(n48365), .ZN(n48367) );
  XOR2HSV0 U52117 ( .A1(n48367), .A2(n48366), .Z(n48368) );
  XNOR2HSV1 U52118 ( .A1(n48369), .A2(n48368), .ZN(n48370) );
  XNOR2HSV1 U52119 ( .A1(n48371), .A2(n48370), .ZN(n48406) );
  NAND2HSV0 U52120 ( .A1(n53717), .A2(n53578), .ZN(n48373) );
  NAND2HSV0 U52121 ( .A1(\pe1/aot [16]), .A2(\pe1/bq[18] ), .ZN(n48372) );
  XOR2HSV0 U52122 ( .A1(n48373), .A2(n48372), .Z(n48377) );
  NAND2HSV0 U52123 ( .A1(\pe1/aot [24]), .A2(n55352), .ZN(n48375) );
  NAND2HSV0 U52124 ( .A1(n42132), .A2(n42092), .ZN(n48374) );
  XOR2HSV0 U52125 ( .A1(n48375), .A2(n48374), .Z(n48376) );
  XOR2HSV0 U52126 ( .A1(n48377), .A2(n48376), .Z(n48386) );
  NAND2HSV0 U52127 ( .A1(\pe1/aot [25]), .A2(\pe1/bq[9] ), .ZN(n48379) );
  NAND2HSV0 U52128 ( .A1(n59985), .A2(n54371), .ZN(n48378) );
  XOR2HSV0 U52129 ( .A1(n48379), .A2(n48378), .Z(n48384) );
  NAND2HSV0 U52130 ( .A1(n54078), .A2(n42373), .ZN(n48382) );
  CLKNHSV0 U52131 ( .I(n44705), .ZN(n54364) );
  NAND2HSV0 U52132 ( .A1(n54364), .A2(n48380), .ZN(n48381) );
  XOR2HSV0 U52133 ( .A1(n48382), .A2(n48381), .Z(n48383) );
  XOR2HSV0 U52134 ( .A1(n48384), .A2(n48383), .Z(n48385) );
  XOR2HSV0 U52135 ( .A1(n48386), .A2(n48385), .Z(n48404) );
  NAND2HSV0 U52136 ( .A1(n59987), .A2(n54179), .ZN(n48388) );
  NAND2HSV0 U52137 ( .A1(n54904), .A2(\pe1/bq[26] ), .ZN(n48387) );
  XOR2HSV0 U52138 ( .A1(n48388), .A2(n48387), .Z(n48392) );
  NAND2HSV0 U52139 ( .A1(n53936), .A2(n54048), .ZN(n48390) );
  NAND2HSV0 U52140 ( .A1(n59990), .A2(\pe1/bq[21] ), .ZN(n48389) );
  XOR2HSV0 U52141 ( .A1(n48390), .A2(n48389), .Z(n48391) );
  XOR2HSV0 U52142 ( .A1(n48392), .A2(n48391), .Z(n48402) );
  NOR2HSV0 U52143 ( .A1(n54672), .A2(n48393), .ZN(n48395) );
  NAND2HSV0 U52144 ( .A1(\pe1/aot [20]), .A2(n53571), .ZN(n48394) );
  XOR2HSV0 U52145 ( .A1(n48395), .A2(n48394), .Z(n48400) );
  NAND2HSV0 U52146 ( .A1(n54978), .A2(n42366), .ZN(n48398) );
  NAND2HSV0 U52147 ( .A1(n48396), .A2(n54995), .ZN(n48397) );
  XOR2HSV0 U52148 ( .A1(n48398), .A2(n48397), .Z(n48399) );
  XOR2HSV0 U52149 ( .A1(n48400), .A2(n48399), .Z(n48401) );
  XOR2HSV0 U52150 ( .A1(n48402), .A2(n48401), .Z(n48403) );
  XOR2HSV0 U52151 ( .A1(n48404), .A2(n48403), .Z(n48405) );
  XOR3HSV2 U52152 ( .A1(n48407), .A2(n48406), .A3(n48405), .Z(n48408) );
  XNOR2HSV1 U52153 ( .A1(n48409), .A2(n48408), .ZN(n48410) );
  XNOR2HSV1 U52154 ( .A1(n48411), .A2(n48410), .ZN(n48413) );
  NAND2HSV0 U52155 ( .A1(n53602), .A2(n55339), .ZN(n48412) );
  XOR2HSV0 U52156 ( .A1(n48413), .A2(n48412), .Z(n48415) );
  NAND2HSV0 U52157 ( .A1(n54265), .A2(\pe1/got [9]), .ZN(n48414) );
  XOR2HSV0 U52158 ( .A1(n48415), .A2(n48414), .Z(n48416) );
  XNOR2HSV1 U52159 ( .A1(n48417), .A2(n48416), .ZN(n48419) );
  NAND2HSV0 U52160 ( .A1(n29773), .A2(n54970), .ZN(n48418) );
  XOR2HSV0 U52161 ( .A1(n48419), .A2(n48418), .Z(n48422) );
  NOR2HSV2 U52162 ( .A1(n41566), .A2(n54453), .ZN(n48421) );
  NAND2HSV0 U52163 ( .A1(n54115), .A2(n54812), .ZN(n48420) );
  XOR3HSV2 U52164 ( .A1(n48422), .A2(n48421), .A3(n48420), .Z(n48423) );
  XNOR2HSV1 U52165 ( .A1(n48424), .A2(n48423), .ZN(n48425) );
  XOR2HSV0 U52166 ( .A1(n48426), .A2(n48425), .Z(n48427) );
  XOR3HSV2 U52167 ( .A1(n48429), .A2(n48428), .A3(n48427), .Z(n48430) );
  XOR2HSV0 U52168 ( .A1(n48431), .A2(n48430), .Z(n48432) );
  XNOR2HSV1 U52169 ( .A1(n48433), .A2(n48432), .ZN(n48434) );
  XNOR2HSV1 U52170 ( .A1(n48435), .A2(n48434), .ZN(n48436) );
  XOR2HSV0 U52171 ( .A1(n48437), .A2(n48436), .Z(n48438) );
  XNOR2HSV1 U52172 ( .A1(n48439), .A2(n48438), .ZN(n48441) );
  CLKNAND2HSV0 U52173 ( .A1(n53768), .A2(n41298), .ZN(n48440) );
  XOR2HSV0 U52174 ( .A1(n48441), .A2(n48440), .Z(n48442) );
  XOR2HSV0 U52175 ( .A1(n48443), .A2(n48442), .Z(n48444) );
  XOR2HSV0 U52176 ( .A1(n48445), .A2(n48444), .Z(n48447) );
  CLKNAND2HSV1 U52177 ( .A1(n54541), .A2(\pe1/got [26]), .ZN(n48446) );
  XNOR2HSV1 U52178 ( .A1(n48447), .A2(n48446), .ZN(n48448) );
  XNOR2HSV4 U52179 ( .A1(n48449), .A2(n48448), .ZN(n48455) );
  NOR2HSV0 U52180 ( .A1(n48451), .A2(n48450), .ZN(n48452) );
  INHSV2 U52181 ( .I(n48452), .ZN(n48454) );
  OAI21HSV4 U52182 ( .A1(n48455), .A2(n48454), .B(n48453), .ZN(n48458) );
  XNOR2HSV4 U52183 ( .A1(n48458), .A2(n48457), .ZN(n48460) );
  CLKNHSV2 U52184 ( .I(n48459), .ZN(n48462) );
  INHSV3 U52185 ( .I(n48460), .ZN(n48461) );
  CLKNHSV0 U52186 ( .I(n54631), .ZN(n59520) );
  CLKNHSV0 U52187 ( .I(n48083), .ZN(n59429) );
  CLKNHSV0 U52188 ( .I(n48083), .ZN(n59430) );
  CLKNHSV0 U52189 ( .I(n48479), .ZN(n59431) );
  CLKNHSV0 U52190 ( .I(n48477), .ZN(n59432) );
  CLKNHSV0 U52191 ( .I(n48083), .ZN(n59435) );
  CLKNHSV0 U52192 ( .I(n48472), .ZN(n59436) );
  CLKNHSV0 U52193 ( .I(n48472), .ZN(n59437) );
  CLKNHSV0 U52194 ( .I(n59660), .ZN(n59438) );
  CLKNHSV0 U52195 ( .I(n48479), .ZN(n59439) );
  CLKNHSV0 U52196 ( .I(n48083), .ZN(n59440) );
  CLKNHSV0 U52197 ( .I(n48478), .ZN(n59442) );
  CLKNHSV0 U52198 ( .I(n48478), .ZN(n59444) );
  CLKNHSV0 U52199 ( .I(n48083), .ZN(n59445) );
  CLKNHSV0 U52200 ( .I(n48472), .ZN(n59446) );
  CLKNHSV0 U52201 ( .I(n48083), .ZN(n59447) );
  CLKNHSV0 U52202 ( .I(n48083), .ZN(n59448) );
  CLKNHSV0 U52203 ( .I(n48476), .ZN(n59449) );
  BUFHSV2 U52204 ( .I(n59397), .Z(n59923) );
  CLKNHSV0 U52205 ( .I(n48472), .ZN(n59476) );
  CLKNHSV0 U52206 ( .I(n48015), .ZN(n59451) );
  CLKNHSV0 U52207 ( .I(n48477), .ZN(n59452) );
  CLKNHSV0 U52208 ( .I(n48015), .ZN(n59453) );
  CLKNHSV0 U52209 ( .I(n59404), .ZN(n48474) );
  CLKNHSV0 U52210 ( .I(n48083), .ZN(n59454) );
  CLKNHSV0 U52211 ( .I(n48479), .ZN(n59455) );
  CLKNHSV0 U52212 ( .I(n48479), .ZN(n59456) );
  CLKNHSV0 U52213 ( .I(n48477), .ZN(n59457) );
  CLKNHSV0 U52214 ( .I(n48478), .ZN(n59458) );
  CLKNHSV0 U52215 ( .I(n59660), .ZN(n59459) );
  CLKNHSV0 U52216 ( .I(n48083), .ZN(n59460) );
  CLKNHSV0 U52217 ( .I(n48015), .ZN(n59461) );
  CLKNHSV0 U52218 ( .I(n48478), .ZN(n59462) );
  CLKNHSV0 U52219 ( .I(n48472), .ZN(n59463) );
  CLKNHSV0 U52220 ( .I(n59660), .ZN(n59464) );
  CLKNHSV0 U52221 ( .I(n48478), .ZN(n59465) );
  CLKNHSV0 U52222 ( .I(n48478), .ZN(n59466) );
  CLKNHSV0 U52223 ( .I(n59660), .ZN(n59467) );
  CLKNHSV0 U52224 ( .I(n48479), .ZN(n59469) );
  CLKNHSV0 U52225 ( .I(n48478), .ZN(n59470) );
  CLKNHSV0 U52226 ( .I(n59660), .ZN(n59471) );
  CLKNHSV0 U52227 ( .I(n48083), .ZN(n59472) );
  CLKNHSV0 U52228 ( .I(n48015), .ZN(n59473) );
  CLKNHSV0 U52229 ( .I(n48474), .ZN(n59474) );
  CLKNHSV0 U52230 ( .I(n48472), .ZN(n59477) );
  CLKNHSV0 U52231 ( .I(n48478), .ZN(n59478) );
  CLKNHSV0 U52232 ( .I(n48478), .ZN(n59479) );
  CLKNHSV0 U52233 ( .I(n48477), .ZN(n59480) );
  CLKNHSV0 U52234 ( .I(n48479), .ZN(n59481) );
  CLKNHSV0 U52235 ( .I(n48479), .ZN(n59482) );
  CLKNHSV0 U52236 ( .I(n48479), .ZN(n59483) );
  CLKNHSV0 U52237 ( .I(n59660), .ZN(n59484) );
  BUFHSV2 U52238 ( .I(n59925), .Z(n59655) );
  INAND2HSV2 U52239 ( .A1(n43873), .B1(n56935), .ZN(n48615) );
  INHSV2 U52240 ( .I(n51118), .ZN(n56339) );
  CLKNAND2HSV1 U52241 ( .A1(n56339), .A2(n55940), .ZN(n48613) );
  CLKNAND2HSV0 U52242 ( .A1(n56780), .A2(n36958), .ZN(n48611) );
  CLKNAND2HSV1 U52243 ( .A1(n48481), .A2(n36955), .ZN(n48609) );
  CLKNAND2HSV0 U52244 ( .A1(n55946), .A2(n46441), .ZN(n48607) );
  CLKNAND2HSV0 U52245 ( .A1(n48482), .A2(n43452), .ZN(n48605) );
  INAND2HSV2 U52246 ( .A1(n48484), .B1(n48483), .ZN(n48603) );
  CLKNAND2HSV0 U52247 ( .A1(n48486), .A2(n48485), .ZN(n48601) );
  NAND2HSV0 U52248 ( .A1(n56265), .A2(n43262), .ZN(n48599) );
  CLKNAND2HSV0 U52249 ( .A1(n59500), .A2(n42996), .ZN(n48597) );
  CLKNAND2HSV0 U52250 ( .A1(n43754), .A2(\pe3/got [18]), .ZN(n48593) );
  NAND2HSV0 U52251 ( .A1(n56178), .A2(n56335), .ZN(n48589) );
  NAND2HSV0 U52252 ( .A1(n43755), .A2(n59967), .ZN(n48579) );
  NAND2HSV0 U52253 ( .A1(n56179), .A2(n59644), .ZN(n48577) );
  NAND2HSV0 U52254 ( .A1(n56180), .A2(n59645), .ZN(n48575) );
  NAND2HSV0 U52255 ( .A1(n56070), .A2(n56241), .ZN(n48571) );
  NAND2HSV0 U52256 ( .A1(n59626), .A2(n48487), .ZN(n48569) );
  NAND2HSV0 U52257 ( .A1(n48488), .A2(n59799), .ZN(n48567) );
  NAND2HSV0 U52258 ( .A1(n37017), .A2(n55950), .ZN(n48510) );
  NAND2HSV0 U52259 ( .A1(\pe3/aot [6]), .A2(\pe3/bq[26] ), .ZN(n48490) );
  NAND2HSV0 U52260 ( .A1(n59808), .A2(\pe3/bq[23] ), .ZN(n48489) );
  XOR2HSV0 U52261 ( .A1(n48490), .A2(n48489), .Z(n48494) );
  NAND2HSV0 U52262 ( .A1(\pe3/aot [16]), .A2(n56640), .ZN(n48492) );
  NAND2HSV0 U52263 ( .A1(n56197), .A2(n56218), .ZN(n48491) );
  XOR2HSV0 U52264 ( .A1(n48492), .A2(n48491), .Z(n48493) );
  XOR2HSV0 U52265 ( .A1(n48494), .A2(n48493), .Z(n48506) );
  NAND2HSV0 U52266 ( .A1(\pe3/aot [22]), .A2(n56187), .ZN(n48498) );
  CLKNHSV0 U52267 ( .I(n48495), .ZN(n56505) );
  NAND2HSV0 U52268 ( .A1(n48496), .A2(n56505), .ZN(n48497) );
  XOR2HSV0 U52269 ( .A1(n48498), .A2(n48497), .Z(n48504) );
  NAND2HSV0 U52270 ( .A1(n56349), .A2(n48499), .ZN(n48502) );
  NAND2HSV0 U52271 ( .A1(n48500), .A2(\pe3/bq[3] ), .ZN(n48501) );
  XOR2HSV0 U52272 ( .A1(n48502), .A2(n48501), .Z(n48503) );
  XOR2HSV0 U52273 ( .A1(n48504), .A2(n48503), .Z(n48505) );
  XOR2HSV0 U52274 ( .A1(n48506), .A2(n48505), .Z(n48508) );
  NAND2HSV0 U52275 ( .A1(n59648), .A2(n56975), .ZN(n48507) );
  XNOR2HSV1 U52276 ( .A1(n48508), .A2(n48507), .ZN(n48509) );
  XNOR2HSV1 U52277 ( .A1(n48510), .A2(n48509), .ZN(n48565) );
  NAND2HSV0 U52278 ( .A1(n48511), .A2(n56823), .ZN(n48562) );
  NAND2HSV0 U52279 ( .A1(n59646), .A2(\pe3/bq[19] ), .ZN(n49282) );
  NOR2HSV0 U52280 ( .A1(n48512), .A2(n49282), .ZN(n48514) );
  AOI22HSV0 U52281 ( .A1(n53249), .A2(\pe3/bq[19] ), .B1(n55867), .B2(n59646), 
        .ZN(n48513) );
  NOR2HSV2 U52282 ( .A1(n48514), .A2(n48513), .ZN(n48519) );
  NAND2HSV0 U52283 ( .A1(n42743), .A2(n55857), .ZN(n55986) );
  NOR2HSV0 U52284 ( .A1(n48515), .A2(n55986), .ZN(n48517) );
  AOI22HSV0 U52285 ( .A1(n43265), .A2(n56971), .B1(\pe3/aot [26]), .B2(n56272), 
        .ZN(n48516) );
  NOR2HSV2 U52286 ( .A1(n48517), .A2(n48516), .ZN(n48518) );
  XNOR2HSV1 U52287 ( .A1(n48519), .A2(n48518), .ZN(n48526) );
  NAND2HSV0 U52288 ( .A1(n59961), .A2(n48520), .ZN(n49420) );
  XNOR2HSV0 U52289 ( .A1(n48524), .A2(n48523), .ZN(n48525) );
  XNOR2HSV1 U52290 ( .A1(n48526), .A2(n48525), .ZN(n48560) );
  NAND2HSV0 U52291 ( .A1(\pe3/aot [5]), .A2(n55960), .ZN(n48529) );
  NAND2HSV0 U52292 ( .A1(n56434), .A2(n48527), .ZN(n48528) );
  XOR2HSV0 U52293 ( .A1(n48529), .A2(n48528), .Z(n48534) );
  NOR2HSV0 U52294 ( .A1(n47447), .A2(n37196), .ZN(n48532) );
  NAND2HSV0 U52295 ( .A1(n48530), .A2(\pe3/bq[7] ), .ZN(n48531) );
  XOR2HSV0 U52296 ( .A1(n48532), .A2(n48531), .Z(n48533) );
  XNOR2HSV1 U52297 ( .A1(n48534), .A2(n48533), .ZN(n48544) );
  NOR2HSV0 U52298 ( .A1(n53229), .A2(n56914), .ZN(n56633) );
  AOI22HSV0 U52299 ( .A1(n55987), .A2(n56428), .B1(n42971), .B2(n56575), .ZN(
        n48535) );
  AOI21HSV0 U52300 ( .A1(n48536), .A2(n56633), .B(n48535), .ZN(n48542) );
  NAND2HSV0 U52301 ( .A1(n56970), .A2(n43052), .ZN(n55651) );
  NOR2HSV0 U52302 ( .A1(n48537), .A2(n55651), .ZN(n48540) );
  AOI22HSV0 U52303 ( .A1(\pe3/aot [8]), .A2(n42530), .B1(n48538), .B2(n56970), 
        .ZN(n48539) );
  NOR2HSV1 U52304 ( .A1(n48540), .A2(n48539), .ZN(n48541) );
  XOR2HSV0 U52305 ( .A1(n48542), .A2(n48541), .Z(n48543) );
  XNOR2HSV1 U52306 ( .A1(n48544), .A2(n48543), .ZN(n48559) );
  NAND2HSV0 U52307 ( .A1(n56204), .A2(n56507), .ZN(n48547) );
  NAND2HSV0 U52308 ( .A1(\pe3/aot [19]), .A2(n55975), .ZN(n48546) );
  XOR2HSV0 U52309 ( .A1(n48547), .A2(n48546), .Z(n48551) );
  NAND2HSV0 U52310 ( .A1(n56087), .A2(n55970), .ZN(n48549) );
  NAND2HSV0 U52311 ( .A1(\pe3/aot [14]), .A2(n55727), .ZN(n48548) );
  XOR2HSV0 U52312 ( .A1(n48549), .A2(n48548), .Z(n48550) );
  XOR2HSV0 U52313 ( .A1(n48551), .A2(n48550), .Z(n48557) );
  NAND2HSV0 U52314 ( .A1(n42818), .A2(n56785), .ZN(n56114) );
  NAND2HSV0 U52315 ( .A1(n55750), .A2(\pe3/bq[4] ), .ZN(n55859) );
  XOR2HSV0 U52316 ( .A1(n56114), .A2(n55859), .Z(n48555) );
  NAND2HSV0 U52317 ( .A1(n55864), .A2(n55616), .ZN(n48552) );
  XOR2HSV0 U52318 ( .A1(n48553), .A2(n48552), .Z(n48554) );
  XOR2HSV0 U52319 ( .A1(n48555), .A2(n48554), .Z(n48556) );
  XOR2HSV0 U52320 ( .A1(n48557), .A2(n48556), .Z(n48558) );
  XOR3HSV2 U52321 ( .A1(n48560), .A2(n48559), .A3(n48558), .Z(n48561) );
  XNOR2HSV1 U52322 ( .A1(n48562), .A2(n48561), .ZN(n48564) );
  NAND2HSV0 U52323 ( .A1(n37316), .A2(n56068), .ZN(n48563) );
  XOR3HSV2 U52324 ( .A1(n48565), .A2(n48564), .A3(n48563), .Z(n48566) );
  XNOR2HSV1 U52325 ( .A1(n48567), .A2(n48566), .ZN(n48568) );
  XNOR2HSV1 U52326 ( .A1(n48569), .A2(n48568), .ZN(n48570) );
  XNOR2HSV1 U52327 ( .A1(n48571), .A2(n48570), .ZN(n48573) );
  NAND2HSV0 U52328 ( .A1(n55895), .A2(n56855), .ZN(n48572) );
  XNOR2HSV1 U52329 ( .A1(n48573), .A2(n48572), .ZN(n48574) );
  XNOR2HSV1 U52330 ( .A1(n48575), .A2(n48574), .ZN(n48576) );
  XNOR2HSV1 U52331 ( .A1(n48577), .A2(n48576), .ZN(n48578) );
  XNOR2HSV1 U52332 ( .A1(n48579), .A2(n48578), .ZN(n48582) );
  NOR2HSV0 U52333 ( .A1(n56391), .A2(n50802), .ZN(n48581) );
  NAND2HSV0 U52334 ( .A1(n56421), .A2(n56392), .ZN(n48580) );
  XOR3HSV1 U52335 ( .A1(n48582), .A2(n48581), .A3(n48580), .Z(n48587) );
  NOR2HSV1 U52336 ( .A1(n48583), .A2(n46042), .ZN(n48586) );
  NAND2HSV0 U52337 ( .A1(n56396), .A2(n48584), .ZN(n48585) );
  XOR3HSV2 U52338 ( .A1(n48587), .A2(n48586), .A3(n48585), .Z(n48588) );
  XNOR2HSV1 U52339 ( .A1(n48589), .A2(n48588), .ZN(n48591) );
  NAND2HSV0 U52340 ( .A1(n55912), .A2(n56065), .ZN(n48590) );
  XNOR2HSV1 U52341 ( .A1(n48591), .A2(n48590), .ZN(n48592) );
  XNOR2HSV1 U52342 ( .A1(n48593), .A2(n48592), .ZN(n48595) );
  NOR2HSV0 U52343 ( .A1(n56406), .A2(n49250), .ZN(n48594) );
  XNOR2HSV1 U52344 ( .A1(n48595), .A2(n48594), .ZN(n48596) );
  XNOR2HSV1 U52345 ( .A1(n48597), .A2(n48596), .ZN(n48598) );
  XNOR2HSV1 U52346 ( .A1(n48599), .A2(n48598), .ZN(n48600) );
  XNOR2HSV1 U52347 ( .A1(n48601), .A2(n48600), .ZN(n48602) );
  XNOR2HSV1 U52348 ( .A1(n48603), .A2(n48602), .ZN(n48604) );
  XNOR2HSV1 U52349 ( .A1(n48605), .A2(n48604), .ZN(n48606) );
  XNOR2HSV1 U52350 ( .A1(n48607), .A2(n48606), .ZN(n48608) );
  XNOR2HSV1 U52351 ( .A1(n48613), .A2(n48612), .ZN(n48614) );
  XOR2HSV0 U52352 ( .A1(n48615), .A2(n48614), .Z(n48618) );
  CLKNAND2HSV2 U52353 ( .A1(n56948), .A2(n42815), .ZN(n48617) );
  CLKAND2HSV1 U52354 ( .A1(n56490), .A2(n29750), .Z(n48616) );
  XOR3HSV2 U52355 ( .A1(n48618), .A2(n48617), .A3(n48616), .Z(\pe3/poht [1])
         );
  NAND2HSV2 U52356 ( .A1(\pe2/aot [2]), .A2(n51803), .ZN(n50917) );
  NAND2HSV2 U52357 ( .A1(n52056), .A2(n51614), .ZN(n51813) );
  CLKNAND2HSV0 U52358 ( .A1(n53291), .A2(n48744), .ZN(n48736) );
  NOR2HSV0 U52359 ( .A1(n51361), .A2(n30686), .ZN(n48731) );
  NAND2HSV0 U52360 ( .A1(n48747), .A2(n51224), .ZN(n48726) );
  NAND2HSV0 U52361 ( .A1(n52572), .A2(n52652), .ZN(n48721) );
  NAND2HSV0 U52362 ( .A1(n51160), .A2(n48167), .ZN(n48717) );
  NAND2HSV0 U52363 ( .A1(n52574), .A2(n51305), .ZN(n48715) );
  NAND2HSV0 U52364 ( .A1(n48748), .A2(n50424), .ZN(n48713) );
  NAND2HSV0 U52365 ( .A1(n29770), .A2(n52641), .ZN(n48711) );
  NAND2HSV0 U52366 ( .A1(n48624), .A2(n50698), .ZN(n48709) );
  NAND2HSV0 U52367 ( .A1(n52580), .A2(n51159), .ZN(n48707) );
  NAND2HSV0 U52368 ( .A1(n48750), .A2(n48841), .ZN(n48703) );
  NAND2HSV0 U52369 ( .A1(n30515), .A2(n51302), .ZN(n48701) );
  NAND2HSV0 U52370 ( .A1(n30255), .A2(n51331), .ZN(n48699) );
  NAND2HSV0 U52371 ( .A1(n30270), .A2(n51362), .ZN(n48697) );
  NAND2HSV0 U52372 ( .A1(n48751), .A2(n51161), .ZN(n48696) );
  NAND2HSV0 U52373 ( .A1(\pe5/aot [13]), .A2(n51167), .ZN(n48627) );
  NAND2HSV0 U52374 ( .A1(\pe5/aot [16]), .A2(n50500), .ZN(n48626) );
  XOR2HSV0 U52375 ( .A1(n48627), .A2(n48626), .Z(n48631) );
  NAND2HSV0 U52376 ( .A1(n52611), .A2(n48237), .ZN(n48629) );
  NAND2HSV0 U52377 ( .A1(\pe5/aot [18]), .A2(n50668), .ZN(n48628) );
  XOR2HSV0 U52378 ( .A1(n48629), .A2(n48628), .Z(n48630) );
  XOR2HSV0 U52379 ( .A1(n48631), .A2(n48630), .Z(n48640) );
  NAND2HSV0 U52380 ( .A1(n40234), .A2(n48764), .ZN(n48633) );
  NAND2HSV0 U52381 ( .A1(\pe5/aot [8]), .A2(n47305), .ZN(n48632) );
  XOR2HSV0 U52382 ( .A1(n48633), .A2(n48632), .Z(n48638) );
  NAND2HSV0 U52383 ( .A1(n48634), .A2(n51191), .ZN(n48636) );
  NAND2HSV0 U52384 ( .A1(n50505), .A2(n52610), .ZN(n48635) );
  XOR2HSV0 U52385 ( .A1(n48636), .A2(n48635), .Z(n48637) );
  XOR2HSV0 U52386 ( .A1(n48638), .A2(n48637), .Z(n48639) );
  XOR2HSV0 U52387 ( .A1(n48640), .A2(n48639), .Z(n48656) );
  NAND2HSV0 U52388 ( .A1(n52607), .A2(n52632), .ZN(n48642) );
  NAND2HSV0 U52389 ( .A1(n51313), .A2(n39445), .ZN(n48641) );
  XOR2HSV0 U52390 ( .A1(n48642), .A2(n48641), .Z(n48646) );
  NAND2HSV0 U52391 ( .A1(n51188), .A2(n48775), .ZN(n48644) );
  NAND2HSV0 U52392 ( .A1(n30788), .A2(\pe5/bq[11] ), .ZN(n48643) );
  XOR2HSV0 U52393 ( .A1(n48644), .A2(n48643), .Z(n48645) );
  XOR2HSV0 U52394 ( .A1(n48646), .A2(n48645), .Z(n48654) );
  NAND2HSV0 U52395 ( .A1(n48829), .A2(n51177), .ZN(n48648) );
  NAND2HSV0 U52396 ( .A1(n48199), .A2(n31045), .ZN(n48647) );
  XOR2HSV0 U52397 ( .A1(n48648), .A2(n48647), .Z(n48652) );
  NAND2HSV0 U52398 ( .A1(n52600), .A2(n48802), .ZN(n48650) );
  NAND2HSV0 U52399 ( .A1(\pe5/aot [23]), .A2(n52672), .ZN(n48649) );
  XOR2HSV0 U52400 ( .A1(n48650), .A2(n48649), .Z(n48651) );
  XOR2HSV0 U52401 ( .A1(n48652), .A2(n48651), .Z(n48653) );
  XOR2HSV0 U52402 ( .A1(n48654), .A2(n48653), .Z(n48655) );
  XOR2HSV0 U52403 ( .A1(n48656), .A2(n48655), .Z(n48694) );
  NAND2HSV0 U52404 ( .A1(n51182), .A2(\pe5/bq[19] ), .ZN(n50516) );
  NOR2HSV0 U52405 ( .A1(n48657), .A2(n50516), .ZN(n48660) );
  AOI22HSV0 U52406 ( .A1(n48658), .A2(n39454), .B1(n48804), .B2(n51182), .ZN(
        n48659) );
  NOR2HSV1 U52407 ( .A1(n48660), .A2(n48659), .ZN(n48673) );
  NOR2HSV0 U52408 ( .A1(n48246), .A2(n45844), .ZN(n48662) );
  INAND2HSV2 U52409 ( .A1(n39123), .B1(\pe5/bq[1] ), .ZN(n48661) );
  XOR2HSV0 U52410 ( .A1(n48662), .A2(n48661), .Z(n48672) );
  NAND2HSV2 U52411 ( .A1(n59944), .A2(\pe5/bq[2] ), .ZN(n52681) );
  NAND2HSV0 U52412 ( .A1(n48663), .A2(\pe5/bq[2] ), .ZN(n48814) );
  OAI21HSV0 U52413 ( .A1(n47230), .A2(n30452), .B(n48814), .ZN(n48664) );
  OAI21HSV0 U52414 ( .A1(n52681), .A2(n48665), .B(n48664), .ZN(n48670) );
  NAND2HSV2 U52415 ( .A1(n48786), .A2(n48778), .ZN(n51289) );
  NOR2HSV0 U52416 ( .A1(n48666), .A2(n51289), .ZN(n48668) );
  AOI22HSV0 U52417 ( .A1(\pe5/aot [21]), .A2(\pe5/bq[10] ), .B1(n48755), .B2(
        n51419), .ZN(n48667) );
  NOR2HSV1 U52418 ( .A1(n48668), .A2(n48667), .ZN(n48669) );
  XOR2HSV0 U52419 ( .A1(n48670), .A2(n48669), .Z(n48671) );
  XOR3HSV2 U52420 ( .A1(n48673), .A2(n48672), .A3(n48671), .Z(n48692) );
  CLKNHSV0 U52421 ( .I(n48674), .ZN(n48678) );
  AOI21HSV0 U52422 ( .A1(n50501), .A2(\pe5/bq[27] ), .B(n48675), .ZN(n48676)
         );
  AOI21HSV2 U52423 ( .A1(n48678), .A2(n48677), .B(n48676), .ZN(n48685) );
  NOR2HSV0 U52424 ( .A1(n48680), .A2(n48679), .ZN(n48683) );
  AOI22HSV0 U52425 ( .A1(n48681), .A2(n51041), .B1(n52585), .B2(n51310), .ZN(
        n48682) );
  NOR2HSV1 U52426 ( .A1(n48683), .A2(n48682), .ZN(n48684) );
  XNOR2HSV1 U52427 ( .A1(n48685), .A2(n48684), .ZN(n48690) );
  NAND2HSV0 U52428 ( .A1(n48796), .A2(n48686), .ZN(n48688) );
  NAND2HSV0 U52429 ( .A1(n37660), .A2(\pe5/bq[7] ), .ZN(n48687) );
  XOR2HSV0 U52430 ( .A1(n48688), .A2(n48687), .Z(n48689) );
  XNOR2HSV1 U52431 ( .A1(n48690), .A2(n48689), .ZN(n48691) );
  XNOR2HSV1 U52432 ( .A1(n48692), .A2(n48691), .ZN(n48693) );
  XNOR2HSV1 U52433 ( .A1(n48694), .A2(n48693), .ZN(n48695) );
  XOR3HSV1 U52434 ( .A1(n48697), .A2(n48696), .A3(n48695), .Z(n48698) );
  XNOR2HSV1 U52435 ( .A1(n48699), .A2(n48698), .ZN(n48700) );
  XNOR2HSV1 U52436 ( .A1(n48701), .A2(n48700), .ZN(n48702) );
  XNOR2HSV1 U52437 ( .A1(n48703), .A2(n48702), .ZN(n48705) );
  NAND2HSV0 U52438 ( .A1(n48848), .A2(n51200), .ZN(n48704) );
  XOR2HSV0 U52439 ( .A1(n48705), .A2(n48704), .Z(n48706) );
  XNOR2HSV1 U52440 ( .A1(n48707), .A2(n48706), .ZN(n48708) );
  XNOR2HSV1 U52441 ( .A1(n48709), .A2(n48708), .ZN(n48710) );
  XNOR2HSV1 U52442 ( .A1(n48711), .A2(n48710), .ZN(n48712) );
  XNOR2HSV1 U52443 ( .A1(n48713), .A2(n48712), .ZN(n48714) );
  XNOR2HSV1 U52444 ( .A1(n48715), .A2(n48714), .ZN(n48716) );
  XNOR2HSV1 U52445 ( .A1(n48717), .A2(n48716), .ZN(n48719) );
  NAND2HSV0 U52446 ( .A1(n44694), .A2(n52568), .ZN(n48718) );
  XOR2HSV0 U52447 ( .A1(n48719), .A2(n48718), .Z(n48720) );
  XNOR2HSV1 U52448 ( .A1(n48721), .A2(n48720), .ZN(n48724) );
  NOR2HSV0 U52449 ( .A1(n50617), .A2(n48722), .ZN(n48723) );
  XNOR2HSV1 U52450 ( .A1(n48724), .A2(n48723), .ZN(n48725) );
  XNOR2HSV1 U52451 ( .A1(n48726), .A2(n48725), .ZN(n48729) );
  CLKNAND2HSV1 U52452 ( .A1(n52569), .A2(n51156), .ZN(n48728) );
  NAND2HSV0 U52453 ( .A1(n51211), .A2(n52566), .ZN(n48727) );
  XOR3HSV2 U52454 ( .A1(n48729), .A2(n48728), .A3(n48727), .Z(n48730) );
  XNOR2HSV1 U52455 ( .A1(n48731), .A2(n48730), .ZN(n48734) );
  NOR2HSV1 U52456 ( .A1(n51217), .A2(n39119), .ZN(n48733) );
  NOR2HSV1 U52457 ( .A1(n52659), .A2(n30516), .ZN(n48732) );
  XOR3HSV2 U52458 ( .A1(n48734), .A2(n48733), .A3(n48732), .Z(n48735) );
  XNOR2HSV1 U52459 ( .A1(n48736), .A2(n48735), .ZN(n48738) );
  NAND2HSV0 U52460 ( .A1(\pe5/got [23]), .A2(n53344), .ZN(n48737) );
  CLKNAND2HSV0 U52461 ( .A1(n51016), .A2(n48743), .ZN(n48882) );
  NOR2HSV0 U52462 ( .A1(n50692), .A2(n39743), .ZN(n48880) );
  NAND2HSV0 U52463 ( .A1(n48745), .A2(n48744), .ZN(n48878) );
  NOR2HSV0 U52464 ( .A1(n51361), .A2(n30516), .ZN(n48876) );
  NAND2HSV0 U52465 ( .A1(n48746), .A2(n51103), .ZN(n48872) );
  NAND2HSV0 U52466 ( .A1(n48747), .A2(n52566), .ZN(n48870) );
  NAND2HSV0 U52467 ( .A1(n51018), .A2(n51224), .ZN(n48866) );
  NAND2HSV0 U52468 ( .A1(n51160), .A2(n52652), .ZN(n48862) );
  NAND2HSV0 U52469 ( .A1(n52574), .A2(n52568), .ZN(n48860) );
  NAND2HSV0 U52470 ( .A1(n48748), .A2(n48167), .ZN(n48858) );
  NAND2HSV0 U52471 ( .A1(n39745), .A2(n48749), .ZN(n48856) );
  NAND2HSV2 U52472 ( .A1(n51162), .A2(n50424), .ZN(n48854) );
  NAND2HSV0 U52473 ( .A1(n52580), .A2(n52641), .ZN(n48852) );
  NAND2HSV0 U52474 ( .A1(n48750), .A2(n51159), .ZN(n48847) );
  NAND2HSV0 U52475 ( .A1(n37659), .A2(n51200), .ZN(n48845) );
  NAND2HSV0 U52476 ( .A1(n48751), .A2(n51302), .ZN(n48840) );
  NAND2HSV0 U52477 ( .A1(n59944), .A2(n30222), .ZN(n48754) );
  NAND2HSV0 U52478 ( .A1(\pe5/got [1]), .A2(n48752), .ZN(n48753) );
  XOR2HSV0 U52479 ( .A1(n48754), .A2(n48753), .Z(n48759) );
  NAND2HSV0 U52480 ( .A1(n51313), .A2(n47305), .ZN(n48757) );
  NAND2HSV0 U52481 ( .A1(\pe5/aot [4]), .A2(n48755), .ZN(n48756) );
  XOR2HSV0 U52482 ( .A1(n48757), .A2(n48756), .Z(n48758) );
  XOR2HSV0 U52483 ( .A1(n48759), .A2(n48758), .Z(n48770) );
  NAND2HSV0 U52484 ( .A1(n48761), .A2(n48760), .ZN(n48763) );
  NAND2HSV0 U52485 ( .A1(n59640), .A2(n51176), .ZN(n48762) );
  XOR2HSV0 U52486 ( .A1(n48763), .A2(n48762), .Z(n48768) );
  NAND2HSV0 U52487 ( .A1(n52675), .A2(n30526), .ZN(n48766) );
  NAND2HSV0 U52488 ( .A1(n59427), .A2(n48764), .ZN(n48765) );
  XOR2HSV0 U52489 ( .A1(n48766), .A2(n48765), .Z(n48767) );
  XOR2HSV0 U52490 ( .A1(n48768), .A2(n48767), .Z(n48769) );
  XOR2HSV0 U52491 ( .A1(n48770), .A2(n48769), .Z(n48772) );
  NAND2HSV0 U52492 ( .A1(n39278), .A2(n51161), .ZN(n48771) );
  XNOR2HSV1 U52493 ( .A1(n48772), .A2(n48771), .ZN(n48774) );
  NAND2HSV0 U52494 ( .A1(n30270), .A2(n51331), .ZN(n48773) );
  XNOR2HSV1 U52495 ( .A1(n48774), .A2(n48773), .ZN(n48839) );
  NAND2HSV0 U52496 ( .A1(n39499), .A2(n48775), .ZN(n48777) );
  NAND2HSV0 U52497 ( .A1(n52584), .A2(n39445), .ZN(n48776) );
  XOR2HSV0 U52498 ( .A1(n48777), .A2(n48776), .Z(n48782) );
  NAND2HSV0 U52499 ( .A1(n30788), .A2(n50668), .ZN(n48780) );
  NAND2HSV0 U52500 ( .A1(\pe5/aot [23]), .A2(n48778), .ZN(n48779) );
  XOR2HSV0 U52501 ( .A1(n48780), .A2(n48779), .Z(n48781) );
  XOR2HSV0 U52502 ( .A1(n48782), .A2(n48781), .Z(n48793) );
  NAND2HSV0 U52503 ( .A1(n51188), .A2(\pe5/bq[11] ), .ZN(n48784) );
  NAND2HSV0 U52504 ( .A1(n59366), .A2(\pe5/bq[1] ), .ZN(n48783) );
  XOR2HSV0 U52505 ( .A1(n48784), .A2(n48783), .Z(n48791) );
  NAND2HSV0 U52506 ( .A1(n48786), .A2(n48785), .ZN(n48789) );
  NAND2HSV0 U52507 ( .A1(n53295), .A2(n48787), .ZN(n48788) );
  XOR2HSV0 U52508 ( .A1(n48789), .A2(n48788), .Z(n48790) );
  XOR2HSV0 U52509 ( .A1(n48791), .A2(n48790), .Z(n48792) );
  XOR2HSV0 U52510 ( .A1(n48793), .A2(n48792), .Z(n48808) );
  NAND2HSV0 U52511 ( .A1(n48077), .A2(\pe5/pq ), .ZN(n48795) );
  NAND2HSV0 U52512 ( .A1(\pe5/aot [13]), .A2(n48237), .ZN(n48794) );
  XOR2HSV0 U52513 ( .A1(n48795), .A2(n48794), .Z(n48800) );
  NAND2HSV0 U52514 ( .A1(n52607), .A2(n52610), .ZN(n48798) );
  NAND2HSV0 U52515 ( .A1(n48796), .A2(\pe5/bq[7] ), .ZN(n48797) );
  XOR2HSV0 U52516 ( .A1(n48798), .A2(n48797), .Z(n48799) );
  XOR2HSV0 U52517 ( .A1(n48800), .A2(n48799), .Z(n48806) );
  NAND2HSV0 U52518 ( .A1(n52623), .A2(n31045), .ZN(n53321) );
  NAND2HSV0 U52519 ( .A1(n52600), .A2(n50500), .ZN(n50584) );
  XNOR2HSV1 U52520 ( .A1(n48806), .A2(n48805), .ZN(n48807) );
  XNOR2HSV1 U52521 ( .A1(n48808), .A2(n48807), .ZN(n48837) );
  CLKNHSV0 U52522 ( .I(n48809), .ZN(n48813) );
  AOI22HSV0 U52523 ( .A1(n59897), .A2(n47291), .B1(n30616), .B2(n48810), .ZN(
        n48811) );
  AOI21HSV0 U52524 ( .A1(n48813), .A2(n48812), .B(n48811), .ZN(n48821) );
  NOR2HSV0 U52525 ( .A1(n48815), .A2(n48814), .ZN(n48819) );
  AOI22HSV0 U52526 ( .A1(n48817), .A2(\pe5/bq[2] ), .B1(n48816), .B2(n53307), 
        .ZN(n48818) );
  NOR2HSV1 U52527 ( .A1(n48819), .A2(n48818), .ZN(n48820) );
  XOR2HSV0 U52528 ( .A1(n48821), .A2(n48820), .Z(n48826) );
  NOR2HSV0 U52529 ( .A1(n48823), .A2(n48822), .ZN(n52621) );
  XOR2HSV0 U52530 ( .A1(n52621), .A2(n48824), .Z(n48825) );
  XNOR2HSV1 U52531 ( .A1(n48826), .A2(n48825), .ZN(n48835) );
  XOR2HSV0 U52532 ( .A1(n48828), .A2(n48827), .Z(n48833) );
  NAND2HSV0 U52533 ( .A1(n48829), .A2(n51191), .ZN(n48831) );
  NAND2HSV0 U52534 ( .A1(n48199), .A2(n52632), .ZN(n48830) );
  XOR2HSV0 U52535 ( .A1(n48831), .A2(n48830), .Z(n48832) );
  XOR2HSV0 U52536 ( .A1(n48833), .A2(n48832), .Z(n48834) );
  XOR2HSV0 U52537 ( .A1(n48835), .A2(n48834), .Z(n48836) );
  XNOR2HSV1 U52538 ( .A1(n48837), .A2(n48836), .ZN(n48838) );
  XOR3HSV2 U52539 ( .A1(n48840), .A2(n48839), .A3(n48838), .Z(n48843) );
  NAND2HSV0 U52540 ( .A1(n30255), .A2(n48841), .ZN(n48842) );
  XOR2HSV0 U52541 ( .A1(n48843), .A2(n48842), .Z(n48844) );
  XNOR2HSV1 U52542 ( .A1(n48845), .A2(n48844), .ZN(n48846) );
  XNOR2HSV1 U52543 ( .A1(n48847), .A2(n48846), .ZN(n48850) );
  NAND2HSV0 U52544 ( .A1(n48848), .A2(n50698), .ZN(n48849) );
  XOR2HSV0 U52545 ( .A1(n48850), .A2(n48849), .Z(n48851) );
  XNOR2HSV1 U52546 ( .A1(n48852), .A2(n48851), .ZN(n48853) );
  XNOR2HSV1 U52547 ( .A1(n48854), .A2(n48853), .ZN(n48855) );
  XNOR2HSV1 U52548 ( .A1(n48856), .A2(n48855), .ZN(n48857) );
  XNOR2HSV1 U52549 ( .A1(n48858), .A2(n48857), .ZN(n48859) );
  XNOR2HSV1 U52550 ( .A1(n48860), .A2(n48859), .ZN(n48861) );
  XNOR2HSV1 U52551 ( .A1(n48862), .A2(n48861), .ZN(n48864) );
  NAND2HSV0 U52552 ( .A1(n30752), .A2(n51157), .ZN(n48863) );
  XOR2HSV0 U52553 ( .A1(n48864), .A2(n48863), .Z(n48865) );
  XNOR2HSV1 U52554 ( .A1(n48866), .A2(n48865), .ZN(n48868) );
  NOR2HSV0 U52555 ( .A1(n50617), .A2(n50422), .ZN(n48867) );
  XNOR2HSV1 U52556 ( .A1(n48868), .A2(n48867), .ZN(n48869) );
  XNOR2HSV1 U52557 ( .A1(n48870), .A2(n48869), .ZN(n48871) );
  XNOR2HSV1 U52558 ( .A1(n48872), .A2(n48871), .ZN(n48874) );
  NAND2HSV0 U52559 ( .A1(n51211), .A2(n45816), .ZN(n48873) );
  XNOR2HSV1 U52560 ( .A1(n48874), .A2(n48873), .ZN(n48875) );
  XNOR2HSV1 U52561 ( .A1(n48876), .A2(n48875), .ZN(n48877) );
  XNOR2HSV1 U52562 ( .A1(n48878), .A2(n48877), .ZN(n48879) );
  XNOR2HSV1 U52563 ( .A1(n48880), .A2(n48879), .ZN(n48881) );
  XNOR2HSV1 U52564 ( .A1(n48882), .A2(n48881), .ZN(n48884) );
  NAND2HSV0 U52565 ( .A1(n59516), .A2(n48739), .ZN(n48883) );
  NOR2HSV4 U52566 ( .A1(n58442), .A2(n58434), .ZN(n48889) );
  INHSV2 U52567 ( .I(n48890), .ZN(n58383) );
  CLKNHSV0 U52568 ( .I(n48477), .ZN(n59502) );
  CLKNHSV0 U52569 ( .I(n48083), .ZN(n59503) );
  CLKNHSV0 U52570 ( .I(n48893), .ZN(n59533) );
  CLKNHSV0 U52571 ( .I(n48083), .ZN(n59510) );
  XOR2HSV0 U52572 ( .A1(n48895), .A2(n48894), .Z(n60084) );
  NAND2HSV2 U52573 ( .A1(n25709), .A2(n52415), .ZN(n48999) );
  CLKNAND2HSV1 U52574 ( .A1(n52854), .A2(n44944), .ZN(n48998) );
  CLKNAND2HSV0 U52575 ( .A1(n25834), .A2(n44711), .ZN(n48996) );
  INHSV2 U52576 ( .I(n44326), .ZN(n53087) );
  CLKNAND2HSV1 U52577 ( .A1(n53087), .A2(n53077), .ZN(n48992) );
  INHSV2 U52578 ( .I(n51894), .ZN(n52919) );
  CLKNAND2HSV0 U52579 ( .A1(n52919), .A2(n38904), .ZN(n48990) );
  NAND2HSV0 U52580 ( .A1(n52920), .A2(n52922), .ZN(n48988) );
  NOR2HSV0 U52581 ( .A1(n52921), .A2(n47570), .ZN(n48986) );
  NAND2HSV0 U52582 ( .A1(n52923), .A2(n52050), .ZN(n48983) );
  NAND2HSV0 U52583 ( .A1(n43926), .A2(n59506), .ZN(n48978) );
  BUFHSV4 U52584 ( .I(n59773), .Z(n52417) );
  NAND2HSV0 U52585 ( .A1(n52417), .A2(n52418), .ZN(n48976) );
  NAND2HSV0 U52586 ( .A1(n51965), .A2(n52172), .ZN(n48973) );
  NAND2HSV0 U52587 ( .A1(n52928), .A2(n52930), .ZN(n48971) );
  NAND2HSV0 U52588 ( .A1(n44714), .A2(n51966), .ZN(n48969) );
  CLKNAND2HSV1 U52589 ( .A1(n52931), .A2(\pe2/got [8]), .ZN(n48966) );
  NAND2HSV0 U52590 ( .A1(n52932), .A2(n53038), .ZN(n48960) );
  NAND2HSV0 U52591 ( .A1(n48896), .A2(n52855), .ZN(n48958) );
  NAND2HSV0 U52592 ( .A1(n59669), .A2(\pe2/got [2]), .ZN(n48954) );
  NAND2HSV0 U52593 ( .A1(n52993), .A2(n52952), .ZN(n48898) );
  NAND2HSV0 U52594 ( .A1(n59358), .A2(n51733), .ZN(n48897) );
  XOR2HSV0 U52595 ( .A1(n48898), .A2(n48897), .Z(n48902) );
  NAND2HSV0 U52596 ( .A1(n59768), .A2(\pe2/bq[21] ), .ZN(n48900) );
  NAND2HSV0 U52597 ( .A1(n59759), .A2(\pe2/bq[2] ), .ZN(n48899) );
  XOR2HSV0 U52598 ( .A1(n48900), .A2(n48899), .Z(n48901) );
  XOR2HSV0 U52599 ( .A1(n48902), .A2(n48901), .Z(n48910) );
  NAND2HSV0 U52600 ( .A1(n52310), .A2(n52484), .ZN(n48904) );
  NAND2HSV0 U52601 ( .A1(\pe2/aot [12]), .A2(n52988), .ZN(n48903) );
  XOR2HSV0 U52602 ( .A1(n48904), .A2(n48903), .Z(n48908) );
  NAND2HSV0 U52603 ( .A1(n44745), .A2(n38803), .ZN(n48906) );
  NAND2HSV0 U52604 ( .A1(\pe2/aot [8]), .A2(n45033), .ZN(n48905) );
  XOR2HSV0 U52605 ( .A1(n48906), .A2(n48905), .Z(n48907) );
  XOR2HSV0 U52606 ( .A1(n48908), .A2(n48907), .Z(n48909) );
  XOR2HSV0 U52607 ( .A1(n48910), .A2(n48909), .Z(n48925) );
  NAND2HSV0 U52608 ( .A1(n59976), .A2(n38792), .ZN(n48912) );
  NAND2HSV0 U52609 ( .A1(n45024), .A2(\pe2/bq[14] ), .ZN(n48911) );
  XOR2HSV0 U52610 ( .A1(n48912), .A2(n48911), .Z(n48916) );
  NAND2HSV0 U52611 ( .A1(\pe2/aot [2]), .A2(n52987), .ZN(n48914) );
  NAND2HSV0 U52612 ( .A1(\pe2/aot [19]), .A2(n52073), .ZN(n48913) );
  XOR2HSV0 U52613 ( .A1(n48914), .A2(n48913), .Z(n48915) );
  XOR2HSV0 U52614 ( .A1(n48916), .A2(n48915), .Z(n48923) );
  NAND2HSV0 U52615 ( .A1(n59974), .A2(n43956), .ZN(n48917) );
  XOR2HSV0 U52616 ( .A1(n52082), .A2(n48917), .Z(n48921) );
  NOR2HSV0 U52617 ( .A1(n51538), .A2(n36530), .ZN(n48919) );
  NAND2HSV0 U52618 ( .A1(n51759), .A2(n52472), .ZN(n48918) );
  XOR2HSV0 U52619 ( .A1(n48919), .A2(n48918), .Z(n48920) );
  XNOR2HSV1 U52620 ( .A1(n48921), .A2(n48920), .ZN(n48922) );
  XNOR2HSV1 U52621 ( .A1(n48923), .A2(n48922), .ZN(n48924) );
  XNOR2HSV1 U52622 ( .A1(n48925), .A2(n48924), .ZN(n48950) );
  NAND2HSV0 U52623 ( .A1(n39052), .A2(\pe2/bq[10] ), .ZN(n48927) );
  NAND2HSV0 U52624 ( .A1(n50930), .A2(n51457), .ZN(n48926) );
  XOR2HSV0 U52625 ( .A1(n48927), .A2(n48926), .Z(n48931) );
  NOR2HSV0 U52626 ( .A1(n38655), .A2(n44718), .ZN(n48929) );
  NAND2HSV0 U52627 ( .A1(n59499), .A2(n52950), .ZN(n48928) );
  XOR2HSV0 U52628 ( .A1(n48929), .A2(n48928), .Z(n48930) );
  XOR2HSV0 U52629 ( .A1(n48931), .A2(n48930), .Z(n48941) );
  NAND2HSV0 U52630 ( .A1(n59977), .A2(n52965), .ZN(n48933) );
  NAND2HSV0 U52631 ( .A1(n59633), .A2(n52179), .ZN(n48932) );
  XOR2HSV0 U52632 ( .A1(n48933), .A2(n48932), .Z(n48939) );
  NOR2HSV0 U52633 ( .A1(n48934), .A2(n51842), .ZN(n52205) );
  NOR2HSV0 U52634 ( .A1(n48935), .A2(n50920), .ZN(n48937) );
  NAND2HSV0 U52635 ( .A1(n59971), .A2(n52851), .ZN(n52207) );
  OAI22HSV0 U52636 ( .A1(n52205), .A2(n48937), .B1(n48936), .B2(n52207), .ZN(
        n48938) );
  XNOR2HSV1 U52637 ( .A1(n48939), .A2(n48938), .ZN(n48940) );
  XNOR2HSV1 U52638 ( .A1(n48941), .A2(n48940), .ZN(n48948) );
  NOR2HSV0 U52639 ( .A1(n38822), .A2(n48621), .ZN(n49607) );
  NOR2HSV0 U52640 ( .A1(n44049), .A2(n48621), .ZN(n52312) );
  AOI21HSV0 U52641 ( .A1(n51921), .A2(\pe2/bq[17] ), .B(n52312), .ZN(n48942)
         );
  AOI21HSV0 U52642 ( .A1(n49607), .A2(n48943), .B(n48942), .ZN(n48944) );
  NOR2HSV0 U52643 ( .A1(n52095), .A2(n36389), .ZN(n52308) );
  XNOR2HSV1 U52644 ( .A1(n48944), .A2(n52308), .ZN(n48946) );
  NAND2HSV0 U52645 ( .A1(n51636), .A2(n45015), .ZN(n52454) );
  NAND2HSV0 U52646 ( .A1(n59758), .A2(n52481), .ZN(n51985) );
  XOR2HSV0 U52647 ( .A1(n52454), .A2(n51985), .Z(n48945) );
  XOR2HSV0 U52648 ( .A1(n48946), .A2(n48945), .Z(n48947) );
  XNOR2HSV1 U52649 ( .A1(n48948), .A2(n48947), .ZN(n48949) );
  XNOR2HSV1 U52650 ( .A1(n48950), .A2(n48949), .ZN(n48952) );
  NAND2HSV0 U52651 ( .A1(n59684), .A2(n59767), .ZN(n48951) );
  XNOR2HSV1 U52652 ( .A1(n48952), .A2(n48951), .ZN(n48953) );
  XNOR2HSV1 U52653 ( .A1(n48954), .A2(n48953), .ZN(n48956) );
  NAND2HSV0 U52654 ( .A1(n59679), .A2(n52239), .ZN(n48955) );
  XNOR2HSV1 U52655 ( .A1(n48956), .A2(n48955), .ZN(n48957) );
  XNOR2HSV1 U52656 ( .A1(n48958), .A2(n48957), .ZN(n48959) );
  XNOR2HSV1 U52657 ( .A1(n48960), .A2(n48959), .ZN(n48962) );
  NAND2HSV0 U52658 ( .A1(n59766), .A2(n53041), .ZN(n48961) );
  XOR2HSV0 U52659 ( .A1(n48962), .A2(n48961), .Z(n48964) );
  CLKNHSV0 U52660 ( .I(n50928), .ZN(n52933) );
  NAND2HSV0 U52661 ( .A1(n52120), .A2(n52933), .ZN(n48963) );
  XNOR2HSV1 U52662 ( .A1(n48964), .A2(n48963), .ZN(n48965) );
  XNOR2HSV1 U52663 ( .A1(n48966), .A2(n48965), .ZN(n48968) );
  NAND2HSV0 U52664 ( .A1(n53056), .A2(\pe2/got [10]), .ZN(n48967) );
  XOR3HSV2 U52665 ( .A1(n48969), .A2(n48968), .A3(n48967), .Z(n48970) );
  XNOR2HSV1 U52666 ( .A1(n48971), .A2(n48970), .ZN(n48972) );
  XNOR2HSV1 U52667 ( .A1(n48973), .A2(n48972), .ZN(n48975) );
  NAND2HSV0 U52668 ( .A1(n59505), .A2(n51608), .ZN(n48974) );
  XOR3HSV2 U52669 ( .A1(n48976), .A2(n48975), .A3(n48974), .Z(n48977) );
  XOR2HSV0 U52670 ( .A1(n48978), .A2(n48977), .Z(n48981) );
  CLKNAND2HSV0 U52671 ( .A1(n52532), .A2(\pe2/got [16]), .ZN(n48980) );
  NAND2HSV0 U52672 ( .A1(n52534), .A2(\pe2/got [17]), .ZN(n48979) );
  XOR3HSV2 U52673 ( .A1(n48981), .A2(n48980), .A3(n48979), .Z(n48982) );
  XNOR2HSV1 U52674 ( .A1(n48983), .A2(n48982), .ZN(n48985) );
  CLKNAND2HSV0 U52675 ( .A1(n53078), .A2(n52042), .ZN(n48984) );
  XOR3HSV2 U52676 ( .A1(n48986), .A2(n48985), .A3(n48984), .Z(n48987) );
  XOR2HSV0 U52677 ( .A1(n48988), .A2(n48987), .Z(n48989) );
  XNOR2HSV1 U52678 ( .A1(n48990), .A2(n48989), .ZN(n48991) );
  XNOR2HSV1 U52679 ( .A1(n48992), .A2(n48991), .ZN(n48994) );
  CLKNAND2HSV0 U52680 ( .A1(n59929), .A2(n52416), .ZN(n48993) );
  XNOR2HSV1 U52681 ( .A1(n48994), .A2(n48993), .ZN(n48995) );
  INHSV2 U52682 ( .I(n49001), .ZN(n59530) );
  INHSV2 U52683 ( .I(ao2[32]), .ZN(n59531) );
  INHSV2 U52684 ( .I(go2[31]), .ZN(n59532) );
  NAND3HSV2 U52685 ( .A1(n46766), .A2(n53102), .A3(n49002), .ZN(n49095) );
  NOR2HSV1 U52686 ( .A1(n53104), .A2(n49003), .ZN(n49004) );
  CLKNAND2HSV1 U52687 ( .A1(n53106), .A2(n49004), .ZN(n49093) );
  CLKNAND2HSV0 U52688 ( .A1(n58712), .A2(n59328), .ZN(n49091) );
  NAND2HSV2 U52689 ( .A1(n58576), .A2(n59176), .ZN(n49089) );
  CLKNAND2HSV0 U52690 ( .A1(n59026), .A2(n58807), .ZN(n49087) );
  CLKNHSV0 U52691 ( .I(n49317), .ZN(n58716) );
  CLKNAND2HSV0 U52692 ( .A1(n58716), .A2(n59178), .ZN(n49085) );
  INHSV1 U52693 ( .I(n49666), .ZN(n59316) );
  CLKNAND2HSV1 U52694 ( .A1(n58717), .A2(n59316), .ZN(n49082) );
  BUFHSV2 U52695 ( .I(n58448), .Z(n58935) );
  CLKNAND2HSV1 U52696 ( .A1(n58935), .A2(n58810), .ZN(n49077) );
  CLKNAND2HSV0 U52697 ( .A1(n58718), .A2(n58811), .ZN(n49075) );
  CLKNHSV2 U52698 ( .I(n53110), .ZN(n58720) );
  CLKNAND2HSV1 U52699 ( .A1(n53111), .A2(n58720), .ZN(n49071) );
  CLKNAND2HSV1 U52700 ( .A1(n59916), .A2(\pe6/got [10]), .ZN(n49069) );
  BUFHSV2 U52701 ( .I(n58658), .Z(n58721) );
  CLKNAND2HSV1 U52702 ( .A1(n53113), .A2(n58721), .ZN(n49067) );
  NOR2HSV0 U52703 ( .A1(n50805), .A2(n58433), .ZN(n49065) );
  CLKNAND2HSV1 U52704 ( .A1(n59032), .A2(n58723), .ZN(n49061) );
  NAND2HSV2 U52705 ( .A1(n59033), .A2(n59292), .ZN(n49059) );
  NAND2HSV0 U52706 ( .A1(n58813), .A2(n58479), .ZN(n49057) );
  NAND2HSV0 U52707 ( .A1(n49743), .A2(n58527), .ZN(n49055) );
  NAND2HSV0 U52708 ( .A1(n49829), .A2(n58724), .ZN(n49053) );
  NAND2HSV0 U52709 ( .A1(n58939), .A2(n58403), .ZN(n49051) );
  CLKNAND2HSV0 U52710 ( .A1(n48038), .A2(n59264), .ZN(n49339) );
  CLKNHSV0 U52711 ( .I(n49339), .ZN(n49006) );
  NOR2HSV0 U52712 ( .A1(n46642), .A2(n32245), .ZN(n49762) );
  AOI22HSV0 U52713 ( .A1(n58975), .A2(n59088), .B1(n49836), .B2(\pe6/bq[4] ), 
        .ZN(n49005) );
  AOI21HSV2 U52714 ( .A1(n49006), .A2(n49762), .B(n49005), .ZN(n49010) );
  NAND2HSV0 U52715 ( .A1(\pe6/bq[8] ), .A2(n46217), .ZN(n49107) );
  NAND2HSV0 U52716 ( .A1(n59066), .A2(\pe6/aot [21]), .ZN(n49008) );
  NAND2HSV0 U52717 ( .A1(\pe6/bq[8] ), .A2(\pe6/aot [21]), .ZN(n59000) );
  CLKNAND2HSV1 U52718 ( .A1(n49205), .A2(n35732), .ZN(n53119) );
  NOR2HSV1 U52719 ( .A1(n59000), .A2(n53119), .ZN(n49007) );
  AOI21HSV2 U52720 ( .A1(n49107), .A2(n49008), .B(n49007), .ZN(n49009) );
  XNOR2HSV1 U52721 ( .A1(n49010), .A2(n49009), .ZN(n49017) );
  BUFHSV2 U52722 ( .I(\pe6/aot [2]), .Z(n58579) );
  CLKNAND2HSV0 U52723 ( .A1(n58356), .A2(n58579), .ZN(n58381) );
  NOR2HSV0 U52724 ( .A1(n49011), .A2(n58381), .ZN(n49013) );
  AOI22HSV0 U52725 ( .A1(n59100), .A2(n58464), .B1(\pe6/aot [19]), .B2(
        \pe6/bq[5] ), .ZN(n49012) );
  NOR2HSV2 U52726 ( .A1(n49013), .A2(n49012), .ZN(n49015) );
  NAND2HSV0 U52727 ( .A1(\pe6/bq[2] ), .A2(n49831), .ZN(n49014) );
  XNOR2HSV1 U52728 ( .A1(n49015), .A2(n49014), .ZN(n49016) );
  XNOR2HSV1 U52729 ( .A1(n49017), .A2(n49016), .ZN(n49049) );
  NAND2HSV0 U52730 ( .A1(\pe6/bq[1] ), .A2(\pe6/aot [23]), .ZN(n49019) );
  NAND2HSV0 U52731 ( .A1(n35750), .A2(\pe6/aot [13]), .ZN(n49018) );
  XOR2HSV0 U52732 ( .A1(n49019), .A2(n49018), .Z(n49023) );
  NAND2HSV0 U52733 ( .A1(n32276), .A2(\pe6/aot [1]), .ZN(n49021) );
  NAND2HSV0 U52734 ( .A1(n36150), .A2(n59266), .ZN(n49020) );
  XOR2HSV0 U52735 ( .A1(n49021), .A2(n49020), .Z(n49022) );
  XOR2HSV0 U52736 ( .A1(n49023), .A2(n49022), .Z(n49032) );
  NAND2HSV0 U52737 ( .A1(\pe6/bq[14] ), .A2(\pe6/aot [10]), .ZN(n49025) );
  NAND2HSV0 U52738 ( .A1(n59075), .A2(\pe6/aot [17]), .ZN(n49024) );
  XOR2HSV0 U52739 ( .A1(n49025), .A2(n49024), .Z(n49030) );
  NAND2HSV0 U52740 ( .A1(n58628), .A2(n58378), .ZN(n58594) );
  NOR2HSV0 U52741 ( .A1(n49026), .A2(n58594), .ZN(n49028) );
  AOI22HSV0 U52742 ( .A1(n50829), .A2(\pe6/aot [5]), .B1(n58842), .B2(n59084), 
        .ZN(n49027) );
  NOR2HSV1 U52743 ( .A1(n49028), .A2(n49027), .ZN(n49029) );
  XNOR2HSV1 U52744 ( .A1(n49030), .A2(n49029), .ZN(n49031) );
  XNOR2HSV1 U52745 ( .A1(n49032), .A2(n49031), .ZN(n49048) );
  NAND2HSV0 U52746 ( .A1(n58833), .A2(n35632), .ZN(n49034) );
  NAND2HSV0 U52747 ( .A1(n58976), .A2(n53115), .ZN(n49033) );
  XOR2HSV0 U52748 ( .A1(n49034), .A2(n49033), .Z(n49038) );
  NAND2HSV0 U52749 ( .A1(n58962), .A2(n49208), .ZN(n49036) );
  NAND2HSV0 U52750 ( .A1(n59045), .A2(n58495), .ZN(n49035) );
  XOR2HSV0 U52751 ( .A1(n49036), .A2(n49035), .Z(n49037) );
  XOR2HSV0 U52752 ( .A1(n49038), .A2(n49037), .Z(n49046) );
  NAND2HSV0 U52753 ( .A1(n59265), .A2(\pe6/aot [11]), .ZN(n49040) );
  NAND2HSV0 U52754 ( .A1(n32982), .A2(\pe6/aot [7]), .ZN(n49039) );
  XOR2HSV0 U52755 ( .A1(n49040), .A2(n49039), .Z(n49044) );
  NOR2HSV0 U52756 ( .A1(n35837), .A2(n58530), .ZN(n49042) );
  CLKNAND2HSV0 U52757 ( .A1(\pe6/bq[21] ), .A2(n58404), .ZN(n49041) );
  XOR2HSV0 U52758 ( .A1(n49042), .A2(n49041), .Z(n49043) );
  XOR2HSV0 U52759 ( .A1(n49044), .A2(n49043), .Z(n49045) );
  XOR2HSV0 U52760 ( .A1(n49046), .A2(n49045), .Z(n49047) );
  XOR3HSV2 U52761 ( .A1(n49049), .A2(n49048), .A3(n49047), .Z(n49050) );
  XNOR2HSV1 U52762 ( .A1(n49051), .A2(n49050), .ZN(n49052) );
  XNOR2HSV1 U52763 ( .A1(n49053), .A2(n49052), .ZN(n49054) );
  XNOR2HSV1 U52764 ( .A1(n49055), .A2(n49054), .ZN(n49056) );
  XNOR2HSV1 U52765 ( .A1(n49057), .A2(n49056), .ZN(n49058) );
  XNOR2HSV1 U52766 ( .A1(n49059), .A2(n49058), .ZN(n49060) );
  XNOR2HSV1 U52767 ( .A1(n49061), .A2(n49060), .ZN(n49063) );
  CLKNAND2HSV0 U52768 ( .A1(n59144), .A2(n36109), .ZN(n49062) );
  XNOR2HSV1 U52769 ( .A1(n49063), .A2(n49062), .ZN(n49064) );
  XNOR2HSV1 U52770 ( .A1(n49065), .A2(n49064), .ZN(n49066) );
  XNOR2HSV1 U52771 ( .A1(n49067), .A2(n49066), .ZN(n49068) );
  XNOR2HSV1 U52772 ( .A1(n49069), .A2(n49068), .ZN(n49070) );
  XNOR2HSV1 U52773 ( .A1(n49071), .A2(n49070), .ZN(n49073) );
  CLKNAND2HSV1 U52774 ( .A1(n59915), .A2(n58719), .ZN(n49072) );
  XNOR2HSV1 U52775 ( .A1(n49073), .A2(n49072), .ZN(n49074) );
  XNOR2HSV1 U52776 ( .A1(n49075), .A2(n49074), .ZN(n49076) );
  XNOR2HSV1 U52777 ( .A1(n49077), .A2(n49076), .ZN(n49080) );
  BUFHSV2 U52778 ( .I(n49078), .Z(n59335) );
  CLKNAND2HSV0 U52779 ( .A1(n59335), .A2(\pe6/got [15]), .ZN(n49079) );
  XOR2HSV0 U52780 ( .A1(n49080), .A2(n49079), .Z(n49081) );
  XNOR2HSV1 U52781 ( .A1(n49082), .A2(n49081), .ZN(n49084) );
  NAND2HSV0 U52782 ( .A1(n59528), .A2(n58715), .ZN(n49083) );
  XOR3HSV2 U52783 ( .A1(n49085), .A2(n49084), .A3(n49083), .Z(n49086) );
  XNOR2HSV1 U52784 ( .A1(n49087), .A2(n49086), .ZN(n49088) );
  XNOR2HSV1 U52785 ( .A1(n49089), .A2(n49088), .ZN(n49090) );
  XNOR2HSV1 U52786 ( .A1(n49091), .A2(n49090), .ZN(n49092) );
  XNOR2HSV1 U52787 ( .A1(n49093), .A2(n49092), .ZN(n49094) );
  XOR2HSV0 U52788 ( .A1(n49095), .A2(n49094), .Z(\pe6/poht [9]) );
  NAND3HSV2 U52789 ( .A1(n46766), .A2(n53102), .A3(n49096), .ZN(n49172) );
  NOR2HSV2 U52790 ( .A1(n53104), .A2(n46270), .ZN(n49097) );
  CLKNAND2HSV1 U52791 ( .A1(n53106), .A2(n49097), .ZN(n49170) );
  NAND2HSV0 U52792 ( .A1(n58712), .A2(n49098), .ZN(n49168) );
  NAND2HSV2 U52793 ( .A1(n53107), .A2(n59031), .ZN(n49166) );
  CLKNAND2HSV1 U52794 ( .A1(n58385), .A2(n32596), .ZN(n49164) );
  CLKNAND2HSV0 U52795 ( .A1(n53109), .A2(n58811), .ZN(n49162) );
  CLKNAND2HSV1 U52796 ( .A1(n59028), .A2(\pe6/got [12]), .ZN(n49159) );
  NAND2HSV0 U52797 ( .A1(n58448), .A2(n44393), .ZN(n49155) );
  CLKNAND2HSV1 U52798 ( .A1(n59680), .A2(n58721), .ZN(n49153) );
  CLKNAND2HSV1 U52799 ( .A1(n53111), .A2(n58709), .ZN(n49149) );
  CLKNAND2HSV0 U52800 ( .A1(n53112), .A2(n58513), .ZN(n49147) );
  NAND2HSV0 U52801 ( .A1(n53113), .A2(n58478), .ZN(n49145) );
  CLKNAND2HSV0 U52802 ( .A1(n59179), .A2(n58479), .ZN(n49143) );
  NAND2HSV0 U52803 ( .A1(n49667), .A2(n59231), .ZN(n49139) );
  NAND2HSV0 U52804 ( .A1(n59379), .A2(n59235), .ZN(n49137) );
  AOI22HSV2 U52805 ( .A1(n58975), .A2(\pe6/aot [14]), .B1(n58842), .B2(n48037), 
        .ZN(n49100) );
  AOI21HSV2 U52806 ( .A1(n53129), .A2(n49101), .B(n49100), .ZN(n49103) );
  XOR2HSV0 U52807 ( .A1(n49103), .A2(n49102), .Z(n49119) );
  CLKNAND2HSV1 U52808 ( .A1(n33023), .A2(n58579), .ZN(n49105) );
  CLKNAND2HSV0 U52809 ( .A1(n58668), .A2(n53134), .ZN(n49104) );
  XOR2HSV0 U52810 ( .A1(n49105), .A2(n49104), .Z(n49111) );
  NOR2HSV0 U52811 ( .A1(n46642), .A2(n46789), .ZN(n49109) );
  NOR2HSV0 U52812 ( .A1(n48042), .A2(n49188), .ZN(n49108) );
  NAND2HSV0 U52813 ( .A1(n49106), .A2(n53115), .ZN(n58677) );
  OAI22HSV1 U52814 ( .A1(n49109), .A2(n49108), .B1(n58677), .B2(n49107), .ZN(
        n49110) );
  XNOR2HSV1 U52815 ( .A1(n49111), .A2(n49110), .ZN(n49118) );
  NAND2HSV0 U52816 ( .A1(n59277), .A2(\pe6/aot [19]), .ZN(n49830) );
  XOR2HSV0 U52817 ( .A1(n49112), .A2(n49830), .Z(n49116) );
  CLKNAND2HSV0 U52818 ( .A1(n32982), .A2(n59252), .ZN(n49114) );
  NAND2HSV0 U52819 ( .A1(n49205), .A2(\pe6/aot [17]), .ZN(n49113) );
  XOR2HSV0 U52820 ( .A1(n49114), .A2(n49113), .Z(n49115) );
  XOR2HSV0 U52821 ( .A1(n49116), .A2(n49115), .Z(n49117) );
  XOR3HSV2 U52822 ( .A1(n49119), .A2(n49118), .A3(n49117), .Z(n49135) );
  NAND2HSV0 U52823 ( .A1(n58976), .A2(\pe6/aot [8]), .ZN(n49121) );
  CLKNHSV0 U52824 ( .I(n48041), .ZN(n59273) );
  NAND2HSV0 U52825 ( .A1(n59273), .A2(\pe6/aot [13]), .ZN(n49120) );
  XOR2HSV0 U52826 ( .A1(n49121), .A2(n49120), .Z(n49125) );
  NAND2HSV0 U52827 ( .A1(n59051), .A2(\pe6/aot [1]), .ZN(n49123) );
  CLKNAND2HSV0 U52828 ( .A1(n35751), .A2(n49847), .ZN(n49122) );
  XOR2HSV0 U52829 ( .A1(n49123), .A2(n49122), .Z(n49124) );
  XOR2HSV0 U52830 ( .A1(n49125), .A2(n49124), .Z(n49133) );
  CLKNAND2HSV0 U52831 ( .A1(n59265), .A2(\pe6/aot [7]), .ZN(n49127) );
  NAND2HSV0 U52832 ( .A1(n59041), .A2(n49760), .ZN(n49126) );
  XOR2HSV0 U52833 ( .A1(n49127), .A2(n49126), .Z(n49131) );
  NOR2HSV0 U52834 ( .A1(n46850), .A2(n59193), .ZN(n49129) );
  CLKNAND2HSV0 U52835 ( .A1(n48044), .A2(\pe6/aot [11]), .ZN(n49128) );
  XOR2HSV0 U52836 ( .A1(n49129), .A2(n49128), .Z(n49130) );
  XOR2HSV0 U52837 ( .A1(n49131), .A2(n49130), .Z(n49132) );
  XOR2HSV0 U52838 ( .A1(n49133), .A2(n49132), .Z(n49134) );
  XNOR2HSV1 U52839 ( .A1(n49135), .A2(n49134), .ZN(n49136) );
  XNOR2HSV1 U52840 ( .A1(n49137), .A2(n49136), .ZN(n49138) );
  XNOR2HSV1 U52841 ( .A1(n49139), .A2(n49138), .ZN(n49141) );
  CLKNAND2HSV0 U52842 ( .A1(n58901), .A2(n48891), .ZN(n49140) );
  XNOR2HSV1 U52843 ( .A1(n49141), .A2(n49140), .ZN(n49142) );
  XOR2HSV0 U52844 ( .A1(n49143), .A2(n49142), .Z(n49144) );
  XNOR2HSV1 U52845 ( .A1(n49145), .A2(n49144), .ZN(n49146) );
  XNOR2HSV1 U52846 ( .A1(n49147), .A2(n49146), .ZN(n49148) );
  XNOR2HSV1 U52847 ( .A1(n49149), .A2(n49148), .ZN(n49151) );
  CLKNAND2HSV1 U52848 ( .A1(n58702), .A2(n59182), .ZN(n49150) );
  XNOR2HSV1 U52849 ( .A1(n49151), .A2(n49150), .ZN(n49152) );
  XNOR2HSV1 U52850 ( .A1(n49153), .A2(n49152), .ZN(n49154) );
  XNOR2HSV1 U52851 ( .A1(n49155), .A2(n49154), .ZN(n49157) );
  NAND2HSV0 U52852 ( .A1(n59677), .A2(n49742), .ZN(n49156) );
  XOR2HSV0 U52853 ( .A1(n49157), .A2(n49156), .Z(n49158) );
  XNOR2HSV1 U52854 ( .A1(n49159), .A2(n49158), .ZN(n49161) );
  XNOR2HSV1 U52855 ( .A1(n49164), .A2(n49163), .ZN(n49165) );
  XNOR2HSV1 U52856 ( .A1(n49166), .A2(n49165), .ZN(n49167) );
  XOR2HSV0 U52857 ( .A1(n49168), .A2(n49167), .Z(n49169) );
  XNOR2HSV1 U52858 ( .A1(n49170), .A2(n49169), .ZN(n49171) );
  XOR2HSV0 U52859 ( .A1(n49172), .A2(n49171), .Z(\pe6/poht [13]) );
  CLKNHSV0 U52860 ( .I(n53104), .ZN(n49175) );
  AND2HSV2 U52861 ( .A1(n49175), .A2(n59316), .Z(n49176) );
  CLKNAND2HSV0 U52862 ( .A1(n49176), .A2(n49177), .ZN(n49180) );
  NAND2HSV0 U52863 ( .A1(n49178), .A2(n59031), .ZN(n49179) );
  NAND2HSV2 U52864 ( .A1(n49180), .A2(n49179), .ZN(n49247) );
  CLKBUFHSV4 U52865 ( .I(n49181), .Z(n58656) );
  CLKNAND2HSV1 U52866 ( .A1(n58656), .A2(n58810), .ZN(n49243) );
  CLKNAND2HSV1 U52867 ( .A1(n58657), .A2(n58654), .ZN(n49241) );
  CLKNAND2HSV0 U52868 ( .A1(n53109), .A2(n49742), .ZN(n49239) );
  CLKNAND2HSV1 U52869 ( .A1(n58611), .A2(n58812), .ZN(n49236) );
  CLKNAND2HSV0 U52870 ( .A1(n58448), .A2(n59182), .ZN(n49232) );
  CLKNAND2HSV1 U52871 ( .A1(n58936), .A2(n58709), .ZN(n49230) );
  NAND2HSV0 U52872 ( .A1(n58662), .A2(n58478), .ZN(n49226) );
  CLKNAND2HSV0 U52873 ( .A1(n53112), .A2(n58479), .ZN(n49224) );
  NAND2HSV0 U52874 ( .A1(n58664), .A2(n58527), .ZN(n49222) );
  NAND2HSV0 U52875 ( .A1(n53114), .A2(n58816), .ZN(n49220) );
  CLKNAND2HSV0 U52876 ( .A1(n58901), .A2(n58403), .ZN(n49218) );
  CLKNAND2HSV0 U52877 ( .A1(n58356), .A2(\pe6/aot [13]), .ZN(n49183) );
  CLKNAND2HSV0 U52878 ( .A1(n58668), .A2(n58459), .ZN(n49182) );
  XOR2HSV0 U52879 ( .A1(n49183), .A2(n49182), .Z(n49187) );
  NAND2HSV0 U52880 ( .A1(n59246), .A2(\pe6/aot [10]), .ZN(n49185) );
  NAND2HSV0 U52881 ( .A1(n58962), .A2(n58449), .ZN(n49184) );
  XOR2HSV0 U52882 ( .A1(n49185), .A2(n49184), .Z(n49186) );
  XOR2HSV0 U52883 ( .A1(n49187), .A2(n49186), .Z(n49198) );
  CLKNAND2HSV1 U52884 ( .A1(n58360), .A2(n58631), .ZN(n58595) );
  CLKNAND2HSV0 U52885 ( .A1(n58405), .A2(n35732), .ZN(n49746) );
  NOR2HSV0 U52886 ( .A1(n58595), .A2(n49746), .ZN(n49190) );
  AOI22HSV0 U52887 ( .A1(n58975), .A2(n32972), .B1(n59189), .B2(n59041), .ZN(
        n49189) );
  NOR2HSV2 U52888 ( .A1(n49190), .A2(n49189), .ZN(n49192) );
  XNOR2HSV1 U52889 ( .A1(n49192), .A2(n49191), .ZN(n49196) );
  NAND2HSV0 U52890 ( .A1(n49844), .A2(n59260), .ZN(n49194) );
  NAND2HSV0 U52891 ( .A1(n58682), .A2(n59252), .ZN(n49193) );
  XOR2HSV0 U52892 ( .A1(n49194), .A2(n49193), .Z(n49195) );
  XOR2HSV0 U52893 ( .A1(n49196), .A2(n49195), .Z(n49197) );
  XOR2HSV0 U52894 ( .A1(n49198), .A2(n49197), .Z(n49216) );
  NAND2HSV0 U52895 ( .A1(n59273), .A2(\pe6/aot [11]), .ZN(n49200) );
  NAND2HSV0 U52896 ( .A1(n58990), .A2(\pe6/aot [17]), .ZN(n49199) );
  XOR2HSV0 U52897 ( .A1(n49200), .A2(n49199), .Z(n49204) );
  CLKNAND2HSV0 U52898 ( .A1(n59240), .A2(n53134), .ZN(n49202) );
  NAND2HSV0 U52899 ( .A1(n35750), .A2(\pe6/aot [7]), .ZN(n49201) );
  XOR2HSV0 U52900 ( .A1(n49202), .A2(n49201), .Z(n49203) );
  XOR2HSV0 U52901 ( .A1(n49204), .A2(n49203), .Z(n49214) );
  NOR2HSV0 U52902 ( .A1(n50847), .A2(n59193), .ZN(n49207) );
  NAND2HSV0 U52903 ( .A1(n49205), .A2(n58842), .ZN(n49206) );
  XOR2HSV0 U52904 ( .A1(n49207), .A2(n49206), .Z(n49212) );
  NAND2HSV0 U52905 ( .A1(n32982), .A2(n49208), .ZN(n59110) );
  CLKNAND2HSV1 U52906 ( .A1(\pe6/bq[4] ), .A2(\pe6/aot [1]), .ZN(n58341) );
  NOR2HSV0 U52907 ( .A1(n59110), .A2(n58341), .ZN(n49210) );
  AOI22HSV0 U52908 ( .A1(\pe6/bq[17] ), .A2(\pe6/aot [1]), .B1(n49208), .B2(
        \pe6/bq[4] ), .ZN(n49209) );
  NOR2HSV2 U52909 ( .A1(n49210), .A2(n49209), .ZN(n49211) );
  XNOR2HSV1 U52910 ( .A1(n49212), .A2(n49211), .ZN(n49213) );
  XNOR2HSV1 U52911 ( .A1(n49214), .A2(n49213), .ZN(n49215) );
  XNOR2HSV1 U52912 ( .A1(n49216), .A2(n49215), .ZN(n49217) );
  XNOR2HSV1 U52913 ( .A1(n49218), .A2(n49217), .ZN(n49219) );
  XNOR2HSV1 U52914 ( .A1(n49220), .A2(n49219), .ZN(n49221) );
  XNOR2HSV1 U52915 ( .A1(n49222), .A2(n49221), .ZN(n49223) );
  XNOR2HSV1 U52916 ( .A1(n49224), .A2(n49223), .ZN(n49225) );
  XNOR2HSV1 U52917 ( .A1(n49226), .A2(n49225), .ZN(n49228) );
  CLKNAND2HSV0 U52918 ( .A1(n58702), .A2(n58513), .ZN(n49227) );
  XNOR2HSV1 U52919 ( .A1(n49228), .A2(n49227), .ZN(n49229) );
  XNOR2HSV1 U52920 ( .A1(n49230), .A2(n49229), .ZN(n49231) );
  XNOR2HSV1 U52921 ( .A1(n49232), .A2(n49231), .ZN(n49234) );
  CLKNAND2HSV0 U52922 ( .A1(n59335), .A2(n58658), .ZN(n49233) );
  XOR2HSV0 U52923 ( .A1(n49234), .A2(n49233), .Z(n49235) );
  XNOR2HSV1 U52924 ( .A1(n49236), .A2(n49235), .ZN(n49238) );
  NAND2HSV0 U52925 ( .A1(n29753), .A2(n58719), .ZN(n49237) );
  XOR3HSV2 U52926 ( .A1(n49239), .A2(n49238), .A3(n49237), .Z(n49240) );
  XNOR2HSV1 U52927 ( .A1(n49241), .A2(n49240), .ZN(n49242) );
  XNOR2HSV1 U52928 ( .A1(n49243), .A2(n49242), .ZN(n49245) );
  AND2HSV2 U52929 ( .A1(n32596), .A2(n58712), .Z(n49244) );
  XNOR2HSV1 U52930 ( .A1(n49245), .A2(n49244), .ZN(n49246) );
  XNOR2HSV1 U52931 ( .A1(n49247), .A2(n49246), .ZN(n49248) );
  XOR2HSV0 U52932 ( .A1(n49249), .A2(n49248), .Z(\pe6/poht [15]) );
  INHSV2 U52933 ( .I(n51118), .ZN(n56907) );
  CLKNAND2HSV0 U52934 ( .A1(n56621), .A2(n56419), .ZN(n49313) );
  INHSV2 U52935 ( .I(n56680), .ZN(n56559) );
  CLKNHSV0 U52936 ( .I(n56936), .ZN(n56541) );
  CLKNHSV0 U52937 ( .I(n56541), .ZN(n49254) );
  INAND2HSV0 U52938 ( .A1(n49254), .B1(n59620), .ZN(n49306) );
  NAND2HSV0 U52939 ( .A1(n49255), .A2(\pe3/got [1]), .ZN(n49304) );
  NAND2HSV0 U52940 ( .A1(\pe3/aot [8]), .A2(n56094), .ZN(n49257) );
  NAND2HSV0 U52941 ( .A1(\pe3/aot [18]), .A2(n56189), .ZN(n49256) );
  XOR2HSV0 U52942 ( .A1(n49257), .A2(n49256), .Z(n49262) );
  NAND2HSV0 U52943 ( .A1(n59344), .A2(n56915), .ZN(n49260) );
  CLKNAND2HSV0 U52944 ( .A1(n42940), .A2(n56348), .ZN(n49259) );
  XOR2HSV0 U52945 ( .A1(n49260), .A2(n49259), .Z(n49261) );
  XOR2HSV0 U52946 ( .A1(n49262), .A2(n49261), .Z(n49271) );
  NAND2HSV0 U52947 ( .A1(n56221), .A2(n43544), .ZN(n49264) );
  CLKNHSV0 U52948 ( .I(n53229), .ZN(n56455) );
  NAND2HSV0 U52949 ( .A1(n56455), .A2(\pe3/bq[11] ), .ZN(n49263) );
  XOR2HSV0 U52950 ( .A1(n49264), .A2(n49263), .Z(n49269) );
  NOR2HSV0 U52951 ( .A1(n37357), .A2(n50722), .ZN(n49267) );
  NAND2HSV0 U52952 ( .A1(\pe3/aot [16]), .A2(n45639), .ZN(n49266) );
  XOR2HSV0 U52953 ( .A1(n49267), .A2(n49266), .Z(n49268) );
  XOR2HSV0 U52954 ( .A1(n49269), .A2(n49268), .Z(n49270) );
  XOR2HSV0 U52955 ( .A1(n49271), .A2(n49270), .Z(n49286) );
  NAND2HSV0 U52956 ( .A1(n56378), .A2(n56454), .ZN(n49274) );
  NAND2HSV0 U52957 ( .A1(n56188), .A2(n56785), .ZN(n49273) );
  XOR2HSV0 U52958 ( .A1(n49274), .A2(n49273), .Z(n49280) );
  CLKNHSV0 U52959 ( .I(n49413), .ZN(n49278) );
  NOR2HSV0 U52960 ( .A1(n56784), .A2(n37196), .ZN(n49277) );
  NAND2HSV2 U52961 ( .A1(n59511), .A2(n56971), .ZN(n52845) );
  OAI22HSV0 U52962 ( .A1(n49278), .A2(n49277), .B1(n49276), .B2(n52845), .ZN(
        n49279) );
  XNOR2HSV1 U52963 ( .A1(n49280), .A2(n49279), .ZN(n49284) );
  NOR2HSV0 U52964 ( .A1(n56567), .A2(n49281), .ZN(n56271) );
  XOR2HSV0 U52965 ( .A1(n56271), .A2(n49282), .Z(n49283) );
  XNOR2HSV1 U52966 ( .A1(n49284), .A2(n49283), .ZN(n49285) );
  XNOR2HSV1 U52967 ( .A1(n49286), .A2(n49285), .ZN(n49302) );
  NAND2HSV0 U52968 ( .A1(n56434), .A2(n42971), .ZN(n49288) );
  NAND2HSV0 U52969 ( .A1(n42728), .A2(\pe3/bq[4] ), .ZN(n49287) );
  XOR2HSV0 U52970 ( .A1(n49288), .A2(n49287), .Z(n49292) );
  NAND2HSV0 U52971 ( .A1(n56439), .A2(\pe3/bq[18] ), .ZN(n49290) );
  NAND2HSV0 U52972 ( .A1(\pe3/aot [10]), .A2(n45534), .ZN(n49289) );
  XOR2HSV0 U52973 ( .A1(n49290), .A2(n49289), .Z(n49291) );
  XOR2HSV0 U52974 ( .A1(n49292), .A2(n49291), .Z(n49300) );
  NAND2HSV0 U52975 ( .A1(n56795), .A2(n56433), .ZN(n49294) );
  NAND2HSV0 U52976 ( .A1(n56354), .A2(n45982), .ZN(n49293) );
  XOR2HSV0 U52977 ( .A1(n49294), .A2(n49293), .Z(n49298) );
  NOR2HSV0 U52978 ( .A1(n56956), .A2(n43039), .ZN(n49296) );
  NAND2HSV0 U52979 ( .A1(n43280), .A2(n56627), .ZN(n49295) );
  XOR2HSV0 U52980 ( .A1(n49296), .A2(n49295), .Z(n49297) );
  XOR2HSV0 U52981 ( .A1(n49298), .A2(n49297), .Z(n49299) );
  XOR2HSV0 U52982 ( .A1(n49300), .A2(n49299), .Z(n49301) );
  XNOR2HSV1 U52983 ( .A1(n49302), .A2(n49301), .ZN(n49303) );
  XNOR2HSV1 U52984 ( .A1(n49304), .A2(n49303), .ZN(n49305) );
  XNOR2HSV1 U52985 ( .A1(n49306), .A2(n49305), .ZN(n49309) );
  NOR2HSV0 U52986 ( .A1(n56391), .A2(n56906), .ZN(n49308) );
  NAND2HSV0 U52987 ( .A1(n56422), .A2(n56781), .ZN(n49307) );
  NOR2HSV0 U52988 ( .A1(n56475), .A2(n56859), .ZN(n49311) );
  NAND2HSV0 U52989 ( .A1(n56396), .A2(n56560), .ZN(n49310) );
  INHSV2 U52990 ( .I(n56778), .ZN(n56266) );
  INHSV2 U52991 ( .I(n49315), .ZN(n59027) );
  BUFHSV2 U52992 ( .I(n46822), .Z(n59172) );
  CLKNHSV0 U52993 ( .I(n49317), .ZN(n58934) );
  CLKNAND2HSV1 U52994 ( .A1(n58935), .A2(n58937), .ZN(n49397) );
  CLKNAND2HSV0 U52995 ( .A1(n58718), .A2(\pe6/got [15]), .ZN(n49395) );
  NAND2HSV0 U52996 ( .A1(n59177), .A2(n58811), .ZN(n49391) );
  NAND2HSV0 U52997 ( .A1(n59916), .A2(n33039), .ZN(n49389) );
  CLKNAND2HSV1 U52998 ( .A1(n58938), .A2(n59181), .ZN(n49387) );
  CLKNAND2HSV1 U52999 ( .A1(n53114), .A2(n58812), .ZN(n49385) );
  NAND2HSV0 U53000 ( .A1(n58722), .A2(n58526), .ZN(n49380) );
  BUFHSV2 U53001 ( .I(\pe6/got [7]), .Z(n58814) );
  CLKNAND2HSV1 U53002 ( .A1(n59033), .A2(n58814), .ZN(n49378) );
  CLKNAND2HSV1 U53003 ( .A1(n59420), .A2(n58398), .ZN(n49376) );
  CLKNAND2HSV1 U53004 ( .A1(n35722), .A2(n59292), .ZN(n49374) );
  CLKNAND2HSV1 U53005 ( .A1(n32165), .A2(n58479), .ZN(n49372) );
  NAND2HSV0 U53006 ( .A1(n49319), .A2(n58527), .ZN(n49370) );
  NAND2HSV0 U53007 ( .A1(n32218), .A2(n58817), .ZN(n49366) );
  NAND2HSV0 U53008 ( .A1(n59050), .A2(n58464), .ZN(n49321) );
  CLKNAND2HSV0 U53009 ( .A1(n59098), .A2(n53134), .ZN(n49320) );
  XOR2HSV0 U53010 ( .A1(n49321), .A2(n49320), .Z(n49326) );
  CLKNAND2HSV0 U53011 ( .A1(n44336), .A2(n49847), .ZN(n58637) );
  OAI21HSV0 U53012 ( .A1(n59205), .A2(n58359), .B(n49322), .ZN(n49323) );
  OAI21HSV0 U53013 ( .A1(n58637), .A2(n49324), .B(n49323), .ZN(n49325) );
  XNOR2HSV1 U53014 ( .A1(n49326), .A2(n49325), .ZN(n49337) );
  NOR2HSV0 U53015 ( .A1(n49327), .A2(n49699), .ZN(n50839) );
  NOR2HSV0 U53016 ( .A1(n58984), .A2(n58463), .ZN(n49329) );
  CLKNAND2HSV1 U53017 ( .A1(n58496), .A2(\pe6/aot [10]), .ZN(n58545) );
  OAI22HSV0 U53018 ( .A1(n50839), .A2(n49329), .B1(n49328), .B2(n58545), .ZN(
        n49335) );
  NOR2HSV0 U53019 ( .A1(n49331), .A2(n49330), .ZN(n49333) );
  AOI22HSV0 U53020 ( .A1(n59054), .A2(n58353), .B1(n58668), .B2(n58631), .ZN(
        n49332) );
  NOR2HSV1 U53021 ( .A1(n49333), .A2(n49332), .ZN(n49334) );
  XOR2HSV0 U53022 ( .A1(n49335), .A2(n49334), .Z(n49336) );
  XNOR2HSV1 U53023 ( .A1(n49337), .A2(n49336), .ZN(n49364) );
  NOR2HSV0 U53024 ( .A1(n48042), .A2(n32373), .ZN(n49683) );
  NOR2HSV0 U53025 ( .A1(n46642), .A2(n32373), .ZN(n49833) );
  NAND2HSV0 U53026 ( .A1(n58990), .A2(n58824), .ZN(n58989) );
  XNOR2HSV1 U53027 ( .A1(n49338), .A2(n58989), .ZN(n49341) );
  NAND2HSV0 U53028 ( .A1(n59089), .A2(\pe6/aot [13]), .ZN(n58985) );
  XOR2HSV0 U53029 ( .A1(n49339), .A2(n58985), .Z(n49340) );
  XOR2HSV0 U53030 ( .A1(n49341), .A2(n49340), .Z(n49347) );
  NAND2HSV0 U53031 ( .A1(\pe6/bq[25] ), .A2(\pe6/aot [1]), .ZN(n50840) );
  XOR2HSV0 U53032 ( .A1(n58863), .A2(n50840), .Z(n49345) );
  NAND2HSV0 U53033 ( .A1(n46210), .A2(n58842), .ZN(n49343) );
  NAND2HSV0 U53034 ( .A1(n59100), .A2(n58459), .ZN(n49342) );
  XOR2HSV0 U53035 ( .A1(n49343), .A2(n49342), .Z(n49344) );
  XNOR2HSV1 U53036 ( .A1(n49345), .A2(n49344), .ZN(n49346) );
  XNOR2HSV1 U53037 ( .A1(n49347), .A2(n49346), .ZN(n49363) );
  NAND2HSV0 U53038 ( .A1(n58682), .A2(\pe6/aot [11]), .ZN(n49349) );
  NAND2HSV0 U53039 ( .A1(n32982), .A2(n59099), .ZN(n49348) );
  XOR2HSV0 U53040 ( .A1(n49349), .A2(n49348), .Z(n49353) );
  NAND2HSV0 U53041 ( .A1(\pe6/bq[2] ), .A2(n59239), .ZN(n49351) );
  NAND2HSV0 U53042 ( .A1(n33023), .A2(n35632), .ZN(n49350) );
  XOR2HSV0 U53043 ( .A1(n49351), .A2(n49350), .Z(n49352) );
  XOR2HSV0 U53044 ( .A1(n49353), .A2(n49352), .Z(n49361) );
  NAND2HSV0 U53045 ( .A1(\pe6/bq[9] ), .A2(\pe6/aot [17]), .ZN(n49355) );
  NAND2HSV0 U53046 ( .A1(n59051), .A2(\pe6/aot [7]), .ZN(n49354) );
  XOR2HSV0 U53047 ( .A1(n49355), .A2(n49354), .Z(n49359) );
  NOR2HSV0 U53048 ( .A1(n48041), .A2(n46637), .ZN(n49357) );
  NAND2HSV0 U53049 ( .A1(n58731), .A2(\pe6/aot [21]), .ZN(n49356) );
  XOR2HSV0 U53050 ( .A1(n49357), .A2(n49356), .Z(n49358) );
  XOR2HSV0 U53051 ( .A1(n49359), .A2(n49358), .Z(n49360) );
  XOR2HSV0 U53052 ( .A1(n49361), .A2(n49360), .Z(n49362) );
  XOR3HSV2 U53053 ( .A1(n49364), .A2(n49363), .A3(n49362), .Z(n49365) );
  XNOR2HSV1 U53054 ( .A1(n49366), .A2(n49365), .ZN(n49368) );
  NAND2HSV0 U53055 ( .A1(n58886), .A2(n58816), .ZN(n49367) );
  XNOR2HSV1 U53056 ( .A1(n49368), .A2(n49367), .ZN(n49369) );
  XNOR2HSV1 U53057 ( .A1(n49370), .A2(n49369), .ZN(n49371) );
  XNOR2HSV1 U53058 ( .A1(n49372), .A2(n49371), .ZN(n49373) );
  XNOR2HSV1 U53059 ( .A1(n49374), .A2(n49373), .ZN(n49375) );
  XNOR2HSV1 U53060 ( .A1(n49376), .A2(n49375), .ZN(n49377) );
  XNOR2HSV1 U53061 ( .A1(n49378), .A2(n49377), .ZN(n49379) );
  XNOR2HSV1 U53062 ( .A1(n49380), .A2(n49379), .ZN(n49383) );
  BUFHSV2 U53063 ( .I(n49381), .Z(n59317) );
  BUFHSV2 U53064 ( .I(\pe6/got [9]), .Z(n59037) );
  CLKNAND2HSV1 U53065 ( .A1(n59317), .A2(n59037), .ZN(n49382) );
  XNOR2HSV1 U53066 ( .A1(n49383), .A2(n49382), .ZN(n49384) );
  XNOR2HSV1 U53067 ( .A1(n49385), .A2(n49384), .ZN(n49386) );
  XNOR2HSV1 U53068 ( .A1(n49387), .A2(n49386), .ZN(n49388) );
  XNOR2HSV1 U53069 ( .A1(n49389), .A2(n49388), .ZN(n49390) );
  XNOR2HSV1 U53070 ( .A1(n49391), .A2(n49390), .ZN(n49393) );
  CLKNAND2HSV1 U53071 ( .A1(n58601), .A2(n58810), .ZN(n49392) );
  XNOR2HSV1 U53072 ( .A1(n49393), .A2(n49392), .ZN(n49394) );
  XNOR2HSV1 U53073 ( .A1(n49395), .A2(n49394), .ZN(n49396) );
  XNOR2HSV1 U53074 ( .A1(n49397), .A2(n49396), .ZN(n49399) );
  CLKNAND2HSV0 U53075 ( .A1(n59161), .A2(n32971), .ZN(n49398) );
  INHSV2 U53076 ( .I(n49739), .ZN(n59029) );
  INHSV2 U53077 ( .I(n49401), .ZN(n59170) );
  INHSV2 U53078 ( .I(n49402), .ZN(n58372) );
  NAND2HSV0 U53079 ( .A1(n56783), .A2(n43374), .ZN(n49490) );
  CLKNAND2HSV0 U53080 ( .A1(n56622), .A2(n56335), .ZN(n49488) );
  NAND2HSV0 U53081 ( .A1(n59920), .A2(n56065), .ZN(n49486) );
  NAND2HSV0 U53082 ( .A1(n56685), .A2(n56174), .ZN(n49484) );
  CLKNAND2HSV1 U53083 ( .A1(n55947), .A2(n56421), .ZN(n49480) );
  CLKNAND2HSV0 U53084 ( .A1(n55824), .A2(n56176), .ZN(n49476) );
  NAND2HSV0 U53085 ( .A1(n56067), .A2(n56683), .ZN(n49467) );
  CLKNAND2HSV0 U53086 ( .A1(n56179), .A2(n56267), .ZN(n49465) );
  NAND2HSV0 U53087 ( .A1(n56180), .A2(n56068), .ZN(n49463) );
  NAND2HSV0 U53088 ( .A1(n56070), .A2(n55950), .ZN(n49459) );
  NAND2HSV0 U53089 ( .A1(n49405), .A2(n56975), .ZN(n49457) );
  NAND2HSV0 U53090 ( .A1(n42950), .A2(\pe3/bq[9] ), .ZN(n49407) );
  NAND2HSV0 U53091 ( .A1(n55858), .A2(n55828), .ZN(n49406) );
  XOR2HSV0 U53092 ( .A1(n49407), .A2(n49406), .Z(n49411) );
  CLKNAND2HSV0 U53093 ( .A1(n56074), .A2(n56213), .ZN(n49409) );
  NAND2HSV0 U53094 ( .A1(n56221), .A2(n42971), .ZN(n49408) );
  XOR2HSV0 U53095 ( .A1(n49409), .A2(n49408), .Z(n49410) );
  XOR2HSV0 U53096 ( .A1(n49411), .A2(n49410), .Z(n49455) );
  OAI21HSV0 U53097 ( .A1(n56914), .A2(n45567), .B(n55986), .ZN(n49412) );
  OAI21HSV1 U53098 ( .A1(n49414), .A2(n49413), .B(n49412), .ZN(n49418) );
  CLKNAND2HSV0 U53099 ( .A1(n56087), .A2(\pe3/bq[4] ), .ZN(n56002) );
  NAND2HSV0 U53100 ( .A1(n42818), .A2(n56529), .ZN(n56115) );
  NOR2HSV0 U53101 ( .A1(n56002), .A2(n56115), .ZN(n49416) );
  AOI22HSV0 U53102 ( .A1(n45695), .A2(n56529), .B1(n42818), .B2(\pe3/bq[4] ), 
        .ZN(n49415) );
  NOR2HSV2 U53103 ( .A1(n49416), .A2(n49415), .ZN(n49417) );
  XNOR2HSV1 U53104 ( .A1(n49418), .A2(n49417), .ZN(n49422) );
  XOR2HSV0 U53105 ( .A1(n49420), .A2(n49419), .Z(n49421) );
  XNOR2HSV1 U53106 ( .A1(n49422), .A2(n49421), .ZN(n49430) );
  NAND2HSV0 U53107 ( .A1(\pe3/aot [14]), .A2(n55975), .ZN(n49425) );
  NAND2HSV0 U53108 ( .A1(n56370), .A2(n56094), .ZN(n49424) );
  XOR2HSV0 U53109 ( .A1(n49425), .A2(n49424), .Z(n49428) );
  CLKNAND2HSV0 U53110 ( .A1(n56378), .A2(n56688), .ZN(n56427) );
  NAND2HSV0 U53111 ( .A1(\pe3/aot [8]), .A2(\pe3/bq[19] ), .ZN(n49426) );
  XOR2HSV0 U53112 ( .A1(n56427), .A2(n49426), .Z(n49427) );
  XOR2HSV0 U53113 ( .A1(n49428), .A2(n49427), .Z(n49429) );
  XNOR2HSV1 U53114 ( .A1(n49430), .A2(n49429), .ZN(n49454) );
  NAND2HSV0 U53115 ( .A1(n56740), .A2(n56433), .ZN(n49432) );
  NAND2HSV0 U53116 ( .A1(n56204), .A2(n56832), .ZN(n49431) );
  XOR2HSV0 U53117 ( .A1(n49432), .A2(n49431), .Z(n49436) );
  NAND2HSV0 U53118 ( .A1(\pe3/aot [16]), .A2(\pe3/bq[11] ), .ZN(n49434) );
  NAND2HSV0 U53119 ( .A1(\pe3/aot [3]), .A2(n55872), .ZN(n49433) );
  XOR2HSV0 U53120 ( .A1(n49434), .A2(n49433), .Z(n49435) );
  XOR2HSV0 U53121 ( .A1(n49436), .A2(n49435), .Z(n49453) );
  NAND2HSV0 U53122 ( .A1(n56439), .A2(n56222), .ZN(n49438) );
  INHSV2 U53123 ( .I(n56567), .ZN(n56520) );
  NAND2HSV0 U53124 ( .A1(n56520), .A2(\pe3/bq[18] ), .ZN(n49437) );
  XOR2HSV0 U53125 ( .A1(n49438), .A2(n49437), .Z(n49443) );
  NAND2HSV0 U53126 ( .A1(n56911), .A2(n49439), .ZN(n49441) );
  NAND2HSV0 U53127 ( .A1(n59511), .A2(\pe3/bq[26] ), .ZN(n49440) );
  XOR2HSV0 U53128 ( .A1(n49441), .A2(n49440), .Z(n49442) );
  XOR2HSV0 U53129 ( .A1(n49443), .A2(n49442), .Z(n49451) );
  NAND2HSV0 U53130 ( .A1(n56113), .A2(n56187), .ZN(n49445) );
  NAND2HSV0 U53131 ( .A1(n56464), .A2(n55970), .ZN(n49444) );
  XOR2HSV0 U53132 ( .A1(n49445), .A2(n49444), .Z(n49449) );
  NAND2HSV0 U53133 ( .A1(n42940), .A2(n56915), .ZN(n49447) );
  NAND2HSV0 U53134 ( .A1(\pe3/aot [11]), .A2(n56640), .ZN(n49446) );
  XOR2HSV0 U53135 ( .A1(n49447), .A2(n49446), .Z(n49448) );
  XOR2HSV0 U53136 ( .A1(n49449), .A2(n49448), .Z(n49450) );
  XOR2HSV0 U53137 ( .A1(n49451), .A2(n49450), .Z(n49452) );
  XOR4HSV1 U53138 ( .A1(n49455), .A2(n49454), .A3(n49453), .A4(n49452), .Z(
        n49456) );
  XNOR2HSV1 U53139 ( .A1(n49457), .A2(n49456), .ZN(n49458) );
  XNOR2HSV1 U53140 ( .A1(n49459), .A2(n49458), .ZN(n49461) );
  NAND2HSV0 U53141 ( .A1(n56127), .A2(n56069), .ZN(n49460) );
  XNOR2HSV1 U53142 ( .A1(n49461), .A2(n49460), .ZN(n49462) );
  XNOR2HSV1 U53143 ( .A1(n49463), .A2(n49462), .ZN(n49464) );
  XNOR2HSV1 U53144 ( .A1(n49465), .A2(n49464), .ZN(n49466) );
  XNOR2HSV1 U53145 ( .A1(n49467), .A2(n49466), .ZN(n49471) );
  NOR2HSV0 U53146 ( .A1(n45728), .A2(n56778), .ZN(n49470) );
  NAND2HSV0 U53147 ( .A1(n56855), .A2(n49468), .ZN(n49469) );
  XOR3HSV1 U53148 ( .A1(n49471), .A2(n49470), .A3(n49469), .Z(n49474) );
  NOR2HSV0 U53149 ( .A1(n56475), .A2(n56680), .ZN(n49473) );
  CLKNAND2HSV0 U53150 ( .A1(n56242), .A2(\pe3/got [10]), .ZN(n49472) );
  XOR3HSV1 U53151 ( .A1(n49474), .A2(n49473), .A3(n49472), .Z(n49475) );
  XNOR2HSV1 U53152 ( .A1(n49476), .A2(n49475), .ZN(n49478) );
  CLKNAND2HSV0 U53153 ( .A1(n46052), .A2(n56247), .ZN(n49477) );
  XNOR2HSV1 U53154 ( .A1(n49478), .A2(n49477), .ZN(n49479) );
  XNOR2HSV1 U53155 ( .A1(n49480), .A2(n49479), .ZN(n49482) );
  NAND2HSV0 U53156 ( .A1(n56662), .A2(n56493), .ZN(n49481) );
  XNOR2HSV1 U53157 ( .A1(n49482), .A2(n49481), .ZN(n49483) );
  XNOR2HSV1 U53158 ( .A1(n49484), .A2(n49483), .ZN(n49485) );
  XNOR2HSV1 U53159 ( .A1(n49486), .A2(n49485), .ZN(n49487) );
  XNOR2HSV1 U53160 ( .A1(n49488), .A2(n49487), .ZN(n49489) );
  XNOR2HSV1 U53161 ( .A1(n49490), .A2(n49489), .ZN(n49491) );
  BUFHSV2 U53162 ( .I(n56260), .Z(n56900) );
  NAND2HSV2 U53163 ( .A1(n25709), .A2(n49492), .ZN(n49602) );
  INAND2HSV2 U53164 ( .A1(n39088), .B1(n52047), .ZN(n49600) );
  NAND2HSV2 U53165 ( .A1(n52048), .A2(n52416), .ZN(n49598) );
  NOR2HSV1 U53166 ( .A1(n52049), .A2(n44327), .ZN(n49590) );
  NAND2HSV0 U53167 ( .A1(n44968), .A2(n51889), .ZN(n49588) );
  NOR2HSV0 U53168 ( .A1(n52921), .A2(n53064), .ZN(n49586) );
  NAND2HSV0 U53169 ( .A1(n52814), .A2(n53055), .ZN(n49578) );
  CLKNAND2HSV0 U53170 ( .A1(n52417), .A2(n49493), .ZN(n49576) );
  NAND2HSV0 U53171 ( .A1(n59634), .A2(\pe2/got [10]), .ZN(n49573) );
  NAND2HSV0 U53172 ( .A1(n52928), .A2(n52052), .ZN(n49571) );
  NAND2HSV0 U53173 ( .A1(n52174), .A2(n52419), .ZN(n49569) );
  NAND2HSV0 U53174 ( .A1(n52287), .A2(\pe2/got [6]), .ZN(n49566) );
  NAND2HSV0 U53175 ( .A1(n45149), .A2(n52239), .ZN(n49560) );
  NAND2HSV0 U53176 ( .A1(n52934), .A2(n51932), .ZN(n49558) );
  NAND2HSV0 U53177 ( .A1(n59679), .A2(n59767), .ZN(n49556) );
  NAND2HSV0 U53178 ( .A1(n39052), .A2(n51825), .ZN(n49496) );
  NAND2HSV0 U53179 ( .A1(\pe2/aot [11]), .A2(\pe2/bq[17] ), .ZN(n49495) );
  XOR2HSV0 U53180 ( .A1(n49496), .A2(n49495), .Z(n49500) );
  NAND2HSV0 U53181 ( .A1(n59768), .A2(n43961), .ZN(n49498) );
  NAND2HSV0 U53182 ( .A1(\pe2/aot [10]), .A2(n52988), .ZN(n49497) );
  XOR2HSV0 U53183 ( .A1(n49498), .A2(n49497), .Z(n49499) );
  XOR2HSV0 U53184 ( .A1(n49500), .A2(n49499), .Z(n49508) );
  NAND2HSV0 U53185 ( .A1(n52974), .A2(n51919), .ZN(n49502) );
  NAND2HSV0 U53186 ( .A1(n51759), .A2(n52073), .ZN(n49501) );
  XOR2HSV0 U53187 ( .A1(n49502), .A2(n49501), .Z(n49506) );
  NAND2HSV0 U53188 ( .A1(n52951), .A2(n51998), .ZN(n49504) );
  NAND2HSV0 U53189 ( .A1(n52184), .A2(n45015), .ZN(n49503) );
  XOR2HSV0 U53190 ( .A1(n49504), .A2(n49503), .Z(n49505) );
  XOR2HSV0 U53191 ( .A1(n49506), .A2(n49505), .Z(n49507) );
  XOR2HSV0 U53192 ( .A1(n49508), .A2(n49507), .Z(n49527) );
  NAND2HSV0 U53193 ( .A1(n51743), .A2(n52438), .ZN(n49510) );
  NAND2HSV0 U53194 ( .A1(n52456), .A2(n45033), .ZN(n49509) );
  XOR2HSV0 U53195 ( .A1(n49510), .A2(n49509), .Z(n49514) );
  NAND2HSV0 U53196 ( .A1(n50930), .A2(n52857), .ZN(n49512) );
  NAND2HSV0 U53197 ( .A1(\pe2/aot [22]), .A2(\pe2/bq[6] ), .ZN(n49511) );
  XOR2HSV0 U53198 ( .A1(n49512), .A2(n49511), .Z(n49513) );
  XOR2HSV0 U53199 ( .A1(n49514), .A2(n49513), .Z(n49525) );
  NAND2HSV0 U53200 ( .A1(n59358), .A2(n51997), .ZN(n49517) );
  NAND2HSV0 U53201 ( .A1(n52294), .A2(n52193), .ZN(n49516) );
  XOR2HSV0 U53202 ( .A1(n49517), .A2(n49516), .Z(n49523) );
  NOR2HSV0 U53203 ( .A1(n51538), .A2(n44854), .ZN(n49521) );
  NOR2HSV0 U53204 ( .A1(n49618), .A2(n49518), .ZN(n49520) );
  NAND2HSV0 U53205 ( .A1(\pe2/aot [2]), .A2(n52950), .ZN(n52091) );
  OAI22HSV1 U53206 ( .A1(n49521), .A2(n49520), .B1(n49519), .B2(n52091), .ZN(
        n49522) );
  XNOR2HSV1 U53207 ( .A1(n49523), .A2(n49522), .ZN(n49524) );
  XNOR2HSV1 U53208 ( .A1(n49525), .A2(n49524), .ZN(n49526) );
  XNOR2HSV1 U53209 ( .A1(n49527), .A2(n49526), .ZN(n49554) );
  CLKNHSV0 U53210 ( .I(n49528), .ZN(n49532) );
  AOI22HSV0 U53211 ( .A1(n49530), .A2(n52851), .B1(n52104), .B2(n51457), .ZN(
        n49531) );
  AOI21HSV1 U53212 ( .A1(n49532), .A2(n52204), .B(n49531), .ZN(n49537) );
  CLKNHSV0 U53213 ( .I(n49533), .ZN(n49535) );
  NOR2HSV0 U53214 ( .A1(n52095), .A2(n47608), .ZN(n51970) );
  AOI22HSV0 U53215 ( .A1(\pe2/aot [7]), .A2(\pe2/bq[21] ), .B1(n39032), .B2(
        \pe2/aot [1]), .ZN(n49534) );
  AOI21HSV0 U53216 ( .A1(n49535), .A2(n51970), .B(n49534), .ZN(n49536) );
  XNOR2HSV1 U53217 ( .A1(n49537), .A2(n49536), .ZN(n49544) );
  NAND2HSV0 U53218 ( .A1(n59972), .A2(\pe2/bq[4] ), .ZN(n52094) );
  NAND2HSV0 U53219 ( .A1(n50956), .A2(n52484), .ZN(n52092) );
  NOR2HSV0 U53220 ( .A1(n49538), .A2(n52092), .ZN(n49539) );
  AOI21HSV0 U53221 ( .A1(n49540), .A2(n52094), .B(n49539), .ZN(n49542) );
  XOR2HSV0 U53222 ( .A1(n49542), .A2(n49541), .Z(n49543) );
  XNOR2HSV1 U53223 ( .A1(n49544), .A2(n49543), .ZN(n49552) );
  NAND2HSV0 U53224 ( .A1(n52070), .A2(n52962), .ZN(n49546) );
  NAND2HSV0 U53225 ( .A1(n52966), .A2(n43956), .ZN(n49545) );
  XOR2HSV0 U53226 ( .A1(n49546), .A2(n49545), .Z(n49550) );
  NAND2HSV0 U53227 ( .A1(n53005), .A2(n38803), .ZN(n49548) );
  NAND2HSV0 U53228 ( .A1(n29736), .A2(n52179), .ZN(n49547) );
  XOR2HSV0 U53229 ( .A1(n49548), .A2(n49547), .Z(n49549) );
  XOR2HSV0 U53230 ( .A1(n49550), .A2(n49549), .Z(n49551) );
  XNOR2HSV1 U53231 ( .A1(n49552), .A2(n49551), .ZN(n49553) );
  XNOR2HSV1 U53232 ( .A1(n49554), .A2(n49553), .ZN(n49555) );
  XNOR2HSV1 U53233 ( .A1(n49556), .A2(n49555), .ZN(n49557) );
  XNOR2HSV1 U53234 ( .A1(n49558), .A2(n49557), .ZN(n49559) );
  XNOR2HSV1 U53235 ( .A1(n49560), .A2(n49559), .ZN(n49562) );
  NAND2HSV0 U53236 ( .A1(n59766), .A2(n51896), .ZN(n49561) );
  XOR2HSV0 U53237 ( .A1(n49562), .A2(n49561), .Z(n49564) );
  NAND2HSV0 U53238 ( .A1(n45218), .A2(n52175), .ZN(n49563) );
  XNOR2HSV1 U53239 ( .A1(n49564), .A2(n49563), .ZN(n49565) );
  XNOR2HSV1 U53240 ( .A1(n49566), .A2(n49565), .ZN(n49568) );
  NAND2HSV0 U53241 ( .A1(n59761), .A2(\pe2/got [8]), .ZN(n49567) );
  XOR3HSV2 U53242 ( .A1(n49569), .A2(n49568), .A3(n49567), .Z(n49570) );
  XNOR2HSV1 U53243 ( .A1(n49571), .A2(n49570), .ZN(n49572) );
  XNOR2HSV1 U53244 ( .A1(n49573), .A2(n49572), .ZN(n49575) );
  NOR2HSV0 U53245 ( .A1(n53065), .A2(n47555), .ZN(n49574) );
  XOR3HSV2 U53246 ( .A1(n49576), .A2(n49575), .A3(n49574), .Z(n49577) );
  XOR2HSV0 U53247 ( .A1(n49578), .A2(n49577), .Z(n49581) );
  CLKNAND2HSV1 U53248 ( .A1(n52532), .A2(n48084), .ZN(n49580) );
  CLKNAND2HSV0 U53249 ( .A1(n52138), .A2(n51964), .ZN(n49579) );
  XOR3HSV2 U53250 ( .A1(n49581), .A2(n49580), .A3(n49579), .Z(n49582) );
  XNOR2HSV1 U53251 ( .A1(n49583), .A2(n49582), .ZN(n49585) );
  CLKNAND2HSV0 U53252 ( .A1(n53078), .A2(n52050), .ZN(n49584) );
  XOR3HSV2 U53253 ( .A1(n49586), .A2(n49585), .A3(n49584), .Z(n49587) );
  XOR2HSV0 U53254 ( .A1(n49588), .A2(n49587), .Z(n49589) );
  XNOR2HSV1 U53255 ( .A1(n49590), .A2(n49589), .ZN(n49594) );
  NAND2HSV2 U53256 ( .A1(n51893), .A2(\pe2/got [21]), .ZN(n49593) );
  CLKNAND2HSV0 U53257 ( .A1(n52399), .A2(n49591), .ZN(n49592) );
  XOR3HSV2 U53258 ( .A1(n49594), .A2(n49593), .A3(n49592), .Z(n49595) );
  XOR2HSV0 U53259 ( .A1(n49596), .A2(n49595), .Z(n49597) );
  XOR2HSV0 U53260 ( .A1(n49598), .A2(n49597), .Z(n49599) );
  XNOR2HSV4 U53261 ( .A1(n49602), .A2(n49601), .ZN(n49605) );
  INAND2HSV2 U53262 ( .A1(n49603), .B1(n52163), .ZN(n49604) );
  XNOR2HSV4 U53263 ( .A1(n49605), .A2(n49604), .ZN(\pe2/poht [5]) );
  CLKNAND2HSV1 U53264 ( .A1(n52047), .A2(n59354), .ZN(n49660) );
  CLKNAND2HSV0 U53265 ( .A1(n51798), .A2(\pe2/got [10]), .ZN(n49655) );
  NOR2HSV1 U53266 ( .A1(n52049), .A2(n51800), .ZN(n49653) );
  CLKNAND2HSV1 U53267 ( .A1(n51799), .A2(\pe2/got [8]), .ZN(n49651) );
  NOR2HSV1 U53268 ( .A1(n47500), .A2(n52018), .ZN(n49649) );
  CLKNAND2HSV1 U53269 ( .A1(n59775), .A2(n59778), .ZN(n49646) );
  NAND2HSV0 U53270 ( .A1(n52895), .A2(n25824), .ZN(n49641) );
  NAND2HSV0 U53271 ( .A1(n59505), .A2(n59767), .ZN(n49639) );
  NOR2HSV0 U53272 ( .A1(n52095), .A2(n48063), .ZN(n52098) );
  NAND2HSV0 U53273 ( .A1(\pe2/aot [8]), .A2(n52193), .ZN(n51453) );
  XOR2HSV0 U53274 ( .A1(n52098), .A2(n51453), .Z(n49609) );
  CLKNAND2HSV0 U53275 ( .A1(n53005), .A2(n52857), .ZN(n51737) );
  XOR2HSV0 U53276 ( .A1(n49607), .A2(n51737), .Z(n49608) );
  XOR2HSV0 U53277 ( .A1(n49609), .A2(n49608), .Z(n49617) );
  NAND2HSV0 U53278 ( .A1(n52056), .A2(\pe2/bq[12] ), .ZN(n49611) );
  NAND2HSV0 U53279 ( .A1(n51636), .A2(n51900), .ZN(n49610) );
  XOR2HSV0 U53280 ( .A1(n49611), .A2(n49610), .Z(n49615) );
  NAND2HSV0 U53281 ( .A1(n44745), .A2(n52905), .ZN(n49613) );
  NAND2HSV0 U53282 ( .A1(n59976), .A2(\pe2/bq[6] ), .ZN(n49612) );
  XOR2HSV0 U53283 ( .A1(n49613), .A2(n49612), .Z(n49614) );
  XOR2HSV0 U53284 ( .A1(n49615), .A2(n49614), .Z(n49616) );
  XOR2HSV0 U53285 ( .A1(n49617), .A2(n49616), .Z(n49637) );
  CLKNAND2HSV1 U53286 ( .A1(\pe2/aot [2]), .A2(n49619), .ZN(n49621) );
  NAND2HSV0 U53287 ( .A1(n51743), .A2(n52851), .ZN(n49620) );
  XOR2HSV0 U53288 ( .A1(n49621), .A2(n49620), .Z(n49625) );
  NAND2HSV0 U53289 ( .A1(\pe2/aot [15]), .A2(n51493), .ZN(n49623) );
  NAND2HSV0 U53290 ( .A1(\pe2/aot [9]), .A2(n51825), .ZN(n49622) );
  XOR2HSV0 U53291 ( .A1(n49623), .A2(n49622), .Z(n49624) );
  XOR2HSV0 U53292 ( .A1(n49625), .A2(n49624), .Z(n49635) );
  NAND2HSV0 U53293 ( .A1(n51460), .A2(n51832), .ZN(n49627) );
  NAND2HSV0 U53294 ( .A1(n59633), .A2(n52063), .ZN(n49626) );
  XOR2HSV0 U53295 ( .A1(n49627), .A2(n49626), .Z(n49633) );
  NOR2HSV0 U53296 ( .A1(n51537), .A2(n49628), .ZN(n49631) );
  NOR2HSV0 U53297 ( .A1(n51538), .A2(n47580), .ZN(n49630) );
  NAND2HSV0 U53298 ( .A1(n52867), .A2(n51839), .ZN(n51924) );
  OAI22HSV2 U53299 ( .A1(n49631), .A2(n49630), .B1(n51924), .B2(n49629), .ZN(
        n49632) );
  XNOR2HSV1 U53300 ( .A1(n49633), .A2(n49632), .ZN(n49634) );
  XNOR2HSV1 U53301 ( .A1(n49635), .A2(n49634), .ZN(n49636) );
  XNOR2HSV1 U53302 ( .A1(n49637), .A2(n49636), .ZN(n49638) );
  XNOR2HSV1 U53303 ( .A1(n49639), .A2(n49638), .ZN(n49640) );
  XNOR2HSV1 U53304 ( .A1(n49641), .A2(n49640), .ZN(n49644) );
  NAND2HSV2 U53305 ( .A1(n51861), .A2(n51933), .ZN(n49643) );
  CLKNAND2HSV1 U53306 ( .A1(n51862), .A2(n51896), .ZN(n49642) );
  XOR3HSV2 U53307 ( .A1(n49644), .A2(n49643), .A3(n49642), .Z(n49645) );
  XNOR2HSV1 U53308 ( .A1(n49646), .A2(n49645), .ZN(n49648) );
  INHSV2 U53309 ( .I(n50928), .ZN(n51895) );
  CLKNAND2HSV0 U53310 ( .A1(n51868), .A2(n51895), .ZN(n49647) );
  XOR3HSV2 U53311 ( .A1(n49649), .A2(n49648), .A3(n49647), .Z(n49650) );
  XOR2HSV0 U53312 ( .A1(n49651), .A2(n49650), .Z(n49652) );
  XNOR2HSV1 U53313 ( .A1(n49653), .A2(n49652), .ZN(n49654) );
  XNOR2HSV1 U53314 ( .A1(n49655), .A2(n49654), .ZN(n49658) );
  INHSV4 U53315 ( .I(n49656), .ZN(n51892) );
  CLKNAND2HSV1 U53316 ( .A1(n51878), .A2(n51892), .ZN(n49657) );
  XNOR2HSV1 U53317 ( .A1(n49658), .A2(n49657), .ZN(n49659) );
  NAND2HSV2 U53318 ( .A1(n52840), .A2(n45289), .ZN(n49662) );
  XNOR2HSV4 U53319 ( .A1(n49664), .A2(n49663), .ZN(\pe2/poht [16]) );
  NAND2HSV0 U53320 ( .A1(n59918), .A2(n59029), .ZN(n49732) );
  NAND2HSV0 U53321 ( .A1(n59680), .A2(n58807), .ZN(n49730) );
  NAND2HSV0 U53322 ( .A1(n59177), .A2(n49098), .ZN(n49725) );
  NAND2HSV0 U53323 ( .A1(n58663), .A2(n58937), .ZN(n49723) );
  CLKNAND2HSV0 U53324 ( .A1(n58938), .A2(\pe6/got [15]), .ZN(n49721) );
  CLKNAND2HSV1 U53325 ( .A1(n59179), .A2(n49741), .ZN(n49719) );
  NAND2HSV0 U53326 ( .A1(n49667), .A2(n33039), .ZN(n49715) );
  NAND2HSV0 U53327 ( .A1(n59050), .A2(n58665), .ZN(n49669) );
  NAND2HSV0 U53328 ( .A1(n58975), .A2(n59239), .ZN(n49668) );
  XOR2HSV0 U53329 ( .A1(n49669), .A2(n49668), .Z(n49673) );
  NAND2HSV0 U53330 ( .A1(n59051), .A2(\pe6/aot [11]), .ZN(n49671) );
  NAND2HSV0 U53331 ( .A1(n48035), .A2(n58459), .ZN(n49670) );
  XOR2HSV0 U53332 ( .A1(n49671), .A2(n49670), .Z(n49672) );
  NAND2HSV0 U53333 ( .A1(n44435), .A2(n58857), .ZN(n49675) );
  NAND2HSV0 U53334 ( .A1(n58976), .A2(n58760), .ZN(n49674) );
  XOR2HSV0 U53335 ( .A1(n49675), .A2(n49674), .Z(n49679) );
  NOR2HSV0 U53336 ( .A1(n59109), .A2(n50840), .ZN(n49677) );
  AOI22HSV0 U53337 ( .A1(n32168), .A2(\pe6/aot [1]), .B1(n59206), .B2(n59250), 
        .ZN(n49676) );
  NOR2HSV2 U53338 ( .A1(n49677), .A2(n49676), .ZN(n49678) );
  CLKNAND2HSV1 U53339 ( .A1(n58962), .A2(n59252), .ZN(n58544) );
  NAND2HSV0 U53340 ( .A1(n58668), .A2(n59044), .ZN(n59188) );
  NAND2HSV0 U53341 ( .A1(n59089), .A2(\pe6/aot [17]), .ZN(n49687) );
  NAND2HSV0 U53342 ( .A1(\pe6/bq[2] ), .A2(n59065), .ZN(n49686) );
  XOR2HSV0 U53343 ( .A1(n49687), .A2(n49686), .Z(n49691) );
  NAND2HSV0 U53344 ( .A1(n59084), .A2(\pe6/aot [21]), .ZN(n49689) );
  NAND2HSV0 U53345 ( .A1(n58990), .A2(n31555), .ZN(n49688) );
  XOR2HSV0 U53346 ( .A1(n49689), .A2(n49688), .Z(n49690) );
  NAND2HSV0 U53347 ( .A1(n59066), .A2(n59061), .ZN(n49693) );
  NAND2HSV0 U53348 ( .A1(n33023), .A2(n32972), .ZN(n49692) );
  XOR2HSV0 U53349 ( .A1(n49693), .A2(n49692), .Z(n49697) );
  NAND2HSV0 U53350 ( .A1(n59045), .A2(n58842), .ZN(n49695) );
  NAND2HSV0 U53351 ( .A1(n58833), .A2(n49208), .ZN(n49694) );
  XOR2HSV0 U53352 ( .A1(n49695), .A2(n49694), .Z(n49696) );
  XOR2HSV0 U53353 ( .A1(n49697), .A2(n49696), .Z(n49698) );
  NAND2HSV0 U53354 ( .A1(n59075), .A2(\pe6/aot [23]), .ZN(n49701) );
  NAND2HSV0 U53355 ( .A1(n59062), .A2(n59272), .ZN(n49700) );
  XOR2HSV0 U53356 ( .A1(n49701), .A2(n49700), .Z(n49705) );
  NAND2HSV0 U53357 ( .A1(n58731), .A2(n58824), .ZN(n49703) );
  NAND2HSV0 U53358 ( .A1(n59251), .A2(n59260), .ZN(n49702) );
  XOR2HSV0 U53359 ( .A1(n49703), .A2(n49702), .Z(n49704) );
  XOR2HSV0 U53360 ( .A1(n49705), .A2(n49704), .Z(n49713) );
  NAND2HSV0 U53361 ( .A1(\pe6/bq[17] ), .A2(\pe6/aot [13]), .ZN(n49707) );
  NAND2HSV0 U53362 ( .A1(n59202), .A2(\pe6/aot [7]), .ZN(n49706) );
  XOR2HSV0 U53363 ( .A1(n49707), .A2(n49706), .Z(n49711) );
  NOR2HSV0 U53364 ( .A1(n46850), .A2(n46637), .ZN(n49709) );
  NAND2HSV0 U53365 ( .A1(n59098), .A2(\pe6/aot [10]), .ZN(n49708) );
  XOR2HSV0 U53366 ( .A1(n49709), .A2(n49708), .Z(n49710) );
  XOR2HSV0 U53367 ( .A1(n49711), .A2(n49710), .Z(n49712) );
  XNOR2HSV1 U53368 ( .A1(n49715), .A2(n49714), .ZN(n49717) );
  CLKNAND2HSV0 U53369 ( .A1(n59144), .A2(n58811), .ZN(n49716) );
  XNOR2HSV1 U53370 ( .A1(n49717), .A2(n49716), .ZN(n49718) );
  XNOR2HSV1 U53371 ( .A1(n49719), .A2(n49718), .ZN(n49720) );
  XNOR2HSV1 U53372 ( .A1(n49721), .A2(n49720), .ZN(n49722) );
  XNOR2HSV1 U53373 ( .A1(n49723), .A2(n49722), .ZN(n49724) );
  XNOR2HSV1 U53374 ( .A1(n49725), .A2(n49724), .ZN(n49728) );
  CLKNAND2HSV1 U53375 ( .A1(n36196), .A2(n36104), .ZN(n49727) );
  XNOR2HSV1 U53376 ( .A1(n49728), .A2(n49727), .ZN(n49729) );
  XNOR2HSV1 U53377 ( .A1(n49730), .A2(n49729), .ZN(n49731) );
  XNOR2HSV1 U53378 ( .A1(n49732), .A2(n49731), .ZN(n49734) );
  CLKNAND2HSV0 U53379 ( .A1(n59335), .A2(n59328), .ZN(n49733) );
  XOR2HSV0 U53380 ( .A1(n49734), .A2(n49733), .Z(n49735) );
  NAND3HSV2 U53381 ( .A1(n46766), .A2(n53102), .A3(n59328), .ZN(n49824) );
  CLKNAND2HSV1 U53382 ( .A1(n49738), .A2(n49737), .ZN(n49828) );
  NOR2HSV1 U53383 ( .A1(n53104), .A2(n49739), .ZN(n49740) );
  CLKNAND2HSV1 U53384 ( .A1(n49828), .A2(n49740), .ZN(n49822) );
  NAND2HSV2 U53385 ( .A1(n53107), .A2(n58715), .ZN(n49818) );
  CLKNAND2HSV0 U53386 ( .A1(n58657), .A2(n59178), .ZN(n49816) );
  CLKNAND2HSV0 U53387 ( .A1(n58716), .A2(\pe6/got [15]), .ZN(n49814) );
  CLKNAND2HSV1 U53388 ( .A1(n58480), .A2(n49741), .ZN(n49811) );
  NAND2HSV0 U53389 ( .A1(n58448), .A2(\pe6/got [12]), .ZN(n49807) );
  CLKNAND2HSV1 U53390 ( .A1(n58936), .A2(n49742), .ZN(n49805) );
  CLKNAND2HSV0 U53391 ( .A1(n53111), .A2(n58658), .ZN(n49801) );
  CLKNAND2HSV1 U53392 ( .A1(n59030), .A2(n58526), .ZN(n49799) );
  CLKNAND2HSV0 U53393 ( .A1(n53113), .A2(n58562), .ZN(n49797) );
  NAND2HSV0 U53394 ( .A1(n59179), .A2(n58513), .ZN(n49795) );
  NAND2HSV0 U53395 ( .A1(n49667), .A2(n58479), .ZN(n49791) );
  CLKNAND2HSV1 U53396 ( .A1(n59379), .A2(\pe6/got [3]), .ZN(n49789) );
  NAND2HSV0 U53397 ( .A1(n58813), .A2(n59231), .ZN(n49787) );
  NAND2HSV0 U53398 ( .A1(n49743), .A2(n59235), .ZN(n49785) );
  NAND2HSV0 U53399 ( .A1(n49844), .A2(n53134), .ZN(n49745) );
  CLKNAND2HSV1 U53400 ( .A1(n58618), .A2(\pe6/aot [6]), .ZN(n58491) );
  NOR2HSV0 U53401 ( .A1(n58986), .A2(n58491), .ZN(n49744) );
  AOI21HSV2 U53402 ( .A1(n49746), .A2(n49745), .B(n49744), .ZN(n49747) );
  NOR2HSV0 U53403 ( .A1(n48887), .A2(n35864), .ZN(n58751) );
  XNOR2HSV1 U53404 ( .A1(n49747), .A2(n58751), .ZN(n49751) );
  NOR2HSV0 U53405 ( .A1(n49680), .A2(n49188), .ZN(n49749) );
  CLKNAND2HSV0 U53406 ( .A1(\pe6/bq[2] ), .A2(n59264), .ZN(n49748) );
  XOR2HSV0 U53407 ( .A1(n49749), .A2(n49748), .Z(n49750) );
  XOR2HSV0 U53408 ( .A1(n49751), .A2(n49750), .Z(n49783) );
  NAND2HSV0 U53409 ( .A1(n32606), .A2(\pe6/aot [2]), .ZN(n49753) );
  NAND2HSV0 U53410 ( .A1(n59051), .A2(n59252), .ZN(n49752) );
  XOR2HSV0 U53411 ( .A1(n49753), .A2(n49752), .Z(n49757) );
  NAND2HSV0 U53412 ( .A1(n59265), .A2(n58495), .ZN(n49755) );
  NAND2HSV0 U53413 ( .A1(n48044), .A2(\pe6/aot [13]), .ZN(n49754) );
  XOR2HSV0 U53414 ( .A1(n49755), .A2(n49754), .Z(n49756) );
  XOR2HSV0 U53415 ( .A1(n49757), .A2(n49756), .Z(n49766) );
  NOR2HSV0 U53416 ( .A1(n48042), .A2(n32858), .ZN(n49759) );
  CLKNAND2HSV0 U53417 ( .A1(n58668), .A2(n58857), .ZN(n49758) );
  XOR2HSV0 U53418 ( .A1(n49759), .A2(n49758), .Z(n49764) );
  NOR2HSV0 U53419 ( .A1(n48047), .A2(n58392), .ZN(n49761) );
  NAND2HSV2 U53420 ( .A1(n59062), .A2(\pe6/aot [7]), .ZN(n58451) );
  NAND2HSV0 U53421 ( .A1(\pe6/bq[15] ), .A2(n49760), .ZN(n59186) );
  OAI22HSV0 U53422 ( .A1(n49762), .A2(n49761), .B1(n58451), .B2(n59186), .ZN(
        n49763) );
  XNOR2HSV1 U53423 ( .A1(n49764), .A2(n49763), .ZN(n49765) );
  XNOR2HSV1 U53424 ( .A1(n49766), .A2(n49765), .ZN(n49782) );
  NAND2HSV0 U53425 ( .A1(n49862), .A2(\pe6/aot [1]), .ZN(n49768) );
  NAND2HSV0 U53426 ( .A1(n35750), .A2(\pe6/aot [11]), .ZN(n49767) );
  XOR2HSV0 U53427 ( .A1(n49768), .A2(n49767), .Z(n49772) );
  CLKNAND2HSV1 U53428 ( .A1(n59066), .A2(\pe6/aot [19]), .ZN(n49770) );
  NAND2HSV0 U53429 ( .A1(n48051), .A2(\pe6/aot [10]), .ZN(n49769) );
  XOR2HSV0 U53430 ( .A1(n49770), .A2(n49769), .Z(n49771) );
  XOR2HSV0 U53431 ( .A1(n49772), .A2(n49771), .Z(n49780) );
  NAND2HSV0 U53432 ( .A1(n59273), .A2(n58842), .ZN(n49774) );
  CLKNAND2HSV0 U53433 ( .A1(n32982), .A2(n49847), .ZN(n49773) );
  XOR2HSV0 U53434 ( .A1(n49774), .A2(n49773), .Z(n49778) );
  NOR2HSV0 U53435 ( .A1(n46146), .A2(n58851), .ZN(n49776) );
  NAND2HSV0 U53436 ( .A1(n36150), .A2(n58459), .ZN(n49775) );
  XOR2HSV0 U53437 ( .A1(n49776), .A2(n49775), .Z(n49777) );
  XOR2HSV0 U53438 ( .A1(n49778), .A2(n49777), .Z(n49779) );
  XOR2HSV0 U53439 ( .A1(n49780), .A2(n49779), .Z(n49781) );
  XOR3HSV2 U53440 ( .A1(n49783), .A2(n49782), .A3(n49781), .Z(n49784) );
  XNOR2HSV1 U53441 ( .A1(n49785), .A2(n49784), .ZN(n49786) );
  XNOR2HSV1 U53442 ( .A1(n49787), .A2(n49786), .ZN(n49788) );
  XNOR2HSV1 U53443 ( .A1(n49789), .A2(n49788), .ZN(n49790) );
  XNOR2HSV1 U53444 ( .A1(n49791), .A2(n49790), .ZN(n49793) );
  NAND2HSV0 U53445 ( .A1(n58901), .A2(n58478), .ZN(n49792) );
  XNOR2HSV1 U53446 ( .A1(n49793), .A2(n49792), .ZN(n49794) );
  XNOR2HSV1 U53447 ( .A1(n49795), .A2(n49794), .ZN(n49796) );
  XNOR2HSV1 U53448 ( .A1(n49797), .A2(n49796), .ZN(n49798) );
  XNOR2HSV1 U53449 ( .A1(n49799), .A2(n49798), .ZN(n49800) );
  XNOR2HSV1 U53450 ( .A1(n49801), .A2(n49800), .ZN(n49803) );
  NAND2HSV0 U53451 ( .A1(n58702), .A2(n58812), .ZN(n49802) );
  XNOR2HSV1 U53452 ( .A1(n49803), .A2(n49802), .ZN(n49804) );
  XNOR2HSV1 U53453 ( .A1(n49805), .A2(n49804), .ZN(n49806) );
  XNOR2HSV1 U53454 ( .A1(n49807), .A2(n49806), .ZN(n49809) );
  NAND2HSV0 U53455 ( .A1(n59161), .A2(n58811), .ZN(n49808) );
  XOR2HSV0 U53456 ( .A1(n49809), .A2(n49808), .Z(n49810) );
  XNOR2HSV1 U53457 ( .A1(n49811), .A2(n49810), .ZN(n49813) );
  NAND2HSV0 U53458 ( .A1(n53172), .A2(n59316), .ZN(n49812) );
  XOR3HSV2 U53459 ( .A1(n49814), .A2(n49813), .A3(n49812), .Z(n49815) );
  XNOR2HSV1 U53460 ( .A1(n49816), .A2(n49815), .ZN(n49817) );
  XOR2HSV0 U53461 ( .A1(n49818), .A2(n49817), .Z(n49820) );
  CLKNAND2HSV0 U53462 ( .A1(n58712), .A2(n58807), .ZN(n49819) );
  XOR2HSV0 U53463 ( .A1(n49820), .A2(n49819), .Z(n49821) );
  XOR2HSV0 U53464 ( .A1(n49822), .A2(n49821), .Z(n49823) );
  XOR2HSV0 U53465 ( .A1(n49824), .A2(n49823), .Z(\pe6/poht [11]) );
  NAND3HSV2 U53466 ( .A1(n46766), .A2(n53102), .A3(n49825), .ZN(n49920) );
  NOR2HSV1 U53467 ( .A1(n53104), .A2(n49826), .ZN(n49827) );
  CLKNAND2HSV1 U53468 ( .A1(n49828), .A2(n49827), .ZN(n49918) );
  CLKNAND2HSV0 U53469 ( .A1(n58712), .A2(n59029), .ZN(n49916) );
  NAND2HSV2 U53470 ( .A1(n53107), .A2(n58807), .ZN(n49914) );
  CLKNAND2HSV0 U53471 ( .A1(n59026), .A2(n58715), .ZN(n49912) );
  CLKNAND2HSV0 U53472 ( .A1(n58716), .A2(n58937), .ZN(n49910) );
  CLKNAND2HSV1 U53473 ( .A1(n58717), .A2(\pe6/got [15]), .ZN(n49907) );
  NAND2HSV0 U53474 ( .A1(n58448), .A2(n58811), .ZN(n49903) );
  CLKNAND2HSV1 U53475 ( .A1(n58936), .A2(n58719), .ZN(n49901) );
  CLKNAND2HSV1 U53476 ( .A1(n53111), .A2(n58812), .ZN(n49897) );
  CLKNAND2HSV1 U53477 ( .A1(n59030), .A2(n58721), .ZN(n49895) );
  CLKNAND2HSV1 U53478 ( .A1(n53113), .A2(n58526), .ZN(n49893) );
  CLKNAND2HSV1 U53479 ( .A1(n59179), .A2(n58814), .ZN(n49891) );
  CLKNAND2HSV1 U53480 ( .A1(n58722), .A2(n58384), .ZN(n49887) );
  CLKNAND2HSV1 U53481 ( .A1(n36105), .A2(\pe6/got [4]), .ZN(n49885) );
  NAND2HSV0 U53482 ( .A1(n58813), .A2(n58527), .ZN(n49883) );
  NAND2HSV0 U53483 ( .A1(n49743), .A2(n58816), .ZN(n49881) );
  NAND2HSV0 U53484 ( .A1(n49829), .A2(n58817), .ZN(n49879) );
  CLKNHSV0 U53485 ( .I(n49830), .ZN(n49834) );
  AOI22HSV0 U53486 ( .A1(n59062), .A2(\pe6/aot [19]), .B1(n49831), .B2(
        \pe6/bq[1] ), .ZN(n49832) );
  AOI21HSV2 U53487 ( .A1(n49834), .A2(n49833), .B(n49832), .ZN(n49840) );
  AOI21HSV0 U53488 ( .A1(n49205), .A2(n49836), .B(n49835), .ZN(n49838) );
  NAND2HSV0 U53489 ( .A1(n59273), .A2(n59264), .ZN(n50836) );
  NOR2HSV0 U53490 ( .A1(n50836), .A2(n53119), .ZN(n49837) );
  NOR2HSV1 U53491 ( .A1(n49838), .A2(n49837), .ZN(n49839) );
  XOR2HSV0 U53492 ( .A1(n49840), .A2(n49839), .Z(n49843) );
  NOR2HSV0 U53493 ( .A1(n46147), .A2(n58851), .ZN(n58978) );
  XOR2HSV0 U53494 ( .A1(n58978), .A2(n49841), .Z(n49842) );
  XNOR2HSV1 U53495 ( .A1(n49843), .A2(n49842), .ZN(n49877) );
  NAND2HSV0 U53496 ( .A1(n49844), .A2(\pe6/aot [7]), .ZN(n49846) );
  NAND2HSV0 U53497 ( .A1(n59089), .A2(\pe6/aot [10]), .ZN(n49845) );
  XOR2HSV0 U53498 ( .A1(n49846), .A2(n49845), .Z(n49851) );
  CLKNAND2HSV0 U53499 ( .A1(n33023), .A2(n49847), .ZN(n49849) );
  CLKNAND2HSV0 U53500 ( .A1(n32982), .A2(n58665), .ZN(n49848) );
  XOR2HSV0 U53501 ( .A1(n49849), .A2(n49848), .Z(n49850) );
  XOR2HSV0 U53502 ( .A1(n49851), .A2(n49850), .Z(n49859) );
  XOR2HSV0 U53503 ( .A1(n49853), .A2(n49852), .Z(n49857) );
  CLKNAND2HSV0 U53504 ( .A1(n58976), .A2(\pe6/aot [11]), .ZN(n49855) );
  NAND2HSV0 U53505 ( .A1(n35750), .A2(n53115), .ZN(n49854) );
  XOR2HSV0 U53506 ( .A1(n49855), .A2(n49854), .Z(n49856) );
  XNOR2HSV1 U53507 ( .A1(n49857), .A2(n49856), .ZN(n49858) );
  XNOR2HSV1 U53508 ( .A1(n49859), .A2(n49858), .ZN(n49876) );
  NAND2HSV0 U53509 ( .A1(\pe6/bq[2] ), .A2(\pe6/aot [21]), .ZN(n49861) );
  NAND2HSV0 U53510 ( .A1(n32606), .A2(n58353), .ZN(n49860) );
  XOR2HSV0 U53511 ( .A1(n49861), .A2(n49860), .Z(n49866) );
  NAND2HSV0 U53512 ( .A1(n59051), .A2(n58459), .ZN(n49864) );
  NAND2HSV0 U53513 ( .A1(n49862), .A2(n59260), .ZN(n49863) );
  XOR2HSV0 U53514 ( .A1(n49864), .A2(n49863), .Z(n49865) );
  XOR2HSV0 U53515 ( .A1(n49866), .A2(n49865), .Z(n49874) );
  NAND2HSV0 U53516 ( .A1(\pe6/bq[8] ), .A2(n58842), .ZN(n49868) );
  NAND2HSV0 U53517 ( .A1(n48044), .A2(n58943), .ZN(n49867) );
  XOR2HSV0 U53518 ( .A1(n49868), .A2(n49867), .Z(n49872) );
  NAND2HSV0 U53519 ( .A1(n58682), .A2(n35632), .ZN(n49870) );
  NAND2HSV0 U53520 ( .A1(n58668), .A2(n58495), .ZN(n49869) );
  XOR2HSV0 U53521 ( .A1(n49870), .A2(n49869), .Z(n49871) );
  XOR2HSV0 U53522 ( .A1(n49872), .A2(n49871), .Z(n49873) );
  XOR2HSV0 U53523 ( .A1(n49874), .A2(n49873), .Z(n49875) );
  XOR3HSV2 U53524 ( .A1(n49877), .A2(n49876), .A3(n49875), .Z(n49878) );
  XNOR2HSV1 U53525 ( .A1(n49879), .A2(n49878), .ZN(n49880) );
  XNOR2HSV1 U53526 ( .A1(n49881), .A2(n49880), .ZN(n49882) );
  XOR2HSV0 U53527 ( .A1(n49883), .A2(n49882), .Z(n49884) );
  XNOR2HSV1 U53528 ( .A1(n49885), .A2(n49884), .ZN(n49886) );
  XNOR2HSV1 U53529 ( .A1(n49887), .A2(n49886), .ZN(n49889) );
  CLKNAND2HSV0 U53530 ( .A1(n59144), .A2(n58659), .ZN(n49888) );
  XNOR2HSV1 U53531 ( .A1(n49889), .A2(n49888), .ZN(n49890) );
  XNOR2HSV1 U53532 ( .A1(n49891), .A2(n49890), .ZN(n49892) );
  XNOR2HSV1 U53533 ( .A1(n49893), .A2(n49892), .ZN(n49894) );
  XNOR2HSV1 U53534 ( .A1(n49895), .A2(n49894), .ZN(n49896) );
  XNOR2HSV1 U53535 ( .A1(n49897), .A2(n49896), .ZN(n49899) );
  CLKNAND2HSV0 U53536 ( .A1(n58702), .A2(n58720), .ZN(n49898) );
  XNOR2HSV1 U53537 ( .A1(n49899), .A2(n49898), .ZN(n49900) );
  XNOR2HSV1 U53538 ( .A1(n49901), .A2(n49900), .ZN(n49902) );
  XNOR2HSV1 U53539 ( .A1(n49903), .A2(n49902), .ZN(n49905) );
  NAND2HSV0 U53540 ( .A1(n58805), .A2(n58810), .ZN(n49904) );
  XOR2HSV0 U53541 ( .A1(n49905), .A2(n49904), .Z(n49906) );
  XNOR2HSV1 U53542 ( .A1(n49907), .A2(n49906), .ZN(n49909) );
  XOR3HSV2 U53543 ( .A1(n49910), .A2(n49909), .A3(n49908), .Z(n49911) );
  XNOR2HSV1 U53544 ( .A1(n49912), .A2(n49911), .ZN(n49913) );
  XNOR2HSV1 U53545 ( .A1(n49914), .A2(n49913), .ZN(n49915) );
  XNOR2HSV1 U53546 ( .A1(n49916), .A2(n49915), .ZN(n49917) );
  XOR2HSV0 U53547 ( .A1(n49918), .A2(n49917), .Z(n49919) );
  XOR2HSV0 U53548 ( .A1(n49920), .A2(n49919), .Z(\pe6/poht [10]) );
  INHSV2 U53549 ( .I(n50042), .ZN(n58052) );
  BUFHSV2 U53550 ( .I(n49921), .Z(n57983) );
  CLKNAND2HSV0 U53551 ( .A1(n57983), .A2(n59663), .ZN(n49953) );
  INHSV2 U53552 ( .I(n49967), .ZN(n58282) );
  NAND2HSV0 U53553 ( .A1(n59683), .A2(n58265), .ZN(n49924) );
  CLKNAND2HSV0 U53554 ( .A1(\pe4/aot [14]), .A2(n58301), .ZN(n49923) );
  XOR2HSV0 U53555 ( .A1(n49924), .A2(n49923), .Z(n49928) );
  NAND2HSV0 U53556 ( .A1(n57234), .A2(n58322), .ZN(n49926) );
  NAND2HSV0 U53557 ( .A1(n59857), .A2(\pe4/bq[4] ), .ZN(n49925) );
  XOR2HSV0 U53558 ( .A1(n49926), .A2(n49925), .Z(n49927) );
  NAND2HSV0 U53559 ( .A1(n59831), .A2(n58077), .ZN(n49931) );
  NAND2HSV0 U53560 ( .A1(\pe4/aot [9]), .A2(n35184), .ZN(n49930) );
  XOR2HSV0 U53561 ( .A1(n49931), .A2(n49930), .Z(n49935) );
  NAND2HSV0 U53562 ( .A1(n47718), .A2(n58003), .ZN(n49933) );
  NAND2HSV0 U53563 ( .A1(n58198), .A2(n58116), .ZN(n49932) );
  XOR2HSV0 U53564 ( .A1(n49933), .A2(n49932), .Z(n49934) );
  XOR2HSV0 U53565 ( .A1(n49935), .A2(n49934), .Z(n49936) );
  NAND2HSV0 U53566 ( .A1(n59953), .A2(\pe4/bq[2] ), .ZN(n49938) );
  NAND2HSV0 U53567 ( .A1(n57993), .A2(\pe4/bq[9] ), .ZN(n49937) );
  XOR2HSV0 U53568 ( .A1(n49938), .A2(n49937), .Z(n49942) );
  CLKNAND2HSV0 U53569 ( .A1(n58070), .A2(\pe4/bq[11] ), .ZN(n49940) );
  NAND2HSV0 U53570 ( .A1(n58199), .A2(\pe4/bq[13] ), .ZN(n49939) );
  XOR2HSV0 U53571 ( .A1(n49940), .A2(n49939), .Z(n49941) );
  XOR2HSV0 U53572 ( .A1(n49942), .A2(n49941), .Z(n49950) );
  NAND2HSV0 U53573 ( .A1(n58283), .A2(n58069), .ZN(n49945) );
  NAND2HSV0 U53574 ( .A1(n58230), .A2(n49943), .ZN(n49944) );
  XOR2HSV0 U53575 ( .A1(n49945), .A2(n49944), .Z(n49948) );
  CLKNAND2HSV0 U53576 ( .A1(n59343), .A2(n57837), .ZN(n49983) );
  CLKNAND2HSV0 U53577 ( .A1(\pe4/aot [2]), .A2(n58084), .ZN(n49946) );
  XOR2HSV0 U53578 ( .A1(n49983), .A2(n49946), .Z(n49947) );
  XOR2HSV0 U53579 ( .A1(n49948), .A2(n49947), .Z(n49949) );
  INHSV2 U53580 ( .I(n47846), .ZN(n58103) );
  XNOR2HSV1 U53581 ( .A1(n49953), .A2(n49952), .ZN(n49957) );
  CLKNAND2HSV0 U53582 ( .A1(n58141), .A2(n58153), .ZN(n49956) );
  INHSV2 U53583 ( .I(n49954), .ZN(n58110) );
  CLKNAND2HSV0 U53584 ( .A1(n57970), .A2(n58110), .ZN(n49955) );
  XOR3HSV2 U53585 ( .A1(n49957), .A2(n49956), .A3(n49955), .Z(n49959) );
  CLKNAND2HSV1 U53586 ( .A1(n58207), .A2(n35400), .ZN(n49958) );
  XNOR2HSV1 U53587 ( .A1(n49959), .A2(n49958), .ZN(n49960) );
  XNOR2HSV1 U53588 ( .A1(n49961), .A2(n49960), .ZN(n49964) );
  NOR2HSV2 U53589 ( .A1(n29774), .A2(n50212), .ZN(n49963) );
  XOR3HSV2 U53590 ( .A1(n49964), .A2(n49963), .A3(n49962), .Z(\pe4/poht [16])
         );
  NAND2HSV2 U53591 ( .A1(n50318), .A2(n59601), .ZN(n50059) );
  CLKNAND2HSV1 U53592 ( .A1(n57673), .A2(n57754), .ZN(n50051) );
  BUFHSV2 U53593 ( .I(n50065), .Z(n58112) );
  CLKNAND2HSV1 U53594 ( .A1(n58112), .A2(n59629), .ZN(n50041) );
  NAND2HSV0 U53595 ( .A1(n57675), .A2(n58102), .ZN(n50031) );
  BUFHSV2 U53596 ( .I(n59835), .Z(n57676) );
  CLKNAND2HSV1 U53597 ( .A1(n57676), .A2(n57677), .ZN(n50029) );
  NAND2HSV0 U53598 ( .A1(n59833), .A2(n58206), .ZN(n50026) );
  NAND2HSV0 U53599 ( .A1(n59682), .A2(n59346), .ZN(n50022) );
  INHSV1 U53600 ( .I(n49967), .ZN(n57680) );
  NAND2HSV0 U53601 ( .A1(n47742), .A2(n57680), .ZN(n50020) );
  NAND2HSV0 U53602 ( .A1(\pe4/aot [22]), .A2(n57798), .ZN(n57353) );
  NOR2HSV0 U53603 ( .A1(n57353), .A2(n49968), .ZN(n49970) );
  AOI22HSV0 U53604 ( .A1(\pe4/aot [22]), .A2(n58301), .B1(n57234), .B2(n57135), 
        .ZN(n49969) );
  NOR2HSV2 U53605 ( .A1(n49970), .A2(n49969), .ZN(n49975) );
  CLKNAND2HSV1 U53606 ( .A1(n58307), .A2(\pe4/bq[10] ), .ZN(n58179) );
  NOR2HSV0 U53607 ( .A1(n49971), .A2(n58179), .ZN(n49973) );
  AOI22HSV0 U53608 ( .A1(n57852), .A2(n58116), .B1(n57505), .B2(n58199), .ZN(
        n49972) );
  NOR2HSV1 U53609 ( .A1(n49973), .A2(n49972), .ZN(n49974) );
  XOR2HSV0 U53610 ( .A1(n49975), .A2(n49974), .Z(n50000) );
  NAND2HSV0 U53611 ( .A1(n57014), .A2(n58130), .ZN(n49977) );
  NAND2HSV0 U53612 ( .A1(\pe4/aot [14]), .A2(\pe4/bq[11] ), .ZN(n49976) );
  XOR2HSV0 U53613 ( .A1(n49977), .A2(n49976), .Z(n49981) );
  NOR2HSV0 U53614 ( .A1(n57025), .A2(n50114), .ZN(n49979) );
  NAND2HSV0 U53615 ( .A1(n57585), .A2(\pe4/bq[12] ), .ZN(n49978) );
  XOR2HSV0 U53616 ( .A1(n49979), .A2(n49978), .Z(n49980) );
  XNOR2HSV1 U53617 ( .A1(n49981), .A2(n49980), .ZN(n49999) );
  NOR2HSV0 U53618 ( .A1(n49982), .A2(n48032), .ZN(n57111) );
  NOR2HSV0 U53619 ( .A1(n34498), .A2(n53219), .ZN(n49984) );
  NAND2HSV0 U53620 ( .A1(n34743), .A2(n58127), .ZN(n57113) );
  OAI22HSV1 U53621 ( .A1(n57111), .A2(n49984), .B1(n57113), .B2(n49983), .ZN(
        n49990) );
  NOR2HSV0 U53622 ( .A1(n49986), .A2(n49985), .ZN(n49988) );
  AOI22HSV0 U53623 ( .A1(n50215), .A2(n57851), .B1(n50250), .B2(n59352), .ZN(
        n49987) );
  NOR2HSV1 U53624 ( .A1(n49988), .A2(n49987), .ZN(n49989) );
  XOR2HSV0 U53625 ( .A1(n49990), .A2(n49989), .Z(n49998) );
  NAND2HSV0 U53626 ( .A1(\pe4/aot [9]), .A2(\pe4/bq[16] ), .ZN(n49992) );
  NAND2HSV0 U53627 ( .A1(n57506), .A2(n57850), .ZN(n49991) );
  XOR2HSV0 U53628 ( .A1(n49992), .A2(n49991), .Z(n49996) );
  NOR2HSV0 U53629 ( .A1(n49929), .A2(n48023), .ZN(n49994) );
  NAND2HSV0 U53630 ( .A1(\pe4/aot [11]), .A2(n58126), .ZN(n49993) );
  XOR2HSV0 U53631 ( .A1(n49994), .A2(n49993), .Z(n49995) );
  XOR2HSV0 U53632 ( .A1(n49996), .A2(n49995), .Z(n49997) );
  XOR4HSV1 U53633 ( .A1(n50000), .A2(n49999), .A3(n49998), .A4(n49997), .Z(
        n50018) );
  NAND2HSV0 U53634 ( .A1(n34022), .A2(\pe4/bq[2] ), .ZN(n50002) );
  NAND2HSV0 U53635 ( .A1(\pe4/aot [7]), .A2(\pe4/bq[18] ), .ZN(n50001) );
  XOR2HSV0 U53636 ( .A1(n50002), .A2(n50001), .Z(n50006) );
  NAND2HSV0 U53637 ( .A1(n57683), .A2(n34879), .ZN(n50004) );
  NAND2HSV0 U53638 ( .A1(\pe4/aot [3]), .A2(\pe4/bq[22] ), .ZN(n50003) );
  XOR2HSV0 U53639 ( .A1(n50004), .A2(n50003), .Z(n50005) );
  XOR2HSV0 U53640 ( .A1(n50006), .A2(n50005), .Z(n50016) );
  NAND2HSV0 U53641 ( .A1(n57692), .A2(n50007), .ZN(n50010) );
  NAND2HSV0 U53642 ( .A1(\pe4/aot [21]), .A2(n57595), .ZN(n50009) );
  XOR2HSV0 U53643 ( .A1(n50010), .A2(n50009), .Z(n50014) );
  NOR2HSV0 U53644 ( .A1(n57326), .A2(n58013), .ZN(n50012) );
  NAND2HSV0 U53645 ( .A1(\pe4/aot [2]), .A2(n57476), .ZN(n50011) );
  XOR2HSV0 U53646 ( .A1(n50012), .A2(n50011), .Z(n50013) );
  XOR2HSV0 U53647 ( .A1(n50014), .A2(n50013), .Z(n50015) );
  XOR2HSV0 U53648 ( .A1(n50016), .A2(n50015), .Z(n50017) );
  XNOR2HSV1 U53649 ( .A1(n50018), .A2(n50017), .ZN(n50019) );
  XNOR2HSV1 U53650 ( .A1(n50020), .A2(n50019), .ZN(n50021) );
  XNOR2HSV1 U53651 ( .A1(n50022), .A2(n50021), .ZN(n50024) );
  NAND2HSV0 U53652 ( .A1(n34405), .A2(n58298), .ZN(n50023) );
  XNOR2HSV1 U53653 ( .A1(n50024), .A2(n50023), .ZN(n50025) );
  XNOR2HSV1 U53654 ( .A1(n50026), .A2(n50025), .ZN(n50028) );
  NAND2HSV0 U53655 ( .A1(n33918), .A2(n58137), .ZN(n50027) );
  XOR3HSV2 U53656 ( .A1(n50029), .A2(n50028), .A3(n50027), .Z(n50030) );
  XNOR2HSV1 U53657 ( .A1(n50031), .A2(n50030), .ZN(n50033) );
  NAND2HSV0 U53658 ( .A1(n57547), .A2(n58111), .ZN(n50032) );
  XNOR2HSV1 U53659 ( .A1(n50033), .A2(n50032), .ZN(n50036) );
  NAND2HSV0 U53660 ( .A1(n34409), .A2(n57818), .ZN(n50035) );
  CLKNAND2HSV1 U53661 ( .A1(n57817), .A2(\pe4/got [10]), .ZN(n50034) );
  XOR3HSV1 U53662 ( .A1(n50036), .A2(n50035), .A3(n50034), .Z(n50039) );
  CLKNAND2HSV1 U53663 ( .A1(n58096), .A2(n50189), .ZN(n50038) );
  CLKNAND2HSV0 U53664 ( .A1(n58097), .A2(\pe4/got [11]), .ZN(n50037) );
  XOR3HSV2 U53665 ( .A1(n50039), .A2(n50038), .A3(n50037), .Z(n50040) );
  XNOR2HSV1 U53666 ( .A1(n50041), .A2(n50040), .ZN(n50045) );
  CLKNAND2HSV1 U53667 ( .A1(n58183), .A2(n57982), .ZN(n50044) );
  INHSV2 U53668 ( .I(n50042), .ZN(n57674) );
  NAND2HSV0 U53669 ( .A1(n58037), .A2(n57674), .ZN(n50043) );
  XOR3HSV2 U53670 ( .A1(n50045), .A2(n50044), .A3(n50043), .Z(n50047) );
  CLKNAND2HSV1 U53671 ( .A1(n58220), .A2(n57189), .ZN(n50046) );
  XNOR2HSV1 U53672 ( .A1(n50047), .A2(n50046), .ZN(n50049) );
  CLKNAND2HSV0 U53673 ( .A1(n57755), .A2(n57457), .ZN(n50048) );
  XNOR2HSV1 U53674 ( .A1(n50049), .A2(n50048), .ZN(n50050) );
  XNOR2HSV1 U53675 ( .A1(n50051), .A2(n50050), .ZN(n50055) );
  INHSV2 U53676 ( .I(n50052), .ZN(n57770) );
  CLKNAND2HSV1 U53677 ( .A1(n58048), .A2(n57770), .ZN(n50054) );
  NAND2HSV0 U53678 ( .A1(n57564), .A2(n50199), .ZN(n50053) );
  XOR3HSV2 U53679 ( .A1(n50055), .A2(n50054), .A3(n50053), .Z(n50057) );
  INHSV2 U53680 ( .I(n50207), .ZN(n57760) );
  CLKNAND2HSV1 U53681 ( .A1(n25843), .A2(n57760), .ZN(n50056) );
  XNOR2HSV1 U53682 ( .A1(n50057), .A2(n50056), .ZN(n50058) );
  XNOR2HSV1 U53683 ( .A1(n50059), .A2(n50058), .ZN(n50063) );
  XOR3HSV2 U53684 ( .A1(n50063), .A2(n50062), .A3(n50061), .Z(\pe4/poht [8])
         );
  INHSV2 U53685 ( .I(n50064), .ZN(n58036) );
  CLKNAND2HSV1 U53686 ( .A1(n58141), .A2(n58036), .ZN(n50101) );
  CLKNAND2HSV0 U53687 ( .A1(n57983), .A2(n58184), .ZN(n50099) );
  NAND2HSV0 U53688 ( .A1(n50065), .A2(n58219), .ZN(n50087) );
  NAND2HSV2 U53689 ( .A1(n58199), .A2(\pe4/bq[9] ), .ZN(n50067) );
  NAND2HSV0 U53690 ( .A1(\pe4/aot [12]), .A2(n58322), .ZN(n50066) );
  XOR2HSV0 U53691 ( .A1(n50067), .A2(n50066), .Z(n50071) );
  CLKNAND2HSV0 U53692 ( .A1(\pe4/aot [2]), .A2(\pe4/bq[11] ), .ZN(n50069) );
  NAND2HSV0 U53693 ( .A1(\pe4/aot [10]), .A2(n58301), .ZN(n50068) );
  XOR2HSV0 U53694 ( .A1(n50069), .A2(n50068), .Z(n50070) );
  XOR2HSV0 U53695 ( .A1(n50071), .A2(n50070), .Z(n50079) );
  NAND2HSV0 U53696 ( .A1(n57692), .A2(n58077), .ZN(n50073) );
  CLKNAND2HSV0 U53697 ( .A1(n58306), .A2(n58130), .ZN(n50072) );
  XOR2HSV0 U53698 ( .A1(n50073), .A2(n50072), .Z(n50077) );
  CLKNAND2HSV1 U53699 ( .A1(n58070), .A2(n58003), .ZN(n50075) );
  NAND2HSV0 U53700 ( .A1(\pe4/aot [9]), .A2(\pe4/bq[4] ), .ZN(n50074) );
  XOR2HSV0 U53701 ( .A1(n50075), .A2(n50074), .Z(n50076) );
  XOR2HSV0 U53702 ( .A1(n50077), .A2(n50076), .Z(n50078) );
  XOR2HSV0 U53703 ( .A1(n50079), .A2(n50078), .Z(n50085) );
  NAND2HSV2 U53704 ( .A1(n58198), .A2(n57784), .ZN(n50349) );
  CLKNAND2HSV1 U53705 ( .A1(\pe4/aot [3]), .A2(n58116), .ZN(n50341) );
  XOR2HSV0 U53706 ( .A1(n50349), .A2(n50341), .Z(n50083) );
  NAND2HSV2 U53707 ( .A1(n57993), .A2(n58010), .ZN(n50081) );
  NAND2HSV0 U53708 ( .A1(n59683), .A2(\pe4/bq[2] ), .ZN(n50080) );
  XOR2HSV0 U53709 ( .A1(n50081), .A2(n50080), .Z(n50082) );
  XOR2HSV0 U53710 ( .A1(n50083), .A2(n50082), .Z(n50084) );
  XNOR2HSV1 U53711 ( .A1(n50085), .A2(n50084), .ZN(n50086) );
  XOR2HSV0 U53712 ( .A1(n50087), .A2(n50086), .Z(n50090) );
  CLKNAND2HSV1 U53713 ( .A1(n57819), .A2(n58298), .ZN(n50089) );
  CLKNAND2HSV0 U53714 ( .A1(n58037), .A2(n59346), .ZN(n50088) );
  XOR3HSV2 U53715 ( .A1(n50090), .A2(n50089), .A3(n50088), .Z(n50093) );
  INHSV2 U53716 ( .I(n50091), .ZN(n58030) );
  CLKNAND2HSV1 U53717 ( .A1(n58103), .A2(n58030), .ZN(n50092) );
  XNOR2HSV1 U53718 ( .A1(n50093), .A2(n50092), .ZN(n50097) );
  INHSV2 U53719 ( .I(n50095), .ZN(n57951) );
  CLKNAND2HSV0 U53720 ( .A1(n58185), .A2(n57951), .ZN(n50096) );
  XNOR2HSV1 U53721 ( .A1(n50097), .A2(n50096), .ZN(n50098) );
  XOR2HSV0 U53722 ( .A1(n50099), .A2(n50098), .Z(n50100) );
  NAND2HSV0 U53723 ( .A1(n58111), .A2(n50199), .ZN(n50102) );
  CLKNHSV0 U53724 ( .I(n57836), .ZN(n57413) );
  CLKNAND2HSV1 U53725 ( .A1(n58207), .A2(n57413), .ZN(n50104) );
  XOR2HSV0 U53726 ( .A1(n50105), .A2(n50104), .Z(n50106) );
  XNOR2HSV1 U53727 ( .A1(n50107), .A2(n50106), .ZN(n50110) );
  NOR2HSV2 U53728 ( .A1(n26761), .A2(n49954), .ZN(n50108) );
  XOR3HSV2 U53729 ( .A1(n50110), .A2(n50109), .A3(n50108), .Z(\pe4/poht [20])
         );
  NAND2HSV0 U53730 ( .A1(n58223), .A2(n57498), .ZN(n50113) );
  CLKNAND2HSV0 U53731 ( .A1(n58070), .A2(n58196), .ZN(n50112) );
  NAND2HSV0 U53732 ( .A1(n58230), .A2(n58130), .ZN(n50116) );
  CLKNHSV0 U53733 ( .I(n50114), .ZN(n57684) );
  NAND2HSV0 U53734 ( .A1(\pe4/aot [2]), .A2(n57684), .ZN(n50115) );
  XOR2HSV0 U53735 ( .A1(n50116), .A2(n50115), .Z(n50117) );
  NAND2HSV0 U53736 ( .A1(n58283), .A2(n58265), .ZN(n50119) );
  NAND2HSV0 U53737 ( .A1(n58199), .A2(n58155), .ZN(n50118) );
  NAND2HSV0 U53738 ( .A1(n50251), .A2(\pe4/bq[1] ), .ZN(n50121) );
  NAND2HSV0 U53739 ( .A1(n58198), .A2(\pe4/bq[2] ), .ZN(n50120) );
  XOR3HSV2 U53740 ( .A1(n50126), .A2(n50125), .A3(n50124), .Z(\pe4/poht [24])
         );
  NAND2HSV2 U53741 ( .A1(n26417), .A2(n57564), .ZN(n50206) );
  CLKNAND2HSV1 U53742 ( .A1(n57673), .A2(n57974), .ZN(n50198) );
  BUFHSV2 U53743 ( .I(n50065), .Z(n58154) );
  CLKNAND2HSV1 U53744 ( .A1(n58154), .A2(\pe4/got [11]), .ZN(n50188) );
  NAND2HSV0 U53745 ( .A1(n59378), .A2(n57677), .ZN(n50178) );
  NAND2HSV0 U53746 ( .A1(n59835), .A2(n58298), .ZN(n50176) );
  NAND2HSV0 U53747 ( .A1(n59833), .A2(n58314), .ZN(n50173) );
  NAND2HSV2 U53748 ( .A1(n57183), .A2(n57680), .ZN(n50171) );
  NAND2HSV0 U53749 ( .A1(\pe4/aot [5]), .A2(\pe4/bq[18] ), .ZN(n50128) );
  NAND2HSV0 U53750 ( .A1(\pe4/aot [6]), .A2(n57926), .ZN(n50127) );
  XOR2HSV0 U53751 ( .A1(n50128), .A2(n50127), .Z(n50133) );
  NAND2HSV2 U53752 ( .A1(n57692), .A2(n58010), .ZN(n58304) );
  NAND2HSV0 U53753 ( .A1(n33867), .A2(n57837), .ZN(n57027) );
  OAI21HSV0 U53754 ( .A1(n47905), .A2(n50129), .B(n57027), .ZN(n50130) );
  OAI21HSV0 U53755 ( .A1(n58304), .A2(n50131), .B(n50130), .ZN(n50132) );
  XNOR2HSV1 U53756 ( .A1(n50133), .A2(n50132), .ZN(n50138) );
  NOR2HSV0 U53757 ( .A1(n50134), .A2(n58013), .ZN(n50136) );
  NAND2HSV0 U53758 ( .A1(n57859), .A2(n57595), .ZN(n50135) );
  XOR2HSV0 U53759 ( .A1(n50136), .A2(n50135), .Z(n50137) );
  XNOR2HSV1 U53760 ( .A1(n50138), .A2(n50137), .ZN(n50169) );
  NAND2HSV0 U53761 ( .A1(n57234), .A2(n57684), .ZN(n50140) );
  NAND2HSV0 U53762 ( .A1(\pe4/aot [9]), .A2(n58126), .ZN(n50139) );
  XOR2HSV0 U53763 ( .A1(n50140), .A2(n50139), .Z(n50144) );
  NAND2HSV0 U53764 ( .A1(n57014), .A2(n57784), .ZN(n50142) );
  NAND2HSV0 U53765 ( .A1(n59839), .A2(n58301), .ZN(n50141) );
  XOR2HSV0 U53766 ( .A1(n50142), .A2(n50141), .Z(n50143) );
  XOR2HSV0 U53767 ( .A1(n50144), .A2(n50143), .Z(n50152) );
  NAND2HSV0 U53768 ( .A1(n59683), .A2(\pe4/bq[12] ), .ZN(n50146) );
  NAND2HSV0 U53769 ( .A1(n59343), .A2(\pe4/bq[11] ), .ZN(n50145) );
  XOR2HSV0 U53770 ( .A1(n50146), .A2(n50145), .Z(n50150) );
  NAND2HSV0 U53771 ( .A1(n35347), .A2(n58130), .ZN(n50148) );
  NAND2HSV0 U53772 ( .A1(\pe4/aot [14]), .A2(n57135), .ZN(n50147) );
  XOR2HSV0 U53773 ( .A1(n50148), .A2(n50147), .Z(n50149) );
  XOR2HSV0 U53774 ( .A1(n50150), .A2(n50149), .Z(n50151) );
  XOR2HSV0 U53775 ( .A1(n50152), .A2(n50151), .Z(n50168) );
  NAND2HSV0 U53776 ( .A1(n57585), .A2(n58116), .ZN(n50154) );
  NAND2HSV0 U53777 ( .A1(\pe4/aot [7]), .A2(n49943), .ZN(n50153) );
  XOR2HSV0 U53778 ( .A1(n50154), .A2(n50153), .Z(n50158) );
  NAND2HSV0 U53779 ( .A1(\pe4/aot [4]), .A2(n50250), .ZN(n50156) );
  NAND2HSV0 U53780 ( .A1(n58283), .A2(n57785), .ZN(n50155) );
  XOR2HSV0 U53781 ( .A1(n50156), .A2(n50155), .Z(n50157) );
  XOR2HSV0 U53782 ( .A1(n50158), .A2(n50157), .Z(n50166) );
  NAND2HSV0 U53783 ( .A1(n57683), .A2(n58127), .ZN(n50160) );
  NAND2HSV0 U53784 ( .A1(n58087), .A2(n34879), .ZN(n50159) );
  XOR2HSV0 U53785 ( .A1(n50160), .A2(n50159), .Z(n50164) );
  NAND2HSV0 U53786 ( .A1(n59951), .A2(\pe4/bq[2] ), .ZN(n50162) );
  NAND2HSV0 U53787 ( .A1(\pe4/aot [2]), .A2(n33969), .ZN(n50161) );
  XOR2HSV0 U53788 ( .A1(n50162), .A2(n50161), .Z(n50163) );
  XOR2HSV0 U53789 ( .A1(n50164), .A2(n50163), .Z(n50165) );
  XOR2HSV0 U53790 ( .A1(n50166), .A2(n50165), .Z(n50167) );
  XOR3HSV2 U53791 ( .A1(n50169), .A2(n50168), .A3(n50167), .Z(n50170) );
  XNOR2HSV1 U53792 ( .A1(n50171), .A2(n50170), .ZN(n50172) );
  XNOR2HSV1 U53793 ( .A1(n50173), .A2(n50172), .ZN(n50175) );
  NAND2HSV0 U53794 ( .A1(n34949), .A2(n58206), .ZN(n50174) );
  XOR3HSV2 U53795 ( .A1(n50176), .A2(n50175), .A3(n50174), .Z(n50177) );
  XNOR2HSV1 U53796 ( .A1(n50178), .A2(n50177), .ZN(n50180) );
  NAND2HSV0 U53797 ( .A1(n59932), .A2(n58184), .ZN(n50179) );
  XNOR2HSV1 U53798 ( .A1(n50180), .A2(n50179), .ZN(n50183) );
  NAND2HSV0 U53799 ( .A1(n57550), .A2(n58102), .ZN(n50182) );
  BUFHSV2 U53800 ( .I(n58060), .Z(n57427) );
  CLKNAND2HSV1 U53801 ( .A1(n57427), .A2(n57177), .ZN(n50181) );
  XOR3HSV1 U53802 ( .A1(n50183), .A2(n50182), .A3(n50181), .Z(n50186) );
  CLKNAND2HSV1 U53803 ( .A1(n58096), .A2(n59663), .ZN(n50185) );
  CLKNAND2HSV0 U53804 ( .A1(n58097), .A2(n57818), .ZN(n50184) );
  XOR3HSV2 U53805 ( .A1(n50186), .A2(n50185), .A3(n50184), .Z(n50187) );
  XNOR2HSV1 U53806 ( .A1(n50188), .A2(n50187), .ZN(n50192) );
  CLKNAND2HSV0 U53807 ( .A1(n58183), .A2(n59629), .ZN(n50191) );
  CLKNAND2HSV0 U53808 ( .A1(n58037), .A2(n50189), .ZN(n50190) );
  XOR3HSV2 U53809 ( .A1(n50192), .A2(n50191), .A3(n50190), .Z(n50194) );
  CLKNAND2HSV0 U53810 ( .A1(n57889), .A2(n58052), .ZN(n50193) );
  XNOR2HSV1 U53811 ( .A1(n50194), .A2(n50193), .ZN(n50196) );
  CLKNAND2HSV0 U53812 ( .A1(n57310), .A2(n57307), .ZN(n50195) );
  XNOR2HSV1 U53813 ( .A1(n50196), .A2(n50195), .ZN(n50197) );
  XNOR2HSV1 U53814 ( .A1(n50198), .A2(n50197), .ZN(n50202) );
  INHSV2 U53815 ( .I(n50211), .ZN(n58217) );
  CLKNAND2HSV1 U53816 ( .A1(n58217), .A2(n34797), .ZN(n50201) );
  NAND2HSV0 U53817 ( .A1(n50199), .A2(n57754), .ZN(n50200) );
  XOR3HSV2 U53818 ( .A1(n50202), .A2(n50201), .A3(n50200), .Z(n50204) );
  NAND2HSV0 U53819 ( .A1(n58186), .A2(n57770), .ZN(n50203) );
  XOR2HSV0 U53820 ( .A1(n50204), .A2(n50203), .Z(n50205) );
  XOR2HSV0 U53821 ( .A1(n50206), .A2(n50205), .Z(n50210) );
  NOR2HSV2 U53822 ( .A1(n26761), .A2(n49965), .ZN(n50208) );
  XOR3HSV2 U53823 ( .A1(n50210), .A2(n50209), .A3(n50208), .Z(\pe4/poht [10])
         );
  NAND2HSV2 U53824 ( .A1(n50318), .A2(n57574), .ZN(n50313) );
  CLKNAND2HSV1 U53825 ( .A1(n58141), .A2(n34594), .ZN(n50307) );
  CLKNAND2HSV0 U53826 ( .A1(n58193), .A2(n33831), .ZN(n50305) );
  NAND2HSV0 U53827 ( .A1(n50213), .A2(n57752), .ZN(n50293) );
  NAND2HSV0 U53828 ( .A1(n57675), .A2(n57413), .ZN(n50282) );
  NAND2HSV0 U53829 ( .A1(n59835), .A2(n58102), .ZN(n50280) );
  BUFHSV2 U53830 ( .I(n59833), .Z(n57678) );
  NAND2HSV0 U53831 ( .A1(n57678), .A2(n58137), .ZN(n50277) );
  NAND2HSV0 U53832 ( .A1(n57458), .A2(n57744), .ZN(n50273) );
  NAND2HSV0 U53833 ( .A1(n50215), .A2(n35184), .ZN(n50217) );
  NAND2HSV0 U53834 ( .A1(n59661), .A2(n57241), .ZN(n50216) );
  XOR2HSV0 U53835 ( .A1(n50217), .A2(n50216), .Z(n50221) );
  NAND2HSV0 U53836 ( .A1(\pe4/aot [11]), .A2(\pe4/bq[16] ), .ZN(n50219) );
  NAND2HSV0 U53837 ( .A1(n34873), .A2(n58084), .ZN(n50218) );
  XOR2HSV0 U53838 ( .A1(n50219), .A2(n50218), .Z(n50220) );
  XOR2HSV0 U53839 ( .A1(n50221), .A2(n50220), .Z(n50229) );
  NAND2HSV0 U53840 ( .A1(n59838), .A2(\pe4/bq[2] ), .ZN(n50223) );
  NAND2HSV0 U53841 ( .A1(\pe4/aot [22]), .A2(n58010), .ZN(n50222) );
  XOR2HSV0 U53842 ( .A1(n50223), .A2(n50222), .Z(n50227) );
  NAND2HSV0 U53843 ( .A1(\pe4/aot [15]), .A2(n58077), .ZN(n50225) );
  NAND2HSV0 U53844 ( .A1(\pe4/aot [14]), .A2(n58127), .ZN(n50224) );
  XOR2HSV0 U53845 ( .A1(n50225), .A2(n50224), .Z(n50226) );
  XOR2HSV0 U53846 ( .A1(n50227), .A2(n50226), .Z(n50228) );
  XOR2HSV0 U53847 ( .A1(n50229), .A2(n50228), .Z(n50245) );
  NAND2HSV0 U53848 ( .A1(\pe4/aot [2]), .A2(n57459), .ZN(n50231) );
  NAND2HSV0 U53849 ( .A1(n33867), .A2(n57798), .ZN(n50230) );
  XOR2HSV0 U53850 ( .A1(n50231), .A2(n50230), .Z(n50235) );
  NAND2HSV0 U53851 ( .A1(\pe4/aot [17]), .A2(n58116), .ZN(n50233) );
  NAND2HSV0 U53852 ( .A1(n58223), .A2(\pe4/bq[22] ), .ZN(n50232) );
  XOR2HSV0 U53853 ( .A1(n50233), .A2(n50232), .Z(n50234) );
  XOR2HSV0 U53854 ( .A1(n50235), .A2(n50234), .Z(n50243) );
  NAND2HSV0 U53855 ( .A1(\pe4/aot [6]), .A2(n57505), .ZN(n50237) );
  NAND2HSV0 U53856 ( .A1(n58198), .A2(n57785), .ZN(n50236) );
  XOR2HSV0 U53857 ( .A1(n50237), .A2(n50236), .Z(n50241) );
  NAND2HSV0 U53858 ( .A1(n57234), .A2(\pe4/bq[11] ), .ZN(n50239) );
  NAND2HSV0 U53859 ( .A1(n47718), .A2(n57850), .ZN(n50238) );
  XOR2HSV0 U53860 ( .A1(n50239), .A2(n50238), .Z(n50240) );
  XOR2HSV0 U53861 ( .A1(n50241), .A2(n50240), .Z(n50242) );
  XOR2HSV0 U53862 ( .A1(n50243), .A2(n50242), .Z(n50244) );
  XOR2HSV0 U53863 ( .A1(n50245), .A2(n50244), .Z(n50265) );
  NAND2HSV0 U53864 ( .A1(n57384), .A2(n57498), .ZN(n50247) );
  NAND2HSV0 U53865 ( .A1(\pe4/aot [24]), .A2(\pe4/bq[3] ), .ZN(n50246) );
  XOR2HSV0 U53866 ( .A1(n50247), .A2(n50246), .Z(n50263) );
  NOR2HSV0 U53867 ( .A1(n57011), .A2(n34276), .ZN(n50340) );
  NOR2HSV0 U53868 ( .A1(n58194), .A2(n50248), .ZN(n57723) );
  AOI22HSV0 U53869 ( .A1(n58307), .A2(n57592), .B1(n33712), .B2(n58283), .ZN(
        n50249) );
  AOI21HSV2 U53870 ( .A1(n50340), .A2(n57723), .B(n50249), .ZN(n50254) );
  NOR2HSV0 U53871 ( .A1(n57775), .A2(n48026), .ZN(n57718) );
  NOR2HSV0 U53872 ( .A1(n57707), .A2(n48022), .ZN(n50364) );
  NOR2HSV0 U53873 ( .A1(n57707), .A2(n48026), .ZN(n57843) );
  AOI21HSV0 U53874 ( .A1(n50251), .A2(n50250), .B(n57843), .ZN(n50252) );
  AOI21HSV1 U53875 ( .A1(n57718), .A2(n50364), .B(n50252), .ZN(n50253) );
  XOR2HSV0 U53876 ( .A1(n50254), .A2(n50253), .Z(n50262) );
  NAND2HSV0 U53877 ( .A1(n57463), .A2(n58126), .ZN(n50256) );
  NAND2HSV0 U53878 ( .A1(\pe4/aot [1]), .A2(n57460), .ZN(n50255) );
  XOR2HSV0 U53879 ( .A1(n50256), .A2(n50255), .Z(n50260) );
  NAND2HSV0 U53880 ( .A1(n59951), .A2(n57851), .ZN(n50258) );
  NAND2HSV0 U53881 ( .A1(n59839), .A2(n58197), .ZN(n50257) );
  XOR2HSV0 U53882 ( .A1(n50258), .A2(n50257), .Z(n50259) );
  XOR2HSV0 U53883 ( .A1(n50260), .A2(n50259), .Z(n50261) );
  XOR3HSV2 U53884 ( .A1(n50263), .A2(n50262), .A3(n50261), .Z(n50264) );
  XNOR2HSV1 U53885 ( .A1(n50265), .A2(n50264), .ZN(n50269) );
  NAND2HSV0 U53886 ( .A1(n50266), .A2(n57680), .ZN(n50268) );
  NAND2HSV0 U53887 ( .A1(n59681), .A2(n59346), .ZN(n50267) );
  XOR3HSV2 U53888 ( .A1(n50269), .A2(n50268), .A3(n50267), .Z(n50271) );
  NAND2HSV0 U53889 ( .A1(n47742), .A2(n57584), .ZN(n50270) );
  XOR2HSV0 U53890 ( .A1(n50271), .A2(n50270), .Z(n50272) );
  XNOR2HSV1 U53891 ( .A1(n50273), .A2(n50272), .ZN(n50275) );
  CLKNAND2HSV1 U53892 ( .A1(n34405), .A2(\pe4/got [5]), .ZN(n50274) );
  XNOR2HSV1 U53893 ( .A1(n50275), .A2(n50274), .ZN(n50276) );
  XNOR2HSV1 U53894 ( .A1(n50277), .A2(n50276), .ZN(n50279) );
  NAND2HSV0 U53895 ( .A1(n59845), .A2(\pe4/got [8]), .ZN(n50278) );
  XOR3HSV2 U53896 ( .A1(n50280), .A2(n50279), .A3(n50278), .Z(n50281) );
  XNOR2HSV1 U53897 ( .A1(n50282), .A2(n50281), .ZN(n50284) );
  NAND2HSV0 U53898 ( .A1(n59932), .A2(n59663), .ZN(n50283) );
  XNOR2HSV1 U53899 ( .A1(n50284), .A2(n50283), .ZN(n50287) );
  NAND2HSV0 U53900 ( .A1(n57550), .A2(n58153), .ZN(n50286) );
  CLKNAND2HSV1 U53901 ( .A1(n58060), .A2(n57888), .ZN(n50285) );
  XOR3HSV1 U53902 ( .A1(n50287), .A2(n50286), .A3(n50285), .Z(n50291) );
  CLKNAND2HSV1 U53903 ( .A1(n57308), .A2(n57674), .ZN(n50290) );
  BUFHSV2 U53904 ( .I(n50288), .Z(n57554) );
  CLKNAND2HSV0 U53905 ( .A1(n57554), .A2(n47657), .ZN(n50289) );
  XOR3HSV2 U53906 ( .A1(n50291), .A2(n50290), .A3(n50289), .Z(n50292) );
  XNOR2HSV1 U53907 ( .A1(n50293), .A2(n50292), .ZN(n50297) );
  INHSV2 U53908 ( .I(n47861), .ZN(n57457) );
  CLKNAND2HSV0 U53909 ( .A1(n47841), .A2(n57457), .ZN(n50296) );
  NAND2HSV0 U53910 ( .A1(n57560), .A2(n59604), .ZN(n50295) );
  XOR3HSV2 U53911 ( .A1(n50297), .A2(n50296), .A3(n50295), .Z(n50300) );
  CLKNAND2HSV0 U53912 ( .A1(n25427), .A2(n57754), .ZN(n50299) );
  XNOR2HSV1 U53913 ( .A1(n50300), .A2(n50299), .ZN(n50303) );
  NAND2HSV0 U53914 ( .A1(n57755), .A2(n57770), .ZN(n50302) );
  XNOR2HSV1 U53915 ( .A1(n50303), .A2(n50302), .ZN(n50304) );
  XNOR2HSV1 U53916 ( .A1(n50305), .A2(n50304), .ZN(n50306) );
  XOR2HSV0 U53917 ( .A1(n50307), .A2(n50306), .Z(n50309) );
  CLKNAND2HSV0 U53918 ( .A1(n57970), .A2(n59601), .ZN(n50308) );
  XNOR2HSV1 U53919 ( .A1(n50309), .A2(n50308), .ZN(n50311) );
  XOR2HSV0 U53920 ( .A1(n50311), .A2(n50310), .Z(n50312) );
  XNOR2HSV1 U53921 ( .A1(n50313), .A2(n50312), .ZN(n50317) );
  NOR2HSV2 U53922 ( .A1(n29774), .A2(n50314), .ZN(n50316) );
  XOR3HSV2 U53923 ( .A1(n50317), .A2(n50316), .A3(n50315), .Z(\pe4/poht [6])
         );
  NAND2HSV2 U53924 ( .A1(n26417), .A2(n35318), .ZN(n50417) );
  CLKNAND2HSV1 U53925 ( .A1(n57673), .A2(n34594), .ZN(n50410) );
  CLKNAND2HSV1 U53926 ( .A1(n50213), .A2(n47656), .ZN(n50399) );
  NAND2HSV0 U53927 ( .A1(n57675), .A2(n57646), .ZN(n50389) );
  NAND2HSV0 U53928 ( .A1(n59835), .A2(\pe4/got [8]), .ZN(n50387) );
  NAND2HSV0 U53929 ( .A1(n57678), .A2(n58102), .ZN(n50383) );
  NAND2HSV0 U53930 ( .A1(n59667), .A2(n59346), .ZN(n50374) );
  NAND2HSV0 U53931 ( .A1(n33498), .A2(n57680), .ZN(n50372) );
  NAND2HSV0 U53932 ( .A1(n57234), .A2(n57986), .ZN(n50320) );
  NAND2HSV0 U53933 ( .A1(n57683), .A2(n57906), .ZN(n50319) );
  XOR2HSV0 U53934 ( .A1(n50320), .A2(n50319), .Z(n50324) );
  NAND2HSV0 U53935 ( .A1(n34743), .A2(\pe4/bq[8] ), .ZN(n50322) );
  NAND2HSV0 U53936 ( .A1(n59951), .A2(n57684), .ZN(n50321) );
  XOR2HSV0 U53937 ( .A1(n50322), .A2(n50321), .Z(n50323) );
  XOR2HSV0 U53938 ( .A1(n50324), .A2(n50323), .Z(n50332) );
  NAND2HSV0 U53939 ( .A1(n34873), .A2(\pe4/bq[16] ), .ZN(n50326) );
  NAND2HSV0 U53940 ( .A1(n57499), .A2(\pe4/bq[3] ), .ZN(n50325) );
  XOR2HSV0 U53941 ( .A1(n50326), .A2(n50325), .Z(n50330) );
  NAND2HSV0 U53942 ( .A1(\pe4/aot [6]), .A2(\pe4/bq[22] ), .ZN(n50328) );
  NAND2HSV0 U53943 ( .A1(n57140), .A2(n57798), .ZN(n50327) );
  XOR2HSV0 U53944 ( .A1(n50328), .A2(n50327), .Z(n50329) );
  XNOR2HSV1 U53945 ( .A1(n50330), .A2(n50329), .ZN(n50331) );
  XNOR2HSV1 U53946 ( .A1(n50332), .A2(n50331), .ZN(n50348) );
  NAND2HSV0 U53947 ( .A1(n59831), .A2(n57592), .ZN(n50334) );
  NAND2HSV0 U53948 ( .A1(\pe4/aot [24]), .A2(n57498), .ZN(n50333) );
  XOR2HSV0 U53949 ( .A1(n50334), .A2(n50333), .Z(n50338) );
  NAND2HSV0 U53950 ( .A1(n57463), .A2(n57348), .ZN(n50336) );
  NAND2HSV0 U53951 ( .A1(\pe4/aot [2]), .A2(n57460), .ZN(n50335) );
  XOR2HSV0 U53952 ( .A1(n50336), .A2(n50335), .Z(n50337) );
  XNOR2HSV1 U53953 ( .A1(n50338), .A2(n50337), .ZN(n50346) );
  NAND2HSV2 U53954 ( .A1(n58307), .A2(n57241), .ZN(n58287) );
  XOR2HSV0 U53955 ( .A1(n50344), .A2(n50343), .Z(n50345) );
  XNOR2HSV1 U53956 ( .A1(n50346), .A2(n50345), .ZN(n50347) );
  XNOR2HSV1 U53957 ( .A1(n50348), .A2(n50347), .ZN(n50370) );
  NOR2HSV0 U53958 ( .A1(n50350), .A2(n50349), .ZN(n50353) );
  CLKNHSV0 U53959 ( .I(n50351), .ZN(n58195) );
  AOI22HSV0 U53960 ( .A1(\pe4/aot [22]), .A2(n58195), .B1(n34636), .B2(n58198), 
        .ZN(n50352) );
  NOR2HSV2 U53961 ( .A1(n50353), .A2(n50352), .ZN(n50359) );
  NOR2HSV0 U53962 ( .A1(n50355), .A2(n50354), .ZN(n50357) );
  AOI22HSV0 U53963 ( .A1(n57327), .A2(\pe4/bq[2] ), .B1(n57014), .B2(
        \pe4/bq[11] ), .ZN(n50356) );
  NOR2HSV2 U53964 ( .A1(n50357), .A2(n50356), .ZN(n50358) );
  XNOR2HSV1 U53965 ( .A1(n50359), .A2(n50358), .ZN(n50362) );
  NAND2HSV0 U53966 ( .A1(\pe4/aot [1]), .A2(n57850), .ZN(n57988) );
  NOR2HSV0 U53967 ( .A1(n57918), .A2(n53219), .ZN(n57016) );
  XNOR2HSV1 U53968 ( .A1(n50362), .A2(n50361), .ZN(n50368) );
  NAND2HSV0 U53969 ( .A1(n57506), .A2(n57785), .ZN(n57717) );
  XOR2HSV0 U53970 ( .A1(n50363), .A2(n57717), .Z(n50366) );
  NAND2HSV0 U53971 ( .A1(n57384), .A2(n57837), .ZN(n57493) );
  XOR2HSV0 U53972 ( .A1(n50364), .A2(n57493), .Z(n50365) );
  XOR2HSV0 U53973 ( .A1(n50366), .A2(n50365), .Z(n50367) );
  XOR2HSV0 U53974 ( .A1(n50368), .A2(n50367), .Z(n50369) );
  XNOR2HSV1 U53975 ( .A1(n50370), .A2(n50369), .ZN(n50371) );
  XNOR2HSV1 U53976 ( .A1(n50372), .A2(n50371), .ZN(n50373) );
  XNOR2HSV1 U53977 ( .A1(n50374), .A2(n50373), .ZN(n50376) );
  NAND2HSV0 U53978 ( .A1(n59681), .A2(n57584), .ZN(n50375) );
  XNOR2HSV1 U53979 ( .A1(n50376), .A2(n50375), .ZN(n50378) );
  NAND2HSV0 U53980 ( .A1(n57679), .A2(n57744), .ZN(n50377) );
  XOR2HSV0 U53981 ( .A1(n50378), .A2(n50377), .Z(n50381) );
  NAND2HSV0 U53982 ( .A1(n59682), .A2(\pe4/got [5]), .ZN(n50380) );
  NAND2HSV0 U53983 ( .A1(n57183), .A2(n58137), .ZN(n50379) );
  XOR3HSV1 U53984 ( .A1(n50381), .A2(n50380), .A3(n50379), .Z(n50382) );
  XNOR2HSV1 U53985 ( .A1(n50383), .A2(n50382), .ZN(n50386) );
  XOR3HSV2 U53986 ( .A1(n50387), .A2(n50386), .A3(n50385), .Z(n50388) );
  XNOR2HSV1 U53987 ( .A1(n50389), .A2(n50388), .ZN(n50391) );
  NAND2HSV0 U53988 ( .A1(n57985), .A2(n58153), .ZN(n50390) );
  XNOR2HSV1 U53989 ( .A1(n50391), .A2(n50390), .ZN(n50394) );
  NAND2HSV0 U53990 ( .A1(n57550), .A2(n50189), .ZN(n50393) );
  CLKNAND2HSV1 U53991 ( .A1(n29758), .A2(n47657), .ZN(n50392) );
  XOR3HSV1 U53992 ( .A1(n50394), .A2(n50393), .A3(n50392), .Z(n50397) );
  CLKNAND2HSV1 U53993 ( .A1(n58029), .A2(n57752), .ZN(n50396) );
  CLKNAND2HSV1 U53994 ( .A1(n59935), .A2(n57674), .ZN(n50395) );
  XOR3HSV2 U53995 ( .A1(n50397), .A2(n50396), .A3(n50395), .Z(n50398) );
  XNOR2HSV1 U53996 ( .A1(n50399), .A2(n50398), .ZN(n50403) );
  NAND2HSV2 U53997 ( .A1(n57819), .A2(\pe4/got [18]), .ZN(n50402) );
  BUFHSV2 U53998 ( .I(n58037), .Z(n57960) );
  CLKNAND2HSV1 U53999 ( .A1(n57960), .A2(n57457), .ZN(n50401) );
  XOR3HSV2 U54000 ( .A1(n50403), .A2(n50402), .A3(n50401), .Z(n50406) );
  CLKNAND2HSV0 U54001 ( .A1(n25427), .A2(n50404), .ZN(n50405) );
  XNOR2HSV1 U54002 ( .A1(n50406), .A2(n50405), .ZN(n50408) );
  CLKNAND2HSV0 U54003 ( .A1(n57755), .A2(n33831), .ZN(n50407) );
  XNOR2HSV1 U54004 ( .A1(n50408), .A2(n50407), .ZN(n50409) );
  XNOR2HSV1 U54005 ( .A1(n50410), .A2(n50409), .ZN(n50413) );
  CLKNAND2HSV1 U54006 ( .A1(n58048), .A2(n59601), .ZN(n50412) );
  XOR3HSV2 U54007 ( .A1(n50413), .A2(n50412), .A3(n50411), .Z(n50415) );
  XNOR2HSV1 U54008 ( .A1(n50415), .A2(n50414), .ZN(n50416) );
  XNOR2HSV1 U54009 ( .A1(n50417), .A2(n50416), .ZN(n50420) );
  NOR2HSV2 U54010 ( .A1(n26761), .A2(n33749), .ZN(n50418) );
  XOR3HSV2 U54011 ( .A1(n50420), .A2(n50419), .A3(n50418), .Z(\pe4/poht [5])
         );
  INHSV2 U54012 ( .I(n50421), .ZN(n50652) );
  NAND2HSV0 U54013 ( .A1(n53359), .A2(n59949), .ZN(n50423) );
  NOR2HSV2 U54014 ( .A1(n50652), .A2(n50423), .ZN(n50491) );
  CLKNAND2HSV1 U54015 ( .A1(n53287), .A2(n50643), .ZN(n50487) );
  CLKNHSV0 U54016 ( .I(n25830), .ZN(n51272) );
  CLKNAND2HSV0 U54017 ( .A1(n51272), .A2(n53285), .ZN(n50485) );
  CLKNAND2HSV0 U54018 ( .A1(n59892), .A2(n48167), .ZN(n50481) );
  CLKNAND2HSV1 U54019 ( .A1(n51016), .A2(n50424), .ZN(n50477) );
  NOR2HSV2 U54020 ( .A1(n48166), .A2(n46978), .ZN(n50472) );
  NAND2HSV0 U54021 ( .A1(n59894), .A2(n52576), .ZN(n50468) );
  CLKNAND2HSV1 U54022 ( .A1(n59882), .A2(\pe5/got [4]), .ZN(n50466) );
  NAND2HSV0 U54023 ( .A1(n59525), .A2(\pe5/got [2]), .ZN(n50462) );
  CLKNAND2HSV0 U54024 ( .A1(n44694), .A2(\pe5/got [1]), .ZN(n50460) );
  NAND2HSV0 U54025 ( .A1(\pe5/aot [4]), .A2(n50500), .ZN(n50498) );
  NAND2HSV0 U54026 ( .A1(n59943), .A2(n51370), .ZN(n50425) );
  XOR2HSV0 U54027 ( .A1(n50498), .A2(n50425), .Z(n50441) );
  NAND2HSV0 U54028 ( .A1(\pe5/aot [18]), .A2(n51276), .ZN(n50427) );
  NAND2HSV0 U54029 ( .A1(n59881), .A2(\pe5/bq[2] ), .ZN(n50426) );
  XOR2HSV0 U54030 ( .A1(n50427), .A2(n50426), .Z(n50432) );
  NOR2HSV0 U54031 ( .A1(n47230), .A2(n50428), .ZN(n50430) );
  NAND2HSV0 U54032 ( .A1(\pe5/aot [10]), .A2(n50533), .ZN(n50429) );
  XOR2HSV0 U54033 ( .A1(n50430), .A2(n50429), .Z(n50431) );
  XNOR2HSV1 U54034 ( .A1(n50432), .A2(n50431), .ZN(n50440) );
  NAND2HSV0 U54035 ( .A1(n51363), .A2(\pe5/bq[14] ), .ZN(n50434) );
  NAND2HSV0 U54036 ( .A1(n53296), .A2(\pe5/bq[11] ), .ZN(n50433) );
  XOR2HSV0 U54037 ( .A1(n50434), .A2(n50433), .Z(n50438) );
  NAND2HSV0 U54038 ( .A1(n51310), .A2(n50668), .ZN(n50436) );
  NAND2HSV0 U54039 ( .A1(\pe5/aot [13]), .A2(n50526), .ZN(n50435) );
  XOR2HSV0 U54040 ( .A1(n50436), .A2(n50435), .Z(n50437) );
  XOR2HSV0 U54041 ( .A1(n50438), .A2(n50437), .Z(n50439) );
  XOR3HSV2 U54042 ( .A1(n50441), .A2(n50440), .A3(n50439), .Z(n50458) );
  NAND2HSV0 U54043 ( .A1(n53299), .A2(\pe5/bq[7] ), .ZN(n50443) );
  NAND2HSV0 U54044 ( .A1(n39490), .A2(n50504), .ZN(n50442) );
  XOR2HSV0 U54045 ( .A1(n50443), .A2(n50442), .Z(n50448) );
  NAND2HSV0 U54046 ( .A1(n59895), .A2(n50444), .ZN(n50446) );
  NAND2HSV0 U54047 ( .A1(n39887), .A2(n53216), .ZN(n50445) );
  XOR2HSV0 U54048 ( .A1(n50446), .A2(n50445), .Z(n50447) );
  XOR2HSV0 U54049 ( .A1(n50448), .A2(n50447), .Z(n50456) );
  CLKNAND2HSV1 U54050 ( .A1(n52611), .A2(n50675), .ZN(n50450) );
  NAND2HSV0 U54051 ( .A1(n59866), .A2(n51176), .ZN(n50449) );
  XOR2HSV0 U54052 ( .A1(n50450), .A2(n50449), .Z(n50454) );
  NOR2HSV0 U54053 ( .A1(n59869), .A2(n39796), .ZN(n50452) );
  NAND2HSV0 U54054 ( .A1(\pe5/aot [16]), .A2(n51281), .ZN(n50451) );
  XOR2HSV0 U54055 ( .A1(n50452), .A2(n50451), .Z(n50453) );
  XOR2HSV0 U54056 ( .A1(n50454), .A2(n50453), .Z(n50455) );
  XOR2HSV0 U54057 ( .A1(n50456), .A2(n50455), .Z(n50457) );
  XNOR2HSV1 U54058 ( .A1(n50458), .A2(n50457), .ZN(n50459) );
  XNOR2HSV1 U54059 ( .A1(n50460), .A2(n50459), .ZN(n50461) );
  XNOR2HSV1 U54060 ( .A1(n50462), .A2(n50461), .ZN(n50464) );
  NOR2HSV0 U54061 ( .A1(n50617), .A2(n51231), .ZN(n50463) );
  XNOR2HSV1 U54062 ( .A1(n50464), .A2(n50463), .ZN(n50465) );
  XNOR2HSV1 U54063 ( .A1(n50466), .A2(n50465), .ZN(n50467) );
  XNOR2HSV1 U54064 ( .A1(n50468), .A2(n50467), .ZN(n50470) );
  NAND2HSV0 U54065 ( .A1(n52653), .A2(n51200), .ZN(n50469) );
  XNOR2HSV1 U54066 ( .A1(n50470), .A2(n50469), .ZN(n50471) );
  XNOR2HSV1 U54067 ( .A1(n50472), .A2(n50471), .ZN(n50475) );
  CLKNAND2HSV0 U54068 ( .A1(n59903), .A2(n50698), .ZN(n50474) );
  NOR2HSV1 U54069 ( .A1(n51360), .A2(n46119), .ZN(n50473) );
  XOR3HSV2 U54070 ( .A1(n50475), .A2(n50474), .A3(n50473), .Z(n50476) );
  XNOR2HSV1 U54071 ( .A1(n50477), .A2(n50476), .ZN(n50479) );
  NAND2HSV0 U54072 ( .A1(n53344), .A2(n51305), .ZN(n50478) );
  XOR2HSV0 U54073 ( .A1(n50479), .A2(n50478), .Z(n50480) );
  XNOR2HSV1 U54074 ( .A1(n50481), .A2(n50480), .ZN(n50483) );
  CLKNAND2HSV0 U54075 ( .A1(n51404), .A2(n53286), .ZN(n50482) );
  XNOR2HSV1 U54076 ( .A1(n50483), .A2(n50482), .ZN(n50484) );
  XNOR2HSV1 U54077 ( .A1(n50485), .A2(n50484), .ZN(n50486) );
  CLKNAND2HSV1 U54078 ( .A1(n29779), .A2(n39881), .ZN(n50488) );
  XOR2HSV0 U54079 ( .A1(n50489), .A2(n50488), .Z(n50490) );
  XNOR2HSV1 U54080 ( .A1(n50491), .A2(n50490), .ZN(n50494) );
  AND2HSV2 U54081 ( .A1(n51108), .A2(n50495), .Z(n50492) );
  CLKNAND2HSV1 U54082 ( .A1(n51109), .A2(n50492), .ZN(n50493) );
  XNOR2HSV1 U54083 ( .A1(n50494), .A2(n50493), .ZN(\pe5/poht [14]) );
  NAND2HSV0 U54084 ( .A1(n53359), .A2(n50495), .ZN(n50496) );
  NOR2HSV2 U54085 ( .A1(n51013), .A2(n50496), .ZN(n50579) );
  NAND2HSV2 U54086 ( .A1(n51155), .A2(n52658), .ZN(n50575) );
  CLKNAND2HSV1 U54087 ( .A1(n52564), .A2(n50643), .ZN(n50573) );
  CLKNAND2HSV1 U54088 ( .A1(n53290), .A2(n50497), .ZN(n50569) );
  CLKNAND2HSV1 U54089 ( .A1(n51016), .A2(n53349), .ZN(n50565) );
  NOR2HSV0 U54090 ( .A1(n53293), .A2(n45901), .ZN(n50560) );
  NAND2HSV0 U54091 ( .A1(n59894), .A2(n51200), .ZN(n50556) );
  CLKNAND2HSV1 U54092 ( .A1(n48747), .A2(n52576), .ZN(n50554) );
  CLKNAND2HSV0 U54093 ( .A1(n51018), .A2(n52579), .ZN(n50549) );
  CLKNAND2HSV1 U54094 ( .A1(n51019), .A2(n51362), .ZN(n50545) );
  NOR2HSV0 U54095 ( .A1(n50499), .A2(n50498), .ZN(n50503) );
  AOI22HSV0 U54096 ( .A1(n50501), .A2(n52610), .B1(n50500), .B2(n52623), .ZN(
        n50502) );
  NOR2HSV2 U54097 ( .A1(n50503), .A2(n50502), .ZN(n50506) );
  NAND2HSV0 U54098 ( .A1(n50505), .A2(n50504), .ZN(n51020) );
  XOR2HSV0 U54099 ( .A1(n50506), .A2(n51020), .Z(n50525) );
  NOR2HSV0 U54100 ( .A1(n50507), .A2(n46916), .ZN(n50509) );
  NAND2HSV0 U54101 ( .A1(n59642), .A2(n48170), .ZN(n50508) );
  XOR2HSV0 U54102 ( .A1(n50509), .A2(n50508), .Z(n50515) );
  NAND2HSV2 U54103 ( .A1(n53296), .A2(n51370), .ZN(n51284) );
  NOR2HSV0 U54104 ( .A1(n50510), .A2(n51284), .ZN(n50513) );
  AOI22HSV0 U54105 ( .A1(\pe5/aot [16]), .A2(n53307), .B1(\pe5/bq[12] ), .B2(
        n50511), .ZN(n50512) );
  NOR2HSV2 U54106 ( .A1(n50513), .A2(n50512), .ZN(n50514) );
  XNOR2HSV1 U54107 ( .A1(n50515), .A2(n50514), .ZN(n50524) );
  XOR2HSV0 U54108 ( .A1(n50517), .A2(n50516), .Z(n50522) );
  NOR2HSV0 U54109 ( .A1(n50518), .A2(n48031), .ZN(n50520) );
  NAND2HSV0 U54110 ( .A1(n40190), .A2(n51276), .ZN(n50519) );
  XOR2HSV0 U54111 ( .A1(n50520), .A2(n50519), .Z(n50521) );
  XOR2HSV0 U54112 ( .A1(n50522), .A2(n50521), .Z(n50523) );
  XOR3HSV2 U54113 ( .A1(n50525), .A2(n50524), .A3(n50523), .Z(n50543) );
  NAND2HSV0 U54114 ( .A1(\pe5/aot [14]), .A2(n50526), .ZN(n50528) );
  NAND2HSV0 U54115 ( .A1(\pe5/aot [13]), .A2(\pe5/bq[7] ), .ZN(n50527) );
  XOR2HSV0 U54116 ( .A1(n50528), .A2(n50527), .Z(n50532) );
  NAND2HSV0 U54117 ( .A1(\pe5/aot [7]), .A2(n50668), .ZN(n50530) );
  NAND2HSV0 U54118 ( .A1(n53295), .A2(\pe5/bq[14] ), .ZN(n50529) );
  XOR2HSV0 U54119 ( .A1(n50530), .A2(n50529), .Z(n50531) );
  XOR2HSV0 U54120 ( .A1(n50532), .A2(n50531), .Z(n50541) );
  NAND2HSV0 U54121 ( .A1(n39887), .A2(\pe5/bq[11] ), .ZN(n50535) );
  NAND2HSV0 U54122 ( .A1(n59897), .A2(n50533), .ZN(n50534) );
  XOR2HSV0 U54123 ( .A1(n50535), .A2(n50534), .Z(n50539) );
  NAND2HSV0 U54124 ( .A1(n52600), .A2(n51176), .ZN(n50537) );
  NAND2HSV0 U54125 ( .A1(n51419), .A2(n52618), .ZN(n50536) );
  XOR2HSV0 U54126 ( .A1(n50537), .A2(n50536), .Z(n50538) );
  XOR2HSV0 U54127 ( .A1(n50539), .A2(n50538), .Z(n50540) );
  XOR2HSV0 U54128 ( .A1(n50541), .A2(n50540), .Z(n50542) );
  XNOR2HSV1 U54129 ( .A1(n50543), .A2(n50542), .ZN(n50544) );
  XNOR2HSV1 U54130 ( .A1(n50545), .A2(n50544), .ZN(n50547) );
  NAND2HSV0 U54131 ( .A1(n44694), .A2(n53197), .ZN(n50546) );
  XOR2HSV0 U54132 ( .A1(n50547), .A2(n50546), .Z(n50548) );
  XNOR2HSV1 U54133 ( .A1(n50549), .A2(n50548), .ZN(n50552) );
  NOR2HSV0 U54134 ( .A1(n50617), .A2(n50550), .ZN(n50551) );
  XNOR2HSV1 U54135 ( .A1(n50552), .A2(n50551), .ZN(n50553) );
  XNOR2HSV1 U54136 ( .A1(n50554), .A2(n50553), .ZN(n50555) );
  XNOR2HSV1 U54137 ( .A1(n50556), .A2(n50555), .ZN(n50558) );
  NAND2HSV0 U54138 ( .A1(n52653), .A2(n51017), .ZN(n50557) );
  XNOR2HSV1 U54139 ( .A1(n50558), .A2(n50557), .ZN(n50559) );
  XNOR2HSV1 U54140 ( .A1(n50560), .A2(n50559), .ZN(n50563) );
  CLKNAND2HSV0 U54141 ( .A1(n40019), .A2(n51358), .ZN(n50562) );
  NOR2HSV1 U54142 ( .A1(n50692), .A2(n46961), .ZN(n50561) );
  XOR3HSV2 U54143 ( .A1(n50563), .A2(n50562), .A3(n50561), .Z(n50564) );
  XNOR2HSV1 U54144 ( .A1(n50565), .A2(n50564), .ZN(n50567) );
  NAND2HSV0 U54145 ( .A1(n53344), .A2(\pe5/got [12]), .ZN(n50566) );
  XOR2HSV0 U54146 ( .A1(n50567), .A2(n50566), .Z(n50568) );
  XNOR2HSV1 U54147 ( .A1(n50569), .A2(n50568), .ZN(n50571) );
  CLKNAND2HSV0 U54148 ( .A1(n51404), .A2(n53285), .ZN(n50570) );
  XNOR2HSV1 U54149 ( .A1(n50571), .A2(n50570), .ZN(n50572) );
  XNOR2HSV1 U54150 ( .A1(n50573), .A2(n50572), .ZN(n50574) );
  XNOR2HSV1 U54151 ( .A1(n50575), .A2(n50574), .ZN(n50577) );
  NAND2HSV2 U54152 ( .A1(n29777), .A2(n59949), .ZN(n50576) );
  XNOR2HSV1 U54153 ( .A1(n50577), .A2(n50576), .ZN(n50578) );
  XOR2HSV2 U54154 ( .A1(n50579), .A2(n50578), .Z(n50582) );
  AND2HSV2 U54155 ( .A1(n53361), .A2(n51103), .Z(n50580) );
  CLKNAND2HSV1 U54156 ( .A1(n51109), .A2(n50580), .ZN(n50581) );
  XNOR2HSV1 U54157 ( .A1(n50582), .A2(n50581), .ZN(\pe5/poht [13]) );
  NAND2HSV0 U54158 ( .A1(n53359), .A2(n39881), .ZN(n50583) );
  NOR2HSV2 U54159 ( .A1(n50652), .A2(n50583), .ZN(n50647) );
  CLKNAND2HSV1 U54160 ( .A1(n53287), .A2(n53285), .ZN(n50642) );
  CLKNAND2HSV0 U54161 ( .A1(n51272), .A2(n53286), .ZN(n50640) );
  CLKNAND2HSV0 U54162 ( .A1(n52670), .A2(n51305), .ZN(n50636) );
  CLKNAND2HSV1 U54163 ( .A1(n51016), .A2(n51358), .ZN(n50632) );
  NOR2HSV0 U54164 ( .A1(n53293), .A2(n45903), .ZN(n50627) );
  NAND2HSV0 U54165 ( .A1(n59894), .A2(n51418), .ZN(n50623) );
  CLKNAND2HSV1 U54166 ( .A1(n52570), .A2(n52579), .ZN(n50621) );
  NAND2HSV0 U54167 ( .A1(n59525), .A2(\pe5/got [1]), .ZN(n50616) );
  XOR2HSV0 U54168 ( .A1(n50585), .A2(n50584), .Z(n50598) );
  NAND2HSV0 U54169 ( .A1(\pe5/aot [13]), .A2(n51373), .ZN(n50587) );
  NAND2HSV0 U54170 ( .A1(n50653), .A2(n51281), .ZN(n50586) );
  XOR2HSV0 U54171 ( .A1(n50587), .A2(n50586), .Z(n50589) );
  NAND2HSV0 U54172 ( .A1(n50588), .A2(n39471), .ZN(n51039) );
  XNOR2HSV1 U54173 ( .A1(n50589), .A2(n51039), .ZN(n50597) );
  NAND2HSV0 U54174 ( .A1(\pe5/aot [4]), .A2(\pe5/bq[14] ), .ZN(n50591) );
  NAND2HSV0 U54175 ( .A1(n39887), .A2(\pe5/bq[9] ), .ZN(n50590) );
  XOR2HSV0 U54176 ( .A1(n50591), .A2(n50590), .Z(n50595) );
  NAND2HSV0 U54177 ( .A1(n59881), .A2(n51276), .ZN(n50593) );
  CLKNAND2HSV0 U54178 ( .A1(\pe5/aot [6]), .A2(n31045), .ZN(n50592) );
  XOR2HSV0 U54179 ( .A1(n50593), .A2(n50592), .Z(n50594) );
  XOR2HSV0 U54180 ( .A1(n50595), .A2(n50594), .Z(n50596) );
  XOR3HSV2 U54181 ( .A1(n50598), .A2(n50597), .A3(n50596), .Z(n50614) );
  CLKNAND2HSV1 U54182 ( .A1(n51313), .A2(n50675), .ZN(n50600) );
  CLKNAND2HSV1 U54183 ( .A1(n51247), .A2(n39592), .ZN(n50599) );
  XOR2HSV0 U54184 ( .A1(n50600), .A2(n50599), .Z(n50604) );
  NAND2HSV0 U54185 ( .A1(n59896), .A2(n50526), .ZN(n50602) );
  NAND2HSV0 U54186 ( .A1(n39490), .A2(n51370), .ZN(n50601) );
  XOR2HSV0 U54187 ( .A1(n50602), .A2(n50601), .Z(n50603) );
  XOR2HSV0 U54188 ( .A1(n50604), .A2(n50603), .Z(n50612) );
  NAND2HSV0 U54189 ( .A1(n59880), .A2(n53216), .ZN(n50606) );
  NAND2HSV0 U54190 ( .A1(n59897), .A2(\pe5/bq[7] ), .ZN(n50605) );
  XOR2HSV0 U54191 ( .A1(n50606), .A2(n50605), .Z(n50610) );
  NOR2HSV0 U54192 ( .A1(n45904), .A2(n45821), .ZN(n50608) );
  NAND2HSV0 U54193 ( .A1(\pe5/aot [16]), .A2(\pe5/bq[2] ), .ZN(n50607) );
  XOR2HSV0 U54194 ( .A1(n50608), .A2(n50607), .Z(n50609) );
  XOR2HSV0 U54195 ( .A1(n50610), .A2(n50609), .Z(n50611) );
  XOR2HSV0 U54196 ( .A1(n50612), .A2(n50611), .Z(n50613) );
  XNOR2HSV1 U54197 ( .A1(n50614), .A2(n50613), .ZN(n50615) );
  XNOR2HSV1 U54198 ( .A1(n50616), .A2(n50615), .ZN(n50619) );
  NOR2HSV0 U54199 ( .A1(n50617), .A2(n51306), .ZN(n50618) );
  XNOR2HSV1 U54200 ( .A1(n50619), .A2(n50618), .ZN(n50620) );
  XNOR2HSV1 U54201 ( .A1(n50621), .A2(n50620), .ZN(n50622) );
  XNOR2HSV1 U54202 ( .A1(n50623), .A2(n50622), .ZN(n50625) );
  NAND2HSV0 U54203 ( .A1(n52653), .A2(n52576), .ZN(n50624) );
  XNOR2HSV1 U54204 ( .A1(n50625), .A2(n50624), .ZN(n50626) );
  XNOR2HSV1 U54205 ( .A1(n50627), .A2(n50626), .ZN(n50630) );
  CLKNAND2HSV0 U54206 ( .A1(n59903), .A2(n51017), .ZN(n50629) );
  NOR2HSV1 U54207 ( .A1(n51218), .A2(n45901), .ZN(n50628) );
  XOR3HSV2 U54208 ( .A1(n50630), .A2(n50629), .A3(n50628), .Z(n50631) );
  XNOR2HSV1 U54209 ( .A1(n50632), .A2(n50631), .ZN(n50634) );
  NAND2HSV0 U54210 ( .A1(n51092), .A2(n53289), .ZN(n50633) );
  XOR2HSV0 U54211 ( .A1(n50634), .A2(n50633), .Z(n50635) );
  XNOR2HSV1 U54212 ( .A1(n50636), .A2(n50635), .ZN(n50638) );
  CLKNAND2HSV1 U54213 ( .A1(n51335), .A2(n48167), .ZN(n50637) );
  XNOR2HSV1 U54214 ( .A1(n50638), .A2(n50637), .ZN(n50639) );
  CLKNAND2HSV1 U54215 ( .A1(n29778), .A2(n50643), .ZN(n50644) );
  XNOR2HSV1 U54216 ( .A1(n50645), .A2(n50644), .ZN(n50646) );
  CLKXOR2HSV4 U54217 ( .A1(n50647), .A2(n50646), .Z(n50650) );
  AND2HSV2 U54218 ( .A1(n53361), .A2(n59949), .Z(n50648) );
  CLKNAND2HSV1 U54219 ( .A1(n53363), .A2(n50648), .ZN(n50649) );
  XNOR2HSV1 U54220 ( .A1(n50650), .A2(n50649), .ZN(\pe5/poht [15]) );
  NAND2HSV0 U54221 ( .A1(n53359), .A2(n40186), .ZN(n50651) );
  NOR2HSV2 U54222 ( .A1(n50652), .A2(n50651), .ZN(n50712) );
  CLKNAND2HSV1 U54223 ( .A1(n53287), .A2(n48167), .ZN(n50708) );
  CLKNAND2HSV0 U54224 ( .A1(n51272), .A2(n51305), .ZN(n50706) );
  CLKNAND2HSV1 U54225 ( .A1(n52565), .A2(n51358), .ZN(n50702) );
  CLKNAND2HSV1 U54226 ( .A1(n51016), .A2(n51017), .ZN(n50697) );
  NOR2HSV2 U54227 ( .A1(n53293), .A2(n50550), .ZN(n50691) );
  NAND2HSV0 U54228 ( .A1(n59894), .A2(\pe5/got [2]), .ZN(n50687) );
  NAND2HSV0 U54229 ( .A1(n59882), .A2(n51362), .ZN(n50685) );
  NAND2HSV0 U54230 ( .A1(n50653), .A2(n51276), .ZN(n50655) );
  NAND2HSV0 U54231 ( .A1(\pe5/aot [13]), .A2(n51281), .ZN(n50654) );
  XOR2HSV0 U54232 ( .A1(n50655), .A2(n50654), .Z(n50659) );
  NAND2HSV0 U54233 ( .A1(n51313), .A2(\pe5/bq[6] ), .ZN(n50657) );
  NAND2HSV0 U54234 ( .A1(n59896), .A2(n51370), .ZN(n50656) );
  XOR2HSV0 U54235 ( .A1(n50657), .A2(n50656), .Z(n50658) );
  XOR2HSV0 U54236 ( .A1(n50659), .A2(n50658), .Z(n50667) );
  NAND2HSV0 U54237 ( .A1(\pe5/aot [6]), .A2(n53216), .ZN(n50661) );
  NAND2HSV0 U54238 ( .A1(n51419), .A2(\pe5/bq[14] ), .ZN(n50660) );
  XOR2HSV0 U54239 ( .A1(n50661), .A2(n50660), .Z(n50665) );
  NAND2HSV0 U54240 ( .A1(n59897), .A2(n51373), .ZN(n50663) );
  CLKNAND2HSV0 U54241 ( .A1(n51363), .A2(\pe5/bq[11] ), .ZN(n50662) );
  XOR2HSV0 U54242 ( .A1(n50663), .A2(n50662), .Z(n50664) );
  XOR2HSV0 U54243 ( .A1(n50665), .A2(n50664), .Z(n50666) );
  XOR2HSV0 U54244 ( .A1(n50667), .A2(n50666), .Z(n50683) );
  NAND2HSV0 U54245 ( .A1(\pe5/aot [3]), .A2(n50668), .ZN(n50670) );
  NAND2HSV0 U54246 ( .A1(n51339), .A2(n39914), .ZN(n50669) );
  XOR2HSV0 U54247 ( .A1(n50670), .A2(n50669), .Z(n50674) );
  NOR2HSV1 U54248 ( .A1(n47230), .A2(n47162), .ZN(n50672) );
  CLKNAND2HSV0 U54249 ( .A1(n39490), .A2(\pe5/bq[2] ), .ZN(n50671) );
  XOR2HSV0 U54250 ( .A1(n50672), .A2(n50671), .Z(n50673) );
  XOR2HSV0 U54251 ( .A1(n50674), .A2(n50673), .Z(n50681) );
  CLKNAND2HSV1 U54252 ( .A1(n53296), .A2(n50675), .ZN(n50677) );
  NAND2HSV0 U54253 ( .A1(\pe5/aot [4]), .A2(n31045), .ZN(n50676) );
  XOR2HSV0 U54254 ( .A1(n50677), .A2(n50676), .Z(n50679) );
  XNOR2HSV1 U54255 ( .A1(n50679), .A2(n50678), .ZN(n50680) );
  XNOR2HSV1 U54256 ( .A1(n50681), .A2(n50680), .ZN(n50682) );
  XNOR2HSV1 U54257 ( .A1(n50683), .A2(n50682), .ZN(n50684) );
  XNOR2HSV1 U54258 ( .A1(n50685), .A2(n50684), .ZN(n50686) );
  XNOR2HSV1 U54259 ( .A1(n50687), .A2(n50686), .ZN(n50689) );
  NAND2HSV0 U54260 ( .A1(n52653), .A2(n51331), .ZN(n50688) );
  XNOR2HSV1 U54261 ( .A1(n50689), .A2(n50688), .ZN(n50690) );
  XNOR2HSV1 U54262 ( .A1(n50691), .A2(n50690), .ZN(n50695) );
  CLKNAND2HSV0 U54263 ( .A1(n59903), .A2(n51334), .ZN(n50694) );
  NOR2HSV1 U54264 ( .A1(n50692), .A2(n45903), .ZN(n50693) );
  XOR3HSV2 U54265 ( .A1(n50695), .A2(n50694), .A3(n50693), .Z(n50696) );
  XNOR2HSV1 U54266 ( .A1(n50697), .A2(n50696), .ZN(n50700) );
  CLKNAND2HSV0 U54267 ( .A1(n51092), .A2(n50698), .ZN(n50699) );
  XOR2HSV0 U54268 ( .A1(n50700), .A2(n50699), .Z(n50701) );
  NAND2HSV0 U54269 ( .A1(n51227), .A2(n52571), .ZN(n50703) );
  XNOR2HSV1 U54270 ( .A1(n50706), .A2(n50705), .ZN(n50707) );
  XNOR2HSV1 U54271 ( .A1(n50708), .A2(n50707), .ZN(n50710) );
  CLKNAND2HSV1 U54272 ( .A1(n29778), .A2(n59367), .ZN(n50709) );
  XNOR2HSV1 U54273 ( .A1(n50710), .A2(n50709), .ZN(n50711) );
  CLKXOR2HSV4 U54274 ( .A1(n50712), .A2(n50711), .Z(n50715) );
  CLKAND2HSV2 U54275 ( .A1(n53361), .A2(n51015), .Z(n50713) );
  CLKNAND2HSV1 U54276 ( .A1(n51109), .A2(n50713), .ZN(n50714) );
  XNOR2HSV1 U54277 ( .A1(n50715), .A2(n50714), .ZN(\pe5/poht [17]) );
  CLKNAND2HSV1 U54278 ( .A1(n56339), .A2(n56771), .ZN(n50749) );
  INHSV2 U54279 ( .I(n56682), .ZN(n56909) );
  INHSV1 U54280 ( .I(n56859), .ZN(n56623) );
  CLKNAND2HSV1 U54281 ( .A1(n56173), .A2(n56623), .ZN(n50745) );
  CLKNHSV0 U54282 ( .I(n50717), .ZN(n56341) );
  CLKNAND2HSV1 U54283 ( .A1(n56341), .A2(n56684), .ZN(n50743) );
  CLKNAND2HSV0 U54284 ( .A1(n55822), .A2(n56735), .ZN(n50741) );
  CLKNHSV0 U54285 ( .I(n56936), .ZN(n56782) );
  NAND2HSV0 U54286 ( .A1(n56175), .A2(n56782), .ZN(n50739) );
  CLKNAND2HSV0 U54287 ( .A1(n48486), .A2(\pe3/got [1]), .ZN(n50737) );
  NAND2HSV0 U54288 ( .A1(n56740), .A2(n56824), .ZN(n56574) );
  NAND2HSV0 U54289 ( .A1(n56221), .A2(\pe3/bq[4] ), .ZN(n50719) );
  XOR2HSV0 U54290 ( .A1(n56574), .A2(n50719), .Z(n50735) );
  CLKNAND2HSV0 U54291 ( .A1(n59961), .A2(n53232), .ZN(n50721) );
  NAND2HSV0 U54292 ( .A1(n59511), .A2(n56627), .ZN(n50720) );
  XOR2HSV0 U54293 ( .A1(n50721), .A2(n50720), .Z(n50726) );
  NOR2HSV1 U54294 ( .A1(n45662), .A2(n49258), .ZN(n50724) );
  NAND2HSV0 U54295 ( .A1(\pe3/aot [8]), .A2(n56529), .ZN(n50723) );
  XOR2HSV0 U54296 ( .A1(n50724), .A2(n50723), .Z(n50725) );
  XNOR2HSV1 U54297 ( .A1(n50726), .A2(n50725), .ZN(n50734) );
  CLKNAND2HSV0 U54298 ( .A1(n56788), .A2(n56832), .ZN(n50728) );
  NAND2HSV0 U54299 ( .A1(n53250), .A2(n56827), .ZN(n50727) );
  XOR2HSV0 U54300 ( .A1(n50728), .A2(n50727), .Z(n50732) );
  NAND2HSV0 U54301 ( .A1(n56423), .A2(n56505), .ZN(n50730) );
  BUFHSV2 U54302 ( .I(\pe3/aot [6]), .Z(n56911) );
  CLKNAND2HSV0 U54303 ( .A1(n56911), .A2(n56867), .ZN(n50729) );
  XOR2HSV0 U54304 ( .A1(n50730), .A2(n50729), .Z(n50731) );
  XOR2HSV0 U54305 ( .A1(n50732), .A2(n50731), .Z(n50733) );
  XOR3HSV2 U54306 ( .A1(n50735), .A2(n50734), .A3(n50733), .Z(n50736) );
  XNOR2HSV1 U54307 ( .A1(n50737), .A2(n50736), .ZN(n50738) );
  XNOR2HSV1 U54308 ( .A1(n50739), .A2(n50738), .ZN(n50740) );
  XNOR2HSV1 U54309 ( .A1(n50741), .A2(n50740), .ZN(n50742) );
  XNOR2HSV1 U54310 ( .A1(n50743), .A2(n50742), .ZN(n50744) );
  XNOR2HSV1 U54311 ( .A1(n50745), .A2(n50744), .ZN(n50746) );
  XOR2HSV0 U54312 ( .A1(n50747), .A2(n50746), .Z(n50748) );
  XOR2HSV0 U54313 ( .A1(n50749), .A2(n50748), .Z(n50751) );
  CLKNAND2HSV1 U54314 ( .A1(n53279), .A2(n56855), .ZN(n50750) );
  INHSV4 U54315 ( .I(n50752), .ZN(n56965) );
  NAND2HSV2 U54316 ( .A1(n56058), .A2(n56558), .ZN(n50754) );
  CLKNAND2HSV1 U54317 ( .A1(n56976), .A2(n56620), .ZN(n50753) );
  XOR3HSV2 U54318 ( .A1(n50755), .A2(n50754), .A3(n50753), .Z(\pe3/poht [22])
         );
  CLKNAND2HSV1 U54319 ( .A1(n56339), .A2(n56495), .ZN(n50798) );
  CLKNAND2HSV0 U54320 ( .A1(n48481), .A2(n56855), .ZN(n50794) );
  CLKNAND2HSV1 U54321 ( .A1(n56341), .A2(n56266), .ZN(n50792) );
  CLKNAND2HSV0 U54322 ( .A1(n55822), .A2(n56779), .ZN(n50790) );
  NAND2HSV0 U54323 ( .A1(n59930), .A2(n56623), .ZN(n50788) );
  CLKNAND2HSV0 U54324 ( .A1(n43869), .A2(n56684), .ZN(n50786) );
  NAND2HSV0 U54325 ( .A1(n46312), .A2(n56735), .ZN(n50784) );
  NAND2HSV0 U54326 ( .A1(n59500), .A2(n56782), .ZN(n50782) );
  NAND2HSV0 U54327 ( .A1(n56662), .A2(\pe3/got [1]), .ZN(n50780) );
  NAND2HSV0 U54328 ( .A1(n56740), .A2(\pe3/bq[4] ), .ZN(n50759) );
  NAND2HSV0 U54329 ( .A1(n56373), .A2(n56937), .ZN(n50758) );
  XOR2HSV0 U54330 ( .A1(n50759), .A2(n50758), .Z(n50763) );
  NAND2HSV0 U54331 ( .A1(n56439), .A2(n53232), .ZN(n50761) );
  NAND2HSV0 U54332 ( .A1(n59961), .A2(n56507), .ZN(n50760) );
  XOR2HSV0 U54333 ( .A1(n50761), .A2(n50760), .Z(n50762) );
  XOR2HSV0 U54334 ( .A1(n50763), .A2(n50762), .Z(n50771) );
  NAND2HSV0 U54335 ( .A1(n53250), .A2(\pe3/bq[11] ), .ZN(n50765) );
  NAND2HSV0 U54336 ( .A1(n56788), .A2(n56627), .ZN(n50764) );
  XOR2HSV0 U54337 ( .A1(n50765), .A2(n50764), .Z(n50769) );
  CLKNAND2HSV0 U54338 ( .A1(n43280), .A2(\pe3/bq[1] ), .ZN(n50767) );
  NAND2HSV0 U54339 ( .A1(\pe3/aot [11]), .A2(n56529), .ZN(n50766) );
  XOR2HSV0 U54340 ( .A1(n50767), .A2(n50766), .Z(n50768) );
  XOR2HSV0 U54341 ( .A1(n50769), .A2(n50768), .Z(n50770) );
  XOR2HSV0 U54342 ( .A1(n50771), .A2(n50770), .Z(n50778) );
  NOR2HSV0 U54343 ( .A1(n53229), .A2(n48495), .ZN(n56577) );
  CLKNAND2HSV1 U54344 ( .A1(n56795), .A2(n55970), .ZN(n56654) );
  CLKNAND2HSV0 U54345 ( .A1(\pe3/aot [8]), .A2(n56835), .ZN(n50772) );
  XNOR2HSV1 U54346 ( .A1(n56654), .A2(n50772), .ZN(n50776) );
  NAND2HSV0 U54347 ( .A1(n59511), .A2(n56644), .ZN(n50774) );
  NAND2HSV0 U54348 ( .A1(n56221), .A2(n45639), .ZN(n50773) );
  XOR2HSV0 U54349 ( .A1(n50774), .A2(n50773), .Z(n50775) );
  XOR3HSV2 U54350 ( .A1(n56577), .A2(n50776), .A3(n50775), .Z(n50777) );
  XNOR2HSV1 U54351 ( .A1(n50778), .A2(n50777), .ZN(n50779) );
  XNOR2HSV1 U54352 ( .A1(n50780), .A2(n50779), .ZN(n50781) );
  XNOR2HSV1 U54353 ( .A1(n50782), .A2(n50781), .ZN(n50783) );
  XNOR2HSV1 U54354 ( .A1(n50784), .A2(n50783), .ZN(n50785) );
  XNOR2HSV1 U54355 ( .A1(n50786), .A2(n50785), .ZN(n50787) );
  XNOR2HSV1 U54356 ( .A1(n50788), .A2(n50787), .ZN(n50789) );
  XNOR2HSV1 U54357 ( .A1(n50790), .A2(n50789), .ZN(n50791) );
  XNOR2HSV1 U54358 ( .A1(n50792), .A2(n50791), .ZN(n50793) );
  XNOR2HSV1 U54359 ( .A1(n50794), .A2(n50793), .ZN(n50795) );
  XOR2HSV0 U54360 ( .A1(n50796), .A2(n50795), .Z(n50797) );
  XOR2HSV0 U54361 ( .A1(n50798), .A2(n50797), .Z(n50801) );
  CLKNAND2HSV0 U54362 ( .A1(n56935), .A2(n56342), .ZN(n50800) );
  NAND2HSV2 U54363 ( .A1(n56948), .A2(n43829), .ZN(n50804) );
  CLKNAND2HSV1 U54364 ( .A1(n56490), .A2(n56176), .ZN(n50803) );
  CLKNAND2HSV2 U54365 ( .A1(n59021), .A2(n59173), .ZN(n50905) );
  CLKNAND2HSV1 U54366 ( .A1(n32970), .A2(n58575), .ZN(n50903) );
  CLKNAND2HSV1 U54367 ( .A1(n59514), .A2(n59027), .ZN(n50901) );
  CLKNAND2HSV1 U54368 ( .A1(n59172), .A2(n49825), .ZN(n50899) );
  CLKNAND2HSV0 U54369 ( .A1(n58934), .A2(n59029), .ZN(n50897) );
  CLKNAND2HSV1 U54370 ( .A1(n58717), .A2(\pe6/got [19]), .ZN(n50894) );
  CLKNAND2HSV1 U54371 ( .A1(n58935), .A2(n32971), .ZN(n50890) );
  NAND2HSV0 U54372 ( .A1(n58718), .A2(n58937), .ZN(n50888) );
  NAND2HSV0 U54373 ( .A1(n59177), .A2(n58810), .ZN(n50884) );
  NAND2HSV0 U54374 ( .A1(n59916), .A2(n58811), .ZN(n50882) );
  NAND2HSV0 U54375 ( .A1(n58938), .A2(n33039), .ZN(n50880) );
  NOR2HSV0 U54376 ( .A1(n50805), .A2(n53110), .ZN(n50878) );
  NAND2HSV0 U54377 ( .A1(n58722), .A2(n59037), .ZN(n50874) );
  CLKNAND2HSV1 U54378 ( .A1(n59033), .A2(n58526), .ZN(n50872) );
  CLKNAND2HSV1 U54379 ( .A1(n44392), .A2(n58814), .ZN(n50870) );
  CLKNAND2HSV1 U54380 ( .A1(n49743), .A2(n58513), .ZN(n50868) );
  CLKNAND2HSV0 U54381 ( .A1(n58815), .A2(n59292), .ZN(n50866) );
  NAND2HSV0 U54382 ( .A1(n58939), .A2(n58479), .ZN(n50864) );
  NAND2HSV0 U54383 ( .A1(n36107), .A2(n58816), .ZN(n50860) );
  NAND2HSV0 U54384 ( .A1(n59183), .A2(n58817), .ZN(n50858) );
  NAND2HSV0 U54385 ( .A1(n59246), .A2(\pe6/aot [19]), .ZN(n50807) );
  NAND2HSV0 U54386 ( .A1(n58833), .A2(\pe6/aot [11]), .ZN(n50806) );
  XOR2HSV0 U54387 ( .A1(n50807), .A2(n50806), .Z(n50811) );
  NAND2HSV0 U54388 ( .A1(n58976), .A2(n58842), .ZN(n50809) );
  NAND2HSV0 U54389 ( .A1(n59089), .A2(n58943), .ZN(n50808) );
  XOR2HSV0 U54390 ( .A1(n50809), .A2(n50808), .Z(n50810) );
  XOR2HSV0 U54391 ( .A1(n50811), .A2(n50810), .Z(n50819) );
  NAND2HSV0 U54392 ( .A1(\pe6/bq[1] ), .A2(n32876), .ZN(n50813) );
  NAND2HSV0 U54393 ( .A1(\pe6/bq[2] ), .A2(n58824), .ZN(n50812) );
  XOR2HSV0 U54394 ( .A1(n50813), .A2(n50812), .Z(n50817) );
  NAND2HSV0 U54395 ( .A1(n44702), .A2(n58459), .ZN(n50815) );
  NAND2HSV0 U54396 ( .A1(n59050), .A2(n58734), .ZN(n50814) );
  XOR2HSV0 U54397 ( .A1(n50815), .A2(n50814), .Z(n50816) );
  XOR2HSV0 U54398 ( .A1(n50817), .A2(n50816), .Z(n50818) );
  XOR2HSV0 U54399 ( .A1(n50819), .A2(n50818), .Z(n50835) );
  CLKNAND2HSV0 U54400 ( .A1(n59098), .A2(\pe6/aot [7]), .ZN(n50821) );
  NAND2HSV0 U54401 ( .A1(\pe6/bq[17] ), .A2(\pe6/aot [10]), .ZN(n50820) );
  XOR2HSV0 U54402 ( .A1(n50821), .A2(n50820), .Z(n50826) );
  NOR2HSV0 U54403 ( .A1(n50822), .A2(n58359), .ZN(n50824) );
  NAND2HSV0 U54404 ( .A1(\pe6/bq[21] ), .A2(n53134), .ZN(n50823) );
  XOR2HSV0 U54405 ( .A1(n50824), .A2(n50823), .Z(n50825) );
  XNOR2HSV1 U54406 ( .A1(n50826), .A2(n50825), .ZN(n50833) );
  NOR2HSV0 U54407 ( .A1(n49680), .A2(n35864), .ZN(n59111) );
  AOI22HSV0 U54408 ( .A1(n58962), .A2(\pe6/aot [17]), .B1(\pe6/aot [21]), .B2(
        n58975), .ZN(n50827) );
  AOI21HSV0 U54409 ( .A1(n58978), .A2(n59111), .B(n50827), .ZN(n50831) );
  CLKNAND2HSV0 U54410 ( .A1(\pe6/bq[11] ), .A2(n58449), .ZN(n53128) );
  XOR2HSV0 U54411 ( .A1(n50831), .A2(n50830), .Z(n50832) );
  XNOR2HSV1 U54412 ( .A1(n50833), .A2(n50832), .ZN(n50834) );
  XNOR2HSV1 U54413 ( .A1(n50835), .A2(n50834), .ZN(n50856) );
  NAND2HSV0 U54414 ( .A1(n33023), .A2(n59099), .ZN(n59195) );
  XOR2HSV0 U54415 ( .A1(n50836), .A2(n59195), .Z(n50854) );
  NOR2HSV0 U54416 ( .A1(n46642), .A2(n50837), .ZN(n58855) );
  AOI22HSV0 U54417 ( .A1(n59062), .A2(\pe6/aot [23]), .B1(n58749), .B2(n58408), 
        .ZN(n50838) );
  AOI21HSV1 U54418 ( .A1(n50839), .A2(n58855), .B(n50838), .ZN(n50844) );
  NAND2HSV0 U54419 ( .A1(n59217), .A2(n58464), .ZN(n59108) );
  NOR2HSV0 U54420 ( .A1(n50840), .A2(n59108), .ZN(n50842) );
  AOI22HSV0 U54421 ( .A1(n48035), .A2(\pe6/aot [1]), .B1(n59206), .B2(
        \pe6/aot [2]), .ZN(n50841) );
  NOR2HSV1 U54422 ( .A1(n50842), .A2(n50841), .ZN(n50843) );
  XOR2HSV0 U54423 ( .A1(n50844), .A2(n50843), .Z(n50853) );
  NAND2HSV0 U54424 ( .A1(n58668), .A2(\pe6/aot [13]), .ZN(n50845) );
  XOR2HSV0 U54425 ( .A1(n50846), .A2(n50845), .Z(n50851) );
  NOR2HSV0 U54426 ( .A1(n50847), .A2(n32245), .ZN(n50849) );
  NAND2HSV0 U54427 ( .A1(\pe6/bq[5] ), .A2(n33004), .ZN(n50848) );
  XOR2HSV0 U54428 ( .A1(n50849), .A2(n50848), .Z(n50850) );
  XOR2HSV0 U54429 ( .A1(n50851), .A2(n50850), .Z(n50852) );
  XOR3HSV2 U54430 ( .A1(n50854), .A2(n50853), .A3(n50852), .Z(n50855) );
  XNOR2HSV1 U54431 ( .A1(n50856), .A2(n50855), .ZN(n50857) );
  XNOR2HSV1 U54432 ( .A1(n50858), .A2(n50857), .ZN(n50859) );
  XNOR2HSV1 U54433 ( .A1(n50860), .A2(n50859), .ZN(n50862) );
  NAND2HSV0 U54434 ( .A1(n58886), .A2(n58527), .ZN(n50861) );
  XNOR2HSV1 U54435 ( .A1(n50862), .A2(n50861), .ZN(n50863) );
  XNOR2HSV1 U54436 ( .A1(n50864), .A2(n50863), .ZN(n50865) );
  XNOR2HSV1 U54437 ( .A1(n50866), .A2(n50865), .ZN(n50867) );
  XNOR2HSV1 U54438 ( .A1(n50868), .A2(n50867), .ZN(n50869) );
  XNOR2HSV1 U54439 ( .A1(n50870), .A2(n50869), .ZN(n50871) );
  XNOR2HSV1 U54440 ( .A1(n50872), .A2(n50871), .ZN(n50873) );
  XNOR2HSV1 U54441 ( .A1(n50874), .A2(n50873), .ZN(n50876) );
  CLKNAND2HSV0 U54442 ( .A1(n59317), .A2(n58812), .ZN(n50875) );
  XNOR2HSV1 U54443 ( .A1(n50876), .A2(n50875), .ZN(n50877) );
  XNOR2HSV1 U54444 ( .A1(n50878), .A2(n50877), .ZN(n50879) );
  XNOR2HSV1 U54445 ( .A1(n50880), .A2(n50879), .ZN(n50881) );
  XNOR2HSV1 U54446 ( .A1(n50882), .A2(n50881), .ZN(n50883) );
  XNOR2HSV1 U54447 ( .A1(n50884), .A2(n50883), .ZN(n50886) );
  CLKNAND2HSV1 U54448 ( .A1(n58601), .A2(\pe6/got [15]), .ZN(n50885) );
  XNOR2HSV1 U54449 ( .A1(n50886), .A2(n50885), .ZN(n50887) );
  XNOR2HSV1 U54450 ( .A1(n50888), .A2(n50887), .ZN(n50889) );
  XNOR2HSV1 U54451 ( .A1(n50890), .A2(n50889), .ZN(n50892) );
  NAND2HSV0 U54452 ( .A1(n58805), .A2(n58715), .ZN(n50891) );
  XOR2HSV0 U54453 ( .A1(n50892), .A2(n50891), .Z(n50893) );
  XNOR2HSV1 U54454 ( .A1(n50894), .A2(n50893), .ZN(n50896) );
  NAND2HSV0 U54455 ( .A1(n59528), .A2(n59328), .ZN(n50895) );
  XOR3HSV2 U54456 ( .A1(n50897), .A2(n50896), .A3(n50895), .Z(n50898) );
  XNOR2HSV1 U54457 ( .A1(n50899), .A2(n50898), .ZN(n50900) );
  XNOR2HSV1 U54458 ( .A1(n50901), .A2(n50900), .ZN(n50902) );
  XNOR2HSV1 U54459 ( .A1(n50903), .A2(n50902), .ZN(n50904) );
  XNOR2HSV4 U54460 ( .A1(n50905), .A2(n50904), .ZN(n50906) );
  XNOR2HSV4 U54461 ( .A1(n50907), .A2(n50906), .ZN(\pe6/poht [6]) );
  INHSV2 U54462 ( .I(n50908), .ZN(n51686) );
  INHSV2 U54463 ( .I(n53032), .ZN(n52900) );
  NAND2HSV2 U54464 ( .A1(n51798), .A2(n51688), .ZN(n50925) );
  NAND2HSV2 U54465 ( .A1(n59499), .A2(n52484), .ZN(n50912) );
  NAND2HSV0 U54466 ( .A1(n59783), .A2(n51832), .ZN(n50911) );
  XOR2HSV0 U54467 ( .A1(n50912), .A2(n50911), .Z(n50916) );
  NOR2HSV0 U54468 ( .A1(n51538), .A2(n51842), .ZN(n50914) );
  CLKNAND2HSV0 U54469 ( .A1(n52456), .A2(n51919), .ZN(n50913) );
  XOR2HSV0 U54470 ( .A1(n50914), .A2(n50913), .Z(n50915) );
  XNOR2HSV1 U54471 ( .A1(n50916), .A2(n50915), .ZN(n50923) );
  NAND2HSV2 U54472 ( .A1(n59978), .A2(\pe2/bq[6] ), .ZN(n51126) );
  NOR2HSV0 U54473 ( .A1(n51126), .A2(n50917), .ZN(n50919) );
  AOI22HSV0 U54474 ( .A1(n59978), .A2(n51803), .B1(n52866), .B2(\pe2/aot [2]), 
        .ZN(n50918) );
  NOR2HSV2 U54475 ( .A1(n50919), .A2(n50918), .ZN(n50921) );
  NAND2HSV2 U54476 ( .A1(n59633), .A2(n52851), .ZN(n52871) );
  XOR2HSV0 U54477 ( .A1(n50921), .A2(n52871), .Z(n50922) );
  XNOR2HSV1 U54478 ( .A1(n50923), .A2(n50922), .ZN(n50924) );
  CLKNAND2HSV1 U54479 ( .A1(n59929), .A2(n51932), .ZN(n50927) );
  NAND2HSV0 U54480 ( .A1(n59790), .A2(n47571), .ZN(n51009) );
  CLKNAND2HSV1 U54481 ( .A1(n44832), .A2(n51726), .ZN(n51007) );
  NOR2HSV0 U54482 ( .A1(n52171), .A2(n47498), .ZN(n51005) );
  NAND2HSV0 U54483 ( .A1(\pe2/got [10]), .A2(n52814), .ZN(n50997) );
  CLKNAND2HSV0 U54484 ( .A1(n52926), .A2(\pe2/got [8]), .ZN(n50995) );
  CLKNAND2HSV0 U54485 ( .A1(n59634), .A2(n52933), .ZN(n50992) );
  CLKNAND2HSV0 U54486 ( .A1(n51609), .A2(n59777), .ZN(n50990) );
  NAND2HSV0 U54487 ( .A1(\pe2/got [4]), .A2(n52929), .ZN(n50988) );
  INHSV2 U54488 ( .I(n53032), .ZN(n52239) );
  NAND2HSV0 U54489 ( .A1(n50929), .A2(n52239), .ZN(n50985) );
  NAND2HSV0 U54490 ( .A1(n52367), .A2(n59767), .ZN(n50981) );
  NAND2HSV0 U54491 ( .A1(\pe2/aot [12]), .A2(n52962), .ZN(n50932) );
  NAND2HSV0 U54492 ( .A1(n50930), .A2(n51805), .ZN(n50931) );
  XOR2HSV0 U54493 ( .A1(n50932), .A2(n50931), .Z(n50936) );
  NAND2HSV0 U54494 ( .A1(n53019), .A2(n51732), .ZN(n50934) );
  NAND2HSV0 U54495 ( .A1(n59358), .A2(n52859), .ZN(n50933) );
  XOR2HSV0 U54496 ( .A1(n50934), .A2(n50933), .Z(n50935) );
  XOR2HSV0 U54497 ( .A1(n50936), .A2(n50935), .Z(n50944) );
  NAND2HSV0 U54498 ( .A1(n51759), .A2(n53223), .ZN(n50938) );
  NAND2HSV0 U54499 ( .A1(n52344), .A2(n52299), .ZN(n50937) );
  XOR2HSV0 U54500 ( .A1(n50938), .A2(n50937), .Z(n50942) );
  CLKNAND2HSV0 U54501 ( .A1(\pe2/aot [6]), .A2(n43961), .ZN(n50940) );
  NAND2HSV0 U54502 ( .A1(n52056), .A2(n52965), .ZN(n50939) );
  XOR2HSV0 U54503 ( .A1(n50940), .A2(n50939), .Z(n50941) );
  XOR2HSV0 U54504 ( .A1(n50942), .A2(n50941), .Z(n50943) );
  XOR2HSV0 U54505 ( .A1(n50944), .A2(n50943), .Z(n50964) );
  NAND2HSV0 U54506 ( .A1(n37801), .A2(n52484), .ZN(n50946) );
  NAND2HSV0 U54507 ( .A1(n39029), .A2(\pe2/bq[4] ), .ZN(n50945) );
  XOR2HSV0 U54508 ( .A1(n50946), .A2(n50945), .Z(n50951) );
  NOR2HSV0 U54509 ( .A1(n50947), .A2(n51842), .ZN(n50949) );
  NAND2HSV0 U54510 ( .A1(\pe2/aot [11]), .A2(\pe2/bq[14] ), .ZN(n50948) );
  XOR2HSV0 U54511 ( .A1(n50949), .A2(n50948), .Z(n50950) );
  XNOR2HSV1 U54512 ( .A1(n50951), .A2(n50950), .ZN(n50962) );
  CLKNHSV0 U54513 ( .I(n50952), .ZN(n50954) );
  NOR2HSV0 U54514 ( .A1(n47503), .A2(n47508), .ZN(n52220) );
  AOI22HSV0 U54515 ( .A1(n52070), .A2(n52448), .B1(n59636), .B2(n51900), .ZN(
        n50953) );
  AOI21HSV2 U54516 ( .A1(n50954), .A2(n52220), .B(n50953), .ZN(n50960) );
  NAND2HSV2 U54517 ( .A1(n52858), .A2(n51614), .ZN(n52898) );
  NOR2HSV0 U54518 ( .A1(n50955), .A2(n52898), .ZN(n50958) );
  CLKNHSV0 U54519 ( .I(n50920), .ZN(n52935) );
  AOI22HSV0 U54520 ( .A1(n50956), .A2(n52935), .B1(\pe2/bq[21] ), .B2(n59978), 
        .ZN(n50957) );
  NOR2HSV1 U54521 ( .A1(n50958), .A2(n50957), .ZN(n50959) );
  XOR2HSV0 U54522 ( .A1(n50960), .A2(n50959), .Z(n50961) );
  XNOR2HSV1 U54523 ( .A1(n50962), .A2(n50961), .ZN(n50963) );
  XNOR2HSV1 U54524 ( .A1(n50964), .A2(n50963), .ZN(n50979) );
  NAND2HSV0 U54525 ( .A1(n52951), .A2(\pe2/bq[17] ), .ZN(n50966) );
  NAND2HSV0 U54526 ( .A1(\pe2/aot [7]), .A2(n52988), .ZN(n50965) );
  XOR2HSV0 U54527 ( .A1(n50966), .A2(n50965), .Z(n50970) );
  NAND2HSV0 U54528 ( .A1(n52966), .A2(n51733), .ZN(n50968) );
  NAND2HSV0 U54529 ( .A1(n59973), .A2(n52481), .ZN(n50967) );
  XOR2HSV0 U54530 ( .A1(n50968), .A2(n50967), .Z(n50969) );
  XOR2HSV0 U54531 ( .A1(n50970), .A2(n50969), .Z(n50977) );
  CLKNAND2HSV0 U54532 ( .A1(\pe2/aot [19]), .A2(\pe2/bq[6] ), .ZN(n52292) );
  XOR2HSV0 U54533 ( .A1(n50971), .A2(n52292), .Z(n50975) );
  NOR2HSV0 U54534 ( .A1(n52095), .A2(n38687), .ZN(n50973) );
  NAND2HSV0 U54535 ( .A1(\pe2/aot [2]), .A2(n52179), .ZN(n50972) );
  XOR2HSV0 U54536 ( .A1(n50973), .A2(n50972), .Z(n50974) );
  XOR2HSV0 U54537 ( .A1(n50975), .A2(n50974), .Z(n50976) );
  XOR2HSV0 U54538 ( .A1(n50977), .A2(n50976), .Z(n50978) );
  XNOR2HSV1 U54539 ( .A1(n50979), .A2(n50978), .ZN(n50980) );
  XNOR2HSV1 U54540 ( .A1(n50981), .A2(n50980), .ZN(n50983) );
  NAND2HSV0 U54541 ( .A1(n44120), .A2(n51932), .ZN(n50982) );
  XOR2HSV0 U54542 ( .A1(n50983), .A2(n50982), .Z(n50984) );
  XNOR2HSV1 U54543 ( .A1(n50985), .A2(n50984), .ZN(n50987) );
  NAND2HSV0 U54544 ( .A1(n59761), .A2(n52175), .ZN(n50986) );
  XOR3HSV2 U54545 ( .A1(n50988), .A2(n50987), .A3(n50986), .Z(n50989) );
  XNOR2HSV1 U54546 ( .A1(n50990), .A2(n50989), .ZN(n50991) );
  XNOR2HSV1 U54547 ( .A1(n50992), .A2(n50991), .ZN(n50994) );
  NAND2HSV0 U54548 ( .A1(n52251), .A2(n44714), .ZN(n50993) );
  XOR3HSV2 U54549 ( .A1(n50995), .A2(n50994), .A3(n50993), .Z(n50996) );
  XNOR2HSV1 U54550 ( .A1(n50997), .A2(n50996), .ZN(n51000) );
  NAND2HSV0 U54551 ( .A1(n59769), .A2(n52930), .ZN(n50999) );
  CLKNAND2HSV0 U54552 ( .A1(n51862), .A2(n52172), .ZN(n50998) );
  XOR3HSV2 U54553 ( .A1(n51000), .A2(n50999), .A3(n50998), .Z(n51001) );
  XNOR2HSV1 U54554 ( .A1(n51002), .A2(n51001), .ZN(n51004) );
  BUFHSV2 U54555 ( .I(n59774), .Z(n53382) );
  NAND2HSV0 U54556 ( .A1(n53382), .A2(n52051), .ZN(n51003) );
  XOR3HSV2 U54557 ( .A1(n51005), .A2(n51004), .A3(n51003), .Z(n51006) );
  XOR2HSV0 U54558 ( .A1(n51007), .A2(n51006), .Z(n51008) );
  CLKNAND2HSV0 U54559 ( .A1(n52399), .A2(n51889), .ZN(n51010) );
  CLKNAND2HSV0 U54560 ( .A1(n53359), .A2(n45816), .ZN(n51012) );
  NOR2HSV2 U54561 ( .A1(n51013), .A2(n51012), .ZN(n51107) );
  NAND2HSV2 U54562 ( .A1(n51155), .A2(n37658), .ZN(n51102) );
  CLKNAND2HSV1 U54563 ( .A1(n52564), .A2(n59949), .ZN(n51100) );
  CLKNAND2HSV0 U54564 ( .A1(n59892), .A2(n51015), .ZN(n51096) );
  CLKNAND2HSV1 U54565 ( .A1(n51016), .A2(n53286), .ZN(n51091) );
  NOR2HSV2 U54566 ( .A1(n48166), .A2(n46961), .ZN(n51086) );
  NAND2HSV0 U54567 ( .A1(n53294), .A2(n50698), .ZN(n51082) );
  CLKNAND2HSV1 U54568 ( .A1(n59882), .A2(n51017), .ZN(n51080) );
  CLKNAND2HSV1 U54569 ( .A1(n51018), .A2(n52576), .ZN(n51076) );
  CLKNAND2HSV0 U54570 ( .A1(n51019), .A2(n53211), .ZN(n51072) );
  NAND2HSV0 U54571 ( .A1(n59392), .A2(n53197), .ZN(n51070) );
  NAND2HSV0 U54572 ( .A1(n59871), .A2(n51362), .ZN(n51068) );
  NAND2HSV0 U54573 ( .A1(n52607), .A2(\pe5/bq[7] ), .ZN(n51173) );
  NOR2HSV0 U54574 ( .A1(n51173), .A2(n51020), .ZN(n51024) );
  AOI22HSV0 U54575 ( .A1(n51022), .A2(n52671), .B1(n50505), .B2(\pe5/bq[7] ), 
        .ZN(n51023) );
  NOR2HSV2 U54576 ( .A1(n51024), .A2(n51023), .ZN(n51026) );
  XNOR2HSV1 U54577 ( .A1(n51026), .A2(n51025), .ZN(n51030) );
  NAND2HSV0 U54578 ( .A1(\pe5/aot [4]), .A2(n52618), .ZN(n51027) );
  XOR2HSV0 U54579 ( .A1(n51028), .A2(n51027), .Z(n51029) );
  XOR2HSV0 U54580 ( .A1(n51030), .A2(n51029), .Z(n51066) );
  NAND2HSV0 U54581 ( .A1(\pe5/aot [16]), .A2(n50526), .ZN(n51032) );
  NAND2HSV0 U54582 ( .A1(n37700), .A2(n51276), .ZN(n51031) );
  XOR2HSV0 U54583 ( .A1(n51032), .A2(n51031), .Z(n51036) );
  CLKNAND2HSV0 U54584 ( .A1(n53323), .A2(n39592), .ZN(n51034) );
  NAND2HSV0 U54585 ( .A1(\pe5/aot [3]), .A2(\pe5/bq[19] ), .ZN(n51033) );
  XOR2HSV0 U54586 ( .A1(n51034), .A2(n51033), .Z(n51035) );
  XOR2HSV0 U54587 ( .A1(n51036), .A2(n51035), .Z(n51047) );
  NAND2HSV0 U54588 ( .A1(n59942), .A2(n53200), .ZN(n51038) );
  NAND2HSV0 U54589 ( .A1(n52591), .A2(\pe5/bq[2] ), .ZN(n51037) );
  XOR2HSV0 U54590 ( .A1(n51038), .A2(n51037), .Z(n51045) );
  NOR2HSV0 U54591 ( .A1(n51040), .A2(n51039), .ZN(n51043) );
  AOI22HSV0 U54592 ( .A1(\pe5/aot [9]), .A2(\pe5/bq[13] ), .B1(n51041), .B2(
        n52623), .ZN(n51042) );
  NOR2HSV2 U54593 ( .A1(n51043), .A2(n51042), .ZN(n51044) );
  XNOR2HSV1 U54594 ( .A1(n51045), .A2(n51044), .ZN(n51046) );
  XNOR2HSV1 U54595 ( .A1(n51047), .A2(n51046), .ZN(n51065) );
  NAND2HSV0 U54596 ( .A1(n53203), .A2(n51048), .ZN(n51050) );
  NAND2HSV0 U54597 ( .A1(n53296), .A2(n39472), .ZN(n51049) );
  XOR2HSV0 U54598 ( .A1(n51050), .A2(n51049), .Z(n51054) );
  NAND2HSV0 U54599 ( .A1(n53295), .A2(n48181), .ZN(n51052) );
  CLKNAND2HSV0 U54600 ( .A1(\pe5/aot [13]), .A2(n51307), .ZN(n51051) );
  XOR2HSV0 U54601 ( .A1(n51052), .A2(n51051), .Z(n51053) );
  XOR2HSV0 U54602 ( .A1(n51054), .A2(n51053), .Z(n51063) );
  NAND2HSV0 U54603 ( .A1(n53299), .A2(n48170), .ZN(n51056) );
  NAND2HSV0 U54604 ( .A1(\pe5/aot [10]), .A2(\pe5/bq[12] ), .ZN(n51055) );
  XOR2HSV0 U54605 ( .A1(n51056), .A2(n51055), .Z(n51061) );
  NOR2HSV0 U54606 ( .A1(n47230), .A2(n51057), .ZN(n51059) );
  NAND2HSV0 U54607 ( .A1(\pe5/aot [18]), .A2(n53307), .ZN(n51058) );
  XOR2HSV0 U54608 ( .A1(n51059), .A2(n51058), .Z(n51060) );
  XOR2HSV0 U54609 ( .A1(n51061), .A2(n51060), .Z(n51062) );
  XOR2HSV0 U54610 ( .A1(n51063), .A2(n51062), .Z(n51064) );
  XOR3HSV2 U54611 ( .A1(n51066), .A2(n51065), .A3(n51064), .Z(n51067) );
  XNOR2HSV1 U54612 ( .A1(n51068), .A2(n51067), .ZN(n51069) );
  XNOR2HSV1 U54613 ( .A1(n51070), .A2(n51069), .ZN(n51071) );
  XNOR2HSV1 U54614 ( .A1(n51072), .A2(n51071), .ZN(n51074) );
  NAND2HSV0 U54615 ( .A1(n44694), .A2(\pe5/got [4]), .ZN(n51073) );
  XOR2HSV0 U54616 ( .A1(n51074), .A2(n51073), .Z(n51075) );
  XNOR2HSV1 U54617 ( .A1(n51076), .A2(n51075), .ZN(n51078) );
  NAND2HSV0 U54618 ( .A1(n59517), .A2(n51200), .ZN(n51077) );
  XNOR2HSV1 U54619 ( .A1(n51078), .A2(n51077), .ZN(n51079) );
  XNOR2HSV1 U54620 ( .A1(n51080), .A2(n51079), .ZN(n51081) );
  XNOR2HSV1 U54621 ( .A1(n51082), .A2(n51081), .ZN(n51084) );
  NAND2HSV0 U54622 ( .A1(n52653), .A2(n51358), .ZN(n51083) );
  XNOR2HSV1 U54623 ( .A1(n51084), .A2(n51083), .ZN(n51085) );
  XNOR2HSV1 U54624 ( .A1(n51086), .A2(n51085), .ZN(n51089) );
  CLKNAND2HSV1 U54625 ( .A1(n53338), .A2(n53349), .ZN(n51088) );
  NOR2HSV1 U54626 ( .A1(n51360), .A2(n46966), .ZN(n51087) );
  XOR3HSV2 U54627 ( .A1(n51089), .A2(n51088), .A3(n51087), .Z(n51090) );
  XNOR2HSV1 U54628 ( .A1(n51091), .A2(n51090), .ZN(n51094) );
  NAND2HSV0 U54629 ( .A1(n51092), .A2(n53285), .ZN(n51093) );
  XOR2HSV0 U54630 ( .A1(n51094), .A2(n51093), .Z(n51095) );
  NAND2HSV0 U54631 ( .A1(n51227), .A2(n52658), .ZN(n51097) );
  XNOR2HSV1 U54632 ( .A1(n51100), .A2(n51099), .ZN(n51101) );
  XNOR2HSV1 U54633 ( .A1(n51102), .A2(n51101), .ZN(n51105) );
  CLKNAND2HSV0 U54634 ( .A1(n29776), .A2(n51103), .ZN(n51104) );
  XNOR2HSV1 U54635 ( .A1(n51105), .A2(n51104), .ZN(n51106) );
  XNOR2HSV1 U54636 ( .A1(n51107), .A2(n51106), .ZN(n51111) );
  NAND3HSV2 U54637 ( .A1(n51109), .A2(n31149), .A3(n51108), .ZN(n51110) );
  XOR2HSV0 U54638 ( .A1(n51111), .A2(n51110), .Z(\pe5/poht [11]) );
  MUX2HSV2 U54639 ( .I0(bo5[31]), .I1(n30344), .S(n48077), .Z(n59540) );
  NAND2HSV2 U54640 ( .A1(n59893), .A2(n52834), .ZN(n51117) );
  CLKNHSV0 U54641 ( .I(n51115), .ZN(n51116) );
  XNOR2HSV1 U54642 ( .A1(n51117), .A2(n51116), .ZN(n60010) );
  INHSV2 U54643 ( .I(n51118), .ZN(n56953) );
  CLKNAND2HSV1 U54644 ( .A1(n51939), .A2(n51120), .ZN(n51149) );
  CLKNAND2HSV1 U54645 ( .A1(n52168), .A2(n51686), .ZN(n51147) );
  CLKNAND2HSV1 U54646 ( .A1(n51893), .A2(n52239), .ZN(n51143) );
  CLKNAND2HSV1 U54647 ( .A1(n59790), .A2(n52895), .ZN(n51141) );
  CLKNAND2HSV0 U54648 ( .A1(n52920), .A2(n51688), .ZN(n51139) );
  NAND2HSV0 U54649 ( .A1(n51547), .A2(n52193), .ZN(n51123) );
  NAND2HSV0 U54650 ( .A1(n51636), .A2(n51623), .ZN(n51564) );
  CLKNAND2HSV1 U54651 ( .A1(n51547), .A2(n52309), .ZN(n52897) );
  NOR2HSV0 U54652 ( .A1(n51564), .A2(n52897), .ZN(n51122) );
  AOI21HSV2 U54653 ( .A1(n51124), .A2(n51123), .B(n51122), .ZN(n51125) );
  CLKNAND2HSV0 U54654 ( .A1(n52951), .A2(n53226), .ZN(n52870) );
  XOR2HSV0 U54655 ( .A1(n51125), .A2(n52870), .Z(n51128) );
  CLKNAND2HSV1 U54656 ( .A1(n52867), .A2(n51457), .ZN(n51539) );
  XOR2HSV0 U54657 ( .A1(n51126), .A2(n51539), .Z(n51127) );
  XOR2HSV0 U54658 ( .A1(n51128), .A2(n51127), .Z(n51137) );
  CLKNAND2HSV1 U54659 ( .A1(n59633), .A2(n52484), .ZN(n51130) );
  NAND2HSV0 U54660 ( .A1(\pe2/aot [2]), .A2(n51825), .ZN(n51129) );
  XOR2HSV0 U54661 ( .A1(n51130), .A2(n51129), .Z(n51135) );
  NOR2HSV1 U54662 ( .A1(n52200), .A2(n50920), .ZN(n51133) );
  CLKNAND2HSV0 U54663 ( .A1(n29736), .A2(n51897), .ZN(n51132) );
  XOR2HSV0 U54664 ( .A1(n51133), .A2(n51132), .Z(n51134) );
  XNOR2HSV1 U54665 ( .A1(n51135), .A2(n51134), .ZN(n51136) );
  XOR2HSV0 U54666 ( .A1(n51137), .A2(n51136), .Z(n51138) );
  XOR2HSV0 U54667 ( .A1(n51139), .A2(n51138), .Z(n51140) );
  XNOR2HSV1 U54668 ( .A1(n51141), .A2(n51140), .ZN(n51142) );
  XNOR2HSV1 U54669 ( .A1(n51143), .A2(n51142), .ZN(n51145) );
  CLKNAND2HSV1 U54670 ( .A1(n51792), .A2(n52855), .ZN(n51144) );
  XNOR2HSV1 U54671 ( .A1(n51145), .A2(n51144), .ZN(n51146) );
  XOR2HSV0 U54672 ( .A1(n51147), .A2(n51146), .Z(n51148) );
  XOR2HSV0 U54673 ( .A1(n51149), .A2(n51148), .Z(n51154) );
  CLKNAND2HSV1 U54674 ( .A1(n52047), .A2(n52890), .ZN(n51152) );
  CLKNAND2HSV1 U54675 ( .A1(n53291), .A2(n51157), .ZN(n51223) );
  NOR2HSV0 U54676 ( .A1(n51361), .A2(n46966), .ZN(n51216) );
  NAND2HSV0 U54677 ( .A1(n51158), .A2(n52641), .ZN(n51209) );
  CLKNAND2HSV1 U54678 ( .A1(n52572), .A2(n51159), .ZN(n51204) );
  NAND2HSV0 U54679 ( .A1(n51160), .A2(n51334), .ZN(n51199) );
  NOR2HSV0 U54680 ( .A1(n51164), .A2(n51163), .ZN(n51166) );
  AOI22HSV0 U54681 ( .A1(\pe5/aot [13]), .A2(\pe5/bq[11] ), .B1(n47291), .B2(
        n51419), .ZN(n51165) );
  NAND2HSV0 U54682 ( .A1(\pe5/aot [14]), .A2(\pe5/bq[10] ), .ZN(n51169) );
  NAND2HSV0 U54683 ( .A1(n52682), .A2(n51167), .ZN(n51168) );
  NAND2HSV0 U54684 ( .A1(n51363), .A2(n39454), .ZN(n51172) );
  CLKNAND2HSV1 U54685 ( .A1(n52623), .A2(\pe5/bq[7] ), .ZN(n51288) );
  NOR2HSV0 U54686 ( .A1(n51170), .A2(n51288), .ZN(n51171) );
  AOI21HSV2 U54687 ( .A1(n51173), .A2(n51172), .B(n51171), .ZN(n51175) );
  NAND2HSV0 U54688 ( .A1(\pe5/aot [7]), .A2(n51176), .ZN(n51179) );
  NAND2HSV0 U54689 ( .A1(\pe5/aot [20]), .A2(n51177), .ZN(n51178) );
  NAND2HSV0 U54690 ( .A1(\pe5/aot [23]), .A2(n53199), .ZN(n51181) );
  CLKNAND2HSV0 U54691 ( .A1(n59942), .A2(n52630), .ZN(n51180) );
  NAND2HSV0 U54692 ( .A1(n51182), .A2(n30607), .ZN(n51184) );
  NAND2HSV0 U54693 ( .A1(\pe5/aot [4]), .A2(n39487), .ZN(n51183) );
  CLKNAND2HSV0 U54694 ( .A1(n50511), .A2(n52610), .ZN(n51186) );
  NAND2HSV0 U54695 ( .A1(n59640), .A2(n52672), .ZN(n51185) );
  NAND2HSV0 U54696 ( .A1(n51187), .A2(n40226), .ZN(n51190) );
  NAND2HSV0 U54697 ( .A1(n51188), .A2(\pe5/bq[2] ), .ZN(n51189) );
  NAND2HSV0 U54698 ( .A1(\pe5/aot [10]), .A2(n52632), .ZN(n51193) );
  NAND2HSV0 U54699 ( .A1(\pe5/aot [18]), .A2(n51191), .ZN(n51192) );
  NAND2HSV0 U54700 ( .A1(\pe5/aot [9]), .A2(n39914), .ZN(n51195) );
  NAND2HSV0 U54701 ( .A1(n52611), .A2(n50668), .ZN(n51194) );
  NAND2HSV0 U54702 ( .A1(n52600), .A2(n31190), .ZN(n51197) );
  NAND2HSV0 U54703 ( .A1(n53299), .A2(\pe5/bq[12] ), .ZN(n51196) );
  XNOR2HSV1 U54704 ( .A1(n51199), .A2(n51198), .ZN(n51202) );
  NAND2HSV0 U54705 ( .A1(n44694), .A2(n51200), .ZN(n51201) );
  XOR2HSV0 U54706 ( .A1(n51202), .A2(n51201), .Z(n51203) );
  XNOR2HSV1 U54707 ( .A1(n51204), .A2(n51203), .ZN(n51207) );
  NAND2HSV0 U54708 ( .A1(n51205), .A2(n47144), .ZN(n51206) );
  XNOR2HSV1 U54709 ( .A1(n51207), .A2(n51206), .ZN(n51208) );
  XNOR2HSV1 U54710 ( .A1(n51209), .A2(n51208), .ZN(n51214) );
  CLKNAND2HSV1 U54711 ( .A1(n52569), .A2(n51210), .ZN(n51213) );
  CLKNAND2HSV0 U54712 ( .A1(n51211), .A2(n59643), .ZN(n51212) );
  XOR3HSV2 U54713 ( .A1(n51214), .A2(n51213), .A3(n51212), .Z(n51215) );
  XNOR2HSV1 U54714 ( .A1(n51216), .A2(n51215), .ZN(n51221) );
  NOR2HSV1 U54715 ( .A1(n51217), .A2(n45817), .ZN(n51220) );
  NOR2HSV1 U54716 ( .A1(n51218), .A2(n31199), .ZN(n51219) );
  XOR3HSV2 U54717 ( .A1(n51221), .A2(n51220), .A3(n51219), .Z(n51222) );
  XNOR2HSV1 U54718 ( .A1(n51223), .A2(n51222), .ZN(n51226) );
  NAND2HSV0 U54719 ( .A1(n53344), .A2(n51224), .ZN(n51225) );
  NAND2HSV2 U54720 ( .A1(n51230), .A2(n51229), .ZN(n52667) );
  INHSV2 U54721 ( .I(n51231), .ZN(n53211) );
  NAND2HSV2 U54722 ( .A1(n52667), .A2(n53211), .ZN(n51245) );
  CLKNAND2HSV1 U54723 ( .A1(n59933), .A2(n51362), .ZN(n51241) );
  CLKNAND2HSV1 U54724 ( .A1(n53203), .A2(n51420), .ZN(n51234) );
  CLKNAND2HSV0 U54725 ( .A1(n51182), .A2(n51336), .ZN(n51233) );
  XOR2HSV0 U54726 ( .A1(n51234), .A2(n51233), .Z(n51239) );
  CLKNAND2HSV1 U54727 ( .A1(\pe5/aot [3]), .A2(\pe5/bq[2] ), .ZN(n51237) );
  CLKNAND2HSV1 U54728 ( .A1(\pe5/aot [4]), .A2(n52581), .ZN(n51236) );
  XOR2HSV0 U54729 ( .A1(n51237), .A2(n51236), .Z(n51238) );
  XOR2HSV0 U54730 ( .A1(n51239), .A2(n51238), .Z(n51240) );
  XNOR2HSV1 U54731 ( .A1(n51241), .A2(n51240), .ZN(n51243) );
  CLKNAND2HSV1 U54732 ( .A1(n29776), .A2(n59357), .ZN(n51242) );
  XNOR2HSV2 U54733 ( .A1(n51243), .A2(n51242), .ZN(n51244) );
  NAND2HSV0 U54734 ( .A1(n29771), .A2(n51418), .ZN(n51246) );
  CLKNAND2HSV1 U54735 ( .A1(n52669), .A2(n51418), .ZN(n51267) );
  INHSV2 U54736 ( .I(n47199), .ZN(n52835) );
  CLKNAND2HSV0 U54737 ( .A1(n52835), .A2(n59355), .ZN(n51265) );
  CLKNAND2HSV1 U54738 ( .A1(n53290), .A2(n51362), .ZN(n51261) );
  NAND2HSV0 U54739 ( .A1(n52682), .A2(\pe5/bq[2] ), .ZN(n51249) );
  CLKNAND2HSV0 U54740 ( .A1(n51247), .A2(n52581), .ZN(n51248) );
  XOR2HSV0 U54741 ( .A1(n51249), .A2(n51248), .Z(n51253) );
  CLKNAND2HSV0 U54742 ( .A1(n59895), .A2(\pe5/bq[7] ), .ZN(n51251) );
  NAND2HSV0 U54743 ( .A1(\pe5/aot [4]), .A2(n51336), .ZN(n51250) );
  XOR2HSV0 U54744 ( .A1(n51251), .A2(n51250), .Z(n51252) );
  XOR2HSV0 U54745 ( .A1(n51253), .A2(n51252), .Z(n51259) );
  CLKNAND2HSV0 U54746 ( .A1(n59945), .A2(n51281), .ZN(n51255) );
  CLKNAND2HSV1 U54747 ( .A1(\pe5/aot [3]), .A2(n51373), .ZN(n51254) );
  XOR2HSV0 U54748 ( .A1(n51255), .A2(n51254), .Z(n51257) );
  NOR2HSV2 U54749 ( .A1(n51232), .A2(n46136), .ZN(n51256) );
  XNOR2HSV1 U54750 ( .A1(n51257), .A2(n51256), .ZN(n51258) );
  XNOR2HSV1 U54751 ( .A1(n51259), .A2(n51258), .ZN(n51260) );
  XNOR2HSV1 U54752 ( .A1(n51261), .A2(n51260), .ZN(n51263) );
  CLKNAND2HSV0 U54753 ( .A1(n52693), .A2(n59357), .ZN(n51262) );
  XNOR2HSV1 U54754 ( .A1(n51263), .A2(n51262), .ZN(n51264) );
  XNOR2HSV1 U54755 ( .A1(n51265), .A2(n51264), .ZN(n51266) );
  NAND2HSV2 U54756 ( .A1(n29779), .A2(\pe5/got [5]), .ZN(n51268) );
  XNOR2HSV1 U54757 ( .A1(n51269), .A2(n51268), .ZN(n51270) );
  NAND2HSV0 U54758 ( .A1(n59893), .A2(n53211), .ZN(n51301) );
  NOR2HSV2 U54759 ( .A1(n51273), .A2(n51306), .ZN(n51299) );
  CLKNAND2HSV0 U54760 ( .A1(n59903), .A2(n51362), .ZN(n51297) );
  CLKNAND2HSV1 U54761 ( .A1(n53295), .A2(\pe5/bq[6] ), .ZN(n51275) );
  NAND2HSV0 U54762 ( .A1(n51339), .A2(\pe5/bq[11] ), .ZN(n51274) );
  XOR2HSV0 U54763 ( .A1(n51275), .A2(n51274), .Z(n51280) );
  CLKNAND2HSV1 U54764 ( .A1(n51313), .A2(\pe5/bq[2] ), .ZN(n51278) );
  NAND2HSV0 U54765 ( .A1(n53323), .A2(n51276), .ZN(n51277) );
  XOR2HSV0 U54766 ( .A1(n51278), .A2(n51277), .Z(n51279) );
  XOR2HSV0 U54767 ( .A1(n51280), .A2(n51279), .Z(n51287) );
  NOR2HSV0 U54768 ( .A1(n59869), .A2(n47162), .ZN(n51283) );
  CLKNAND2HSV0 U54769 ( .A1(\pe5/aot [9]), .A2(n51281), .ZN(n51282) );
  XOR2HSV0 U54770 ( .A1(n51283), .A2(n51282), .Z(n51285) );
  XNOR2HSV1 U54771 ( .A1(n51285), .A2(n51284), .ZN(n51286) );
  XNOR2HSV1 U54772 ( .A1(n51287), .A2(n51286), .ZN(n51295) );
  XOR2HSV0 U54773 ( .A1(n51289), .A2(n51288), .Z(n51293) );
  NOR2HSV0 U54774 ( .A1(n47230), .A2(n51021), .ZN(n51291) );
  NAND2HSV0 U54775 ( .A1(\pe5/aot [4]), .A2(n50675), .ZN(n51290) );
  XOR2HSV0 U54776 ( .A1(n51291), .A2(n51290), .Z(n51292) );
  XOR2HSV0 U54777 ( .A1(n51293), .A2(n51292), .Z(n51294) );
  XNOR2HSV1 U54778 ( .A1(n51295), .A2(n51294), .ZN(n51296) );
  XNOR2HSV1 U54779 ( .A1(n51297), .A2(n51296), .ZN(n51298) );
  XNOR2HSV1 U54780 ( .A1(n51299), .A2(n51298), .ZN(n51300) );
  XNOR2HSV1 U54781 ( .A1(n51301), .A2(n51300), .ZN(n51304) );
  CLKNAND2HSV0 U54782 ( .A1(n51092), .A2(n51302), .ZN(n51303) );
  INHSV2 U54783 ( .I(n51306), .ZN(n53197) );
  NAND2HSV0 U54784 ( .A1(n59893), .A2(n53197), .ZN(n51330) );
  NOR2HSV1 U54785 ( .A1(n51360), .A2(n48625), .ZN(n51328) );
  NAND2HSV0 U54786 ( .A1(n51247), .A2(n51336), .ZN(n51309) );
  NAND2HSV0 U54787 ( .A1(n53203), .A2(n51307), .ZN(n51308) );
  XOR2HSV0 U54788 ( .A1(n51309), .A2(n51308), .Z(n51326) );
  NAND2HSV0 U54789 ( .A1(n51310), .A2(n52671), .ZN(n51312) );
  CLKNAND2HSV0 U54790 ( .A1(n59895), .A2(n53216), .ZN(n51311) );
  XOR2HSV0 U54791 ( .A1(n51312), .A2(n51311), .Z(n51317) );
  NOR2HSV1 U54792 ( .A1(n47409), .A2(n46136), .ZN(n51315) );
  NAND2HSV0 U54793 ( .A1(n51313), .A2(n52581), .ZN(n51314) );
  XOR2HSV0 U54794 ( .A1(n51315), .A2(n51314), .Z(n51316) );
  XNOR2HSV1 U54795 ( .A1(n51317), .A2(n51316), .ZN(n51325) );
  CLKNAND2HSV1 U54796 ( .A1(n39887), .A2(\pe5/bq[2] ), .ZN(n51319) );
  NAND2HSV0 U54797 ( .A1(n59880), .A2(n51420), .ZN(n51318) );
  XOR2HSV0 U54798 ( .A1(n51319), .A2(n51318), .Z(n51323) );
  NOR2HSV0 U54799 ( .A1(n59869), .A2(n46916), .ZN(n51321) );
  NAND2HSV0 U54800 ( .A1(n50501), .A2(\pe5/bq[7] ), .ZN(n51320) );
  XOR2HSV0 U54801 ( .A1(n51321), .A2(n51320), .Z(n51322) );
  XOR2HSV0 U54802 ( .A1(n51323), .A2(n51322), .Z(n51324) );
  XOR3HSV2 U54803 ( .A1(n51326), .A2(n51325), .A3(n51324), .Z(n51327) );
  XOR2HSV0 U54804 ( .A1(n51328), .A2(n51327), .Z(n51329) );
  XNOR2HSV1 U54805 ( .A1(n51330), .A2(n51329), .ZN(n51333) );
  NAND2HSV0 U54806 ( .A1(n51399), .A2(n51331), .ZN(n51332) );
  NAND2HSV2 U54807 ( .A1(n52667), .A2(n52576), .ZN(n51356) );
  CLKNAND2HSV1 U54808 ( .A1(n52564), .A2(n59357), .ZN(n51351) );
  NAND2HSV2 U54809 ( .A1(n51335), .A2(\pe5/got [1]), .ZN(n51349) );
  CLKNAND2HSV0 U54810 ( .A1(\pe5/aot [3]), .A2(n51336), .ZN(n51338) );
  CLKNAND2HSV0 U54811 ( .A1(\pe5/aot [4]), .A2(n51281), .ZN(n51337) );
  XOR2HSV0 U54812 ( .A1(n51338), .A2(n51337), .Z(n51343) );
  CLKNAND2HSV1 U54813 ( .A1(n53203), .A2(n52671), .ZN(n51341) );
  CLKNAND2HSV1 U54814 ( .A1(n51339), .A2(\pe5/bq[6] ), .ZN(n51340) );
  XOR2HSV0 U54815 ( .A1(n51341), .A2(n51340), .Z(n51342) );
  XNOR2HSV1 U54816 ( .A1(n51343), .A2(n51342), .ZN(n51347) );
  CLKNAND2HSV0 U54817 ( .A1(n59945), .A2(\pe5/bq[2] ), .ZN(n51345) );
  CLKNAND2HSV1 U54818 ( .A1(n52682), .A2(n51276), .ZN(n51344) );
  XOR2HSV0 U54819 ( .A1(n51345), .A2(n51344), .Z(n51346) );
  XNOR2HSV1 U54820 ( .A1(n51347), .A2(n51346), .ZN(n51348) );
  XNOR2HSV1 U54821 ( .A1(n51349), .A2(n51348), .ZN(n51350) );
  XNOR2HSV1 U54822 ( .A1(n51351), .A2(n51350), .ZN(n51354) );
  CLKNAND2HSV1 U54823 ( .A1(n52669), .A2(n52579), .ZN(n51353) );
  NAND2HSV2 U54824 ( .A1(n29775), .A2(n52577), .ZN(n51352) );
  XOR3HSV2 U54825 ( .A1(n51354), .A2(n51353), .A3(n51352), .Z(n51355) );
  NAND2HSV0 U54826 ( .A1(n53210), .A2(\pe5/got [6]), .ZN(n51357) );
  NAND2HSV2 U54827 ( .A1(n52668), .A2(n48167), .ZN(n51415) );
  CLKNAND2HSV1 U54828 ( .A1(n51014), .A2(n51358), .ZN(n51408) );
  CLKNAND2HSV0 U54829 ( .A1(n59892), .A2(n51359), .ZN(n51403) );
  NAND2HSV0 U54830 ( .A1(n59893), .A2(n51334), .ZN(n51398) );
  NOR2HSV1 U54831 ( .A1(n51360), .A2(n50550), .ZN(n51396) );
  NAND2HSV0 U54832 ( .A1(n59903), .A2(n59355), .ZN(n51394) );
  NOR2HSV0 U54833 ( .A1(n51361), .A2(n51306), .ZN(n51392) );
  NAND2HSV0 U54834 ( .A1(n52653), .A2(n51362), .ZN(n51390) );
  NAND2HSV0 U54835 ( .A1(\pe5/aot [13]), .A2(n53199), .ZN(n51365) );
  NAND2HSV0 U54836 ( .A1(n51363), .A2(n50533), .ZN(n51364) );
  XOR2HSV0 U54837 ( .A1(n51365), .A2(n51364), .Z(n51369) );
  NAND2HSV0 U54838 ( .A1(\pe5/aot [4]), .A2(n53216), .ZN(n51367) );
  NAND2HSV0 U54839 ( .A1(n51339), .A2(\pe5/bq[13] ), .ZN(n51366) );
  XOR2HSV0 U54840 ( .A1(n51367), .A2(n51366), .Z(n51368) );
  XOR2HSV0 U54841 ( .A1(n51369), .A2(n51368), .Z(n51379) );
  CLKNAND2HSV0 U54842 ( .A1(\pe5/aot [2]), .A2(n39615), .ZN(n51372) );
  CLKNAND2HSV0 U54843 ( .A1(n51313), .A2(n51370), .ZN(n51371) );
  XOR2HSV0 U54844 ( .A1(n51372), .A2(n51371), .Z(n51377) );
  NAND2HSV0 U54845 ( .A1(n39887), .A2(n51373), .ZN(n51375) );
  NAND2HSV0 U54846 ( .A1(n52675), .A2(n50526), .ZN(n51374) );
  XOR2HSV0 U54847 ( .A1(n51375), .A2(n51374), .Z(n51376) );
  XOR2HSV0 U54848 ( .A1(n51377), .A2(n51376), .Z(n51378) );
  XOR2HSV0 U54849 ( .A1(n51379), .A2(n51378), .Z(n51388) );
  CLKNAND2HSV1 U54850 ( .A1(\pe5/aot [3]), .A2(\pe5/bq[11] ), .ZN(n51381) );
  NAND2HSV0 U54851 ( .A1(n59896), .A2(\pe5/bq[2] ), .ZN(n51380) );
  XOR2HSV0 U54852 ( .A1(n51381), .A2(n51380), .Z(n51385) );
  XOR2HSV0 U54853 ( .A1(n51383), .A2(n51382), .Z(n51384) );
  XOR3HSV2 U54854 ( .A1(n51386), .A2(n51385), .A3(n51384), .Z(n51387) );
  XNOR2HSV1 U54855 ( .A1(n51388), .A2(n51387), .ZN(n51389) );
  XOR2HSV0 U54856 ( .A1(n51390), .A2(n51389), .Z(n51391) );
  XOR2HSV0 U54857 ( .A1(n51392), .A2(n51391), .Z(n51393) );
  XNOR2HSV1 U54858 ( .A1(n51394), .A2(n51393), .ZN(n51395) );
  XNOR2HSV1 U54859 ( .A1(n51396), .A2(n51395), .ZN(n51397) );
  XNOR2HSV1 U54860 ( .A1(n51398), .A2(n51397), .ZN(n51401) );
  CLKNAND2HSV0 U54861 ( .A1(n51399), .A2(\pe5/got [6]), .ZN(n51400) );
  XNOR2HSV1 U54862 ( .A1(n51401), .A2(n51400), .ZN(n51402) );
  XNOR2HSV1 U54863 ( .A1(n51403), .A2(n51402), .ZN(n51406) );
  CLKNAND2HSV0 U54864 ( .A1(n51404), .A2(n47144), .ZN(n51405) );
  XNOR2HSV1 U54865 ( .A1(n51406), .A2(n51405), .ZN(n51407) );
  XNOR2HSV1 U54866 ( .A1(n51408), .A2(n51407), .ZN(n51410) );
  NOR2HSV1 U54867 ( .A1(n47139), .A2(n46961), .ZN(n51409) );
  XOR2HSV0 U54868 ( .A1(n51410), .A2(n51409), .Z(n51413) );
  NAND2HSV0 U54869 ( .A1(n51411), .A2(n59643), .ZN(n51412) );
  XOR2HSV0 U54870 ( .A1(n51413), .A2(n51412), .Z(n51414) );
  XNOR2HSV1 U54871 ( .A1(n51417), .A2(n51416), .ZN(\pe5/poht [19]) );
  NAND2HSV0 U54872 ( .A1(n51014), .A2(n51362), .ZN(n51429) );
  NOR2HSV0 U54873 ( .A1(n45904), .A2(n51021), .ZN(n51427) );
  NAND2HSV2 U54874 ( .A1(n51419), .A2(n53307), .ZN(n51422) );
  CLKNAND2HSV1 U54875 ( .A1(\pe5/aot [3]), .A2(n51420), .ZN(n51421) );
  XOR2HSV0 U54876 ( .A1(n51422), .A2(n51421), .Z(n51426) );
  CLKNAND2HSV0 U54877 ( .A1(n59945), .A2(n53199), .ZN(n51424) );
  CLKNAND2HSV0 U54878 ( .A1(\pe5/aot [4]), .A2(\pe5/bq[2] ), .ZN(n51423) );
  XOR2HSV0 U54879 ( .A1(n51424), .A2(n51423), .Z(n51425) );
  XOR3HSV2 U54880 ( .A1(n51427), .A2(n51426), .A3(n51425), .Z(n51428) );
  XNOR2HSV1 U54881 ( .A1(n51429), .A2(n51428), .ZN(n51432) );
  CLKNAND2HSV1 U54882 ( .A1(n59933), .A2(n53197), .ZN(n51431) );
  CLKNAND2HSV1 U54883 ( .A1(n29778), .A2(n53211), .ZN(n51430) );
  XOR3HSV2 U54884 ( .A1(n51432), .A2(n51431), .A3(n51430), .Z(n51433) );
  NAND2HSV0 U54885 ( .A1(n53210), .A2(n52576), .ZN(n51435) );
  XNOR2HSV1 U54886 ( .A1(n51436), .A2(n51435), .ZN(\pe5/poht [27]) );
  BUFHSV2 U54887 ( .I(n51437), .Z(n51440) );
  NOR2HSV0 U54888 ( .A1(n51441), .A2(n52710), .ZN(n51442) );
  XOR2HSV0 U54889 ( .A1(n51442), .A2(poh6[9]), .Z(po[10]) );
  NOR2HSV0 U54890 ( .A1(n51443), .A2(n52701), .ZN(n51444) );
  XOR2HSV0 U54891 ( .A1(n51444), .A2(poh6[11]), .Z(po[12]) );
  NOR2HSV2 U54892 ( .A1(n29748), .A2(n32793), .ZN(n51446) );
  XOR2HSV0 U54893 ( .A1(n51446), .A2(poh6[12]), .Z(po[13]) );
  XOR2HSV0 U54894 ( .A1(n51447), .A2(poh6[18]), .Z(po[19]) );
  OAI21HSV0 U54895 ( .A1(n51450), .A2(n51449), .B(n51448), .ZN(n60061) );
  CLKNAND2HSV1 U54896 ( .A1(n53087), .A2(n52175), .ZN(n51483) );
  CLKNAND2HSV0 U54897 ( .A1(n52919), .A2(n52855), .ZN(n51481) );
  NAND2HSV0 U54898 ( .A1(n44968), .A2(n52900), .ZN(n51479) );
  CLKNAND2HSV0 U54899 ( .A1(n51868), .A2(n51932), .ZN(n51477) );
  NAND2HSV0 U54900 ( .A1(n60002), .A2(n51688), .ZN(n51475) );
  NOR2HSV0 U54901 ( .A1(n51453), .A2(n51452), .ZN(n51455) );
  AOI22HSV0 U54902 ( .A1(n52951), .A2(n51803), .B1(n52322), .B2(n52344), .ZN(
        n51454) );
  NOR2HSV2 U54903 ( .A1(n51455), .A2(n51454), .ZN(n51456) );
  XOR2HSV0 U54904 ( .A1(n51456), .A2(n51540), .Z(n51473) );
  NAND2HSV0 U54905 ( .A1(n59633), .A2(n51897), .ZN(n51459) );
  NAND2HSV0 U54906 ( .A1(n52056), .A2(n51457), .ZN(n51458) );
  XOR2HSV0 U54907 ( .A1(n51459), .A2(n51458), .Z(n51464) );
  NOR2HSV2 U54908 ( .A1(n52095), .A2(n47508), .ZN(n51462) );
  NAND2HSV0 U54909 ( .A1(n51460), .A2(n51493), .ZN(n51461) );
  XOR2HSV0 U54910 ( .A1(n51462), .A2(n51461), .Z(n51463) );
  XNOR2HSV1 U54911 ( .A1(n51464), .A2(n51463), .ZN(n51472) );
  NAND2HSV0 U54912 ( .A1(\pe2/aot [2]), .A2(n52448), .ZN(n51466) );
  NAND2HSV0 U54913 ( .A1(n52456), .A2(n52866), .ZN(n51465) );
  XOR2HSV0 U54914 ( .A1(n51466), .A2(n51465), .Z(n51470) );
  CLKNAND2HSV0 U54915 ( .A1(n59768), .A2(n52484), .ZN(n51468) );
  NAND2HSV0 U54916 ( .A1(n59976), .A2(\pe2/bq[1] ), .ZN(n51467) );
  XOR2HSV0 U54917 ( .A1(n51468), .A2(n51467), .Z(n51469) );
  XOR2HSV0 U54918 ( .A1(n51470), .A2(n51469), .Z(n51471) );
  XOR3HSV2 U54919 ( .A1(n51473), .A2(n51472), .A3(n51471), .Z(n51474) );
  XNOR2HSV1 U54920 ( .A1(n51475), .A2(n51474), .ZN(n51476) );
  XNOR2HSV1 U54921 ( .A1(n51477), .A2(n51476), .ZN(n51478) );
  XOR2HSV0 U54922 ( .A1(n51479), .A2(n51478), .Z(n51480) );
  XOR2HSV0 U54923 ( .A1(n51481), .A2(n51480), .Z(n51482) );
  CLKNAND2HSV1 U54924 ( .A1(n51792), .A2(n51939), .ZN(n51484) );
  CLKNAND2HSV1 U54925 ( .A1(n52047), .A2(\pe2/got [10]), .ZN(n51527) );
  CLKNAND2HSV0 U54926 ( .A1(n59475), .A2(n52052), .ZN(n51525) );
  CLKNAND2HSV1 U54927 ( .A1(n53087), .A2(n51939), .ZN(n51519) );
  CLKNAND2HSV0 U54928 ( .A1(n59790), .A2(n51686), .ZN(n51517) );
  NAND2HSV0 U54929 ( .A1(n51799), .A2(n52855), .ZN(n51515) );
  NAND2HSV0 U54930 ( .A1(n60002), .A2(n51932), .ZN(n51513) );
  NAND2HSV0 U54931 ( .A1(n51485), .A2(n51688), .ZN(n51510) );
  NAND2HSV0 U54932 ( .A1(n51486), .A2(n52322), .ZN(n51488) );
  NAND2HSV0 U54933 ( .A1(n53019), .A2(n51803), .ZN(n51487) );
  XOR2HSV0 U54934 ( .A1(n51488), .A2(n51487), .Z(n51492) );
  CLKNAND2HSV0 U54935 ( .A1(\pe2/aot [7]), .A2(\pe2/bq[6] ), .ZN(n51490) );
  CLKNAND2HSV0 U54936 ( .A1(n52951), .A2(n51897), .ZN(n51489) );
  XOR2HSV0 U54937 ( .A1(n51490), .A2(n51489), .Z(n51491) );
  XOR2HSV0 U54938 ( .A1(n51492), .A2(n51491), .Z(n51501) );
  NAND2HSV0 U54939 ( .A1(n59976), .A2(n51493), .ZN(n51495) );
  NAND2HSV0 U54940 ( .A1(n52456), .A2(n51832), .ZN(n51494) );
  XOR2HSV0 U54941 ( .A1(n51495), .A2(n51494), .Z(n51499) );
  NAND2HSV0 U54942 ( .A1(n51547), .A2(n51733), .ZN(n51497) );
  NAND2HSV0 U54943 ( .A1(\pe2/aot [2]), .A2(n52073), .ZN(n51496) );
  XOR2HSV0 U54944 ( .A1(n51497), .A2(n51496), .Z(n51498) );
  XOR2HSV0 U54945 ( .A1(n51499), .A2(n51498), .Z(n51500) );
  XOR2HSV0 U54946 ( .A1(n51501), .A2(n51500), .Z(n51508) );
  CLKNAND2HSV0 U54947 ( .A1(n59977), .A2(n52484), .ZN(n51503) );
  NAND2HSV0 U54948 ( .A1(n52056), .A2(n51825), .ZN(n51502) );
  XOR2HSV0 U54949 ( .A1(n51503), .A2(n51502), .Z(n51506) );
  NAND2HSV0 U54950 ( .A1(\pe2/aot [12]), .A2(n51532), .ZN(n51703) );
  NAND2HSV0 U54951 ( .A1(n52867), .A2(n51997), .ZN(n51504) );
  XOR2HSV0 U54952 ( .A1(n51703), .A2(n51504), .Z(n51505) );
  XOR2HSV0 U54953 ( .A1(n51506), .A2(n51505), .Z(n51507) );
  XNOR2HSV1 U54954 ( .A1(n51508), .A2(n51507), .ZN(n51509) );
  XNOR2HSV1 U54955 ( .A1(n51510), .A2(n51509), .ZN(n51512) );
  CLKNAND2HSV0 U54956 ( .A1(n51868), .A2(n52900), .ZN(n51511) );
  XOR3HSV2 U54957 ( .A1(n51513), .A2(n51512), .A3(n51511), .Z(n51514) );
  XOR2HSV0 U54958 ( .A1(n51515), .A2(n51514), .Z(n51516) );
  XOR2HSV0 U54959 ( .A1(n51517), .A2(n51516), .Z(n51518) );
  XNOR2HSV1 U54960 ( .A1(n51519), .A2(n51518), .ZN(n51521) );
  CLKNAND2HSV1 U54961 ( .A1(n25828), .A2(n52890), .ZN(n51520) );
  XNOR2HSV1 U54962 ( .A1(n51521), .A2(n51520), .ZN(n51522) );
  XOR2HSV0 U54963 ( .A1(n51523), .A2(n51522), .Z(n51524) );
  XOR2HSV0 U54964 ( .A1(n51525), .A2(n51524), .Z(n51526) );
  NAND2HSV2 U54965 ( .A1(n25709), .A2(n51892), .ZN(n51528) );
  XNOR2HSV4 U54966 ( .A1(n51529), .A2(n51528), .ZN(n51531) );
  CLKNAND2HSV0 U54967 ( .A1(n59794), .A2(\pe2/got [12]), .ZN(n51530) );
  XNOR2HSV4 U54968 ( .A1(n51531), .A2(n51530), .ZN(\pe2/poht [20]) );
  CLKNAND2HSV0 U54969 ( .A1(n52919), .A2(n52900), .ZN(n51560) );
  NAND2HSV0 U54970 ( .A1(n59522), .A2(n51932), .ZN(n51558) );
  CLKNAND2HSV1 U54971 ( .A1(n51782), .A2(n51688), .ZN(n51556) );
  NAND2HSV0 U54972 ( .A1(n59633), .A2(n52309), .ZN(n51534) );
  NAND2HSV0 U54973 ( .A1(n59977), .A2(n51532), .ZN(n51533) );
  XOR2HSV0 U54974 ( .A1(n51534), .A2(n51533), .Z(n51554) );
  NAND2HSV0 U54975 ( .A1(n59768), .A2(n53226), .ZN(n51536) );
  NAND2HSV0 U54976 ( .A1(n52951), .A2(n52484), .ZN(n51535) );
  XOR2HSV0 U54977 ( .A1(n51536), .A2(n51535), .Z(n51544) );
  NOR2HSV0 U54978 ( .A1(n51537), .A2(n49529), .ZN(n51542) );
  NOR2HSV0 U54979 ( .A1(n51538), .A2(n51567), .ZN(n51541) );
  OAI22HSV2 U54980 ( .A1(n51542), .A2(n51541), .B1(n51540), .B2(n51539), .ZN(
        n51543) );
  XNOR2HSV1 U54981 ( .A1(n51544), .A2(n51543), .ZN(n51553) );
  NAND2HSV0 U54982 ( .A1(n52456), .A2(n51897), .ZN(n51546) );
  NAND2HSV0 U54983 ( .A1(n52056), .A2(n52866), .ZN(n51545) );
  XOR2HSV0 U54984 ( .A1(n51546), .A2(n51545), .Z(n51551) );
  NOR2HSV1 U54985 ( .A1(n49618), .A2(n47511), .ZN(n51549) );
  NAND2HSV0 U54986 ( .A1(n51547), .A2(n51997), .ZN(n51548) );
  XOR2HSV0 U54987 ( .A1(n51549), .A2(n51548), .Z(n51550) );
  XOR2HSV0 U54988 ( .A1(n51551), .A2(n51550), .Z(n51552) );
  XOR3HSV2 U54989 ( .A1(n51554), .A2(n51553), .A3(n51552), .Z(n51555) );
  XNOR2HSV1 U54990 ( .A1(n51556), .A2(n51555), .ZN(n51557) );
  XOR2HSV0 U54991 ( .A1(n51558), .A2(n51557), .Z(n51559) );
  XOR2HSV0 U54992 ( .A1(n51560), .A2(n51559), .Z(n51562) );
  CLKNAND2HSV1 U54993 ( .A1(n51878), .A2(n51686), .ZN(n51561) );
  CLKNAND2HSV1 U54994 ( .A1(n52902), .A2(\pe2/got [12]), .ZN(n51606) );
  CLKNAND2HSV0 U54995 ( .A1(n59475), .A2(n51892), .ZN(n51605) );
  CLKNAND2HSV1 U54996 ( .A1(n51797), .A2(\pe2/got [10]), .ZN(n51603) );
  CLKNAND2HSV1 U54997 ( .A1(n51893), .A2(n59371), .ZN(n51599) );
  CLKNAND2HSV0 U54998 ( .A1(n59790), .A2(n51895), .ZN(n51597) );
  NAND2HSV0 U54999 ( .A1(n59522), .A2(n51939), .ZN(n51595) );
  NOR2HSV1 U55000 ( .A1(n52171), .A2(n50909), .ZN(n51593) );
  CLKNAND2HSV1 U55001 ( .A1(n52923), .A2(n51933), .ZN(n51590) );
  NAND2HSV0 U55002 ( .A1(n59792), .A2(n51733), .ZN(n52436) );
  XOR2HSV0 U55003 ( .A1(n51563), .A2(n52436), .Z(n51566) );
  CLKNAND2HSV1 U55004 ( .A1(n51921), .A2(n51919), .ZN(n51704) );
  XOR2HSV0 U55005 ( .A1(n51564), .A2(n51704), .Z(n51565) );
  XOR2HSV0 U55006 ( .A1(n51566), .A2(n51565), .Z(n51575) );
  CLKNAND2HSV0 U55007 ( .A1(n51460), .A2(n51897), .ZN(n51569) );
  INHSV2 U55008 ( .I(n51567), .ZN(n53223) );
  NAND2HSV0 U55009 ( .A1(n59633), .A2(n53223), .ZN(n51568) );
  XOR2HSV0 U55010 ( .A1(n51569), .A2(n51568), .Z(n51573) );
  NAND2HSV0 U55011 ( .A1(\pe2/aot [2]), .A2(n52472), .ZN(n51571) );
  NAND2HSV0 U55012 ( .A1(n59783), .A2(\pe2/bq[14] ), .ZN(n51570) );
  XOR2HSV0 U55013 ( .A1(n51571), .A2(n51570), .Z(n51572) );
  XNOR2HSV1 U55014 ( .A1(n51573), .A2(n51572), .ZN(n51574) );
  XNOR2HSV1 U55015 ( .A1(n51575), .A2(n51574), .ZN(n51585) );
  NAND2HSV0 U55016 ( .A1(n51824), .A2(n51900), .ZN(n51577) );
  NAND2HSV0 U55017 ( .A1(n53019), .A2(\pe2/bq[6] ), .ZN(n51576) );
  XOR2HSV0 U55018 ( .A1(n51577), .A2(n51576), .Z(n51581) );
  NAND2HSV0 U55019 ( .A1(n52951), .A2(n51832), .ZN(n51579) );
  NAND2HSV0 U55020 ( .A1(n53005), .A2(n52905), .ZN(n51578) );
  XOR2HSV0 U55021 ( .A1(n51579), .A2(n51578), .Z(n51580) );
  XNOR2HSV1 U55022 ( .A1(n51581), .A2(n51580), .ZN(n51583) );
  NOR2HSV0 U55023 ( .A1(n45165), .A2(n50920), .ZN(n52937) );
  CLKNAND2HSV0 U55024 ( .A1(n59976), .A2(n51803), .ZN(n52939) );
  XOR2HSV0 U55025 ( .A1(n52937), .A2(n52939), .Z(n51582) );
  XNOR2HSV1 U55026 ( .A1(n51583), .A2(n51582), .ZN(n51584) );
  XNOR2HSV1 U55027 ( .A1(n51585), .A2(n51584), .ZN(n51588) );
  NAND2HSV0 U55028 ( .A1(n59769), .A2(n52896), .ZN(n51587) );
  CLKNAND2HSV0 U55029 ( .A1(n52534), .A2(n52895), .ZN(n51586) );
  XOR3HSV2 U55030 ( .A1(n51588), .A2(n51587), .A3(n51586), .Z(n51589) );
  XNOR2HSV1 U55031 ( .A1(n51590), .A2(n51589), .ZN(n51592) );
  CLKNAND2HSV0 U55032 ( .A1(n51868), .A2(n51686), .ZN(n51591) );
  XOR3HSV2 U55033 ( .A1(n51593), .A2(n51592), .A3(n51591), .Z(n51594) );
  XOR2HSV0 U55034 ( .A1(n51595), .A2(n51594), .Z(n51596) );
  XOR2HSV0 U55035 ( .A1(n51597), .A2(n51596), .Z(n51598) );
  XNOR2HSV1 U55036 ( .A1(n51599), .A2(n51598), .ZN(n51601) );
  CLKNAND2HSV1 U55037 ( .A1(n51878), .A2(n52052), .ZN(n51600) );
  XNOR2HSV1 U55038 ( .A1(n51601), .A2(n51600), .ZN(n51602) );
  XOR2HSV0 U55039 ( .A1(n51603), .A2(n51602), .Z(n51604) );
  INAND2HSV2 U55040 ( .A1(n52169), .B1(n52047), .ZN(n51681) );
  CLKNAND2HSV1 U55041 ( .A1(n52048), .A2(n47571), .ZN(n51679) );
  CLKNAND2HSV1 U55042 ( .A1(n25835), .A2(n51726), .ZN(n51677) );
  CLKNAND2HSV1 U55043 ( .A1(n51798), .A2(n51608), .ZN(n51673) );
  NOR2HSV1 U55044 ( .A1(n52170), .A2(n51607), .ZN(n51671) );
  CLKNAND2HSV0 U55045 ( .A1(n51799), .A2(n52172), .ZN(n51669) );
  NOR2HSV1 U55046 ( .A1(n52171), .A2(n44045), .ZN(n51667) );
  NAND2HSV0 U55047 ( .A1(n59775), .A2(n52052), .ZN(n51664) );
  NAND2HSV0 U55048 ( .A1(n59506), .A2(n59777), .ZN(n51659) );
  CLKNAND2HSV0 U55049 ( .A1(n52417), .A2(n51896), .ZN(n51657) );
  BUFHSV2 U55050 ( .I(n51965), .Z(n52927) );
  CLKNAND2HSV1 U55051 ( .A1(n52927), .A2(n51933), .ZN(n51654) );
  NAND2HSV0 U55052 ( .A1(n51609), .A2(n52895), .ZN(n51652) );
  NAND2HSV0 U55053 ( .A1(n51610), .A2(n52901), .ZN(n51650) );
  CLKNAND2HSV1 U55054 ( .A1(n51920), .A2(n52859), .ZN(n51738) );
  NAND2HSV0 U55055 ( .A1(n59976), .A2(n52063), .ZN(n51613) );
  NAND2HSV0 U55056 ( .A1(\pe2/aot [2]), .A2(n38792), .ZN(n51612) );
  XOR2HSV0 U55057 ( .A1(n51613), .A2(n51612), .Z(n51618) );
  NAND2HSV0 U55058 ( .A1(n59783), .A2(n44197), .ZN(n51616) );
  NAND2HSV0 U55059 ( .A1(\pe2/aot [20]), .A2(n51614), .ZN(n51615) );
  XOR2HSV0 U55060 ( .A1(n51616), .A2(n51615), .Z(n51617) );
  XOR2HSV0 U55061 ( .A1(n51618), .A2(n51617), .Z(n51629) );
  NAND2HSV0 U55062 ( .A1(n51824), .A2(\pe2/bq[17] ), .ZN(n51620) );
  NAND2HSV0 U55063 ( .A1(n59792), .A2(\pe2/bq[18] ), .ZN(n51619) );
  XOR2HSV0 U55064 ( .A1(n51620), .A2(n51619), .Z(n51627) );
  NOR2HSV0 U55065 ( .A1(n51622), .A2(n51621), .ZN(n51625) );
  AOI22HSV0 U55066 ( .A1(n52070), .A2(n52866), .B1(\pe2/aot [12]), .B2(n51623), 
        .ZN(n51624) );
  NOR2HSV2 U55067 ( .A1(n51625), .A2(n51624), .ZN(n51626) );
  XNOR2HSV1 U55068 ( .A1(n51627), .A2(n51626), .ZN(n51628) );
  XNOR2HSV1 U55069 ( .A1(n51629), .A2(n51628), .ZN(n51647) );
  NAND2HSV0 U55070 ( .A1(n59973), .A2(n51897), .ZN(n51631) );
  NAND2HSV0 U55071 ( .A1(n51460), .A2(n51900), .ZN(n51630) );
  XOR2HSV0 U55072 ( .A1(n51631), .A2(n51630), .Z(n51635) );
  NAND2HSV0 U55073 ( .A1(n59633), .A2(\pe2/bq[14] ), .ZN(n51633) );
  NAND2HSV0 U55074 ( .A1(n52056), .A2(\pe2/bq[16] ), .ZN(n51632) );
  XOR2HSV0 U55075 ( .A1(n51633), .A2(n51632), .Z(n51634) );
  XOR2HSV0 U55076 ( .A1(n51635), .A2(n51634), .Z(n51645) );
  NAND2HSV0 U55077 ( .A1(n51636), .A2(n49619), .ZN(n51638) );
  NAND2HSV0 U55078 ( .A1(\pe2/aot [19]), .A2(n51919), .ZN(n51637) );
  XOR2HSV0 U55079 ( .A1(n51638), .A2(n51637), .Z(n51643) );
  NAND2HSV0 U55080 ( .A1(n59975), .A2(n53223), .ZN(n51641) );
  NAND2HSV0 U55081 ( .A1(n51639), .A2(\pe2/bq[3] ), .ZN(n51640) );
  XOR2HSV0 U55082 ( .A1(n51641), .A2(n51640), .Z(n51642) );
  XOR2HSV0 U55083 ( .A1(n51643), .A2(n51642), .Z(n51644) );
  XOR2HSV0 U55084 ( .A1(n51645), .A2(n51644), .Z(n51646) );
  XOR3HSV2 U55085 ( .A1(n51648), .A2(n51647), .A3(n51646), .Z(n51649) );
  XNOR2HSV1 U55086 ( .A1(n51650), .A2(n51649), .ZN(n51651) );
  XNOR2HSV1 U55087 ( .A1(n51652), .A2(n51651), .ZN(n51653) );
  XNOR2HSV1 U55088 ( .A1(n51654), .A2(n51653), .ZN(n51656) );
  NOR2HSV0 U55089 ( .A1(n45071), .A2(n50908), .ZN(n51655) );
  XOR3HSV2 U55090 ( .A1(n51657), .A2(n51656), .A3(n51655), .Z(n51658) );
  XOR2HSV0 U55091 ( .A1(n51659), .A2(n51658), .Z(n51662) );
  CLKNAND2HSV1 U55092 ( .A1(n59769), .A2(n51895), .ZN(n51661) );
  CLKNAND2HSV1 U55093 ( .A1(n52138), .A2(n59371), .ZN(n51660) );
  XOR3HSV2 U55094 ( .A1(n51662), .A2(n51661), .A3(n51660), .Z(n51663) );
  XNOR2HSV1 U55095 ( .A1(n51664), .A2(n51663), .ZN(n51666) );
  CLKNAND2HSV1 U55096 ( .A1(n51782), .A2(n49493), .ZN(n51665) );
  XOR3HSV2 U55097 ( .A1(n51667), .A2(n51666), .A3(n51665), .Z(n51668) );
  XOR2HSV0 U55098 ( .A1(n51669), .A2(n51668), .Z(n51670) );
  XNOR2HSV1 U55099 ( .A1(n51671), .A2(n51670), .ZN(n51672) );
  XNOR2HSV1 U55100 ( .A1(n51673), .A2(n51672), .ZN(n51675) );
  CLKNAND2HSV1 U55101 ( .A1(n51792), .A2(n52051), .ZN(n51674) );
  XNOR2HSV1 U55102 ( .A1(n51675), .A2(n51674), .ZN(n51676) );
  XOR2HSV0 U55103 ( .A1(n51677), .A2(n51676), .Z(n51678) );
  XOR2HSV0 U55104 ( .A1(n51679), .A2(n51678), .Z(n51680) );
  XOR2HSV0 U55105 ( .A1(n51681), .A2(n51680), .Z(n51683) );
  XNOR2HSV4 U55106 ( .A1(n51683), .A2(n51682), .ZN(n51685) );
  CLKNAND2HSV0 U55107 ( .A1(n59790), .A2(n51939), .ZN(n51723) );
  NAND2HSV0 U55108 ( .A1(n59522), .A2(n51686), .ZN(n51721) );
  NOR2HSV0 U55109 ( .A1(n52171), .A2(n53032), .ZN(n51719) );
  NAND2HSV0 U55110 ( .A1(n51485), .A2(n51932), .ZN(n51716) );
  CLKNAND2HSV0 U55111 ( .A1(n52534), .A2(n51688), .ZN(n51714) );
  NAND2HSV0 U55112 ( .A1(n59976), .A2(n52484), .ZN(n51690) );
  NAND2HSV0 U55113 ( .A1(n59768), .A2(n51897), .ZN(n51689) );
  XOR2HSV0 U55114 ( .A1(n51690), .A2(n51689), .Z(n51694) );
  NAND2HSV0 U55115 ( .A1(n59977), .A2(n51803), .ZN(n51692) );
  NAND2HSV0 U55116 ( .A1(n52456), .A2(n53223), .ZN(n51691) );
  XOR2HSV0 U55117 ( .A1(n51692), .A2(n51691), .Z(n51693) );
  XOR2HSV0 U55118 ( .A1(n51694), .A2(n51693), .Z(n51702) );
  NAND2HSV0 U55119 ( .A1(\pe2/aot [8]), .A2(\pe2/bq[6] ), .ZN(n51696) );
  NAND2HSV0 U55120 ( .A1(n51824), .A2(n52448), .ZN(n51695) );
  XOR2HSV0 U55121 ( .A1(n51696), .A2(n51695), .Z(n51700) );
  CLKNAND2HSV0 U55122 ( .A1(n52056), .A2(n52322), .ZN(n51698) );
  NAND2HSV0 U55123 ( .A1(\pe2/aot [7]), .A2(n51832), .ZN(n51697) );
  XOR2HSV0 U55124 ( .A1(n51698), .A2(n51697), .Z(n51699) );
  XOR2HSV0 U55125 ( .A1(n51700), .A2(n51699), .Z(n51701) );
  XOR2HSV0 U55126 ( .A1(n51702), .A2(n51701), .Z(n51712) );
  NAND2HSV2 U55127 ( .A1(n52966), .A2(n51614), .ZN(n51984) );
  NAND2HSV0 U55128 ( .A1(n52867), .A2(n51900), .ZN(n51705) );
  XNOR2HSV1 U55129 ( .A1(n51706), .A2(n51705), .ZN(n51710) );
  NOR2HSV0 U55130 ( .A1(n52095), .A2(n49628), .ZN(n51708) );
  NAND2HSV0 U55131 ( .A1(\pe2/aot [2]), .A2(n51733), .ZN(n51707) );
  XOR2HSV0 U55132 ( .A1(n51708), .A2(n51707), .Z(n51709) );
  XOR2HSV0 U55133 ( .A1(n51710), .A2(n51709), .Z(n51711) );
  XNOR2HSV1 U55134 ( .A1(n51712), .A2(n51711), .ZN(n51713) );
  XNOR2HSV1 U55135 ( .A1(n51714), .A2(n51713), .ZN(n51715) );
  XNOR2HSV1 U55136 ( .A1(n51716), .A2(n51715), .ZN(n51718) );
  CLKNAND2HSV0 U55137 ( .A1(n51868), .A2(n52855), .ZN(n51717) );
  XOR3HSV2 U55138 ( .A1(n51719), .A2(n51718), .A3(n51717), .Z(n51720) );
  XOR2HSV0 U55139 ( .A1(n51721), .A2(n51720), .Z(n51722) );
  XOR2HSV0 U55140 ( .A1(n51723), .A2(n51722), .Z(n51725) );
  CLKNAND2HSV1 U55141 ( .A1(n25828), .A2(\pe2/got [8]), .ZN(n51724) );
  INHSV2 U55142 ( .I(n51727), .ZN(n53093) );
  CLKNAND2HSV1 U55143 ( .A1(n51728), .A2(n52172), .ZN(n51791) );
  NOR2HSV1 U55144 ( .A1(n52170), .A2(n49656), .ZN(n51789) );
  CLKNAND2HSV1 U55145 ( .A1(n51799), .A2(\pe2/got [10]), .ZN(n51787) );
  NOR2HSV1 U55146 ( .A1(n52921), .A2(n44188), .ZN(n51785) );
  NAND2HSV0 U55147 ( .A1(n59775), .A2(n51895), .ZN(n51781) );
  NAND2HSV0 U55148 ( .A1(n59984), .A2(n52173), .ZN(n51776) );
  CLKNAND2HSV1 U55149 ( .A1(n52926), .A2(\pe2/got [2]), .ZN(n51774) );
  CLKNAND2HSV1 U55150 ( .A1(n59634), .A2(n52896), .ZN(n51771) );
  NAND2HSV0 U55151 ( .A1(n52056), .A2(\pe2/bq[14] ), .ZN(n51731) );
  NAND2HSV0 U55152 ( .A1(\pe2/aot [6]), .A2(n51729), .ZN(n51730) );
  XOR2HSV0 U55153 ( .A1(n51731), .A2(n51730), .Z(n51752) );
  NAND2HSV0 U55154 ( .A1(n59792), .A2(n51732), .ZN(n51735) );
  NAND2HSV0 U55155 ( .A1(n59633), .A2(n51733), .ZN(n51734) );
  XOR2HSV0 U55156 ( .A1(n51735), .A2(n51734), .Z(n51742) );
  NOR2HSV0 U55157 ( .A1(n45165), .A2(n51842), .ZN(n51740) );
  NOR2HSV0 U55158 ( .A1(n51736), .A2(n49529), .ZN(n51739) );
  OAI22HSV2 U55159 ( .A1(n51740), .A2(n51739), .B1(n51738), .B2(n51737), .ZN(
        n51741) );
  XNOR2HSV1 U55160 ( .A1(n51742), .A2(n51741), .ZN(n51751) );
  NAND2HSV0 U55161 ( .A1(n52966), .A2(\pe2/bq[6] ), .ZN(n51745) );
  NAND2HSV0 U55162 ( .A1(n51743), .A2(\pe2/bq[3] ), .ZN(n51744) );
  XOR2HSV0 U55163 ( .A1(n51745), .A2(n51744), .Z(n51749) );
  NAND2HSV0 U55164 ( .A1(n59974), .A2(n51803), .ZN(n51747) );
  NAND2HSV0 U55165 ( .A1(n59976), .A2(n53223), .ZN(n51746) );
  XOR2HSV0 U55166 ( .A1(n51747), .A2(n51746), .Z(n51748) );
  XOR2HSV0 U55167 ( .A1(n51749), .A2(n51748), .Z(n51750) );
  XOR3HSV2 U55168 ( .A1(n51752), .A2(n51751), .A3(n51750), .Z(n51769) );
  NAND2HSV0 U55169 ( .A1(n52951), .A2(\pe2/bq[11] ), .ZN(n51754) );
  NAND2HSV0 U55170 ( .A1(\pe2/aot [9]), .A2(n52063), .ZN(n51753) );
  XOR2HSV0 U55171 ( .A1(n51754), .A2(n51753), .Z(n51758) );
  NAND2HSV0 U55172 ( .A1(\pe2/aot [2]), .A2(\pe2/bq[17] ), .ZN(n51756) );
  NAND2HSV0 U55173 ( .A1(n59783), .A2(n52988), .ZN(n51755) );
  XOR2HSV0 U55174 ( .A1(n51756), .A2(n51755), .Z(n51757) );
  XOR2HSV0 U55175 ( .A1(n51758), .A2(n51757), .Z(n51767) );
  NAND2HSV0 U55176 ( .A1(n51759), .A2(n51919), .ZN(n51761) );
  NAND2HSV0 U55177 ( .A1(n51824), .A2(n49619), .ZN(n51760) );
  XOR2HSV0 U55178 ( .A1(n51761), .A2(n51760), .Z(n51765) );
  NOR2HSV0 U55179 ( .A1(n52103), .A2(n50920), .ZN(n51763) );
  NAND2HSV0 U55180 ( .A1(\pe2/aot [10]), .A2(n52193), .ZN(n51762) );
  XOR2HSV0 U55181 ( .A1(n51763), .A2(n51762), .Z(n51764) );
  XOR2HSV0 U55182 ( .A1(n51765), .A2(n51764), .Z(n51766) );
  XOR2HSV0 U55183 ( .A1(n51767), .A2(n51766), .Z(n51768) );
  XNOR2HSV1 U55184 ( .A1(n51769), .A2(n51768), .ZN(n51770) );
  XNOR2HSV1 U55185 ( .A1(n51771), .A2(n51770), .ZN(n51773) );
  NOR2HSV0 U55186 ( .A1(n53065), .A2(n53032), .ZN(n51772) );
  XOR3HSV2 U55187 ( .A1(n51774), .A2(n51773), .A3(n51772), .Z(n51775) );
  XOR2HSV0 U55188 ( .A1(n51776), .A2(n51775), .Z(n51779) );
  CLKNAND2HSV1 U55189 ( .A1(n59769), .A2(n52175), .ZN(n51778) );
  CLKNAND2HSV1 U55190 ( .A1(n52138), .A2(n51939), .ZN(n51777) );
  XOR3HSV2 U55191 ( .A1(n51779), .A2(n51778), .A3(n51777), .Z(n51780) );
  XNOR2HSV1 U55192 ( .A1(n51781), .A2(n51780), .ZN(n51784) );
  CLKNAND2HSV1 U55193 ( .A1(n51782), .A2(n52052), .ZN(n51783) );
  XOR3HSV2 U55194 ( .A1(n51785), .A2(n51784), .A3(n51783), .Z(n51786) );
  XOR2HSV0 U55195 ( .A1(n51787), .A2(n51786), .Z(n51788) );
  XNOR2HSV1 U55196 ( .A1(n51789), .A2(n51788), .ZN(n51790) );
  XNOR2HSV1 U55197 ( .A1(n51791), .A2(n51790), .ZN(n51794) );
  CLKNAND2HSV1 U55198 ( .A1(n51792), .A2(n59375), .ZN(n51793) );
  CLKNHSV0 U55199 ( .I(n59983), .ZN(n51795) );
  INAND2HSV2 U55200 ( .A1(n51795), .B1(n53093), .ZN(n51886) );
  CLKNAND2HSV1 U55201 ( .A1(n51120), .A2(n51796), .ZN(n51884) );
  CLKNAND2HSV1 U55202 ( .A1(n52918), .A2(n52051), .ZN(n51882) );
  CLKNAND2HSV1 U55203 ( .A1(n51798), .A2(n52418), .ZN(n51877) );
  NOR2HSV1 U55204 ( .A1(n52170), .A2(n47555), .ZN(n51875) );
  CLKNAND2HSV0 U55205 ( .A1(n51799), .A2(n49493), .ZN(n51873) );
  NOR2HSV0 U55206 ( .A1(n52171), .A2(n51800), .ZN(n51871) );
  NAND2HSV0 U55207 ( .A1(n51485), .A2(\pe2/got [8]), .ZN(n51867) );
  NAND2HSV0 U55208 ( .A1(n51801), .A2(n59778), .ZN(n51860) );
  CLKNAND2HSV0 U55209 ( .A1(n52926), .A2(n51933), .ZN(n51858) );
  NAND2HSV0 U55210 ( .A1(n51965), .A2(\pe2/got [2]), .ZN(n51855) );
  NAND2HSV0 U55211 ( .A1(n51802), .A2(n52896), .ZN(n51853) );
  NAND2HSV0 U55212 ( .A1(n59358), .A2(n51803), .ZN(n51971) );
  NOR2HSV0 U55213 ( .A1(n51971), .A2(n51804), .ZN(n51807) );
  AOI22HSV0 U55214 ( .A1(n59358), .A2(n51805), .B1(n59973), .B2(n52309), .ZN(
        n51806) );
  NOR2HSV2 U55215 ( .A1(n51807), .A2(n51806), .ZN(n51812) );
  NAND2HSV0 U55216 ( .A1(n52951), .A2(\pe2/bq[14] ), .ZN(n51975) );
  NOR2HSV0 U55217 ( .A1(n51975), .A2(n51808), .ZN(n51810) );
  AOI22HSV0 U55218 ( .A1(\pe2/aot [8]), .A2(n52438), .B1(\pe2/bq[14] ), .B2(
        n52456), .ZN(n51809) );
  NOR2HSV1 U55219 ( .A1(n51810), .A2(n51809), .ZN(n51811) );
  XNOR2HSV1 U55220 ( .A1(n51812), .A2(n51811), .ZN(n51821) );
  NAND2HSV0 U55221 ( .A1(n52056), .A2(n52337), .ZN(n51816) );
  NOR2HSV0 U55222 ( .A1(n51814), .A2(n51813), .ZN(n51815) );
  AOI21HSV2 U55223 ( .A1(n51817), .A2(n51816), .B(n51815), .ZN(n51819) );
  NAND2HSV0 U55224 ( .A1(n51920), .A2(\pe2/bq[6] ), .ZN(n51818) );
  XNOR2HSV1 U55225 ( .A1(n51819), .A2(n51818), .ZN(n51820) );
  XNOR2HSV1 U55226 ( .A1(n51821), .A2(n51820), .ZN(n51831) );
  NAND2HSV0 U55227 ( .A1(\pe2/aot [9]), .A2(n51900), .ZN(n51823) );
  NAND2HSV0 U55228 ( .A1(\pe2/aot [17]), .A2(n52905), .ZN(n51822) );
  XOR2HSV0 U55229 ( .A1(n51823), .A2(n51822), .Z(n51829) );
  NAND2HSV0 U55230 ( .A1(n51824), .A2(\pe2/bq[16] ), .ZN(n51827) );
  NAND2HSV0 U55231 ( .A1(n53005), .A2(n51825), .ZN(n51826) );
  XOR2HSV0 U55232 ( .A1(n51827), .A2(n51826), .Z(n51828) );
  XOR2HSV0 U55233 ( .A1(n51829), .A2(n51828), .Z(n51830) );
  XOR2HSV0 U55234 ( .A1(n51831), .A2(n51830), .Z(n51851) );
  NAND2HSV0 U55235 ( .A1(n51921), .A2(n51832), .ZN(n51834) );
  NAND2HSV0 U55236 ( .A1(\pe2/aot [2]), .A2(n52988), .ZN(n51833) );
  XOR2HSV0 U55237 ( .A1(n51834), .A2(n51833), .Z(n51838) );
  NOR2HSV0 U55238 ( .A1(n52431), .A2(n49515), .ZN(n51836) );
  NAND2HSV0 U55239 ( .A1(n59976), .A2(n52193), .ZN(n51835) );
  XOR2HSV0 U55240 ( .A1(n51836), .A2(n51835), .Z(n51837) );
  XNOR2HSV1 U55241 ( .A1(n51838), .A2(n51837), .ZN(n51849) );
  NAND2HSV0 U55242 ( .A1(n59792), .A2(n44074), .ZN(n51841) );
  NAND2HSV0 U55243 ( .A1(n59633), .A2(n51839), .ZN(n51840) );
  XOR2HSV0 U55244 ( .A1(n51841), .A2(n51840), .Z(n51847) );
  NOR2HSV0 U55245 ( .A1(n47503), .A2(n51842), .ZN(n51845) );
  NOR2HSV0 U55246 ( .A1(n52095), .A2(n52429), .ZN(n51844) );
  OAI22HSV0 U55247 ( .A1(n51845), .A2(n51844), .B1(n51843), .B2(n51967), .ZN(
        n51846) );
  XNOR2HSV1 U55248 ( .A1(n51847), .A2(n51846), .ZN(n51848) );
  XNOR2HSV1 U55249 ( .A1(n51849), .A2(n51848), .ZN(n51850) );
  XNOR2HSV1 U55250 ( .A1(n51851), .A2(n51850), .ZN(n51852) );
  XNOR2HSV1 U55251 ( .A1(n51853), .A2(n51852), .ZN(n51854) );
  XNOR2HSV1 U55252 ( .A1(n51855), .A2(n51854), .ZN(n51857) );
  NOR2HSV0 U55253 ( .A1(n53065), .A2(n50909), .ZN(n51856) );
  XOR3HSV2 U55254 ( .A1(n51858), .A2(n51857), .A3(n51856), .Z(n51859) );
  XOR2HSV0 U55255 ( .A1(n51860), .A2(n51859), .Z(n51865) );
  NAND2HSV2 U55256 ( .A1(n51861), .A2(n59777), .ZN(n51864) );
  CLKNAND2HSV0 U55257 ( .A1(n51862), .A2(n51895), .ZN(n51863) );
  XOR3HSV2 U55258 ( .A1(n51865), .A2(n51864), .A3(n51863), .Z(n51866) );
  XNOR2HSV1 U55259 ( .A1(n51867), .A2(n51866), .ZN(n51870) );
  CLKNAND2HSV0 U55260 ( .A1(n51868), .A2(\pe2/got [10]), .ZN(n51869) );
  XOR3HSV2 U55261 ( .A1(n51871), .A2(n51870), .A3(n51869), .Z(n51872) );
  XOR2HSV0 U55262 ( .A1(n51873), .A2(n51872), .Z(n51874) );
  XNOR2HSV1 U55263 ( .A1(n51875), .A2(n51874), .ZN(n51876) );
  XNOR2HSV1 U55264 ( .A1(n51877), .A2(n51876), .ZN(n51880) );
  CLKNAND2HSV1 U55265 ( .A1(n51878), .A2(n59354), .ZN(n51879) );
  XNOR2HSV1 U55266 ( .A1(n51880), .A2(n51879), .ZN(n51881) );
  XOR2HSV0 U55267 ( .A1(n51882), .A2(n51881), .Z(n51883) );
  XOR2HSV0 U55268 ( .A1(n51884), .A2(n51883), .Z(n51885) );
  XOR2HSV0 U55269 ( .A1(n51886), .A2(n51885), .Z(n51888) );
  NAND2HSV2 U55270 ( .A1(n25709), .A2(n44712), .ZN(n51887) );
  XNOR2HSV4 U55271 ( .A1(n51888), .A2(n51887), .ZN(n51891) );
  CLKNAND2HSV0 U55272 ( .A1(n51889), .A2(n51961), .ZN(n51890) );
  XNOR2HSV4 U55273 ( .A1(n51891), .A2(n51890), .ZN(\pe2/poht [13]) );
  CLKNAND2HSV1 U55274 ( .A1(n52414), .A2(n52418), .ZN(n51957) );
  CLKNAND2HSV0 U55275 ( .A1(n59475), .A2(\pe2/got [12]), .ZN(n51955) );
  CLKNAND2HSV1 U55276 ( .A1(n52918), .A2(n51892), .ZN(n51953) );
  CLKNAND2HSV1 U55277 ( .A1(n51893), .A2(\pe2/got [9]), .ZN(n51948) );
  NOR2HSV0 U55278 ( .A1(n51894), .A2(n44188), .ZN(n51946) );
  NAND2HSV0 U55279 ( .A1(n59522), .A2(n51895), .ZN(n51944) );
  NOR2HSV0 U55280 ( .A1(n52171), .A2(n50908), .ZN(n51942) );
  CLKNAND2HSV1 U55281 ( .A1(n51485), .A2(n51896), .ZN(n51938) );
  NAND2HSV0 U55282 ( .A1(n52896), .A2(n52814), .ZN(n51931) );
  NAND2HSV0 U55283 ( .A1(n59976), .A2(n51897), .ZN(n51899) );
  NAND2HSV0 U55284 ( .A1(\pe2/aot [9]), .A2(n51832), .ZN(n51898) );
  XOR2HSV0 U55285 ( .A1(n51899), .A2(n51898), .Z(n51904) );
  NAND2HSV0 U55286 ( .A1(n51824), .A2(n52438), .ZN(n51902) );
  NAND2HSV0 U55287 ( .A1(n29736), .A2(n51900), .ZN(n51901) );
  XOR2HSV0 U55288 ( .A1(n51902), .A2(n51901), .Z(n51903) );
  XOR2HSV0 U55289 ( .A1(n51904), .A2(n51903), .Z(n51912) );
  NAND2HSV0 U55290 ( .A1(\pe2/aot [15]), .A2(\pe2/bq[1] ), .ZN(n51906) );
  NAND2HSV0 U55291 ( .A1(\pe2/aot [2]), .A2(\pe2/bq[14] ), .ZN(n51905) );
  XOR2HSV0 U55292 ( .A1(n51906), .A2(n51905), .Z(n51910) );
  CLKNAND2HSV1 U55293 ( .A1(n51636), .A2(n52063), .ZN(n51908) );
  NAND2HSV0 U55294 ( .A1(n52951), .A2(n53223), .ZN(n51907) );
  XOR2HSV0 U55295 ( .A1(n51908), .A2(n51907), .Z(n51909) );
  XOR2HSV0 U55296 ( .A1(n51910), .A2(n51909), .Z(n51911) );
  XOR2HSV0 U55297 ( .A1(n51912), .A2(n51911), .Z(n51929) );
  NAND2HSV0 U55298 ( .A1(n53005), .A2(n51803), .ZN(n51914) );
  NAND2HSV0 U55299 ( .A1(n59783), .A2(\pe2/bq[15] ), .ZN(n51913) );
  XOR2HSV0 U55300 ( .A1(n51914), .A2(n51913), .Z(n51918) );
  NAND2HSV0 U55301 ( .A1(\pe2/aot [7]), .A2(n51623), .ZN(n51916) );
  NAND2HSV0 U55302 ( .A1(n51460), .A2(\pe2/bq[6] ), .ZN(n51915) );
  XOR2HSV0 U55303 ( .A1(n51916), .A2(n51915), .Z(n51917) );
  XOR2HSV0 U55304 ( .A1(n51918), .A2(n51917), .Z(n51927) );
  NAND2HSV0 U55305 ( .A1(n51920), .A2(n51919), .ZN(n51923) );
  NAND2HSV0 U55306 ( .A1(n51921), .A2(\pe2/bq[3] ), .ZN(n51922) );
  XOR2HSV0 U55307 ( .A1(n51923), .A2(n51922), .Z(n51925) );
  XNOR2HSV1 U55308 ( .A1(n51925), .A2(n51924), .ZN(n51926) );
  XNOR2HSV1 U55309 ( .A1(n51927), .A2(n51926), .ZN(n51928) );
  XNOR2HSV1 U55310 ( .A1(n51929), .A2(n51928), .ZN(n51930) );
  XNOR2HSV1 U55311 ( .A1(n51931), .A2(n51930), .ZN(n51936) );
  NAND2HSV0 U55312 ( .A1(n59769), .A2(n51932), .ZN(n51935) );
  CLKNAND2HSV0 U55313 ( .A1(n51862), .A2(n51933), .ZN(n51934) );
  XOR3HSV2 U55314 ( .A1(n51936), .A2(n51935), .A3(n51934), .Z(n51937) );
  XNOR2HSV1 U55315 ( .A1(n51938), .A2(n51937), .ZN(n51941) );
  CLKNAND2HSV1 U55316 ( .A1(n53078), .A2(n51939), .ZN(n51940) );
  XOR3HSV2 U55317 ( .A1(n51942), .A2(n51941), .A3(n51940), .Z(n51943) );
  XOR2HSV0 U55318 ( .A1(n51944), .A2(n51943), .Z(n51945) );
  XNOR2HSV1 U55319 ( .A1(n51946), .A2(n51945), .ZN(n51947) );
  XNOR2HSV1 U55320 ( .A1(n51948), .A2(n51947), .ZN(n51951) );
  CLKNAND2HSV0 U55321 ( .A1(n51949), .A2(\pe2/got [10]), .ZN(n51950) );
  XNOR2HSV1 U55322 ( .A1(n51951), .A2(n51950), .ZN(n51952) );
  XOR2HSV0 U55323 ( .A1(n51953), .A2(n51952), .Z(n51954) );
  XOR2HSV0 U55324 ( .A1(n51955), .A2(n51954), .Z(n51956) );
  XNOR2HSV4 U55325 ( .A1(n51960), .A2(n51959), .ZN(n51963) );
  CLKNAND2HSV0 U55326 ( .A1(n45289), .A2(n51961), .ZN(n51962) );
  XNOR2HSV4 U55327 ( .A1(n51963), .A2(n51962), .ZN(\pe2/poht [17]) );
  CLKNAND2HSV1 U55328 ( .A1(n52047), .A2(n52533), .ZN(n52041) );
  CLKNAND2HSV1 U55329 ( .A1(n53087), .A2(n51964), .ZN(n52037) );
  NOR2HSV1 U55330 ( .A1(n52170), .A2(n47498), .ZN(n52035) );
  CLKNAND2HSV0 U55331 ( .A1(n44968), .A2(n53055), .ZN(n52033) );
  NOR2HSV2 U55332 ( .A1(n52921), .A2(n49656), .ZN(n52031) );
  CLKNAND2HSV0 U55333 ( .A1(n52923), .A2(\pe2/got [10]), .ZN(n52028) );
  NAND2HSV0 U55334 ( .A1(n52174), .A2(n59506), .ZN(n52023) );
  CLKNAND2HSV0 U55335 ( .A1(n52417), .A2(n53038), .ZN(n52021) );
  NAND2HSV0 U55336 ( .A1(n51965), .A2(n51896), .ZN(n52017) );
  NAND2HSV0 U55337 ( .A1(n51609), .A2(\pe2/got [3]), .ZN(n52015) );
  NAND2HSV0 U55338 ( .A1(n59761), .A2(n51932), .ZN(n52013) );
  NAND2HSV0 U55339 ( .A1(n59767), .A2(n51966), .ZN(n52011) );
  NOR2HSV0 U55340 ( .A1(n38946), .A2(n51842), .ZN(n51969) );
  OAI22HSV0 U55341 ( .A1(n51970), .A2(n51969), .B1(n51968), .B2(n51967), .ZN(
        n51974) );
  XOR2HSV0 U55342 ( .A1(n51972), .A2(n51971), .Z(n51973) );
  XOR3HSV1 U55343 ( .A1(n51975), .A2(n51974), .A3(n51973), .Z(n52009) );
  NAND2HSV0 U55344 ( .A1(n52294), .A2(\pe2/bq[3] ), .ZN(n51977) );
  NAND2HSV0 U55345 ( .A1(n52456), .A2(n38803), .ZN(n51976) );
  XOR2HSV0 U55346 ( .A1(n51977), .A2(n51976), .Z(n51981) );
  NAND2HSV0 U55347 ( .A1(\pe2/bq[17] ), .A2(n29736), .ZN(n51979) );
  NAND2HSV0 U55348 ( .A1(\pe2/aot [10]), .A2(n51733), .ZN(n51978) );
  XOR2HSV0 U55349 ( .A1(n51979), .A2(n51978), .Z(n51980) );
  XOR2HSV0 U55350 ( .A1(n51981), .A2(n51980), .Z(n51990) );
  NOR2HSV0 U55351 ( .A1(n51538), .A2(n52429), .ZN(n51983) );
  NAND2HSV0 U55352 ( .A1(n52993), .A2(n52988), .ZN(n51982) );
  XOR2HSV0 U55353 ( .A1(n51983), .A2(n51982), .Z(n51988) );
  NOR2HSV0 U55354 ( .A1(n38822), .A2(n47511), .ZN(n51986) );
  OAI22HSV2 U55355 ( .A1(n52204), .A2(n51986), .B1(n51985), .B2(n51984), .ZN(
        n51987) );
  XNOR2HSV1 U55356 ( .A1(n51988), .A2(n51987), .ZN(n51989) );
  XNOR2HSV1 U55357 ( .A1(n51990), .A2(n51989), .ZN(n52008) );
  NAND2HSV0 U55358 ( .A1(n59768), .A2(n52962), .ZN(n51992) );
  NAND2HSV0 U55359 ( .A1(n39019), .A2(n52073), .ZN(n51991) );
  XOR2HSV0 U55360 ( .A1(n51992), .A2(n51991), .Z(n51996) );
  CLKNAND2HSV0 U55361 ( .A1(\pe2/aot [20]), .A2(n51805), .ZN(n51994) );
  NAND2HSV0 U55362 ( .A1(\pe2/aot [7]), .A2(n43956), .ZN(n51993) );
  XOR2HSV0 U55363 ( .A1(n51994), .A2(n51993), .Z(n51995) );
  XOR2HSV0 U55364 ( .A1(n51996), .A2(n51995), .Z(n52006) );
  NAND2HSV0 U55365 ( .A1(n53005), .A2(n51997), .ZN(n52000) );
  NAND2HSV0 U55366 ( .A1(\pe2/aot [2]), .A2(n51998), .ZN(n51999) );
  XOR2HSV0 U55367 ( .A1(n52000), .A2(n51999), .Z(n52004) );
  NAND2HSV0 U55368 ( .A1(n52070), .A2(n52859), .ZN(n52002) );
  NAND2HSV0 U55369 ( .A1(n59636), .A2(n53223), .ZN(n52001) );
  XOR2HSV0 U55370 ( .A1(n52002), .A2(n52001), .Z(n52003) );
  XOR2HSV0 U55371 ( .A1(n52004), .A2(n52003), .Z(n52005) );
  XOR2HSV0 U55372 ( .A1(n52006), .A2(n52005), .Z(n52007) );
  XOR3HSV2 U55373 ( .A1(n52009), .A2(n52008), .A3(n52007), .Z(n52010) );
  XNOR2HSV1 U55374 ( .A1(n52011), .A2(n52010), .ZN(n52012) );
  XOR2HSV0 U55375 ( .A1(n52013), .A2(n52012), .Z(n52014) );
  XNOR2HSV1 U55376 ( .A1(n52015), .A2(n52014), .ZN(n52016) );
  XNOR2HSV1 U55377 ( .A1(n52017), .A2(n52016), .ZN(n52020) );
  NOR2HSV0 U55378 ( .A1(n53065), .A2(n52018), .ZN(n52019) );
  XOR3HSV2 U55379 ( .A1(n52021), .A2(n52020), .A3(n52019), .Z(n52022) );
  XOR2HSV0 U55380 ( .A1(n52023), .A2(n52022), .Z(n52026) );
  CLKNAND2HSV0 U55381 ( .A1(n52532), .A2(n59371), .ZN(n52025) );
  NAND2HSV0 U55382 ( .A1(n52534), .A2(n52052), .ZN(n52024) );
  XOR3HSV2 U55383 ( .A1(n52026), .A2(n52025), .A3(n52024), .Z(n52027) );
  XNOR2HSV1 U55384 ( .A1(n52028), .A2(n52027), .ZN(n52030) );
  CLKNAND2HSV0 U55385 ( .A1(n53078), .A2(n52172), .ZN(n52029) );
  XOR3HSV2 U55386 ( .A1(n52031), .A2(n52030), .A3(n52029), .Z(n52032) );
  XOR2HSV0 U55387 ( .A1(n52033), .A2(n52032), .Z(n52034) );
  XNOR2HSV1 U55388 ( .A1(n52035), .A2(n52034), .ZN(n52036) );
  XNOR2HSV1 U55389 ( .A1(n52037), .A2(n52036), .ZN(n52039) );
  CLKNAND2HSV0 U55390 ( .A1(n52399), .A2(n51796), .ZN(n52038) );
  XNOR2HSV1 U55391 ( .A1(n52039), .A2(n52038), .ZN(n52040) );
  NAND2HSV2 U55392 ( .A1(n25709), .A2(n52042), .ZN(n52043) );
  XNOR2HSV4 U55393 ( .A1(n52044), .A2(n52043), .ZN(n52046) );
  INAND2HSV2 U55394 ( .A1(n38711), .B1(n53097), .ZN(n52045) );
  XNOR2HSV4 U55395 ( .A1(n52046), .A2(n52045), .ZN(\pe2/poht [11]) );
  CLKNAND2HSV1 U55396 ( .A1(n52047), .A2(\pe2/got [24]), .ZN(n52160) );
  CLKNAND2HSV1 U55397 ( .A1(n52048), .A2(n43924), .ZN(n52158) );
  CLKNAND2HSV0 U55398 ( .A1(n59927), .A2(n59685), .ZN(n52152) );
  NOR2HSV1 U55399 ( .A1(n52049), .A2(n47570), .ZN(n52150) );
  CLKNAND2HSV0 U55400 ( .A1(n44968), .A2(n52050), .ZN(n52148) );
  NOR2HSV0 U55401 ( .A1(n52921), .A2(n52526), .ZN(n52146) );
  NAND2HSV0 U55402 ( .A1(n52814), .A2(n52172), .ZN(n52137) );
  NAND2HSV0 U55403 ( .A1(n52417), .A2(\pe2/got [10]), .ZN(n52135) );
  NAND2HSV0 U55404 ( .A1(n52927), .A2(n52052), .ZN(n52132) );
  NAND2HSV0 U55405 ( .A1(n51609), .A2(\pe2/got [8]), .ZN(n52130) );
  NAND2HSV0 U55406 ( .A1(\pe2/got [6]), .A2(n52419), .ZN(n52128) );
  NAND2HSV0 U55407 ( .A1(n52176), .A2(n52175), .ZN(n52124) );
  NAND2HSV0 U55408 ( .A1(n39011), .A2(n51932), .ZN(n52117) );
  NAND2HSV0 U55409 ( .A1(n52053), .A2(n59767), .ZN(n52115) );
  NAND2HSV0 U55410 ( .A1(n52998), .A2(n51493), .ZN(n52055) );
  NAND2HSV0 U55411 ( .A1(n52184), .A2(n52179), .ZN(n52054) );
  XOR2HSV0 U55412 ( .A1(n52055), .A2(n52054), .Z(n52060) );
  NAND2HSV0 U55413 ( .A1(\pe2/aot [5]), .A2(n52299), .ZN(n52058) );
  NAND2HSV0 U55414 ( .A1(n52456), .A2(\pe2/bq[21] ), .ZN(n52057) );
  XOR2HSV0 U55415 ( .A1(n52058), .A2(n52057), .Z(n52059) );
  XOR2HSV0 U55416 ( .A1(n52060), .A2(n52059), .Z(n52069) );
  NAND2HSV0 U55417 ( .A1(n53005), .A2(n43956), .ZN(n52062) );
  NAND2HSV0 U55418 ( .A1(n59768), .A2(n52988), .ZN(n52061) );
  XOR2HSV0 U55419 ( .A1(n52062), .A2(n52061), .Z(n52067) );
  NAND2HSV0 U55420 ( .A1(n52951), .A2(n43961), .ZN(n52065) );
  NAND2HSV0 U55421 ( .A1(\pe2/aot [17]), .A2(n52063), .ZN(n52064) );
  XOR2HSV0 U55422 ( .A1(n52065), .A2(n52064), .Z(n52066) );
  XOR2HSV0 U55423 ( .A1(n52067), .A2(n52066), .Z(n52068) );
  XOR2HSV0 U55424 ( .A1(n52069), .A2(n52068), .Z(n52090) );
  NAND2HSV0 U55425 ( .A1(n52070), .A2(n51733), .ZN(n52072) );
  NAND2HSV0 U55426 ( .A1(n52974), .A2(n51614), .ZN(n52071) );
  XOR2HSV0 U55427 ( .A1(n52072), .A2(n52071), .Z(n52077) );
  NAND2HSV0 U55428 ( .A1(n51743), .A2(n52073), .ZN(n52075) );
  NAND2HSV0 U55429 ( .A1(n59975), .A2(\pe2/bq[14] ), .ZN(n52074) );
  XOR2HSV0 U55430 ( .A1(n52075), .A2(n52074), .Z(n52076) );
  XOR2HSV0 U55431 ( .A1(n52077), .A2(n52076), .Z(n52088) );
  NAND2HSV0 U55432 ( .A1(\pe2/aot [7]), .A2(n52965), .ZN(n52079) );
  NAND2HSV0 U55433 ( .A1(\pe2/aot [10]), .A2(\pe2/bq[17] ), .ZN(n52078) );
  XOR2HSV0 U55434 ( .A1(n52079), .A2(n52078), .Z(n52086) );
  NOR2HSV0 U55435 ( .A1(n44871), .A2(n51131), .ZN(n52084) );
  NOR2HSV0 U55436 ( .A1(n52080), .A2(n51567), .ZN(n52083) );
  OAI22HSV0 U55437 ( .A1(n52084), .A2(n52083), .B1(n52082), .B2(n52081), .ZN(
        n52085) );
  XNOR2HSV1 U55438 ( .A1(n52086), .A2(n52085), .ZN(n52087) );
  XNOR2HSV1 U55439 ( .A1(n52088), .A2(n52087), .ZN(n52089) );
  XNOR2HSV1 U55440 ( .A1(n52090), .A2(n52089), .ZN(n52113) );
  NOR2HSV0 U55441 ( .A1(n51538), .A2(n38687), .ZN(n53022) );
  XOR2HSV0 U55442 ( .A1(n53022), .A2(n52091), .Z(n52111) );
  OAI21HSV0 U55443 ( .A1(n48621), .A2(n47574), .B(n52092), .ZN(n52093) );
  OAI21HSV1 U55444 ( .A1(n52094), .A2(n52223), .B(n52093), .ZN(n52100) );
  INHSV2 U55445 ( .I(n52095), .ZN(n53016) );
  AOI22HSV0 U55446 ( .A1(n59976), .A2(\pe2/bq[16] ), .B1(\pe2/bq[26] ), .B2(
        n53016), .ZN(n52096) );
  AOI21HSV0 U55447 ( .A1(n52098), .A2(n52097), .B(n52096), .ZN(n52099) );
  XNOR2HSV1 U55448 ( .A1(n52100), .A2(n52099), .ZN(n52110) );
  NAND2HSV0 U55449 ( .A1(n59587), .A2(n52859), .ZN(n52101) );
  XOR2HSV0 U55450 ( .A1(n52102), .A2(n52101), .Z(n52108) );
  NOR2HSV0 U55451 ( .A1(n52103), .A2(n47511), .ZN(n52106) );
  NAND2HSV0 U55452 ( .A1(n52104), .A2(\pe2/bq[6] ), .ZN(n52105) );
  XOR2HSV0 U55453 ( .A1(n52106), .A2(n52105), .Z(n52107) );
  XOR2HSV0 U55454 ( .A1(n52108), .A2(n52107), .Z(n52109) );
  XOR3HSV2 U55455 ( .A1(n52111), .A2(n52110), .A3(n52109), .Z(n52112) );
  XNOR2HSV1 U55456 ( .A1(n52113), .A2(n52112), .ZN(n52114) );
  XNOR2HSV1 U55457 ( .A1(n52115), .A2(n52114), .ZN(n52116) );
  XNOR2HSV1 U55458 ( .A1(n52117), .A2(n52116), .ZN(n52119) );
  NAND2HSV0 U55459 ( .A1(n59766), .A2(n52239), .ZN(n52118) );
  XOR2HSV0 U55460 ( .A1(n52119), .A2(n52118), .Z(n52122) );
  NAND2HSV0 U55461 ( .A1(n52120), .A2(n51896), .ZN(n52121) );
  XNOR2HSV1 U55462 ( .A1(n52122), .A2(n52121), .ZN(n52123) );
  XNOR2HSV1 U55463 ( .A1(n52124), .A2(n52123), .ZN(n52127) );
  NAND2HSV0 U55464 ( .A1(n59761), .A2(n52125), .ZN(n52126) );
  XOR3HSV2 U55465 ( .A1(n52128), .A2(n52127), .A3(n52126), .Z(n52129) );
  XNOR2HSV1 U55466 ( .A1(n52130), .A2(n52129), .ZN(n52131) );
  XNOR2HSV1 U55467 ( .A1(n52132), .A2(n52131), .ZN(n52134) );
  NOR2HSV0 U55468 ( .A1(n53065), .A2(n49656), .ZN(n52133) );
  XOR3HSV2 U55469 ( .A1(n52135), .A2(n52134), .A3(n52133), .Z(n52136) );
  XOR2HSV0 U55470 ( .A1(n52137), .A2(n52136), .Z(n52141) );
  CLKNAND2HSV0 U55471 ( .A1(n52532), .A2(n53055), .ZN(n52140) );
  CLKNAND2HSV0 U55472 ( .A1(n52138), .A2(n51958), .ZN(n52139) );
  XOR3HSV2 U55473 ( .A1(n52141), .A2(n52140), .A3(n52139), .Z(n52142) );
  XNOR2HSV1 U55474 ( .A1(n52143), .A2(n52142), .ZN(n52145) );
  NAND2HSV0 U55475 ( .A1(n53382), .A2(n38782), .ZN(n52144) );
  XOR3HSV2 U55476 ( .A1(n52146), .A2(n52145), .A3(n52144), .Z(n52147) );
  XOR2HSV0 U55477 ( .A1(n52148), .A2(n52147), .Z(n52149) );
  XNOR2HSV1 U55478 ( .A1(n52150), .A2(n52149), .ZN(n52151) );
  XNOR2HSV1 U55479 ( .A1(n52152), .A2(n52151), .ZN(n52154) );
  CLKNAND2HSV0 U55480 ( .A1(n52399), .A2(n52167), .ZN(n52153) );
  XNOR2HSV1 U55481 ( .A1(n52154), .A2(n52153), .ZN(n52155) );
  XOR2HSV0 U55482 ( .A1(n52156), .A2(n52155), .Z(n52157) );
  XOR2HSV0 U55483 ( .A1(n52158), .A2(n52157), .Z(n52159) );
  XOR2HSV0 U55484 ( .A1(n52160), .A2(n52159), .Z(n52162) );
  NAND2HSV2 U55485 ( .A1(n52910), .A2(n44711), .ZN(n52161) );
  XNOR2HSV4 U55486 ( .A1(n52162), .A2(n52161), .ZN(n52166) );
  INAND2HSV2 U55487 ( .A1(n52164), .B1(n52163), .ZN(n52165) );
  XNOR2HSV4 U55488 ( .A1(n52166), .A2(n52165), .ZN(\pe2/poht [6]) );
  NAND2HSV2 U55489 ( .A1(n25709), .A2(n52416), .ZN(n52282) );
  CLKNAND2HSV1 U55490 ( .A1(n52854), .A2(n45249), .ZN(n52280) );
  CLKNAND2HSV1 U55491 ( .A1(n45389), .A2(n52167), .ZN(n52275) );
  CLKNAND2HSV1 U55492 ( .A1(n59929), .A2(n59685), .ZN(n52273) );
  CLKNAND2HSV1 U55493 ( .A1(n59927), .A2(n59982), .ZN(n52271) );
  NOR2HSV1 U55494 ( .A1(n52170), .A2(n52169), .ZN(n52269) );
  CLKNAND2HSV0 U55495 ( .A1(n52920), .A2(n38782), .ZN(n52267) );
  NOR2HSV0 U55496 ( .A1(n52171), .A2(n47573), .ZN(n52265) );
  NAND2HSV0 U55497 ( .A1(n59769), .A2(n52172), .ZN(n52258) );
  NAND2HSV0 U55498 ( .A1(n52930), .A2(n25824), .ZN(n52256) );
  CLKNAND2HSV0 U55499 ( .A1(n52417), .A2(n44714), .ZN(n52254) );
  NAND2HSV0 U55500 ( .A1(n52927), .A2(\pe2/got [8]), .ZN(n52250) );
  NAND2HSV0 U55501 ( .A1(n51609), .A2(n52174), .ZN(n52248) );
  NAND2HSV0 U55502 ( .A1(n52175), .A2(n52419), .ZN(n52246) );
  NAND2HSV0 U55503 ( .A1(n51896), .A2(n52176), .ZN(n52243) );
  NAND2HSV0 U55504 ( .A1(n52932), .A2(n52896), .ZN(n52236) );
  CLKNAND2HSV0 U55505 ( .A1(n52456), .A2(n52965), .ZN(n52178) );
  NAND2HSV0 U55506 ( .A1(\pe2/aot [8]), .A2(n52988), .ZN(n52177) );
  XOR2HSV0 U55507 ( .A1(n52178), .A2(n52177), .Z(n52183) );
  NAND2HSV0 U55508 ( .A1(n52344), .A2(n52179), .ZN(n52181) );
  NAND2HSV0 U55509 ( .A1(\pe2/aot [2]), .A2(n38053), .ZN(n52180) );
  XOR2HSV0 U55510 ( .A1(n52181), .A2(n52180), .Z(n52182) );
  XOR2HSV0 U55511 ( .A1(n52183), .A2(n52182), .Z(n52192) );
  NAND2HSV0 U55512 ( .A1(n59499), .A2(\pe2/bq[21] ), .ZN(n52186) );
  NAND2HSV0 U55513 ( .A1(n52184), .A2(n52299), .ZN(n52185) );
  XOR2HSV0 U55514 ( .A1(n52186), .A2(n52185), .Z(n52190) );
  NAND2HSV0 U55515 ( .A1(n59636), .A2(n51733), .ZN(n52188) );
  NAND2HSV0 U55516 ( .A1(n53005), .A2(\pe2/bq[14] ), .ZN(n52187) );
  XOR2HSV0 U55517 ( .A1(n52188), .A2(n52187), .Z(n52189) );
  XOR2HSV0 U55518 ( .A1(n52190), .A2(n52189), .Z(n52191) );
  XOR2HSV0 U55519 ( .A1(n52192), .A2(n52191), .Z(n52213) );
  NAND2HSV0 U55520 ( .A1(\pe2/aot [17]), .A2(n52193), .ZN(n52195) );
  NAND2HSV0 U55521 ( .A1(\pe2/aot [7]), .A2(n43961), .ZN(n52194) );
  XOR2HSV0 U55522 ( .A1(n52195), .A2(n52194), .Z(n52199) );
  NAND2HSV0 U55523 ( .A1(n59975), .A2(n52962), .ZN(n52197) );
  NAND2HSV0 U55524 ( .A1(\pe2/aot [10]), .A2(\pe2/bq[16] ), .ZN(n52196) );
  XOR2HSV0 U55525 ( .A1(n52197), .A2(n52196), .Z(n52198) );
  XNOR2HSV1 U55526 ( .A1(n52199), .A2(n52198), .ZN(n52211) );
  NOR2HSV0 U55527 ( .A1(n52095), .A2(n44854), .ZN(n52445) );
  NOR2HSV0 U55528 ( .A1(n52200), .A2(n44844), .ZN(n52203) );
  OAI22HSV0 U55529 ( .A1(n52445), .A2(n52203), .B1(n52202), .B2(n52201), .ZN(
        n52209) );
  NAND2HSV0 U55530 ( .A1(n59758), .A2(n52857), .ZN(n52206) );
  AOI22HSV1 U55531 ( .A1(n52207), .A2(n52206), .B1(n52205), .B2(n52204), .ZN(
        n52208) );
  XOR2HSV0 U55532 ( .A1(n52209), .A2(n52208), .Z(n52210) );
  XNOR2HSV1 U55533 ( .A1(n52211), .A2(n52210), .ZN(n52212) );
  XNOR2HSV1 U55534 ( .A1(n52213), .A2(n52212), .ZN(n52234) );
  CLKNHSV0 U55535 ( .I(n52939), .ZN(n52218) );
  AOI21HSV0 U55536 ( .A1(n59976), .A2(n52215), .B(n52214), .ZN(n52216) );
  AOI21HSV0 U55537 ( .A1(n52218), .A2(n52217), .B(n52216), .ZN(n52222) );
  XOR2HSV0 U55538 ( .A1(n52220), .A2(n52219), .Z(n52221) );
  XOR3HSV2 U55539 ( .A1(n52223), .A2(n52222), .A3(n52221), .Z(n52232) );
  NAND2HSV0 U55540 ( .A1(n59587), .A2(\pe2/bq[6] ), .ZN(n52224) );
  XOR2HSV0 U55541 ( .A1(n52225), .A2(n52224), .Z(n52230) );
  NOR2HSV0 U55542 ( .A1(n52226), .A2(n49515), .ZN(n52228) );
  NAND2HSV0 U55543 ( .A1(n52294), .A2(n52859), .ZN(n52227) );
  XOR2HSV0 U55544 ( .A1(n52228), .A2(n52227), .Z(n52229) );
  XOR2HSV0 U55545 ( .A1(n52230), .A2(n52229), .Z(n52231) );
  XOR2HSV0 U55546 ( .A1(n52232), .A2(n52231), .Z(n52233) );
  XNOR2HSV1 U55547 ( .A1(n52234), .A2(n52233), .ZN(n52235) );
  XNOR2HSV1 U55548 ( .A1(n52236), .A2(n52235), .ZN(n52238) );
  NAND2HSV0 U55549 ( .A1(n59766), .A2(n51932), .ZN(n52237) );
  XOR2HSV0 U55550 ( .A1(n52238), .A2(n52237), .Z(n52241) );
  NAND2HSV0 U55551 ( .A1(n44120), .A2(n52239), .ZN(n52240) );
  XNOR2HSV1 U55552 ( .A1(n52241), .A2(n52240), .ZN(n52242) );
  XNOR2HSV1 U55553 ( .A1(n52243), .A2(n52242), .ZN(n52245) );
  NAND2HSV0 U55554 ( .A1(n59761), .A2(\pe2/got [6]), .ZN(n52244) );
  XOR3HSV2 U55555 ( .A1(n52246), .A2(n52245), .A3(n52244), .Z(n52247) );
  XNOR2HSV1 U55556 ( .A1(n52248), .A2(n52247), .ZN(n52249) );
  XNOR2HSV1 U55557 ( .A1(n52250), .A2(n52249), .ZN(n52253) );
  NAND2HSV0 U55558 ( .A1(n52251), .A2(\pe2/got [10]), .ZN(n52252) );
  XOR3HSV2 U55559 ( .A1(n52254), .A2(n52253), .A3(n52252), .Z(n52255) );
  XNOR2HSV1 U55560 ( .A1(n52256), .A2(n52255), .ZN(n52257) );
  XNOR2HSV1 U55561 ( .A1(n52258), .A2(n52257), .ZN(n52260) );
  CLKNAND2HSV0 U55562 ( .A1(n51862), .A2(n53055), .ZN(n52259) );
  XNOR2HSV1 U55563 ( .A1(n52260), .A2(n52259), .ZN(n52261) );
  XNOR2HSV1 U55564 ( .A1(n52262), .A2(n52261), .ZN(n52264) );
  CLKNAND2HSV0 U55565 ( .A1(n53382), .A2(n51796), .ZN(n52263) );
  XOR3HSV2 U55566 ( .A1(n52265), .A2(n52264), .A3(n52263), .Z(n52266) );
  XOR2HSV0 U55567 ( .A1(n52267), .A2(n52266), .Z(n52268) );
  XNOR2HSV1 U55568 ( .A1(n52269), .A2(n52268), .ZN(n52270) );
  XNOR2HSV1 U55569 ( .A1(n52271), .A2(n52270), .ZN(n52272) );
  XNOR2HSV1 U55570 ( .A1(n52273), .A2(n52272), .ZN(n52274) );
  XNOR2HSV1 U55571 ( .A1(n52275), .A2(n52274), .ZN(n52278) );
  XNOR2HSV1 U55572 ( .A1(n52278), .A2(n52277), .ZN(n52279) );
  XOR2HSV0 U55573 ( .A1(n52280), .A2(n52279), .Z(n52281) );
  XNOR2HSV4 U55574 ( .A1(n52282), .A2(n52281), .ZN(n52284) );
  INAND2HSV2 U55575 ( .A1(n39088), .B1(n52558), .ZN(n52283) );
  XNOR2HSV4 U55576 ( .A1(n52284), .A2(n52283), .ZN(\pe2/poht [7]) );
  CLKNAND2HSV1 U55577 ( .A1(n52047), .A2(n38327), .ZN(n52408) );
  CLKNAND2HSV1 U55578 ( .A1(n51120), .A2(n59981), .ZN(n52406) );
  INAND2HSV0 U55579 ( .A1(n52285), .B1(n52918), .ZN(n52404) );
  CLKNAND2HSV0 U55580 ( .A1(n52919), .A2(n53077), .ZN(n52398) );
  NAND2HSV0 U55581 ( .A1(n59522), .A2(n38904), .ZN(n52396) );
  NOR2HSV0 U55582 ( .A1(n52921), .A2(n44327), .ZN(n52394) );
  CLKNAND2HSV1 U55583 ( .A1(n52923), .A2(n39075), .ZN(n52391) );
  NAND2HSV0 U55584 ( .A1(n59506), .A2(\pe2/got [16]), .ZN(n52386) );
  NAND2HSV0 U55585 ( .A1(n52286), .A2(n51608), .ZN(n52384) );
  CLKNAND2HSV0 U55586 ( .A1(n52927), .A2(n53055), .ZN(n52381) );
  NAND2HSV0 U55587 ( .A1(n52928), .A2(n52172), .ZN(n52379) );
  NAND2HSV0 U55588 ( .A1(\pe2/got [10]), .A2(n52929), .ZN(n52377) );
  NAND2HSV0 U55589 ( .A1(n52287), .A2(\pe2/got [9]), .ZN(n52373) );
  NAND2HSV0 U55590 ( .A1(n52932), .A2(n53041), .ZN(n52366) );
  NAND2HSV0 U55591 ( .A1(n52288), .A2(n53038), .ZN(n52364) );
  NOR2HSV0 U55592 ( .A1(n53033), .A2(n50910), .ZN(n52360) );
  AOI22HSV0 U55593 ( .A1(n52289), .A2(n52935), .B1(n59759), .B2(n52484), .ZN(
        n52290) );
  AOI21HSV0 U55594 ( .A1(n52947), .A2(n52291), .B(n52290), .ZN(n52298) );
  NOR2HSV0 U55595 ( .A1(n52293), .A2(n52292), .ZN(n52296) );
  AOI22HSV0 U55596 ( .A1(n52998), .A2(n52866), .B1(n52294), .B2(n52438), .ZN(
        n52295) );
  NOR2HSV1 U55597 ( .A1(n52296), .A2(n52295), .ZN(n52297) );
  XOR2HSV0 U55598 ( .A1(n52298), .A2(n52297), .Z(n52321) );
  NAND2HSV0 U55599 ( .A1(n59768), .A2(n52299), .ZN(n52302) );
  NAND2HSV0 U55600 ( .A1(n52951), .A2(n52300), .ZN(n52301) );
  XOR2HSV0 U55601 ( .A1(n52302), .A2(n52301), .Z(n52306) );
  NAND2HSV0 U55602 ( .A1(n39029), .A2(n51997), .ZN(n52304) );
  NAND2HSV0 U55603 ( .A1(n39052), .A2(n52073), .ZN(n52303) );
  XOR2HSV0 U55604 ( .A1(n52304), .A2(n52303), .Z(n52305) );
  XOR2HSV0 U55605 ( .A1(n52306), .A2(n52305), .Z(n52320) );
  NOR2HSV0 U55606 ( .A1(n49618), .A2(n44699), .ZN(n52460) );
  AOI22HSV0 U55607 ( .A1(\pe2/aot [2]), .A2(n36608), .B1(n38393), .B2(n53016), 
        .ZN(n52307) );
  AOI21HSV2 U55608 ( .A1(n52308), .A2(n52460), .B(n52307), .ZN(n52314) );
  NOR2HSV0 U55609 ( .A1(n44095), .A2(n51842), .ZN(n52491) );
  AOI22HSV0 U55610 ( .A1(n52974), .A2(n52994), .B1(n52310), .B2(n52309), .ZN(
        n52311) );
  AOI21HSV2 U55611 ( .A1(n52312), .A2(n52491), .B(n52311), .ZN(n52313) );
  XNOR2HSV1 U55612 ( .A1(n52314), .A2(n52313), .ZN(n52318) );
  NAND2HSV0 U55613 ( .A1(n52955), .A2(n52962), .ZN(n52316) );
  NAND2HSV0 U55614 ( .A1(n51759), .A2(\pe2/bq[14] ), .ZN(n52315) );
  XOR2HSV0 U55615 ( .A1(n52316), .A2(n52315), .Z(n52317) );
  XNOR2HSV1 U55616 ( .A1(n52318), .A2(n52317), .ZN(n52319) );
  XOR3HSV2 U55617 ( .A1(n52321), .A2(n52320), .A3(n52319), .Z(n52357) );
  NAND2HSV0 U55618 ( .A1(n37801), .A2(n52322), .ZN(n52324) );
  NAND2HSV0 U55619 ( .A1(n52485), .A2(\pe2/bq[2] ), .ZN(n52323) );
  XOR2HSV0 U55620 ( .A1(n52324), .A2(n52323), .Z(n52328) );
  NAND2HSV0 U55621 ( .A1(n59636), .A2(\pe2/bq[17] ), .ZN(n52326) );
  NAND2HSV0 U55622 ( .A1(n59974), .A2(n51732), .ZN(n52325) );
  XOR2HSV0 U55623 ( .A1(n52326), .A2(n52325), .Z(n52327) );
  XOR2HSV0 U55624 ( .A1(n52328), .A2(n52327), .Z(n52336) );
  NAND2HSV0 U55625 ( .A1(n59976), .A2(n52965), .ZN(n52330) );
  NAND2HSV0 U55626 ( .A1(n53005), .A2(n38792), .ZN(n52329) );
  XOR2HSV0 U55627 ( .A1(n52330), .A2(n52329), .Z(n52334) );
  NAND2HSV0 U55628 ( .A1(n59499), .A2(n38064), .ZN(n52332) );
  NAND2HSV0 U55629 ( .A1(n52456), .A2(n44987), .ZN(n52331) );
  XOR2HSV0 U55630 ( .A1(n52332), .A2(n52331), .Z(n52333) );
  XOR2HSV0 U55631 ( .A1(n52334), .A2(n52333), .Z(n52335) );
  XOR2HSV0 U55632 ( .A1(n52336), .A2(n52335), .Z(n52354) );
  NAND2HSV0 U55633 ( .A1(n52966), .A2(n52988), .ZN(n52339) );
  NAND2HSV0 U55634 ( .A1(n59973), .A2(n52337), .ZN(n52338) );
  XOR2HSV0 U55635 ( .A1(n52339), .A2(n52338), .Z(n52343) );
  NAND2HSV0 U55636 ( .A1(n53009), .A2(\pe2/bq[21] ), .ZN(n52341) );
  NAND2HSV0 U55637 ( .A1(n59633), .A2(n38053), .ZN(n52340) );
  XOR2HSV0 U55638 ( .A1(n52341), .A2(n52340), .Z(n52342) );
  XOR2HSV0 U55639 ( .A1(n52343), .A2(n52342), .Z(n52352) );
  NAND2HSV0 U55640 ( .A1(n52993), .A2(n52973), .ZN(n52346) );
  NAND2HSV0 U55641 ( .A1(n52344), .A2(n52987), .ZN(n52345) );
  XOR2HSV0 U55642 ( .A1(n52346), .A2(n52345), .Z(n52350) );
  NOR2HSV0 U55643 ( .A1(n47574), .A2(n51567), .ZN(n52348) );
  NAND2HSV0 U55644 ( .A1(n50956), .A2(n51457), .ZN(n52347) );
  XOR2HSV0 U55645 ( .A1(n52348), .A2(n52347), .Z(n52349) );
  XOR2HSV0 U55646 ( .A1(n52350), .A2(n52349), .Z(n52351) );
  XOR2HSV0 U55647 ( .A1(n52352), .A2(n52351), .Z(n52353) );
  XOR2HSV0 U55648 ( .A1(n52354), .A2(n52353), .Z(n52356) );
  NAND2HSV0 U55649 ( .A1(n38539), .A2(n52895), .ZN(n52355) );
  XOR3HSV2 U55650 ( .A1(n52357), .A2(n52356), .A3(n52355), .Z(n52359) );
  NAND2HSV0 U55651 ( .A1(n59669), .A2(n52239), .ZN(n52358) );
  XOR3HSV2 U55652 ( .A1(n52360), .A2(n52359), .A3(n52358), .Z(n52362) );
  NAND2HSV0 U55653 ( .A1(n38702), .A2(n59984), .ZN(n52361) );
  XNOR2HSV1 U55654 ( .A1(n52362), .A2(n52361), .ZN(n52363) );
  XNOR2HSV1 U55655 ( .A1(n52364), .A2(n52363), .ZN(n52365) );
  XNOR2HSV1 U55656 ( .A1(n52366), .A2(n52365), .ZN(n52369) );
  NAND2HSV0 U55657 ( .A1(n52367), .A2(n59757), .ZN(n52368) );
  XOR2HSV0 U55658 ( .A1(n52369), .A2(n52368), .Z(n52371) );
  NAND2HSV0 U55659 ( .A1(n53050), .A2(\pe2/got [8]), .ZN(n52370) );
  XNOR2HSV1 U55660 ( .A1(n52371), .A2(n52370), .ZN(n52372) );
  XNOR2HSV1 U55661 ( .A1(n52373), .A2(n52372), .ZN(n52376) );
  NAND2HSV0 U55662 ( .A1(n53056), .A2(n52374), .ZN(n52375) );
  XOR3HSV2 U55663 ( .A1(n52377), .A2(n52376), .A3(n52375), .Z(n52378) );
  XNOR2HSV1 U55664 ( .A1(n52379), .A2(n52378), .ZN(n52380) );
  XNOR2HSV1 U55665 ( .A1(n52381), .A2(n52380), .ZN(n52383) );
  NOR2HSV0 U55666 ( .A1(n53065), .A2(n47573), .ZN(n52382) );
  XOR3HSV2 U55667 ( .A1(n52384), .A2(n52383), .A3(n52382), .Z(n52385) );
  XNOR2HSV1 U55668 ( .A1(n52386), .A2(n52385), .ZN(n52389) );
  NAND2HSV0 U55669 ( .A1(n52924), .A2(\pe2/got [17]), .ZN(n52388) );
  NAND2HSV0 U55670 ( .A1(n59361), .A2(n52925), .ZN(n52387) );
  XOR3HSV2 U55671 ( .A1(n52389), .A2(n52388), .A3(n52387), .Z(n52390) );
  XNOR2HSV1 U55672 ( .A1(n52391), .A2(n52390), .ZN(n52393) );
  NAND2HSV0 U55673 ( .A1(n53382), .A2(n52922), .ZN(n52392) );
  XOR3HSV2 U55674 ( .A1(n52394), .A2(n52393), .A3(n52392), .Z(n52395) );
  XOR2HSV0 U55675 ( .A1(n52396), .A2(n52395), .Z(n52397) );
  XNOR2HSV1 U55676 ( .A1(n52398), .A2(n52397), .ZN(n52402) );
  NAND2HSV0 U55677 ( .A1(n59927), .A2(n59584), .ZN(n52401) );
  CLKNAND2HSV0 U55678 ( .A1(n52399), .A2(\pe2/got [25]), .ZN(n52400) );
  XOR3HSV2 U55679 ( .A1(n52402), .A2(n52401), .A3(n52400), .Z(n52403) );
  XOR2HSV0 U55680 ( .A1(n52404), .A2(n52403), .Z(n52405) );
  XOR2HSV0 U55681 ( .A1(n52408), .A2(n52407), .Z(n52410) );
  NAND2HSV2 U55682 ( .A1(n52910), .A2(n59635), .ZN(n52409) );
  XNOR2HSV4 U55683 ( .A1(n52410), .A2(n52409), .ZN(n52413) );
  INAND2HSV2 U55684 ( .A1(n52411), .B1(n52558), .ZN(n52412) );
  XNOR2HSV4 U55685 ( .A1(n52413), .A2(n52412), .ZN(\pe2/poht [2]) );
  CLKNAND2HSV1 U55686 ( .A1(n52414), .A2(n52916), .ZN(n52555) );
  CLKNAND2HSV0 U55687 ( .A1(n52918), .A2(n44944), .ZN(n52551) );
  CLKNAND2HSV0 U55688 ( .A1(n52919), .A2(n52416), .ZN(n52546) );
  NAND2HSV0 U55689 ( .A1(n52920), .A2(n53077), .ZN(n52544) );
  NOR2HSV0 U55690 ( .A1(n52921), .A2(n38711), .ZN(n52542) );
  CLKNAND2HSV0 U55691 ( .A1(n52923), .A2(\pe2/got [20]), .ZN(n52539) );
  NAND2HSV0 U55692 ( .A1(n52814), .A2(\pe2/got [17]), .ZN(n52531) );
  CLKNAND2HSV0 U55693 ( .A1(n52417), .A2(n51964), .ZN(n52529) );
  CLKNAND2HSV1 U55694 ( .A1(n52927), .A2(n51958), .ZN(n52525) );
  NAND2HSV0 U55695 ( .A1(n52928), .A2(n52418), .ZN(n52523) );
  NAND2HSV0 U55696 ( .A1(n52930), .A2(n52419), .ZN(n52521) );
  CLKNAND2HSV0 U55697 ( .A1(n52931), .A2(\pe2/got [10]), .ZN(n52518) );
  NAND2HSV0 U55698 ( .A1(n52932), .A2(n52933), .ZN(n52512) );
  NAND2HSV0 U55699 ( .A1(n48896), .A2(n53041), .ZN(n52510) );
  NAND2HSV0 U55700 ( .A1(n43928), .A2(n59984), .ZN(n52506) );
  NAND2HSV0 U55701 ( .A1(n59684), .A2(n52239), .ZN(n52422) );
  NOR2HSV0 U55702 ( .A1(n52420), .A2(n50926), .ZN(n52421) );
  XNOR2HSV1 U55703 ( .A1(n52422), .A2(n52421), .ZN(n52504) );
  NOR2HSV0 U55704 ( .A1(n38907), .A2(n50910), .ZN(n52502) );
  NAND2HSV0 U55705 ( .A1(\pe2/aot [12]), .A2(n52965), .ZN(n52424) );
  NAND2HSV0 U55706 ( .A1(n44745), .A2(n52988), .ZN(n52423) );
  XOR2HSV0 U55707 ( .A1(n52424), .A2(n52423), .Z(n52428) );
  NAND2HSV0 U55708 ( .A1(n59974), .A2(\pe2/bq[17] ), .ZN(n52426) );
  NAND2HSV0 U55709 ( .A1(n51759), .A2(n49619), .ZN(n52425) );
  XOR2HSV0 U55710 ( .A1(n52426), .A2(n52425), .Z(n52427) );
  XOR2HSV0 U55711 ( .A1(n52428), .A2(n52427), .Z(n52442) );
  NOR2HSV0 U55712 ( .A1(n38822), .A2(n52429), .ZN(n52435) );
  NOR2HSV0 U55713 ( .A1(n52431), .A2(n52430), .ZN(n52434) );
  OAI22HSV0 U55714 ( .A1(n52435), .A2(n52434), .B1(n52433), .B2(n52432), .ZN(
        n52440) );
  XNOR2HSV1 U55715 ( .A1(n52440), .A2(n52439), .ZN(n52441) );
  XNOR2HSV1 U55716 ( .A1(n52442), .A2(n52441), .ZN(n52465) );
  NOR2HSV0 U55717 ( .A1(n52447), .A2(n52446), .ZN(n52451) );
  AOI22HSV0 U55718 ( .A1(n52449), .A2(n52935), .B1(\pe2/aot [22]), .B2(n52448), 
        .ZN(n52450) );
  NOR2HSV1 U55719 ( .A1(n52451), .A2(n52450), .ZN(n52452) );
  XOR2HSV0 U55720 ( .A1(n52453), .A2(n52452), .Z(n52463) );
  NOR2HSV0 U55721 ( .A1(n52455), .A2(n52454), .ZN(n52459) );
  AOI22HSV0 U55722 ( .A1(n52457), .A2(n45015), .B1(n38064), .B2(n52456), .ZN(
        n52458) );
  NOR2HSV2 U55723 ( .A1(n52459), .A2(n52458), .ZN(n52461) );
  XNOR2HSV1 U55724 ( .A1(n52461), .A2(n52460), .ZN(n52462) );
  XNOR2HSV1 U55725 ( .A1(n52463), .A2(n52462), .ZN(n52464) );
  XNOR2HSV1 U55726 ( .A1(n52465), .A2(n52464), .ZN(n52501) );
  NAND2HSV0 U55727 ( .A1(n59976), .A2(\pe2/bq[21] ), .ZN(n52467) );
  NAND2HSV0 U55728 ( .A1(n59768), .A2(n52179), .ZN(n52466) );
  XOR2HSV0 U55729 ( .A1(n52467), .A2(n52466), .Z(n52471) );
  NAND2HSV0 U55730 ( .A1(n59969), .A2(\pe2/bq[2] ), .ZN(n52469) );
  NAND2HSV0 U55731 ( .A1(n59971), .A2(n51457), .ZN(n52468) );
  XOR2HSV0 U55732 ( .A1(n52469), .A2(n52468), .Z(n52470) );
  XOR2HSV0 U55733 ( .A1(n52471), .A2(n52470), .Z(n52480) );
  NAND2HSV0 U55734 ( .A1(\pe2/aot [19]), .A2(n52472), .ZN(n52474) );
  NAND2HSV0 U55735 ( .A1(n52993), .A2(n52987), .ZN(n52473) );
  XOR2HSV0 U55736 ( .A1(n52474), .A2(n52473), .Z(n52478) );
  NAND2HSV0 U55737 ( .A1(n59973), .A2(n52984), .ZN(n52476) );
  NAND2HSV0 U55738 ( .A1(n59499), .A2(n39032), .ZN(n52475) );
  XOR2HSV0 U55739 ( .A1(n52476), .A2(n52475), .Z(n52477) );
  XOR2HSV0 U55740 ( .A1(n52478), .A2(n52477), .Z(n52479) );
  XOR2HSV0 U55741 ( .A1(n52480), .A2(n52479), .Z(n52499) );
  NAND2HSV0 U55742 ( .A1(n59758), .A2(n52073), .ZN(n52483) );
  NAND2HSV0 U55743 ( .A1(\pe2/aot [23]), .A2(n52481), .ZN(n52482) );
  XOR2HSV0 U55744 ( .A1(n52483), .A2(n52482), .Z(n52489) );
  NAND2HSV0 U55745 ( .A1(n52485), .A2(n52484), .ZN(n52487) );
  NAND2HSV0 U55746 ( .A1(n52955), .A2(\pe2/bq[14] ), .ZN(n52486) );
  XOR2HSV0 U55747 ( .A1(n52487), .A2(n52486), .Z(n52488) );
  XOR2HSV0 U55748 ( .A1(n52489), .A2(n52488), .Z(n52497) );
  XOR2HSV0 U55749 ( .A1(n52491), .A2(n52490), .Z(n52495) );
  NOR2HSV0 U55750 ( .A1(n38655), .A2(n51567), .ZN(n52493) );
  NAND2HSV0 U55751 ( .A1(n52974), .A2(\pe2/bq[6] ), .ZN(n52492) );
  XOR2HSV0 U55752 ( .A1(n52493), .A2(n52492), .Z(n52494) );
  XOR2HSV0 U55753 ( .A1(n52495), .A2(n52494), .Z(n52496) );
  XOR2HSV0 U55754 ( .A1(n52497), .A2(n52496), .Z(n52498) );
  XOR2HSV0 U55755 ( .A1(n52499), .A2(n52498), .Z(n52500) );
  XOR3HSV2 U55756 ( .A1(n52502), .A2(n52501), .A3(n52500), .Z(n52503) );
  XNOR2HSV1 U55757 ( .A1(n52504), .A2(n52503), .ZN(n52505) );
  XNOR2HSV1 U55758 ( .A1(n52506), .A2(n52505), .ZN(n52508) );
  NAND2HSV0 U55759 ( .A1(n38702), .A2(n53038), .ZN(n52507) );
  XNOR2HSV1 U55760 ( .A1(n52508), .A2(n52507), .ZN(n52509) );
  XNOR2HSV1 U55761 ( .A1(n52510), .A2(n52509), .ZN(n52511) );
  XNOR2HSV1 U55762 ( .A1(n52512), .A2(n52511), .ZN(n52514) );
  NAND2HSV0 U55763 ( .A1(n59766), .A2(\pe2/got [8]), .ZN(n52513) );
  XOR2HSV0 U55764 ( .A1(n52514), .A2(n52513), .Z(n52516) );
  NAND2HSV0 U55765 ( .A1(n53050), .A2(\pe2/got [9]), .ZN(n52515) );
  XNOR2HSV1 U55766 ( .A1(n52516), .A2(n52515), .ZN(n52517) );
  XNOR2HSV1 U55767 ( .A1(n52518), .A2(n52517), .ZN(n52520) );
  NAND2HSV0 U55768 ( .A1(n53056), .A2(n52172), .ZN(n52519) );
  XOR3HSV2 U55769 ( .A1(n52521), .A2(n52520), .A3(n52519), .Z(n52522) );
  XNOR2HSV1 U55770 ( .A1(n52523), .A2(n52522), .ZN(n52524) );
  XNOR2HSV1 U55771 ( .A1(n52525), .A2(n52524), .ZN(n52528) );
  NOR2HSV0 U55772 ( .A1(n53065), .A2(n52526), .ZN(n52527) );
  XOR3HSV2 U55773 ( .A1(n52529), .A2(n52528), .A3(n52527), .Z(n52530) );
  XOR2HSV0 U55774 ( .A1(n52531), .A2(n52530), .Z(n52537) );
  CLKNAND2HSV0 U55775 ( .A1(n52532), .A2(n52925), .ZN(n52536) );
  NAND2HSV0 U55776 ( .A1(n52534), .A2(n52533), .ZN(n52535) );
  XOR3HSV2 U55777 ( .A1(n52537), .A2(n52536), .A3(n52535), .Z(n52538) );
  XNOR2HSV1 U55778 ( .A1(n52539), .A2(n52538), .ZN(n52541) );
  CLKNAND2HSV0 U55779 ( .A1(n53078), .A2(n52276), .ZN(n52540) );
  XOR3HSV2 U55780 ( .A1(n52542), .A2(n52541), .A3(n52540), .Z(n52543) );
  XOR2HSV0 U55781 ( .A1(n52544), .A2(n52543), .Z(n52545) );
  XOR2HSV0 U55782 ( .A1(n52546), .A2(n52545), .Z(n52549) );
  CLKNAND2HSV1 U55783 ( .A1(n53087), .A2(\pe2/got [25]), .ZN(n52548) );
  CLKNAND2HSV0 U55784 ( .A1(n59929), .A2(n53086), .ZN(n52547) );
  XOR3HSV2 U55785 ( .A1(n52549), .A2(n52548), .A3(n52547), .Z(n52550) );
  XOR2HSV0 U55786 ( .A1(n52551), .A2(n52550), .Z(n52552) );
  XOR2HSV0 U55787 ( .A1(n52553), .A2(n52552), .Z(n52554) );
  XOR2HSV0 U55788 ( .A1(n52555), .A2(n52554), .Z(n52557) );
  NAND2HSV2 U55789 ( .A1(n52910), .A2(n38873), .ZN(n52556) );
  INAND2HSV2 U55790 ( .A1(n52559), .B1(n52558), .ZN(n52560) );
  XNOR2HSV4 U55791 ( .A1(n52561), .A2(n52560), .ZN(\pe2/poht [1]) );
  CLKNAND2HSV1 U55792 ( .A1(n51016), .A2(n52566), .ZN(n52664) );
  NOR2HSV0 U55793 ( .A1(n52567), .A2(n48722), .ZN(n52657) );
  CLKNAND2HSV1 U55794 ( .A1(n52569), .A2(n52568), .ZN(n52651) );
  NAND2HSV0 U55795 ( .A1(n52570), .A2(n48167), .ZN(n52649) );
  NAND2HSV0 U55796 ( .A1(n52572), .A2(n52571), .ZN(n52645) );
  NAND2HSV0 U55797 ( .A1(n59878), .A2(n50698), .ZN(n52640) );
  NAND2HSV0 U55798 ( .A1(n48681), .A2(n39471), .ZN(n52583) );
  NAND2HSV0 U55799 ( .A1(n59879), .A2(n52581), .ZN(n52582) );
  XOR2HSV0 U55800 ( .A1(n52583), .A2(n52582), .Z(n52589) );
  NAND2HSV0 U55801 ( .A1(n52584), .A2(n39914), .ZN(n52587) );
  NAND2HSV0 U55802 ( .A1(n59866), .A2(n52585), .ZN(n52586) );
  XOR2HSV0 U55803 ( .A1(n52587), .A2(n52586), .Z(n52588) );
  NAND2HSV0 U55804 ( .A1(n52590), .A2(\pe5/bq[2] ), .ZN(n52593) );
  NAND2HSV0 U55805 ( .A1(n52591), .A2(\pe5/bq[7] ), .ZN(n52592) );
  XOR2HSV0 U55806 ( .A1(n52593), .A2(n52592), .Z(n52599) );
  NAND2HSV0 U55807 ( .A1(n59895), .A2(n52594), .ZN(n52597) );
  NAND2HSV0 U55808 ( .A1(n51313), .A2(n52595), .ZN(n52596) );
  XOR2HSV0 U55809 ( .A1(n52597), .A2(n52596), .Z(n52598) );
  NAND2HSV0 U55810 ( .A1(n52600), .A2(n30891), .ZN(n52602) );
  NAND2HSV0 U55811 ( .A1(n53295), .A2(n46933), .ZN(n52601) );
  XOR2HSV0 U55812 ( .A1(n52602), .A2(n52601), .Z(n52606) );
  NAND2HSV0 U55813 ( .A1(n50501), .A2(n30607), .ZN(n52604) );
  NAND2HSV0 U55814 ( .A1(\pe5/aot [18]), .A2(n48775), .ZN(n52603) );
  XOR2HSV0 U55815 ( .A1(n52604), .A2(n52603), .Z(n52605) );
  NAND2HSV0 U55816 ( .A1(n52607), .A2(n48778), .ZN(n52609) );
  NAND2HSV0 U55817 ( .A1(n59640), .A2(\pe5/bq[11] ), .ZN(n52608) );
  XOR2HSV0 U55818 ( .A1(n52609), .A2(n52608), .Z(n52615) );
  NAND2HSV0 U55819 ( .A1(n52611), .A2(n52610), .ZN(n52613) );
  NAND2HSV0 U55820 ( .A1(n51187), .A2(n50526), .ZN(n52612) );
  XOR2HSV0 U55821 ( .A1(n52613), .A2(n52612), .Z(n52614) );
  NAND2HSV0 U55822 ( .A1(n39499), .A2(n53200), .ZN(n52617) );
  NAND2HSV0 U55823 ( .A1(n40190), .A2(\pe5/bq[8] ), .ZN(n52616) );
  AOI22HSV0 U55824 ( .A1(n50505), .A2(n52619), .B1(n52618), .B2(\pe5/aot [9]), 
        .ZN(n52620) );
  AOI21HSV0 U55825 ( .A1(n52622), .A2(n52621), .B(n52620), .ZN(n52629) );
  NAND2HSV0 U55826 ( .A1(\pe5/aot [23]), .A2(n51370), .ZN(n52626) );
  CLKNAND2HSV1 U55827 ( .A1(n52623), .A2(n51370), .ZN(n52680) );
  NOR2HSV0 U55828 ( .A1(n52624), .A2(n52680), .ZN(n52625) );
  AOI21HSV2 U55829 ( .A1(n52627), .A2(n52626), .B(n52625), .ZN(n52628) );
  NAND2HSV0 U55830 ( .A1(n52631), .A2(n52630), .ZN(n52634) );
  NAND2HSV0 U55831 ( .A1(\pe5/aot [13]), .A2(n52632), .ZN(n52633) );
  XOR2HSV0 U55832 ( .A1(n52634), .A2(n52633), .Z(n52638) );
  NAND2HSV0 U55833 ( .A1(n53304), .A2(n39487), .ZN(n52636) );
  NAND2HSV0 U55834 ( .A1(n59880), .A2(n39454), .ZN(n52635) );
  XOR2HSV0 U55835 ( .A1(n52636), .A2(n52635), .Z(n52637) );
  XNOR2HSV1 U55836 ( .A1(n52640), .A2(n52639), .ZN(n52643) );
  NAND2HSV0 U55837 ( .A1(n44694), .A2(n52641), .ZN(n52642) );
  XOR2HSV0 U55838 ( .A1(n52643), .A2(n52642), .Z(n52644) );
  XNOR2HSV1 U55839 ( .A1(n52645), .A2(n52644), .ZN(n52647) );
  NAND2HSV0 U55840 ( .A1(n59517), .A2(n53349), .ZN(n52646) );
  XNOR2HSV1 U55841 ( .A1(n52647), .A2(n52646), .ZN(n52648) );
  XNOR2HSV1 U55842 ( .A1(n52649), .A2(n52648), .ZN(n52650) );
  XNOR2HSV1 U55843 ( .A1(n52651), .A2(n52650), .ZN(n52655) );
  NAND2HSV0 U55844 ( .A1(n52653), .A2(n52652), .ZN(n52654) );
  XNOR2HSV1 U55845 ( .A1(n52655), .A2(n52654), .ZN(n52656) );
  XNOR2HSV1 U55846 ( .A1(n52657), .A2(n52656), .ZN(n52662) );
  CLKNAND2HSV1 U55847 ( .A1(n53338), .A2(n52658), .ZN(n52661) );
  NOR2HSV2 U55848 ( .A1(n52659), .A2(n50422), .ZN(n52660) );
  XOR3HSV2 U55849 ( .A1(n52662), .A2(n52661), .A3(n52660), .Z(n52663) );
  XNOR2HSV1 U55850 ( .A1(n52664), .A2(n52663), .ZN(n52666) );
  NAND2HSV0 U55851 ( .A1(n59516), .A2(n37556), .ZN(n52665) );
  CLKNAND2HSV1 U55852 ( .A1(n52670), .A2(\pe5/got [2]), .ZN(n52692) );
  NAND2HSV0 U55853 ( .A1(n53344), .A2(\pe5/got [1]), .ZN(n52690) );
  CLKNAND2HSV0 U55854 ( .A1(n50501), .A2(n52671), .ZN(n52674) );
  NAND2HSV0 U55855 ( .A1(n51339), .A2(n52672), .ZN(n52673) );
  XOR2HSV0 U55856 ( .A1(n52674), .A2(n52673), .Z(n52679) );
  NAND2HSV0 U55857 ( .A1(n52675), .A2(n52581), .ZN(n52677) );
  CLKNAND2HSV0 U55858 ( .A1(\pe5/aot [3]), .A2(\pe5/bq[6] ), .ZN(n52676) );
  XOR2HSV0 U55859 ( .A1(n52677), .A2(n52676), .Z(n52678) );
  XOR2HSV0 U55860 ( .A1(n52679), .A2(n52678), .Z(n52688) );
  XOR2HSV0 U55861 ( .A1(n52681), .A2(n52680), .Z(n52686) );
  NOR2HSV1 U55862 ( .A1(n51232), .A2(n47207), .ZN(n52684) );
  NAND2HSV0 U55863 ( .A1(n52682), .A2(n51281), .ZN(n52683) );
  XOR2HSV0 U55864 ( .A1(n52684), .A2(n52683), .Z(n52685) );
  XOR2HSV0 U55865 ( .A1(n52686), .A2(n52685), .Z(n52687) );
  XOR2HSV0 U55866 ( .A1(n52688), .A2(n52687), .Z(n52689) );
  XNOR2HSV1 U55867 ( .A1(n52690), .A2(n52689), .ZN(n52691) );
  BUFHSV2 U55868 ( .I(n59407), .Z(n59652) );
  BUFHSV2 U55869 ( .I(n59429), .Z(n59651) );
  BUFHSV2 U55870 ( .I(n59925), .Z(n59657) );
  BUFHSV2 U55871 ( .I(n59925), .Z(n59654) );
  BUFHSV2 U55872 ( .I(n59925), .Z(n59653) );
  BUFHSV2 U55873 ( .I(n59925), .Z(n59650) );
  BUFHSV2 U55874 ( .I(n59484), .Z(n59922) );
  BUFHSV2 U55875 ( .I(n59925), .Z(n59658) );
  BUFHSV2 U55876 ( .I(n59397), .Z(n59921) );
  BUFHSV2 U55877 ( .I(n59651), .Z(n59649) );
  INAND2HSV0 U55878 ( .A1(n52701), .B1(n52700), .ZN(n52702) );
  INHSV2 U55879 ( .I(n52702), .ZN(n52703) );
  XOR2HSV0 U55880 ( .A1(n52703), .A2(poh6[2]), .Z(po[3]) );
  CLKNHSV0 U55881 ( .I(n52704), .ZN(n52708) );
  NOR2HSV0 U55882 ( .A1(n52706), .A2(n52705), .ZN(n52707) );
  XOR3HSV0 U55883 ( .A1(n52709), .A2(n52708), .A3(n52707), .Z(n52711) );
  NOR2HSV0 U55884 ( .A1(n52711), .A2(n52710), .ZN(n52712) );
  XOR2HSV0 U55885 ( .A1(n52712), .A2(poh6[3]), .Z(po[4]) );
  NAND2HSV0 U55886 ( .A1(n59669), .A2(n47997), .ZN(n52722) );
  CLKNHSV2 U55887 ( .I(n52718), .ZN(n52720) );
  XOR2HSV0 U55888 ( .A1(n52720), .A2(n29743), .Z(n52721) );
  XNOR2HSV1 U55889 ( .A1(n52722), .A2(n52721), .ZN(n60100) );
  NAND2HSV0 U55890 ( .A1(n59662), .A2(n52723), .ZN(n52724) );
  XOR2HSV0 U55891 ( .A1(n33300), .A2(n52724), .Z(n60081) );
  NAND2HSV0 U55892 ( .A1(n52727), .A2(n52726), .ZN(n52728) );
  XOR2HSV0 U55893 ( .A1(n52733), .A2(n52732), .Z(n60073) );
  XOR2HSV0 U55894 ( .A1(n52735), .A2(n52734), .Z(n60072) );
  NAND2HSV0 U55895 ( .A1(n54456), .A2(n53650), .ZN(n52737) );
  XNOR2HSV1 U55896 ( .A1(n52737), .A2(n25398), .ZN(n60017) );
  NAND2HSV0 U55897 ( .A1(n52738), .A2(n36924), .ZN(n52740) );
  XNOR2HSV0 U55898 ( .A1(n52740), .A2(n52739), .ZN(n52742) );
  NAND2HSV0 U55899 ( .A1(n56070), .A2(n52726), .ZN(n52741) );
  XOR2HSV0 U55900 ( .A1(n52742), .A2(n52741), .Z(n60048) );
  NOR2HSV0 U55901 ( .A1(n41802), .A2(n44522), .ZN(n52744) );
  XOR2HSV0 U55902 ( .A1(n52744), .A2(n52743), .Z(pov1[11]) );
  NAND2HSV0 U55903 ( .A1(n59725), .A2(n52831), .ZN(n52764) );
  XOR2HSV0 U55904 ( .A1(n52764), .A2(n52763), .Z(pov1[14]) );
  NOR2HSV0 U55905 ( .A1(n52765), .A2(n32793), .ZN(n52766) );
  XOR2HSV0 U55906 ( .A1(n52766), .A2(poh6[14]), .Z(po[15]) );
  NAND2HSV0 U55907 ( .A1(n59878), .A2(n52767), .ZN(n52770) );
  CLKNHSV0 U55908 ( .I(n52768), .ZN(n52769) );
  XNOR2HSV1 U55909 ( .A1(n52770), .A2(n52769), .ZN(n60033) );
  CLKNHSV0 U55910 ( .I(n29751), .ZN(n52782) );
  NAND2HSV0 U55911 ( .A1(n29742), .A2(n52780), .ZN(n52781) );
  XNOR2HSV1 U55912 ( .A1(n52782), .A2(n52781), .ZN(n52783) );
  NOR2HSV1 U55913 ( .A1(n52783), .A2(n32685), .ZN(n52784) );
  XOR2HSV0 U55914 ( .A1(n52784), .A2(poh6[16]), .Z(po[17]) );
  CLKNHSV0 U55915 ( .I(n52793), .ZN(n52794) );
  NAND3HSV1 U55916 ( .A1(n52796), .A2(n52795), .A3(n52794), .ZN(n52798) );
  XOR2HSV0 U55917 ( .A1(n52798), .A2(n52797), .Z(n60011) );
  NAND2HSV0 U55918 ( .A1(n59525), .A2(n52799), .ZN(n52801) );
  XNOR2HSV1 U55919 ( .A1(n52801), .A2(n52800), .ZN(n52807) );
  AND2HSV2 U55920 ( .A1(n52803), .A2(n52802), .Z(n52805) );
  AND2HSV2 U55921 ( .A1(n52805), .A2(n52804), .Z(n52806) );
  XNOR2HSV1 U55922 ( .A1(n52807), .A2(n52806), .ZN(n60069) );
  XNOR2HSV1 U55923 ( .A1(n52821), .A2(n25878), .ZN(n60066) );
  XOR2HSV0 U55924 ( .A1(n52826), .A2(n35439), .Z(n60057) );
  CLKNAND2HSV0 U55925 ( .A1(n44968), .A2(n38264), .ZN(n52828) );
  XOR2HSV0 U55926 ( .A1(n52828), .A2(n29769), .Z(n60093) );
  CLKNHSV0 U55927 ( .I(n52829), .ZN(n52830) );
  INHSV2 U55928 ( .I(n52830), .ZN(n52833) );
  CLKNAND2HSV1 U55929 ( .A1(n59751), .A2(n52831), .ZN(n52832) );
  XOR2HSV0 U55930 ( .A1(n52833), .A2(n52832), .Z(pov1[25]) );
  NAND2HSV2 U55931 ( .A1(n51014), .A2(n52834), .ZN(n52837) );
  XOR2HSV0 U55932 ( .A1(n52837), .A2(n52836), .Z(n60000) );
  XOR2HSV0 U55933 ( .A1(n52839), .A2(n52838), .Z(n60006) );
  CLKNAND2HSV1 U55934 ( .A1(n52840), .A2(n47997), .ZN(n52842) );
  XOR2HSV0 U55935 ( .A1(n52842), .A2(n52841), .Z(n60014) );
  CLKBUFHSV4 U55936 ( .I(n54553), .Z(n55569) );
  CLKNAND2HSV1 U55937 ( .A1(n55569), .A2(n53367), .ZN(n52844) );
  CLKNHSV0 U55938 ( .I(n48470), .ZN(n52843) );
  XOR2HSV0 U55939 ( .A1(n52844), .A2(n52843), .Z(n60044) );
  CLKNAND2HSV0 U55940 ( .A1(n56817), .A2(n56975), .ZN(n52846) );
  XOR2HSV0 U55941 ( .A1(n52846), .A2(n52845), .Z(\pe3/poht [31]) );
  NOR2HSV2 U55942 ( .A1(n29752), .A2(n46581), .ZN(n52850) );
  XOR2HSV0 U55943 ( .A1(n52847), .A2(n52848), .Z(n52849) );
  XOR2HSV0 U55944 ( .A1(n52850), .A2(n52849), .Z(pov4[31]) );
  CLKNAND2HSV1 U55945 ( .A1(n51688), .A2(n52558), .ZN(n52853) );
  NAND2HSV2 U55946 ( .A1(n53016), .A2(n52851), .ZN(n52852) );
  XOR2HSV0 U55947 ( .A1(n52853), .A2(n52852), .Z(\pe2/poht [31]) );
  CLKNAND2HSV1 U55948 ( .A1(n52854), .A2(n59777), .ZN(n52889) );
  CLKNAND2HSV1 U55949 ( .A1(n25831), .A2(n51686), .ZN(n52887) );
  CLKNAND2HSV0 U55950 ( .A1(n52918), .A2(n52855), .ZN(n52885) );
  INAND2HSV2 U55951 ( .A1(n47554), .B1(n52900), .ZN(n52883) );
  CLKNAND2HSV1 U55952 ( .A1(n52919), .A2(n52901), .ZN(n52879) );
  CLKNAND2HSV1 U55953 ( .A1(n52858), .A2(n52857), .ZN(n52861) );
  CLKNAND2HSV0 U55954 ( .A1(\pe2/aot [2]), .A2(n52859), .ZN(n52860) );
  XOR2HSV0 U55955 ( .A1(n52861), .A2(n52860), .Z(n52865) );
  CLKNAND2HSV1 U55956 ( .A1(n51803), .A2(n29736), .ZN(n52863) );
  NAND2HSV0 U55957 ( .A1(n52456), .A2(n52905), .ZN(n52862) );
  XOR2HSV0 U55958 ( .A1(n52863), .A2(n52862), .Z(n52864) );
  XOR2HSV0 U55959 ( .A1(n52865), .A2(n52864), .Z(n52877) );
  NAND2HSV0 U55960 ( .A1(n52867), .A2(n52866), .ZN(n52869) );
  NAND2HSV0 U55961 ( .A1(n59783), .A2(n53223), .ZN(n52868) );
  XOR2HSV0 U55962 ( .A1(n52869), .A2(n52868), .Z(n52875) );
  NOR2HSV0 U55963 ( .A1(n52871), .A2(n52870), .ZN(n52873) );
  AOI22HSV0 U55964 ( .A1(\pe2/aot [7]), .A2(n53226), .B1(n52951), .B2(n51532), 
        .ZN(n52872) );
  NOR2HSV2 U55965 ( .A1(n52873), .A2(n52872), .ZN(n52874) );
  XNOR2HSV1 U55966 ( .A1(n52875), .A2(n52874), .ZN(n52876) );
  XNOR2HSV1 U55967 ( .A1(n52877), .A2(n52876), .ZN(n52878) );
  XNOR2HSV1 U55968 ( .A1(n52879), .A2(n52878), .ZN(n52880) );
  XNOR2HSV1 U55969 ( .A1(n52881), .A2(n52880), .ZN(n52882) );
  XNOR2HSV1 U55970 ( .A1(n52883), .A2(n52882), .ZN(n52884) );
  XOR2HSV0 U55971 ( .A1(n52885), .A2(n52884), .Z(n52886) );
  XOR2HSV0 U55972 ( .A1(n52887), .A2(n52886), .Z(n52888) );
  XOR2HSV0 U55973 ( .A1(n52889), .A2(n52888), .Z(n52892) );
  NAND2HSV2 U55974 ( .A1(n52910), .A2(n52890), .ZN(n52891) );
  NAND2HSV0 U55975 ( .A1(n59794), .A2(\pe2/got [8]), .ZN(n52893) );
  XOR2HSV0 U55976 ( .A1(n52894), .A2(n52893), .Z(\pe2/poht [24]) );
  CLKNAND2HSV0 U55977 ( .A1(n59792), .A2(n53226), .ZN(n52899) );
  NAND2HSV2 U55978 ( .A1(n52902), .A2(n52901), .ZN(n52909) );
  CLKNAND2HSV1 U55979 ( .A1(\pe2/aot [2]), .A2(n53226), .ZN(n52904) );
  CLKNAND2HSV0 U55980 ( .A1(\pe2/aot [3]), .A2(n51532), .ZN(n52903) );
  XOR2HSV0 U55981 ( .A1(n52904), .A2(n52903), .Z(n52907) );
  CLKNAND2HSV1 U55982 ( .A1(n51547), .A2(n52905), .ZN(n52906) );
  XNOR2HSV1 U55983 ( .A1(n52907), .A2(n52906), .ZN(n52908) );
  XOR2HSV0 U55984 ( .A1(n52909), .A2(n52908), .Z(n52911) );
  CLKNAND2HSV0 U55985 ( .A1(n59351), .A2(n52558), .ZN(n52912) );
  XOR2HSV0 U55986 ( .A1(n52913), .A2(n52912), .Z(\pe2/poht [29]) );
  NAND2HSV2 U55987 ( .A1(n58655), .A2(n59235), .ZN(n52915) );
  NAND2HSV2 U55988 ( .A1(n58336), .A2(\pe6/aot [1]), .ZN(n52914) );
  XOR2HSV0 U55989 ( .A1(n52915), .A2(n52914), .Z(\pe6/poht [31]) );
  CLKNAND2HSV0 U55990 ( .A1(n52919), .A2(n44711), .ZN(n53085) );
  NAND2HSV0 U55991 ( .A1(n52920), .A2(n52416), .ZN(n53083) );
  NOR2HSV0 U55992 ( .A1(n52921), .A2(n45248), .ZN(n53081) );
  NAND2HSV0 U55993 ( .A1(n52923), .A2(n52922), .ZN(n53076) );
  NAND2HSV0 U55994 ( .A1(n52924), .A2(n39075), .ZN(n53072) );
  NAND2HSV0 U55995 ( .A1(n59506), .A2(n52925), .ZN(n53070) );
  CLKNAND2HSV0 U55996 ( .A1(n52926), .A2(n51796), .ZN(n53068) );
  CLKNAND2HSV1 U55997 ( .A1(n52927), .A2(n51964), .ZN(n53063) );
  NAND2HSV0 U55998 ( .A1(n52928), .A2(n51608), .ZN(n53061) );
  NAND2HSV0 U55999 ( .A1(n52172), .A2(n52929), .ZN(n53059) );
  NAND2HSV0 U56000 ( .A1(n52931), .A2(n52930), .ZN(n53054) );
  NAND2HSV0 U56001 ( .A1(n52932), .A2(\pe2/got [8]), .ZN(n53047) );
  NAND2HSV0 U56002 ( .A1(n52934), .A2(n52933), .ZN(n53045) );
  AOI22HSV0 U56003 ( .A1(n38558), .A2(n52935), .B1(n43961), .B2(n59636), .ZN(
        n52936) );
  AOI21HSV0 U56004 ( .A1(n52938), .A2(n52937), .B(n52936), .ZN(n52945) );
  NOR2HSV0 U56005 ( .A1(n52940), .A2(n52939), .ZN(n52943) );
  AOI22HSV0 U56006 ( .A1(n52941), .A2(n51803), .B1(n45033), .B2(n59976), .ZN(
        n52942) );
  NOR2HSV1 U56007 ( .A1(n52943), .A2(n52942), .ZN(n52944) );
  XOR2HSV0 U56008 ( .A1(n52945), .A2(n52944), .Z(n52949) );
  XOR2HSV0 U56009 ( .A1(n52947), .A2(n52946), .Z(n52948) );
  XNOR2HSV1 U56010 ( .A1(n52949), .A2(n52948), .ZN(n52961) );
  NAND2HSV0 U56011 ( .A1(n52951), .A2(n52950), .ZN(n52954) );
  NAND2HSV0 U56012 ( .A1(n59633), .A2(n52952), .ZN(n52953) );
  XOR2HSV0 U56013 ( .A1(n52954), .A2(n52953), .Z(n52959) );
  NAND2HSV0 U56014 ( .A1(n45295), .A2(\pe2/bq[6] ), .ZN(n52957) );
  NAND2HSV0 U56015 ( .A1(n52955), .A2(n43956), .ZN(n52956) );
  XOR2HSV0 U56016 ( .A1(n52957), .A2(n52956), .Z(n52958) );
  XOR2HSV0 U56017 ( .A1(n52959), .A2(n52958), .Z(n52960) );
  XOR2HSV0 U56018 ( .A1(n52961), .A2(n52960), .Z(n53031) );
  NAND2HSV0 U56019 ( .A1(n39052), .A2(n52962), .ZN(n52964) );
  NAND2HSV0 U56020 ( .A1(\pe2/aot [23]), .A2(n51997), .ZN(n52963) );
  XOR2HSV0 U56021 ( .A1(n52964), .A2(n52963), .Z(n52970) );
  NAND2HSV0 U56022 ( .A1(n52966), .A2(n52965), .ZN(n52968) );
  NAND2HSV0 U56023 ( .A1(\pe2/aot [19]), .A2(\pe2/bq[14] ), .ZN(n52967) );
  XOR2HSV0 U56024 ( .A1(n52968), .A2(n52967), .Z(n52969) );
  XOR2HSV0 U56025 ( .A1(n52970), .A2(n52969), .Z(n52980) );
  NAND2HSV0 U56026 ( .A1(n59968), .A2(n51805), .ZN(n52972) );
  NAND2HSV0 U56027 ( .A1(\pe2/got [1]), .A2(n36602), .ZN(n52971) );
  XOR2HSV0 U56028 ( .A1(n52972), .A2(n52971), .Z(n52978) );
  NAND2HSV0 U56029 ( .A1(n52456), .A2(n52973), .ZN(n52976) );
  NAND2HSV0 U56030 ( .A1(n52974), .A2(n52859), .ZN(n52975) );
  XOR2HSV0 U56031 ( .A1(n52976), .A2(n52975), .Z(n52977) );
  XOR2HSV0 U56032 ( .A1(n52978), .A2(n52977), .Z(n52979) );
  XOR2HSV0 U56033 ( .A1(n52980), .A2(n52979), .Z(n52983) );
  NAND2HSV2 U56034 ( .A1(n52981), .A2(n51932), .ZN(n52982) );
  XNOR2HSV1 U56035 ( .A1(n52983), .A2(n52982), .ZN(n53030) );
  NAND2HSV0 U56036 ( .A1(n51743), .A2(\pe2/bq[17] ), .ZN(n52986) );
  NAND2HSV0 U56037 ( .A1(n51759), .A2(n52984), .ZN(n52985) );
  XOR2HSV0 U56038 ( .A1(n52986), .A2(n52985), .Z(n52992) );
  NAND2HSV0 U56039 ( .A1(n59499), .A2(n52987), .ZN(n52990) );
  NAND2HSV0 U56040 ( .A1(n59974), .A2(n52988), .ZN(n52989) );
  XOR2HSV0 U56041 ( .A1(n52990), .A2(n52989), .Z(n52991) );
  XOR2HSV0 U56042 ( .A1(n52992), .A2(n52991), .Z(n53004) );
  NAND2HSV0 U56043 ( .A1(n52993), .A2(n36608), .ZN(n52997) );
  NAND2HSV0 U56044 ( .A1(n52995), .A2(n52994), .ZN(n52996) );
  XOR2HSV0 U56045 ( .A1(n52997), .A2(n52996), .Z(n53002) );
  NAND2HSV0 U56046 ( .A1(n52998), .A2(\pe2/bq[8] ), .ZN(n53000) );
  NAND2HSV0 U56047 ( .A1(\pe2/aot [22]), .A2(n52073), .ZN(n52999) );
  XOR2HSV0 U56048 ( .A1(n53000), .A2(n52999), .Z(n53001) );
  XOR2HSV0 U56049 ( .A1(n53002), .A2(n53001), .Z(n53003) );
  XOR2HSV0 U56050 ( .A1(n53004), .A2(n53003), .Z(n53028) );
  NAND2HSV0 U56051 ( .A1(n53005), .A2(\pe2/bq[21] ), .ZN(n53008) );
  NAND2HSV0 U56052 ( .A1(n59758), .A2(n53006), .ZN(n53007) );
  XOR2HSV0 U56053 ( .A1(n53008), .A2(n53007), .Z(n53013) );
  NOR2HSV0 U56054 ( .A1(n38655), .A2(n47511), .ZN(n53011) );
  NAND2HSV0 U56055 ( .A1(n53009), .A2(n52179), .ZN(n53010) );
  XOR2HSV0 U56056 ( .A1(n53011), .A2(n53010), .Z(n53012) );
  XOR2HSV0 U56057 ( .A1(n53013), .A2(n53012), .Z(n53026) );
  NAND2HSV0 U56058 ( .A1(\pe2/pq ), .A2(n53014), .ZN(n53018) );
  NAND2HSV0 U56059 ( .A1(n53016), .A2(n53015), .ZN(n53017) );
  XOR2HSV0 U56060 ( .A1(n53018), .A2(n53017), .Z(n53024) );
  AOI22HSV0 U56061 ( .A1(n53019), .A2(n45015), .B1(n38393), .B2(n52344), .ZN(
        n53020) );
  AOI21HSV0 U56062 ( .A1(n53022), .A2(n53021), .B(n53020), .ZN(n53023) );
  XNOR2HSV1 U56063 ( .A1(n53024), .A2(n53023), .ZN(n53025) );
  XNOR2HSV1 U56064 ( .A1(n53026), .A2(n53025), .ZN(n53027) );
  XNOR2HSV1 U56065 ( .A1(n53028), .A2(n53027), .ZN(n53029) );
  XOR3HSV2 U56066 ( .A1(n53031), .A2(n53030), .A3(n53029), .Z(n53037) );
  NAND2HSV0 U56067 ( .A1(n59684), .A2(n59984), .ZN(n53035) );
  NOR2HSV0 U56068 ( .A1(n53033), .A2(n53032), .ZN(n53034) );
  XNOR2HSV1 U56069 ( .A1(n53035), .A2(n53034), .ZN(n53036) );
  XOR2HSV0 U56070 ( .A1(n53037), .A2(n53036), .Z(n53040) );
  NAND2HSV0 U56071 ( .A1(n43928), .A2(n53038), .ZN(n53039) );
  XOR2HSV0 U56072 ( .A1(n53040), .A2(n53039), .Z(n53043) );
  NAND2HSV0 U56073 ( .A1(n44254), .A2(n53041), .ZN(n53042) );
  XNOR2HSV1 U56074 ( .A1(n53043), .A2(n53042), .ZN(n53044) );
  XNOR2HSV1 U56075 ( .A1(n53045), .A2(n53044), .ZN(n53046) );
  XNOR2HSV1 U56076 ( .A1(n53047), .A2(n53046), .ZN(n53049) );
  NAND2HSV0 U56077 ( .A1(n59766), .A2(\pe2/got [9]), .ZN(n53048) );
  XOR2HSV0 U56078 ( .A1(n53049), .A2(n53048), .Z(n53052) );
  NAND2HSV0 U56079 ( .A1(n53050), .A2(\pe2/got [10]), .ZN(n53051) );
  XNOR2HSV1 U56080 ( .A1(n53052), .A2(n53051), .ZN(n53053) );
  XNOR2HSV1 U56081 ( .A1(n53054), .A2(n53053), .ZN(n53058) );
  NAND2HSV0 U56082 ( .A1(n53056), .A2(n53055), .ZN(n53057) );
  XOR3HSV2 U56083 ( .A1(n53059), .A2(n53058), .A3(n53057), .Z(n53060) );
  XNOR2HSV1 U56084 ( .A1(n53061), .A2(n53060), .ZN(n53062) );
  XNOR2HSV1 U56085 ( .A1(n53063), .A2(n53062), .ZN(n53067) );
  NOR2HSV0 U56086 ( .A1(n53065), .A2(n53064), .ZN(n53066) );
  XOR3HSV2 U56087 ( .A1(n53068), .A2(n53067), .A3(n53066), .Z(n53069) );
  XNOR2HSV1 U56088 ( .A1(n53070), .A2(n53069), .ZN(n53071) );
  XNOR2HSV1 U56089 ( .A1(n53072), .A2(n53071), .ZN(n53074) );
  NAND2HSV0 U56090 ( .A1(n59361), .A2(n52042), .ZN(n53073) );
  XNOR2HSV1 U56091 ( .A1(n53074), .A2(n53073), .ZN(n53075) );
  XNOR2HSV1 U56092 ( .A1(n53076), .A2(n53075), .ZN(n53080) );
  CLKNAND2HSV0 U56093 ( .A1(n53078), .A2(n53077), .ZN(n53079) );
  XOR3HSV2 U56094 ( .A1(n53081), .A2(n53080), .A3(n53079), .Z(n53082) );
  XOR2HSV0 U56095 ( .A1(n53083), .A2(n53082), .Z(n53084) );
  XNOR2HSV1 U56096 ( .A1(n53085), .A2(n53084), .ZN(n53090) );
  NAND2HSV2 U56097 ( .A1(n53087), .A2(n53086), .ZN(n53089) );
  CLKNAND2HSV0 U56098 ( .A1(n59929), .A2(n44944), .ZN(n53088) );
  XOR3HSV2 U56099 ( .A1(n53090), .A2(n53089), .A3(n53088), .Z(n53091) );
  INAND2HSV0 U56100 ( .A1(n53098), .B1(n53097), .ZN(n53099) );
  XOR2HSV0 U56101 ( .A1(n53100), .A2(n53099), .Z(po2) );
  NOR2HSV1 U56102 ( .A1(n53104), .A2(n53103), .ZN(n53105) );
  CLKNAND2HSV1 U56103 ( .A1(n53106), .A2(n53105), .ZN(n53183) );
  CLKNAND2HSV0 U56104 ( .A1(n59031), .A2(n59024), .ZN(n53181) );
  CLKNHSV0 U56105 ( .I(n32596), .ZN(n53108) );
  INAND2HSV2 U56106 ( .A1(n53108), .B1(n53107), .ZN(n53179) );
  CLKNAND2HSV1 U56107 ( .A1(n58385), .A2(n58810), .ZN(n53177) );
  CLKNAND2HSV0 U56108 ( .A1(n53109), .A2(n59180), .ZN(n53175) );
  CLKNAND2HSV1 U56109 ( .A1(n58480), .A2(n49742), .ZN(n53171) );
  CLKNAND2HSV0 U56110 ( .A1(n58448), .A2(n58658), .ZN(n53167) );
  CLKNAND2HSV1 U56111 ( .A1(n59680), .A2(n59182), .ZN(n53165) );
  CLKNAND2HSV0 U56112 ( .A1(n53111), .A2(n58513), .ZN(n53161) );
  NAND2HSV0 U56113 ( .A1(n53112), .A2(n58478), .ZN(n53159) );
  CLKNAND2HSV0 U56114 ( .A1(n53113), .A2(n58479), .ZN(n53157) );
  NAND2HSV0 U56115 ( .A1(n53114), .A2(n58527), .ZN(n53155) );
  NAND2HSV0 U56116 ( .A1(n49667), .A2(n58403), .ZN(n53151) );
  NAND2HSV0 U56117 ( .A1(n59273), .A2(n53115), .ZN(n53117) );
  NAND2HSV0 U56118 ( .A1(n59277), .A2(n59088), .ZN(n53116) );
  XOR2HSV0 U56119 ( .A1(n53117), .A2(n53116), .Z(n53121) );
  NAND2HSV0 U56120 ( .A1(\pe6/bq[14] ), .A2(\pe6/aot [5]), .ZN(n53118) );
  XOR2HSV0 U56121 ( .A1(n53119), .A2(n53118), .Z(n53120) );
  XOR2HSV0 U56122 ( .A1(n53121), .A2(n53120), .Z(n53149) );
  NOR2HSV0 U56123 ( .A1(n48047), .A2(n58530), .ZN(n53123) );
  CLKNAND2HSV0 U56124 ( .A1(n59041), .A2(\pe6/aot [17]), .ZN(n53122) );
  XOR2HSV0 U56125 ( .A1(n53123), .A2(n53122), .Z(n53127) );
  CLKNHSV0 U56126 ( .I(n58382), .ZN(n53125) );
  NOR2HSV0 U56127 ( .A1(n58984), .A2(n44396), .ZN(n59106) );
  AOI22HSV1 U56128 ( .A1(n58833), .A2(\pe6/aot [3]), .B1(n58842), .B2(n59062), 
        .ZN(n53124) );
  AOI21HSV2 U56129 ( .A1(n53125), .A2(n59106), .B(n53124), .ZN(n53126) );
  XNOR2HSV1 U56130 ( .A1(n53127), .A2(n53126), .ZN(n53131) );
  XOR2HSV0 U56131 ( .A1(n53129), .A2(n53128), .Z(n53130) );
  XNOR2HSV1 U56132 ( .A1(n53131), .A2(n53130), .ZN(n53148) );
  NAND2HSV0 U56133 ( .A1(n58976), .A2(\pe6/aot [7]), .ZN(n53133) );
  NAND2HSV0 U56134 ( .A1(n59246), .A2(\pe6/aot [11]), .ZN(n53132) );
  XOR2HSV0 U56135 ( .A1(n53133), .A2(n53132), .Z(n53138) );
  CLKNAND2HSV0 U56136 ( .A1(n59265), .A2(n53134), .ZN(n53136) );
  NAND2HSV0 U56137 ( .A1(n44336), .A2(n58495), .ZN(n53135) );
  XOR2HSV0 U56138 ( .A1(n53136), .A2(n53135), .Z(n53137) );
  XOR2HSV0 U56139 ( .A1(n53138), .A2(n53137), .Z(n53146) );
  NAND2HSV0 U56140 ( .A1(n48044), .A2(\pe6/aot [10]), .ZN(n53140) );
  NAND2HSV0 U56141 ( .A1(n33023), .A2(\pe6/aot [1]), .ZN(n53139) );
  XOR2HSV0 U56142 ( .A1(n53140), .A2(n53139), .Z(n53144) );
  NAND2HSV0 U56143 ( .A1(n32982), .A2(n59260), .ZN(n53142) );
  NAND2HSV0 U56144 ( .A1(n48038), .A2(\pe6/aot [13]), .ZN(n53141) );
  XOR2HSV0 U56145 ( .A1(n53142), .A2(n53141), .Z(n53143) );
  XOR2HSV0 U56146 ( .A1(n53144), .A2(n53143), .Z(n53145) );
  XOR2HSV0 U56147 ( .A1(n53146), .A2(n53145), .Z(n53147) );
  XOR3HSV2 U56148 ( .A1(n53149), .A2(n53148), .A3(n53147), .Z(n53150) );
  XNOR2HSV1 U56149 ( .A1(n53151), .A2(n53150), .ZN(n53153) );
  NAND2HSV0 U56150 ( .A1(n58901), .A2(n58724), .ZN(n53152) );
  XNOR2HSV1 U56151 ( .A1(n53153), .A2(n53152), .ZN(n53154) );
  XOR2HSV0 U56152 ( .A1(n53155), .A2(n53154), .Z(n53156) );
  XNOR2HSV1 U56153 ( .A1(n53157), .A2(n53156), .ZN(n53158) );
  XNOR2HSV1 U56154 ( .A1(n53159), .A2(n53158), .ZN(n53160) );
  XNOR2HSV1 U56155 ( .A1(n53161), .A2(n53160), .ZN(n53163) );
  CLKNAND2HSV0 U56156 ( .A1(n59915), .A2(n58709), .ZN(n53162) );
  XNOR2HSV1 U56157 ( .A1(n53163), .A2(n53162), .ZN(n53164) );
  XNOR2HSV1 U56158 ( .A1(n53165), .A2(n53164), .ZN(n53166) );
  XNOR2HSV1 U56159 ( .A1(n53167), .A2(n53166), .ZN(n53169) );
  NAND2HSV0 U56160 ( .A1(n59677), .A2(n44393), .ZN(n53168) );
  XOR2HSV0 U56161 ( .A1(n53169), .A2(n53168), .Z(n53170) );
  XNOR2HSV1 U56162 ( .A1(n53171), .A2(n53170), .ZN(n53174) );
  NAND2HSV0 U56163 ( .A1(n53172), .A2(n58711), .ZN(n53173) );
  XOR3HSV2 U56164 ( .A1(n53175), .A2(n53174), .A3(n53173), .Z(n53176) );
  XNOR2HSV1 U56165 ( .A1(n53177), .A2(n53176), .ZN(n53178) );
  XNOR2HSV1 U56166 ( .A1(n53179), .A2(n53178), .ZN(n53180) );
  XOR2HSV0 U56167 ( .A1(n53181), .A2(n53180), .Z(n53182) );
  XNOR2HSV1 U56168 ( .A1(n53183), .A2(n53182), .ZN(n53184) );
  XOR2HSV0 U56169 ( .A1(n53185), .A2(n53184), .Z(\pe6/poht [14]) );
  INHSV2 U56170 ( .I(n55185), .ZN(n54988) );
  NAND2HSV2 U56171 ( .A1(n59373), .A2(n54988), .ZN(n53186) );
  XOR2HSV0 U56172 ( .A1(n53187), .A2(n53186), .Z(\pe1/poht [31]) );
  AOI21HSV1 U56173 ( .A1(n53188), .A2(n39239), .B(n48625), .ZN(n53189) );
  OAI21HSV0 U56174 ( .A1(n29761), .A2(n53190), .B(n53189), .ZN(n53194) );
  NAND2HSV2 U56175 ( .A1(n51182), .A2(\pe5/bq[2] ), .ZN(n53192) );
  CLKNAND2HSV1 U56176 ( .A1(n59866), .A2(n53199), .ZN(n53191) );
  XOR2HSV0 U56177 ( .A1(n53192), .A2(n53191), .Z(n53193) );
  XOR2HSV0 U56178 ( .A1(n53194), .A2(n53193), .Z(n53196) );
  NAND2HSV0 U56179 ( .A1(n53197), .A2(n53210), .ZN(n53195) );
  XOR2HSV0 U56180 ( .A1(n53196), .A2(n53195), .Z(\pe5/poht [30]) );
  NAND2HSV2 U56181 ( .A1(n29779), .A2(n51362), .ZN(n53207) );
  CLKNAND2HSV1 U56182 ( .A1(\pe5/aot [3]), .A2(n53199), .ZN(n53202) );
  CLKNAND2HSV1 U56183 ( .A1(n51339), .A2(n53200), .ZN(n53201) );
  XOR2HSV0 U56184 ( .A1(n53202), .A2(n53201), .Z(n53205) );
  NAND2HSV2 U56185 ( .A1(n53203), .A2(\pe5/bq[2] ), .ZN(n53204) );
  XNOR2HSV1 U56186 ( .A1(n53205), .A2(n53204), .ZN(n53206) );
  XOR2HSV0 U56187 ( .A1(n53207), .A2(n53206), .Z(n53208) );
  NAND2HSV0 U56188 ( .A1(n53211), .A2(n53210), .ZN(n53212) );
  XOR2HSV0 U56189 ( .A1(n53213), .A2(n53212), .Z(\pe5/poht [29]) );
  MUX2HSV2 U56190 ( .I0(bo6[2]), .I1(\pe6/bq[2] ), .S(n53214), .Z(n59539) );
  MUX2HSV2 U56191 ( .I0(bo5[11]), .I1(\pe5/bq[11] ), .S(n53215), .Z(n59541) );
  MUX2HSV2 U56192 ( .I0(bo5[10]), .I1(n53216), .S(n53215), .Z(n59542) );
  MUX2HSV2 U56193 ( .I0(bo5[2]), .I1(\pe5/bq[2] ), .S(n53215), .Z(n59544) );
  MUX2HSV2 U56194 ( .I0(bo4[21]), .I1(n33969), .S(n34496), .Z(n59545) );
  MUX2HSV2 U56195 ( .I0(bo4[17]), .I1(n57926), .S(n48073), .Z(n59546) );
  MUX2HSV2 U56196 ( .I0(bo4[14]), .I1(n58069), .S(n48073), .Z(n59547) );
  MUX2HSV2 U56197 ( .I0(bo4[13]), .I1(n58127), .S(n53220), .Z(n59548) );
  MUX2HSV2 U56198 ( .I0(bo4[11]), .I1(\pe4/bq[11] ), .S(n48082), .Z(n59549) );
  MUX2HSV2 U56199 ( .I0(bo4[10]), .I1(n58116), .S(n48073), .Z(n59550) );
  MUX2HSV2 U56200 ( .I0(bo4[9]), .I1(n58113), .S(n48073), .Z(n59551) );
  MUX2HSV2 U56201 ( .I0(bo4[4]), .I1(n57498), .S(n47659), .Z(n59552) );
  MUX2HSV2 U56202 ( .I0(bo4[2]), .I1(\pe4/bq[2] ), .S(n34054), .Z(n59553) );
  MUX2HSV2 U56203 ( .I0(bo3[24]), .I1(n55872), .S(n46124), .Z(n59557) );
  MUX2HSV2 U56204 ( .I0(bo3[7]), .I1(\pe3/bq[7] ), .S(n53221), .Z(n59560) );
  MUX2HSV2 U56205 ( .I0(bo2[12]), .I1(\pe2/bq[12] ), .S(n46619), .Z(n59564) );
  MUX2HSV2 U56206 ( .I0(bo2[8]), .I1(n53223), .S(n53222), .Z(n59565) );
  MUX2HSV2 U56207 ( .I0(bo2[5]), .I1(n52857), .S(n53224), .Z(n59566) );
  MUX2HSV2 U56208 ( .I0(bo2[2]), .I1(n53226), .S(n53225), .Z(n59567) );
  CLKNAND2HSV1 U56209 ( .A1(n56341), .A2(n56177), .ZN(n53274) );
  CLKNAND2HSV0 U56210 ( .A1(n55822), .A2(n56855), .ZN(n53272) );
  CLKNHSV0 U56211 ( .I(n53227), .ZN(n56736) );
  CLKNAND2HSV0 U56212 ( .A1(n56736), .A2(n56266), .ZN(n53270) );
  CLKNAND2HSV0 U56213 ( .A1(n56622), .A2(n56779), .ZN(n53268) );
  NAND2HSV0 U56214 ( .A1(n56737), .A2(n56623), .ZN(n53266) );
  CLKNAND2HSV0 U56215 ( .A1(n56684), .A2(n59500), .ZN(n53264) );
  CLKNAND2HSV0 U56216 ( .A1(n56624), .A2(n56782), .ZN(n53260) );
  NAND2HSV0 U56217 ( .A1(n59821), .A2(\pe3/got [1]), .ZN(n53258) );
  CLKNAND2HSV0 U56218 ( .A1(n56378), .A2(n55857), .ZN(n53231) );
  CLKNHSV0 U56219 ( .I(n53229), .ZN(n56695) );
  NAND2HSV0 U56220 ( .A1(n56695), .A2(\pe3/bq[4] ), .ZN(n53230) );
  XOR2HSV0 U56221 ( .A1(n53231), .A2(n53230), .Z(n53236) );
  NAND2HSV0 U56222 ( .A1(n56221), .A2(n53232), .ZN(n53234) );
  NAND2HSV0 U56223 ( .A1(n59511), .A2(n56094), .ZN(n53233) );
  XOR2HSV0 U56224 ( .A1(n53234), .A2(n53233), .Z(n53235) );
  XOR2HSV0 U56225 ( .A1(n53236), .A2(n53235), .Z(n53244) );
  NAND2HSV0 U56226 ( .A1(n56423), .A2(n56832), .ZN(n53238) );
  NAND2HSV0 U56227 ( .A1(n56911), .A2(n56627), .ZN(n53237) );
  XOR2HSV0 U56228 ( .A1(n53238), .A2(n53237), .Z(n53242) );
  NOR2HSV0 U56229 ( .A1(n47447), .A2(n49258), .ZN(n53240) );
  CLKNAND2HSV0 U56230 ( .A1(\pe3/aot [2]), .A2(n48499), .ZN(n53239) );
  XOR2HSV0 U56231 ( .A1(n53240), .A2(n53239), .Z(n53241) );
  XOR2HSV0 U56232 ( .A1(n53242), .A2(n53241), .Z(n53243) );
  XOR2HSV0 U56233 ( .A1(n53244), .A2(n53243), .Z(n53256) );
  NAND2HSV0 U56234 ( .A1(n56074), .A2(\pe3/bq[11] ), .ZN(n56563) );
  NAND2HSV0 U56235 ( .A1(n56439), .A2(n56507), .ZN(n56635) );
  NOR2HSV0 U56236 ( .A1(n56563), .A2(n56635), .ZN(n53246) );
  AOI22HSV0 U56237 ( .A1(n56788), .A2(n56507), .B1(\pe3/bq[11] ), .B2(n59816), 
        .ZN(n53245) );
  NOR2HSV1 U56238 ( .A1(n53246), .A2(n53245), .ZN(n53254) );
  NAND2HSV0 U56239 ( .A1(n56197), .A2(n56867), .ZN(n53248) );
  NAND2HSV0 U56240 ( .A1(\pe3/aot [8]), .A2(\pe3/bq[8] ), .ZN(n53247) );
  XOR2HSV0 U56241 ( .A1(n53248), .A2(n53247), .Z(n53253) );
  NOR2HSV0 U56242 ( .A1(n56382), .A2(n50722), .ZN(n56578) );
  NAND2HSV0 U56243 ( .A1(n53249), .A2(n55975), .ZN(n56116) );
  CLKNAND2HSV1 U56244 ( .A1(n53250), .A2(n56529), .ZN(n56940) );
  CLKNAND2HSV0 U56245 ( .A1(n56188), .A2(n56505), .ZN(n56649) );
  XOR2HSV0 U56246 ( .A1(n53251), .A2(n56649), .Z(n53252) );
  XOR3HSV2 U56247 ( .A1(n53254), .A2(n53253), .A3(n53252), .Z(n53255) );
  XNOR2HSV1 U56248 ( .A1(n53256), .A2(n53255), .ZN(n53257) );
  XNOR2HSV1 U56249 ( .A1(n53258), .A2(n53257), .ZN(n53259) );
  XNOR2HSV1 U56250 ( .A1(n53260), .A2(n53259), .ZN(n53262) );
  NAND2HSV0 U56251 ( .A1(n43463), .A2(n56735), .ZN(n53261) );
  XNOR2HSV1 U56252 ( .A1(n53262), .A2(n53261), .ZN(n53263) );
  XNOR2HSV1 U56253 ( .A1(n53264), .A2(n53263), .ZN(n53265) );
  XNOR2HSV1 U56254 ( .A1(n53266), .A2(n53265), .ZN(n53267) );
  XNOR2HSV1 U56255 ( .A1(n53268), .A2(n53267), .ZN(n53269) );
  XNOR2HSV1 U56256 ( .A1(n53270), .A2(n53269), .ZN(n53271) );
  XNOR2HSV1 U56257 ( .A1(n53272), .A2(n53271), .ZN(n53273) );
  XNOR2HSV1 U56258 ( .A1(n53274), .A2(n53273), .ZN(n53275) );
  XNOR2HSV1 U56259 ( .A1(n53278), .A2(n53277), .ZN(n53281) );
  NAND2HSV2 U56260 ( .A1(n56907), .A2(n56618), .ZN(n53280) );
  NAND2HSV2 U56261 ( .A1(n56058), .A2(n56419), .ZN(n53283) );
  CLKNAND2HSV1 U56262 ( .A1(n56900), .A2(\pe3/got [14]), .ZN(n53282) );
  XOR3HSV2 U56263 ( .A1(n53284), .A2(n53283), .A3(n53282), .Z(\pe3/poht [17])
         );
  CLKNAND2HSV1 U56264 ( .A1(n29778), .A2(n53285), .ZN(n53357) );
  CLKNAND2HSV1 U56265 ( .A1(n53287), .A2(n53286), .ZN(n53355) );
  CLKNAND2HSV1 U56266 ( .A1(n53288), .A2(n48167), .ZN(n53353) );
  CLKNAND2HSV0 U56267 ( .A1(n53290), .A2(n53289), .ZN(n53348) );
  CLKNAND2HSV0 U56268 ( .A1(n53291), .A2(n50698), .ZN(n53343) );
  NOR2HSV0 U56269 ( .A1(n53293), .A2(n53292), .ZN(n53337) );
  CLKNAND2HSV1 U56270 ( .A1(n53294), .A2(n52579), .ZN(n53333) );
  CLKNAND2HSV1 U56271 ( .A1(n59882), .A2(\pe5/got [2]), .ZN(n53331) );
  NAND2HSV0 U56272 ( .A1(n59517), .A2(n51362), .ZN(n53329) );
  CLKNAND2HSV0 U56273 ( .A1(n53295), .A2(\pe5/bq[11] ), .ZN(n53298) );
  CLKNAND2HSV1 U56274 ( .A1(n53296), .A2(n51307), .ZN(n53297) );
  XOR2HSV0 U56275 ( .A1(n53298), .A2(n53297), .Z(n53303) );
  NAND2HSV2 U56276 ( .A1(\pe5/aot [4]), .A2(\pe5/bq[13] ), .ZN(n53301) );
  NAND2HSV0 U56277 ( .A1(n53299), .A2(n51373), .ZN(n53300) );
  XOR2HSV0 U56278 ( .A1(n53301), .A2(n53300), .Z(n53302) );
  XOR2HSV0 U56279 ( .A1(n53303), .A2(n53302), .Z(n53313) );
  CLKNAND2HSV0 U56280 ( .A1(n51313), .A2(\pe5/bq[7] ), .ZN(n53306) );
  NAND2HSV0 U56281 ( .A1(n53304), .A2(n53216), .ZN(n53305) );
  XOR2HSV0 U56282 ( .A1(n53306), .A2(n53305), .Z(n53311) );
  NAND2HSV0 U56283 ( .A1(\pe5/aot [13]), .A2(n53307), .ZN(n53309) );
  NAND2HSV0 U56284 ( .A1(n59943), .A2(\pe5/bq[2] ), .ZN(n53308) );
  XOR2HSV0 U56285 ( .A1(n53309), .A2(n53308), .Z(n53310) );
  XOR2HSV0 U56286 ( .A1(n53311), .A2(n53310), .Z(n53312) );
  XOR2HSV0 U56287 ( .A1(n53313), .A2(n53312), .Z(n53327) );
  CLKNAND2HSV1 U56288 ( .A1(\pe5/aot [14]), .A2(n40226), .ZN(n53316) );
  NAND2HSV0 U56289 ( .A1(n51419), .A2(n53314), .ZN(n53315) );
  XOR2HSV0 U56290 ( .A1(n53316), .A2(n53315), .Z(n53320) );
  NAND2HSV0 U56291 ( .A1(n39887), .A2(n48760), .ZN(n53318) );
  NAND2HSV0 U56292 ( .A1(\pe5/aot [16]), .A2(n53199), .ZN(n53317) );
  XOR2HSV0 U56293 ( .A1(n53318), .A2(n53317), .Z(n53319) );
  XOR2HSV0 U56294 ( .A1(n53320), .A2(n53319), .Z(n53325) );
  XOR2HSV0 U56295 ( .A1(n53325), .A2(n53324), .Z(n53326) );
  XOR2HSV0 U56296 ( .A1(n53327), .A2(n53326), .Z(n53328) );
  XNOR2HSV1 U56297 ( .A1(n53329), .A2(n53328), .ZN(n53330) );
  XNOR2HSV1 U56298 ( .A1(n53331), .A2(n53330), .ZN(n53332) );
  XNOR2HSV1 U56299 ( .A1(n53333), .A2(n53332), .ZN(n53335) );
  CLKNAND2HSV0 U56300 ( .A1(n52653), .A2(n51418), .ZN(n53334) );
  XNOR2HSV1 U56301 ( .A1(n53335), .A2(n53334), .ZN(n53336) );
  XNOR2HSV1 U56302 ( .A1(n53337), .A2(n53336), .ZN(n53341) );
  CLKNAND2HSV1 U56303 ( .A1(n53338), .A2(n51200), .ZN(n53340) );
  NOR2HSV2 U56304 ( .A1(n51360), .A2(n46978), .ZN(n53339) );
  XOR3HSV2 U56305 ( .A1(n53341), .A2(n53340), .A3(n53339), .Z(n53342) );
  XNOR2HSV1 U56306 ( .A1(n53343), .A2(n53342), .ZN(n53346) );
  CLKNAND2HSV0 U56307 ( .A1(n53344), .A2(n59891), .ZN(n53345) );
  XNOR2HSV1 U56308 ( .A1(n53346), .A2(n53345), .ZN(n53347) );
  XNOR2HSV1 U56309 ( .A1(n53348), .A2(n53347), .ZN(n53351) );
  CLKNAND2HSV0 U56310 ( .A1(n59535), .A2(n53349), .ZN(n53350) );
  XNOR2HSV1 U56311 ( .A1(n53351), .A2(n53350), .ZN(n53352) );
  XNOR2HSV1 U56312 ( .A1(n53353), .A2(n53352), .ZN(n53354) );
  XNOR2HSV1 U56313 ( .A1(n53355), .A2(n53354), .ZN(n53356) );
  XOR2HSV0 U56314 ( .A1(n53357), .A2(n53356), .Z(n53366) );
  NAND2HSV2 U56315 ( .A1(n53359), .A2(n51015), .ZN(n53360) );
  NOR2HSV2 U56316 ( .A1(n51013), .A2(n53360), .ZN(n53365) );
  AND2HSV2 U56317 ( .A1(n53361), .A2(n39881), .Z(n53362) );
  CLKNAND2HSV1 U56318 ( .A1(n53363), .A2(n53362), .ZN(n53364) );
  XOR3HSV2 U56319 ( .A1(n53366), .A2(n53365), .A3(n53364), .Z(\pe5/poht [16])
         );
  NAND2HSV0 U56320 ( .A1(n56180), .A2(n46107), .ZN(n53370) );
  XOR2HSV0 U56321 ( .A1(n53370), .A2(n53369), .Z(n53371) );
  XOR2HSV0 U56322 ( .A1(n53372), .A2(n53371), .Z(n60089) );
  XNOR2HSV0 U56323 ( .A1(n53377), .A2(n53376), .ZN(n53379) );
  XOR2HSV0 U56324 ( .A1(n53379), .A2(n53378), .Z(n60087) );
  NAND2HSV0 U56325 ( .A1(n52934), .A2(n44709), .ZN(n53380) );
  XOR2HSV0 U56326 ( .A1(n53380), .A2(n53381), .Z(n60099) );
  CLKNAND2HSV1 U56327 ( .A1(n53382), .A2(n47997), .ZN(n53383) );
  XOR2HSV0 U56328 ( .A1(n53383), .A2(n39113), .Z(n60094) );
  XOR2HSV0 U56329 ( .A1(n53388), .A2(n53387), .Z(pov2[28]) );
  INHSV2 U56330 ( .I(n53791), .ZN(n55541) );
  CLKNAND2HSV0 U56331 ( .A1(n55541), .A2(n40873), .ZN(n53510) );
  CLKNAND2HSV0 U56332 ( .A1(n59489), .A2(n59374), .ZN(n53508) );
  CLKNAND2HSV0 U56333 ( .A1(n53792), .A2(n53520), .ZN(n53502) );
  CLKNAND2HSV1 U56334 ( .A1(n53656), .A2(n53655), .ZN(n55341) );
  CLKNAND2HSV0 U56335 ( .A1(n55341), .A2(n53390), .ZN(n53498) );
  NAND2HSV0 U56336 ( .A1(n55229), .A2(\pe1/got [21]), .ZN(n53496) );
  NAND2HSV0 U56337 ( .A1(n53521), .A2(\pe1/got [19]), .ZN(n53492) );
  NOR2HSV0 U56338 ( .A1(n53391), .A2(n54248), .ZN(n53490) );
  NAND2HSV0 U56339 ( .A1(n53522), .A2(n54135), .ZN(n53488) );
  NAND2HSV0 U56340 ( .A1(n53392), .A2(n54161), .ZN(n53486) );
  NOR2HSV0 U56341 ( .A1(n54454), .A2(n54039), .ZN(n53484) );
  CLKNHSV0 U56342 ( .I(n53393), .ZN(n53794) );
  INHSV2 U56343 ( .I(n53794), .ZN(n54731) );
  NOR2HSV0 U56344 ( .A1(n54731), .A2(n54957), .ZN(n53482) );
  NAND2HSV0 U56345 ( .A1(n54557), .A2(n55087), .ZN(n53479) );
  NAND2HSV0 U56346 ( .A1(n54041), .A2(n54970), .ZN(n53477) );
  NOR2HSV0 U56347 ( .A1(n41301), .A2(n55163), .ZN(n53472) );
  CLKNHSV1 U56348 ( .I(n55019), .ZN(n54894) );
  NAND2HSV0 U56349 ( .A1(n41332), .A2(n54894), .ZN(n53468) );
  NAND2HSV0 U56350 ( .A1(n42360), .A2(n53863), .ZN(n53462) );
  NAND2HSV0 U56351 ( .A1(n53979), .A2(n54104), .ZN(n53460) );
  NAND2HSV0 U56352 ( .A1(\pe1/aot [16]), .A2(n48380), .ZN(n53395) );
  NAND2HSV0 U56353 ( .A1(n59619), .A2(\pe1/bq[27] ), .ZN(n53394) );
  XOR2HSV0 U56354 ( .A1(n53395), .A2(n53394), .Z(n53399) );
  NAND2HSV0 U56355 ( .A1(n54303), .A2(n40557), .ZN(n53397) );
  NAND2HSV0 U56356 ( .A1(n59987), .A2(n55352), .ZN(n53396) );
  XOR2HSV0 U56357 ( .A1(n53397), .A2(n53396), .Z(n53398) );
  XOR2HSV0 U56358 ( .A1(n53399), .A2(n53398), .Z(n53407) );
  NAND2HSV0 U56359 ( .A1(n41768), .A2(\pe1/bq[11] ), .ZN(n53401) );
  NAND2HSV0 U56360 ( .A1(n53812), .A2(n42092), .ZN(n53400) );
  XOR2HSV0 U56361 ( .A1(n53401), .A2(n53400), .Z(n53405) );
  BUFHSV2 U56362 ( .I(n53936), .Z(n54662) );
  NAND2HSV0 U56363 ( .A1(n54662), .A2(n54565), .ZN(n53403) );
  NAND2HSV0 U56364 ( .A1(n54500), .A2(n54179), .ZN(n53402) );
  XOR2HSV0 U56365 ( .A1(n53403), .A2(n53402), .Z(n53404) );
  XOR2HSV0 U56366 ( .A1(n53405), .A2(n53404), .Z(n53406) );
  XOR2HSV0 U56367 ( .A1(n53407), .A2(n53406), .Z(n53428) );
  NAND2HSV0 U56368 ( .A1(n54364), .A2(n42373), .ZN(n53408) );
  XOR2HSV0 U56369 ( .A1(n53409), .A2(n53408), .Z(n53426) );
  NOR2HSV0 U56370 ( .A1(n55504), .A2(n41622), .ZN(n53659) );
  NOR2HSV0 U56371 ( .A1(n55524), .A2(n53410), .ZN(n53971) );
  NOR2HSV0 U56372 ( .A1(n55504), .A2(n53410), .ZN(n53661) );
  AOI21HSV0 U56373 ( .A1(n59373), .A2(n53411), .B(n53661), .ZN(n53412) );
  AOI21HSV1 U56374 ( .A1(n53659), .A2(n53971), .B(n53412), .ZN(n53417) );
  CLKNHSV0 U56375 ( .I(n55185), .ZN(n54063) );
  NAND2HSV0 U56376 ( .A1(\pe1/aot [22]), .A2(n54063), .ZN(n54641) );
  NOR2HSV0 U56377 ( .A1(n53413), .A2(n54641), .ZN(n53415) );
  CLKNHSV0 U56378 ( .I(n55185), .ZN(n54292) );
  AOI22HSV0 U56379 ( .A1(n59985), .A2(n54292), .B1(n54078), .B2(\pe1/bq[9] ), 
        .ZN(n53414) );
  NOR2HSV1 U56380 ( .A1(n53415), .A2(n53414), .ZN(n53416) );
  XOR2HSV0 U56381 ( .A1(n53417), .A2(n53416), .Z(n53425) );
  CLKNHSV0 U56382 ( .I(n54829), .ZN(n54497) );
  NAND2HSV0 U56383 ( .A1(n54497), .A2(n53571), .ZN(n53419) );
  NAND2HSV0 U56384 ( .A1(n55496), .A2(n41623), .ZN(n53418) );
  XOR2HSV0 U56385 ( .A1(n53419), .A2(n53418), .Z(n53423) );
  NAND2HSV0 U56386 ( .A1(n53954), .A2(n53798), .ZN(n53421) );
  NAND2HSV0 U56387 ( .A1(n54307), .A2(n55394), .ZN(n53420) );
  XOR2HSV0 U56388 ( .A1(n53421), .A2(n53420), .Z(n53422) );
  XOR2HSV0 U56389 ( .A1(n53423), .A2(n53422), .Z(n53424) );
  XOR3HSV2 U56390 ( .A1(n53426), .A2(n53425), .A3(n53424), .Z(n53427) );
  XOR2HSV0 U56391 ( .A1(n53428), .A2(n53427), .Z(n53457) );
  NAND2HSV0 U56392 ( .A1(\pe1/aot [15]), .A2(n54836), .ZN(n53430) );
  NAND2HSV0 U56393 ( .A1(n53538), .A2(n55110), .ZN(n53429) );
  XOR2HSV0 U56394 ( .A1(n53430), .A2(n53429), .Z(n53434) );
  NAND2HSV0 U56395 ( .A1(\pe1/aot [14]), .A2(n54995), .ZN(n53432) );
  NAND2HSV0 U56396 ( .A1(n55452), .A2(n54048), .ZN(n53431) );
  XOR2HSV0 U56397 ( .A1(n53432), .A2(n53431), .Z(n53433) );
  XOR2HSV0 U56398 ( .A1(n53434), .A2(n53433), .Z(n53442) );
  NAND2HSV2 U56399 ( .A1(n59986), .A2(n55544), .ZN(n53436) );
  NAND2HSV0 U56400 ( .A1(n53717), .A2(\pe1/bq[21] ), .ZN(n53435) );
  XOR2HSV0 U56401 ( .A1(n53436), .A2(n53435), .Z(n53440) );
  NAND2HSV0 U56402 ( .A1(n54578), .A2(n53578), .ZN(n53438) );
  NAND2HSV0 U56403 ( .A1(n59990), .A2(\pe1/bq[18] ), .ZN(n53437) );
  XOR2HSV0 U56404 ( .A1(n53438), .A2(n53437), .Z(n53439) );
  XNOR2HSV1 U56405 ( .A1(n53440), .A2(n53439), .ZN(n53441) );
  XNOR2HSV1 U56406 ( .A1(n53442), .A2(n53441), .ZN(n53455) );
  NAND2HSV0 U56407 ( .A1(n59590), .A2(n59755), .ZN(n53453) );
  NAND2HSV2 U56408 ( .A1(n54978), .A2(n54289), .ZN(n55306) );
  NOR2HSV0 U56409 ( .A1(n53443), .A2(n55306), .ZN(n53445) );
  AOI22HSV0 U56410 ( .A1(n53931), .A2(n54289), .B1(n54465), .B2(n59495), .ZN(
        n53444) );
  NOR2HSV2 U56411 ( .A1(n53445), .A2(n53444), .ZN(n53451) );
  NAND2HSV0 U56412 ( .A1(n53848), .A2(n55518), .ZN(n54306) );
  NOR2HSV0 U56413 ( .A1(n53446), .A2(n54306), .ZN(n53449) );
  AOI22HSV0 U56414 ( .A1(n40683), .A2(n55491), .B1(n59589), .B2(n55231), .ZN(
        n53448) );
  NOR2HSV1 U56415 ( .A1(n53449), .A2(n53448), .ZN(n53450) );
  XOR2HSV0 U56416 ( .A1(n53451), .A2(n53450), .Z(n53452) );
  XOR2HSV0 U56417 ( .A1(n53453), .A2(n53452), .Z(n53454) );
  XNOR2HSV1 U56418 ( .A1(n53455), .A2(n53454), .ZN(n53456) );
  XNOR2HSV1 U56419 ( .A1(n53457), .A2(n53456), .ZN(n53459) );
  NAND2HSV0 U56420 ( .A1(n53795), .A2(n55319), .ZN(n53458) );
  XOR3HSV2 U56421 ( .A1(n53460), .A2(n53459), .A3(n53458), .Z(n53461) );
  XNOR2HSV1 U56422 ( .A1(n53462), .A2(n53461), .ZN(n53464) );
  NAND2HSV0 U56423 ( .A1(n53602), .A2(n55475), .ZN(n53463) );
  XOR2HSV0 U56424 ( .A1(n53464), .A2(n53463), .Z(n53466) );
  NAND2HSV0 U56425 ( .A1(n54265), .A2(n53523), .ZN(n53465) );
  XOR2HSV0 U56426 ( .A1(n53466), .A2(n53465), .Z(n53467) );
  XNOR2HSV1 U56427 ( .A1(n53468), .A2(n53467), .ZN(n53470) );
  NAND2HSV0 U56428 ( .A1(n29762), .A2(\pe1/got [8]), .ZN(n53469) );
  XOR2HSV0 U56429 ( .A1(n53470), .A2(n53469), .Z(n53471) );
  XNOR2HSV1 U56430 ( .A1(n53472), .A2(n53471), .ZN(n53475) );
  NAND2HSV0 U56431 ( .A1(n54115), .A2(n53473), .ZN(n53474) );
  XOR2HSV0 U56432 ( .A1(n53475), .A2(n53474), .Z(n53476) );
  XNOR2HSV1 U56433 ( .A1(n53477), .A2(n53476), .ZN(n53478) );
  XNOR2HSV1 U56434 ( .A1(n53479), .A2(n53478), .ZN(n53481) );
  NAND2HSV0 U56435 ( .A1(n54521), .A2(\pe1/got [14]), .ZN(n53480) );
  XOR3HSV2 U56436 ( .A1(n53482), .A2(n53481), .A3(n53480), .Z(n53483) );
  XNOR2HSV1 U56437 ( .A1(n53484), .A2(n53483), .ZN(n53485) );
  XNOR2HSV1 U56438 ( .A1(n53486), .A2(n53485), .ZN(n53487) );
  XNOR2HSV1 U56439 ( .A1(n53488), .A2(n53487), .ZN(n53489) );
  XNOR2HSV1 U56440 ( .A1(n53490), .A2(n53489), .ZN(n53491) );
  XNOR2HSV1 U56441 ( .A1(n53492), .A2(n53491), .ZN(n53494) );
  NAND2HSV0 U56442 ( .A1(n53768), .A2(n44530), .ZN(n53493) );
  XOR2HSV0 U56443 ( .A1(n53494), .A2(n53493), .Z(n53495) );
  XNOR2HSV1 U56444 ( .A1(n53496), .A2(n53495), .ZN(n53497) );
  XNOR2HSV1 U56445 ( .A1(n53498), .A2(n53497), .ZN(n53500) );
  BUFHSV2 U56446 ( .I(n55144), .Z(n54711) );
  INAND2HSV2 U56447 ( .A1(n54711), .B1(\pe1/got [23]), .ZN(n53499) );
  XNOR2HSV1 U56448 ( .A1(n53500), .A2(n53499), .ZN(n53501) );
  XNOR2HSV1 U56449 ( .A1(n53502), .A2(n53501), .ZN(n53506) );
  INAND2HSV2 U56450 ( .A1(n55529), .B1(\pe1/got [25]), .ZN(n53505) );
  CLKNAND2HSV0 U56451 ( .A1(n55213), .A2(n41689), .ZN(n53504) );
  XOR3HSV2 U56452 ( .A1(n53506), .A2(n53505), .A3(n53504), .Z(n53507) );
  XOR2HSV0 U56453 ( .A1(n53508), .A2(n53507), .Z(n53509) );
  XOR2HSV0 U56454 ( .A1(n53510), .A2(n53509), .Z(n53517) );
  NAND2HSV2 U56455 ( .A1(n25840), .A2(n53512), .ZN(n53516) );
  NAND2HSV2 U56456 ( .A1(n53514), .A2(n53513), .ZN(n53515) );
  XOR3HSV2 U56457 ( .A1(n53517), .A2(n53516), .A3(n53515), .Z(\pe1/poht [2])
         );
  INHSV2 U56458 ( .I(n53791), .ZN(n55574) );
  CLKNAND2HSV0 U56459 ( .A1(n55574), .A2(n53518), .ZN(n53648) );
  NAND2HSV2 U56460 ( .A1(n29654), .A2(n53519), .ZN(n53654) );
  INHSV2 U56461 ( .I(n53654), .ZN(n54635) );
  CLKNAND2HSV0 U56462 ( .A1(n55489), .A2(n54033), .ZN(n53646) );
  CLKNAND2HSV0 U56463 ( .A1(n53792), .A2(n41689), .ZN(n53641) );
  CLKNAND2HSV0 U56464 ( .A1(n55341), .A2(n53520), .ZN(n53637) );
  NAND2HSV0 U56465 ( .A1(n55229), .A2(\pe1/got [23]), .ZN(n53635) );
  NAND2HSV0 U56466 ( .A1(n53521), .A2(n54724), .ZN(n53631) );
  CLKNHSV0 U56467 ( .I(n59360), .ZN(n53912) );
  NOR2HSV0 U56468 ( .A1(n53912), .A2(n48338), .ZN(n53629) );
  NAND2HSV0 U56469 ( .A1(n53522), .A2(n59995), .ZN(n53627) );
  CLKNAND2HSV0 U56470 ( .A1(n41508), .A2(n54716), .ZN(n53625) );
  NOR2HSV0 U56471 ( .A1(n54040), .A2(n53911), .ZN(n53623) );
  NOR2HSV0 U56472 ( .A1(n54731), .A2(n54039), .ZN(n53621) );
  NAND2HSV0 U56473 ( .A1(n54557), .A2(n54969), .ZN(n53618) );
  NAND2HSV0 U56474 ( .A1(n54264), .A2(n54812), .ZN(n53616) );
  NOR2HSV0 U56475 ( .A1(n41566), .A2(n55082), .ZN(n53612) );
  NAND2HSV0 U56476 ( .A1(n54456), .A2(\pe1/got [9]), .ZN(n53608) );
  NAND2HSV2 U56477 ( .A1(n53524), .A2(n53523), .ZN(n53601) );
  NAND2HSV0 U56478 ( .A1(n59529), .A2(n53863), .ZN(n53599) );
  NAND2HSV0 U56479 ( .A1(n53795), .A2(n55475), .ZN(n53598) );
  NAND2HSV0 U56480 ( .A1(n59373), .A2(n25179), .ZN(n53676) );
  NOR2HSV0 U56481 ( .A1(n53525), .A2(n53676), .ZN(n53528) );
  AOI22HSV0 U56482 ( .A1(n55595), .A2(n25179), .B1(n40684), .B2(n59373), .ZN(
        n53527) );
  NOR2HSV2 U56483 ( .A1(n53528), .A2(n53527), .ZN(n53534) );
  NAND2HSV0 U56484 ( .A1(\pe1/aot [25]), .A2(n54988), .ZN(n54184) );
  NOR2HSV0 U56485 ( .A1(n53529), .A2(n54184), .ZN(n53532) );
  AOI22HSV0 U56486 ( .A1(n25226), .A2(n54292), .B1(\pe1/aot [25]), .B2(n55501), 
        .ZN(n53531) );
  NOR2HSV1 U56487 ( .A1(n53532), .A2(n53531), .ZN(n53533) );
  XNOR2HSV1 U56488 ( .A1(n53534), .A2(n53533), .ZN(n53537) );
  NAND2HSV0 U56489 ( .A1(\pe1/aot [3]), .A2(n53411), .ZN(n53658) );
  XOR2HSV0 U56490 ( .A1(n53535), .A2(n53658), .Z(n53536) );
  XNOR2HSV1 U56491 ( .A1(n53537), .A2(n53536), .ZN(n53562) );
  NAND2HSV0 U56492 ( .A1(n53673), .A2(\pe1/bq[2] ), .ZN(n53540) );
  NAND2HSV0 U56493 ( .A1(n53538), .A2(\pe1/bq[4] ), .ZN(n53539) );
  XOR2HSV0 U56494 ( .A1(n53540), .A2(n53539), .Z(n53542) );
  NAND2HSV0 U56495 ( .A1(n59675), .A2(n54104), .ZN(n53541) );
  XOR2HSV0 U56496 ( .A1(n53542), .A2(n53541), .Z(n53544) );
  NAND2HSV0 U56497 ( .A1(n41248), .A2(\pe1/got [3]), .ZN(n53543) );
  XNOR2HSV1 U56498 ( .A1(n53544), .A2(n53543), .ZN(n53561) );
  NAND2HSV0 U56499 ( .A1(\pe1/aot [15]), .A2(\pe1/bq[18] ), .ZN(n53546) );
  NAND2HSV0 U56500 ( .A1(\pe1/aot [14]), .A2(n42092), .ZN(n53545) );
  XOR2HSV0 U56501 ( .A1(n53546), .A2(n53545), .Z(n53550) );
  NAND2HSV0 U56502 ( .A1(n53954), .A2(n55352), .ZN(n53548) );
  NAND2HSV0 U56503 ( .A1(n54307), .A2(\pe1/bq[9] ), .ZN(n53547) );
  XOR2HSV0 U56504 ( .A1(n53548), .A2(n53547), .Z(n53549) );
  XOR2HSV0 U56505 ( .A1(n53550), .A2(n53549), .Z(n53559) );
  NAND2HSV0 U56506 ( .A1(n59990), .A2(n54565), .ZN(n53552) );
  NAND2HSV0 U56507 ( .A1(n59987), .A2(n42373), .ZN(n53551) );
  XOR2HSV0 U56508 ( .A1(n53552), .A2(n53551), .Z(n53557) );
  NOR2HSV0 U56509 ( .A1(n55307), .A2(n53553), .ZN(n53555) );
  NAND2HSV0 U56510 ( .A1(n42093), .A2(n54179), .ZN(n53554) );
  XOR2HSV0 U56511 ( .A1(n53555), .A2(n53554), .Z(n53556) );
  XOR2HSV0 U56512 ( .A1(n53557), .A2(n53556), .Z(n53558) );
  XOR2HSV0 U56513 ( .A1(n53559), .A2(n53558), .Z(n53560) );
  XOR3HSV2 U56514 ( .A1(n53562), .A2(n53561), .A3(n53560), .Z(n53596) );
  NAND2HSV0 U56515 ( .A1(n53717), .A2(n54048), .ZN(n53564) );
  NAND2HSV0 U56516 ( .A1(n59985), .A2(n54668), .ZN(n53563) );
  XOR2HSV0 U56517 ( .A1(n53564), .A2(n53563), .Z(n53568) );
  INHSV1 U56518 ( .I(n54093), .ZN(n54274) );
  NAND2HSV0 U56519 ( .A1(n53931), .A2(n54274), .ZN(n53566) );
  NAND2HSV0 U56520 ( .A1(n54500), .A2(n48380), .ZN(n53565) );
  XOR2HSV0 U56521 ( .A1(n53566), .A2(n53565), .Z(n53567) );
  XOR2HSV0 U56522 ( .A1(n53568), .A2(n53567), .Z(n53577) );
  NAND2HSV0 U56523 ( .A1(n54497), .A2(n54836), .ZN(n53570) );
  NAND2HSV0 U56524 ( .A1(n41169), .A2(\pe1/bq[11] ), .ZN(n53569) );
  XOR2HSV0 U56525 ( .A1(n53570), .A2(n53569), .Z(n53575) );
  NAND2HSV0 U56526 ( .A1(n54364), .A2(n53571), .ZN(n53573) );
  NAND2HSV0 U56527 ( .A1(n40683), .A2(n54289), .ZN(n53572) );
  XOR2HSV0 U56528 ( .A1(n53573), .A2(n53572), .Z(n53574) );
  XOR2HSV0 U56529 ( .A1(n53575), .A2(n53574), .Z(n53576) );
  XOR2HSV0 U56530 ( .A1(n53577), .A2(n53576), .Z(n53594) );
  NAND2HSV0 U56531 ( .A1(n54662), .A2(n42106), .ZN(n53580) );
  NAND2HSV0 U56532 ( .A1(n54188), .A2(n53578), .ZN(n53579) );
  XOR2HSV0 U56533 ( .A1(n53580), .A2(n53579), .Z(n53584) );
  NAND2HSV2 U56534 ( .A1(n59986), .A2(n55231), .ZN(n53582) );
  NAND2HSV0 U56535 ( .A1(\pe1/aot [16]), .A2(n54995), .ZN(n53581) );
  XOR2HSV0 U56536 ( .A1(n53582), .A2(n53581), .Z(n53583) );
  XOR2HSV0 U56537 ( .A1(n53584), .A2(n53583), .Z(n53592) );
  NAND2HSV0 U56538 ( .A1(n53812), .A2(\pe1/bq[21] ), .ZN(n53586) );
  NAND2HSV0 U56539 ( .A1(\pe1/aot [5]), .A2(n53805), .ZN(n53585) );
  XOR2HSV0 U56540 ( .A1(n53586), .A2(n53585), .Z(n53590) );
  NAND2HSV0 U56541 ( .A1(n59619), .A2(n40553), .ZN(n53588) );
  NAND2HSV0 U56542 ( .A1(n59992), .A2(n41771), .ZN(n53587) );
  XOR2HSV0 U56543 ( .A1(n53588), .A2(n53587), .Z(n53589) );
  XOR2HSV0 U56544 ( .A1(n53590), .A2(n53589), .Z(n53591) );
  XOR2HSV0 U56545 ( .A1(n53592), .A2(n53591), .Z(n53593) );
  XOR2HSV0 U56546 ( .A1(n53594), .A2(n53593), .Z(n53595) );
  XNOR2HSV1 U56547 ( .A1(n53596), .A2(n53595), .ZN(n53597) );
  XOR3HSV1 U56548 ( .A1(n53599), .A2(n53598), .A3(n53597), .Z(n53600) );
  XNOR2HSV1 U56549 ( .A1(n53601), .A2(n53600), .ZN(n53604) );
  NAND2HSV0 U56550 ( .A1(n53602), .A2(n55570), .ZN(n53603) );
  XOR2HSV0 U56551 ( .A1(n53604), .A2(n53603), .Z(n53606) );
  NAND2HSV0 U56552 ( .A1(n59919), .A2(n55339), .ZN(n53605) );
  XOR2HSV0 U56553 ( .A1(n53606), .A2(n53605), .Z(n53607) );
  XNOR2HSV1 U56554 ( .A1(n53608), .A2(n53607), .ZN(n53610) );
  NAND2HSV0 U56555 ( .A1(n29773), .A2(n55088), .ZN(n53609) );
  XOR2HSV0 U56556 ( .A1(n53610), .A2(n53609), .Z(n53611) );
  XNOR2HSV1 U56557 ( .A1(n53612), .A2(n53611), .ZN(n53614) );
  NAND2HSV0 U56558 ( .A1(n53996), .A2(n55337), .ZN(n53613) );
  XOR2HSV0 U56559 ( .A1(n53614), .A2(n53613), .Z(n53615) );
  XNOR2HSV1 U56560 ( .A1(n53616), .A2(n53615), .ZN(n53617) );
  XNOR2HSV1 U56561 ( .A1(n53618), .A2(n53617), .ZN(n53620) );
  NAND2HSV0 U56562 ( .A1(n41850), .A2(n54161), .ZN(n53619) );
  XOR3HSV2 U56563 ( .A1(n53621), .A2(n53620), .A3(n53619), .Z(n53622) );
  XNOR2HSV1 U56564 ( .A1(n53623), .A2(n53622), .ZN(n53624) );
  XNOR2HSV1 U56565 ( .A1(n53625), .A2(n53624), .ZN(n53626) );
  XNOR2HSV1 U56566 ( .A1(n53627), .A2(n53626), .ZN(n53628) );
  XNOR2HSV1 U56567 ( .A1(n53629), .A2(n53628), .ZN(n53630) );
  XNOR2HSV1 U56568 ( .A1(n53631), .A2(n53630), .ZN(n53633) );
  NAND2HSV0 U56569 ( .A1(n53768), .A2(n54160), .ZN(n53632) );
  XOR2HSV0 U56570 ( .A1(n53633), .A2(n53632), .Z(n53634) );
  XNOR2HSV1 U56571 ( .A1(n53635), .A2(n53634), .ZN(n53636) );
  XNOR2HSV1 U56572 ( .A1(n53637), .A2(n53636), .ZN(n53639) );
  INAND2HSV2 U56573 ( .A1(n54711), .B1(\pe1/got [25]), .ZN(n53638) );
  XNOR2HSV1 U56574 ( .A1(n53639), .A2(n53638), .ZN(n53640) );
  XNOR2HSV1 U56575 ( .A1(n53641), .A2(n53640), .ZN(n53644) );
  INHSV2 U56576 ( .I(n54146), .ZN(n55330) );
  INAND2HSV2 U56577 ( .A1(n55330), .B1(n59374), .ZN(n53643) );
  CLKNAND2HSV0 U56578 ( .A1(n55476), .A2(n40873), .ZN(n53642) );
  XOR3HSV2 U56579 ( .A1(n53644), .A2(n53643), .A3(n53642), .Z(n53645) );
  XOR2HSV0 U56580 ( .A1(n53646), .A2(n53645), .Z(n53647) );
  XOR2HSV0 U56581 ( .A1(n53648), .A2(n53647), .Z(n53653) );
  NAND2HSV2 U56582 ( .A1(n59428), .A2(n53649), .ZN(n53652) );
  INHSV2 U56583 ( .I(n54154), .ZN(n55158) );
  XOR3HSV2 U56584 ( .A1(n53653), .A2(n53652), .A3(n53651), .Z(po1) );
  INHSV2 U56585 ( .I(n53791), .ZN(n55488) );
  CLKNAND2HSV0 U56586 ( .A1(n55488), .A2(n53512), .ZN(n53785) );
  BUFHSV2 U56587 ( .I(n53654), .Z(n55289) );
  CLKNAND2HSV1 U56588 ( .A1(n55289), .A2(\pe1/got [28]), .ZN(n53783) );
  CLKNAND2HSV0 U56589 ( .A1(n53792), .A2(\pe1/got [25]), .ZN(n53778) );
  CLKNAND2HSV1 U56590 ( .A1(n53656), .A2(n53655), .ZN(n55450) );
  CLKNAND2HSV0 U56591 ( .A1(\pe1/got [23]), .A2(n55450), .ZN(n53774) );
  NAND2HSV0 U56592 ( .A1(n55229), .A2(n54160), .ZN(n53772) );
  BUFHSV2 U56593 ( .I(n59391), .Z(n54038) );
  CLKNAND2HSV1 U56594 ( .A1(n54038), .A2(n44530), .ZN(n53767) );
  NOR2HSV1 U56595 ( .A1(n53912), .A2(n41928), .ZN(n53765) );
  CLKNAND2HSV0 U56596 ( .A1(n29741), .A2(n54716), .ZN(n53763) );
  CLKNAND2HSV0 U56597 ( .A1(n54814), .A2(n54135), .ZN(n53761) );
  INHSV2 U56598 ( .I(n53657), .ZN(n54040) );
  NOR2HSV0 U56599 ( .A1(n54040), .A2(n53793), .ZN(n53759) );
  NOR2HSV0 U56600 ( .A1(n54731), .A2(n54884), .ZN(n53757) );
  NAND2HSV0 U56601 ( .A1(n53913), .A2(n54812), .ZN(n53754) );
  NAND2HSV0 U56602 ( .A1(n54264), .A2(n55087), .ZN(n53752) );
  NOR2HSV0 U56603 ( .A1(n42438), .A2(n54636), .ZN(n53748) );
  NAND2HSV0 U56604 ( .A1(n54456), .A2(n55339), .ZN(n53744) );
  NAND2HSV0 U56605 ( .A1(n42360), .A2(n55475), .ZN(n53738) );
  NAND2HSV0 U56606 ( .A1(n59529), .A2(n55514), .ZN(n53736) );
  NAND2HSV0 U56607 ( .A1(n26833), .A2(n54104), .ZN(n53670) );
  CLKNHSV0 U56608 ( .I(n53658), .ZN(n53662) );
  AOI21HSV0 U56609 ( .A1(n59389), .A2(n40553), .B(n53659), .ZN(n53660) );
  AOI21HSV2 U56610 ( .A1(n53662), .A2(n53661), .B(n53660), .ZN(n53668) );
  INHSV2 U56611 ( .I(n54399), .ZN(n54083) );
  NAND2HSV0 U56612 ( .A1(n59385), .A2(n54083), .ZN(n53665) );
  NAND2HSV0 U56613 ( .A1(n53812), .A2(n54083), .ZN(n55240) );
  NOR2HSV0 U56614 ( .A1(n53663), .A2(n55240), .ZN(n53664) );
  AOI21HSV0 U56615 ( .A1(n53666), .A2(n53665), .B(n53664), .ZN(n53667) );
  XOR2HSV0 U56616 ( .A1(n53668), .A2(n53667), .Z(n53669) );
  XNOR2HSV1 U56617 ( .A1(n53670), .A2(n53669), .ZN(n53682) );
  NAND2HSV2 U56618 ( .A1(n54912), .A2(n54063), .ZN(n55312) );
  NOR2HSV0 U56619 ( .A1(n53671), .A2(n55312), .ZN(n53675) );
  CLKNHSV0 U56620 ( .I(n55185), .ZN(n55392) );
  AOI22HSV0 U56621 ( .A1(n53673), .A2(n55392), .B1(n42092), .B2(n55103), .ZN(
        n53674) );
  NOR2HSV2 U56622 ( .A1(n53675), .A2(n53674), .ZN(n53677) );
  XOR2HSV0 U56623 ( .A1(n53677), .A2(n53676), .Z(n53680) );
  NOR2HSV0 U56624 ( .A1(n46629), .A2(n54735), .ZN(n54295) );
  NAND2HSV0 U56625 ( .A1(n59992), .A2(n41644), .ZN(n53678) );
  XOR2HSV0 U56626 ( .A1(n54295), .A2(n53678), .Z(n53679) );
  XNOR2HSV1 U56627 ( .A1(n53680), .A2(n53679), .ZN(n53681) );
  XNOR2HSV1 U56628 ( .A1(n53682), .A2(n53681), .ZN(n53699) );
  NAND2HSV0 U56629 ( .A1(n54662), .A2(\pe1/bq[21] ), .ZN(n53684) );
  NAND2HSV2 U56630 ( .A1(n59986), .A2(n54289), .ZN(n53683) );
  XOR2HSV0 U56631 ( .A1(n53684), .A2(n53683), .Z(n53688) );
  NAND2HSV0 U56632 ( .A1(n54497), .A2(n41424), .ZN(n53686) );
  NAND2HSV0 U56633 ( .A1(n59619), .A2(n53805), .ZN(n53685) );
  XOR2HSV0 U56634 ( .A1(n53686), .A2(n53685), .Z(n53687) );
  XOR2HSV0 U56635 ( .A1(n53688), .A2(n53687), .Z(n53697) );
  NAND2HSV0 U56636 ( .A1(\pe1/aot [16]), .A2(n54836), .ZN(n53690) );
  NAND2HSV0 U56637 ( .A1(n53954), .A2(\pe1/bq[9] ), .ZN(n53689) );
  XOR2HSV0 U56638 ( .A1(n53690), .A2(n53689), .Z(n53695) );
  NAND2HSV0 U56639 ( .A1(n41768), .A2(n42373), .ZN(n53693) );
  NAND2HSV0 U56640 ( .A1(\pe1/aot [21]), .A2(\pe1/bq[11] ), .ZN(n53692) );
  XOR2HSV0 U56641 ( .A1(n53693), .A2(n53692), .Z(n53694) );
  XOR2HSV0 U56642 ( .A1(n53695), .A2(n53694), .Z(n53696) );
  XOR2HSV0 U56643 ( .A1(n53697), .A2(n53696), .Z(n53698) );
  XOR2HSV0 U56644 ( .A1(n53699), .A2(n53698), .Z(n53733) );
  NAND2HSV0 U56645 ( .A1(n54500), .A2(n54999), .ZN(n53701) );
  NAND2HSV0 U56646 ( .A1(\pe1/aot [15]), .A2(n54995), .ZN(n53700) );
  XOR2HSV0 U56647 ( .A1(n53701), .A2(n53700), .Z(n53705) );
  NAND2HSV0 U56648 ( .A1(n59993), .A2(n41771), .ZN(n53703) );
  NAND2HSV0 U56649 ( .A1(n40683), .A2(\pe1/bq[4] ), .ZN(n53702) );
  XOR2HSV0 U56650 ( .A1(n53703), .A2(n53702), .Z(n53704) );
  XOR2HSV0 U56651 ( .A1(n53705), .A2(n53704), .Z(n53714) );
  NAND2HSV0 U56652 ( .A1(n54904), .A2(n53949), .ZN(n53707) );
  NAND2HSV0 U56653 ( .A1(n54188), .A2(n54048), .ZN(n53706) );
  XOR2HSV0 U56654 ( .A1(n53707), .A2(n53706), .Z(n53712) );
  NAND2HSV0 U56655 ( .A1(\pe1/aot [24]), .A2(n53708), .ZN(n53710) );
  NAND2HSV0 U56656 ( .A1(\pe1/aot [14]), .A2(\pe1/bq[18] ), .ZN(n53709) );
  XOR2HSV0 U56657 ( .A1(n53710), .A2(n53709), .Z(n53711) );
  XOR2HSV0 U56658 ( .A1(n53712), .A2(n53711), .Z(n53713) );
  XOR2HSV0 U56659 ( .A1(n53714), .A2(n53713), .Z(n53731) );
  NAND2HSV0 U56660 ( .A1(\pe1/aot [25]), .A2(n54274), .ZN(n53716) );
  NAND2HSV0 U56661 ( .A1(n59985), .A2(\pe1/bq[2] ), .ZN(n53715) );
  XOR2HSV0 U56662 ( .A1(n53716), .A2(n53715), .Z(n53722) );
  NAND2HSV0 U56663 ( .A1(n53717), .A2(n54465), .ZN(n53720) );
  NAND2HSV0 U56664 ( .A1(n54578), .A2(n53718), .ZN(n53719) );
  XOR2HSV0 U56665 ( .A1(n53720), .A2(n53719), .Z(n53721) );
  XOR2HSV0 U56666 ( .A1(n53722), .A2(n53721), .Z(n53729) );
  NOR2HSV0 U56667 ( .A1(n41885), .A2(n53723), .ZN(n53725) );
  NAND2HSV0 U56668 ( .A1(n54364), .A2(n54179), .ZN(n53724) );
  XOR2HSV0 U56669 ( .A1(n53725), .A2(n53724), .Z(n53727) );
  NAND2HSV0 U56670 ( .A1(n59675), .A2(\pe1/got [1]), .ZN(n53726) );
  XOR2HSV0 U56671 ( .A1(n53727), .A2(n53726), .Z(n53728) );
  XNOR2HSV1 U56672 ( .A1(n53729), .A2(n53728), .ZN(n53730) );
  XNOR2HSV1 U56673 ( .A1(n53731), .A2(n53730), .ZN(n53732) );
  XNOR2HSV1 U56674 ( .A1(n53733), .A2(n53732), .ZN(n53735) );
  NAND2HSV0 U56675 ( .A1(n53795), .A2(n53863), .ZN(n53734) );
  XOR3HSV2 U56676 ( .A1(n53736), .A2(n53735), .A3(n53734), .Z(n53737) );
  XNOR2HSV1 U56677 ( .A1(n53738), .A2(n53737), .ZN(n53740) );
  NAND2HSV0 U56678 ( .A1(n59686), .A2(n55448), .ZN(n53739) );
  XOR2HSV0 U56679 ( .A1(n53740), .A2(n53739), .Z(n53742) );
  NAND2HSV0 U56680 ( .A1(n54265), .A2(n54894), .ZN(n53741) );
  XOR2HSV0 U56681 ( .A1(n53742), .A2(n53741), .Z(n53743) );
  XNOR2HSV1 U56682 ( .A1(n53744), .A2(n53743), .ZN(n53746) );
  NAND2HSV0 U56683 ( .A1(n29763), .A2(n55145), .ZN(n53745) );
  XOR2HSV0 U56684 ( .A1(n53746), .A2(n53745), .Z(n53747) );
  XNOR2HSV1 U56685 ( .A1(n53748), .A2(n53747), .ZN(n53750) );
  NAND2HSV0 U56686 ( .A1(n53996), .A2(n54970), .ZN(n53749) );
  XOR2HSV0 U56687 ( .A1(n53750), .A2(n53749), .Z(n53751) );
  XNOR2HSV1 U56688 ( .A1(n53752), .A2(n53751), .ZN(n53753) );
  XNOR2HSV1 U56689 ( .A1(n53754), .A2(n53753), .ZN(n53756) );
  BUFHSV2 U56690 ( .I(n41312), .Z(n53877) );
  NOR2HSV2 U56691 ( .A1(n53877), .A2(n54039), .ZN(n53755) );
  XOR3HSV2 U56692 ( .A1(n53757), .A2(n53756), .A3(n53755), .Z(n53758) );
  XNOR2HSV1 U56693 ( .A1(n53759), .A2(n53758), .ZN(n53760) );
  XNOR2HSV1 U56694 ( .A1(n53761), .A2(n53760), .ZN(n53762) );
  XNOR2HSV1 U56695 ( .A1(n53763), .A2(n53762), .ZN(n53764) );
  XOR2HSV0 U56696 ( .A1(n53765), .A2(n53764), .Z(n53766) );
  XNOR2HSV1 U56697 ( .A1(n53767), .A2(n53766), .ZN(n53770) );
  NAND2HSV0 U56698 ( .A1(n53768), .A2(\pe1/got [21]), .ZN(n53769) );
  XOR2HSV0 U56699 ( .A1(n53770), .A2(n53769), .Z(n53771) );
  XNOR2HSV1 U56700 ( .A1(n53772), .A2(n53771), .ZN(n53773) );
  XNOR2HSV1 U56701 ( .A1(n53774), .A2(n53773), .ZN(n53776) );
  INHSV2 U56702 ( .I(n54711), .ZN(n55069) );
  CLKNAND2HSV0 U56703 ( .A1(n55069), .A2(n53520), .ZN(n53775) );
  XNOR2HSV1 U56704 ( .A1(n53776), .A2(n53775), .ZN(n53777) );
  XNOR2HSV1 U56705 ( .A1(n53778), .A2(n53777), .ZN(n53781) );
  INAND2HSV2 U56706 ( .A1(n55330), .B1(n41689), .ZN(n53780) );
  CLKNAND2HSV0 U56707 ( .A1(n55213), .A2(n59374), .ZN(n53779) );
  XOR3HSV2 U56708 ( .A1(n53781), .A2(n53780), .A3(n53779), .Z(n53782) );
  XOR2HSV0 U56709 ( .A1(n53783), .A2(n53782), .Z(n53784) );
  XOR2HSV0 U56710 ( .A1(n53785), .A2(n53784), .Z(n53790) );
  NAND2HSV2 U56711 ( .A1(n53786), .A2(n59428), .ZN(n53789) );
  NAND2HSV0 U56712 ( .A1(n59520), .A2(n53787), .ZN(n53788) );
  XOR3HSV2 U56713 ( .A1(n53790), .A2(n53789), .A3(n53788), .Z(\pe1/poht [1])
         );
  CLKNAND2HSV0 U56714 ( .A1(n55593), .A2(\pe1/got [26]), .ZN(n53907) );
  CLKNAND2HSV1 U56715 ( .A1(n55489), .A2(\pe1/got [25]), .ZN(n53905) );
  INHSV2 U56716 ( .I(n53792), .ZN(n55162) );
  CLKNAND2HSV1 U56717 ( .A1(n55449), .A2(n54160), .ZN(n53900) );
  NAND2HSV0 U56718 ( .A1(n59521), .A2(n44530), .ZN(n53896) );
  NAND2HSV0 U56719 ( .A1(n59422), .A2(\pe1/got [19]), .ZN(n53894) );
  CLKNAND2HSV1 U56720 ( .A1(n54038), .A2(n54135), .ZN(n53890) );
  NOR2HSV1 U56721 ( .A1(n53912), .A2(n53793), .ZN(n53888) );
  CLKNAND2HSV1 U56722 ( .A1(n29741), .A2(n54241), .ZN(n53886) );
  CLKNAND2HSV0 U56723 ( .A1(n41508), .A2(n54969), .ZN(n53884) );
  NOR2HSV1 U56724 ( .A1(n54040), .A2(n54957), .ZN(n53882) );
  INHSV2 U56725 ( .I(n53794), .ZN(n54815) );
  NOR2HSV0 U56726 ( .A1(n54815), .A2(n55082), .ZN(n53880) );
  NAND2HSV0 U56727 ( .A1(n53913), .A2(n55088), .ZN(n53876) );
  CLKNAND2HSV0 U56728 ( .A1(n54162), .A2(n55145), .ZN(n53874) );
  NAND2HSV0 U56729 ( .A1(n54456), .A2(\pe1/got [5]), .ZN(n53867) );
  NAND2HSV0 U56730 ( .A1(n42360), .A2(n54104), .ZN(n53860) );
  NAND2HSV0 U56731 ( .A1(n53795), .A2(n54455), .ZN(n53858) );
  NAND2HSV0 U56732 ( .A1(n54662), .A2(\pe1/bq[18] ), .ZN(n53797) );
  NAND2HSV0 U56733 ( .A1(\pe1/aot [15]), .A2(n41641), .ZN(n53796) );
  XOR2HSV0 U56734 ( .A1(n53797), .A2(n53796), .Z(n53802) );
  NAND2HSV0 U56735 ( .A1(n59987), .A2(n53798), .ZN(n53800) );
  NAND2HSV0 U56736 ( .A1(\pe1/aot [14]), .A2(\pe1/bq[15] ), .ZN(n53799) );
  XOR2HSV0 U56737 ( .A1(n53800), .A2(n53799), .Z(n53801) );
  XOR2HSV0 U56738 ( .A1(n53802), .A2(n53801), .Z(n53811) );
  NAND2HSV0 U56739 ( .A1(\pe1/aot [24]), .A2(n54289), .ZN(n53804) );
  NAND2HSV0 U56740 ( .A1(n53954), .A2(n55231), .ZN(n53803) );
  XOR2HSV0 U56741 ( .A1(n53804), .A2(n53803), .Z(n53809) );
  CLKNHSV0 U56742 ( .I(n55524), .ZN(n54743) );
  NAND2HSV0 U56743 ( .A1(n54743), .A2(n53805), .ZN(n53807) );
  NAND2HSV0 U56744 ( .A1(n55496), .A2(n41644), .ZN(n53806) );
  XOR2HSV0 U56745 ( .A1(n53807), .A2(n53806), .Z(n53808) );
  XOR2HSV0 U56746 ( .A1(n53809), .A2(n53808), .Z(n53810) );
  XOR2HSV0 U56747 ( .A1(n53811), .A2(n53810), .Z(n53830) );
  NAND2HSV0 U56748 ( .A1(n44541), .A2(\pe1/bq[16] ), .ZN(n53814) );
  NAND2HSV0 U56749 ( .A1(n53812), .A2(\pe1/bq[17] ), .ZN(n53813) );
  XOR2HSV0 U56750 ( .A1(n53814), .A2(n53813), .Z(n53818) );
  NAND2HSV0 U56751 ( .A1(n55553), .A2(n53949), .ZN(n53816) );
  NAND2HSV0 U56752 ( .A1(n54364), .A2(n55352), .ZN(n53815) );
  XOR2HSV0 U56753 ( .A1(n53816), .A2(n53815), .Z(n53817) );
  XOR2HSV0 U56754 ( .A1(n53818), .A2(n53817), .Z(n53828) );
  NOR2HSV0 U56755 ( .A1(n54901), .A2(n53819), .ZN(n53821) );
  NAND2HSV0 U56756 ( .A1(n54904), .A2(\pe1/bq[21] ), .ZN(n53820) );
  XOR2HSV0 U56757 ( .A1(n53821), .A2(n53820), .Z(n53826) );
  NAND2HSV0 U56758 ( .A1(n59619), .A2(n54274), .ZN(n55354) );
  NOR2HSV0 U56759 ( .A1(n53822), .A2(n55354), .ZN(n53824) );
  AOI22HSV0 U56760 ( .A1(n54078), .A2(n55394), .B1(n41173), .B2(n55433), .ZN(
        n53823) );
  NOR2HSV2 U56761 ( .A1(n53824), .A2(n53823), .ZN(n53825) );
  XNOR2HSV1 U56762 ( .A1(n53826), .A2(n53825), .ZN(n53827) );
  XNOR2HSV1 U56763 ( .A1(n53828), .A2(n53827), .ZN(n53829) );
  XNOR2HSV1 U56764 ( .A1(n53830), .A2(n53829), .ZN(n53856) );
  NOR2HSV1 U56765 ( .A1(n54846), .A2(n55185), .ZN(n55343) );
  CLKNHSV0 U56766 ( .I(n54846), .ZN(n55093) );
  AOI22HSV0 U56767 ( .A1(n40683), .A2(n54292), .B1(n42092), .B2(n55093), .ZN(
        n53831) );
  AOI21HSV0 U56768 ( .A1(n53832), .A2(n55343), .B(n53831), .ZN(n53837) );
  NOR2HSV0 U56769 ( .A1(n46629), .A2(n53834), .ZN(n54076) );
  NOR2HSV0 U56770 ( .A1(n53833), .A2(n54399), .ZN(n53968) );
  INHSV1 U56771 ( .I(n53834), .ZN(n55451) );
  AOI22HSV0 U56772 ( .A1(n54293), .A2(n55491), .B1(n40898), .B2(n55451), .ZN(
        n53835) );
  AOI21HSV1 U56773 ( .A1(n54076), .A2(n53968), .B(n53835), .ZN(n53836) );
  XOR2HSV0 U56774 ( .A1(n53837), .A2(n53836), .Z(n53845) );
  NOR2HSV0 U56775 ( .A1(n54829), .A2(n48059), .ZN(n53970) );
  NOR2HSV0 U56776 ( .A1(n54673), .A2(n53691), .ZN(n54087) );
  NOR2HSV0 U56777 ( .A1(n54673), .A2(n48059), .ZN(n54313) );
  AOI21HSV0 U56778 ( .A1(n42373), .A2(n54900), .B(n54313), .ZN(n53838) );
  AOI21HSV1 U56779 ( .A1(n53970), .A2(n54087), .B(n53838), .ZN(n53843) );
  NAND2HSV0 U56780 ( .A1(n55578), .A2(n54565), .ZN(n54734) );
  NOR2HSV0 U56781 ( .A1(n53839), .A2(n54734), .ZN(n53841) );
  AOI22HSV0 U56782 ( .A1(n55380), .A2(n54565), .B1(n41771), .B2(n59730), .ZN(
        n53840) );
  NOR2HSV2 U56783 ( .A1(n53841), .A2(n53840), .ZN(n53842) );
  XNOR2HSV1 U56784 ( .A1(n53843), .A2(n53842), .ZN(n53844) );
  XNOR2HSV1 U56785 ( .A1(n53845), .A2(n53844), .ZN(n53854) );
  NAND2HSV0 U56786 ( .A1(n54578), .A2(n54302), .ZN(n53847) );
  NAND2HSV0 U56787 ( .A1(n54500), .A2(\pe1/bq[11] ), .ZN(n53846) );
  XOR2HSV0 U56788 ( .A1(n53847), .A2(n53846), .Z(n53852) );
  NAND2HSV0 U56789 ( .A1(n42093), .A2(\pe1/bq[9] ), .ZN(n53850) );
  NAND2HSV0 U56790 ( .A1(n53848), .A2(n54371), .ZN(n53849) );
  XOR2HSV0 U56791 ( .A1(n53850), .A2(n53849), .Z(n53851) );
  XOR2HSV0 U56792 ( .A1(n53852), .A2(n53851), .Z(n53853) );
  XNOR2HSV1 U56793 ( .A1(n53854), .A2(n53853), .ZN(n53855) );
  XNOR2HSV1 U56794 ( .A1(n53856), .A2(n53855), .ZN(n53857) );
  XNOR2HSV1 U56795 ( .A1(n53858), .A2(n53857), .ZN(n53859) );
  XNOR2HSV1 U56796 ( .A1(n53860), .A2(n53859), .ZN(n53862) );
  NAND2HSV0 U56797 ( .A1(n59686), .A2(n55319), .ZN(n53861) );
  XOR2HSV0 U56798 ( .A1(n53862), .A2(n53861), .Z(n53865) );
  NAND2HSV0 U56799 ( .A1(n54265), .A2(n53863), .ZN(n53864) );
  XOR2HSV0 U56800 ( .A1(n53865), .A2(n53864), .Z(n53866) );
  XNOR2HSV1 U56801 ( .A1(n53867), .A2(n53866), .ZN(n53869) );
  NAND2HSV0 U56802 ( .A1(n29762), .A2(\pe1/got [6]), .ZN(n53868) );
  XOR2HSV0 U56803 ( .A1(n53869), .A2(n53868), .Z(n53872) );
  NOR2HSV0 U56804 ( .A1(n41301), .A2(n55019), .ZN(n53871) );
  NAND2HSV0 U56805 ( .A1(n53996), .A2(\pe1/got [8]), .ZN(n53870) );
  XOR3HSV1 U56806 ( .A1(n53872), .A2(n53871), .A3(n53870), .Z(n53873) );
  XNOR2HSV1 U56807 ( .A1(n53874), .A2(n53873), .ZN(n53875) );
  XNOR2HSV1 U56808 ( .A1(n53876), .A2(n53875), .ZN(n53879) );
  BUFHSV2 U56809 ( .I(n54879), .Z(n54453) );
  NOR2HSV2 U56810 ( .A1(n53877), .A2(n54453), .ZN(n53878) );
  XOR3HSV2 U56811 ( .A1(n53880), .A2(n53879), .A3(n53878), .Z(n53881) );
  XNOR2HSV1 U56812 ( .A1(n53882), .A2(n53881), .ZN(n53883) );
  XNOR2HSV1 U56813 ( .A1(n53884), .A2(n53883), .ZN(n53885) );
  XNOR2HSV1 U56814 ( .A1(n53886), .A2(n53885), .ZN(n53887) );
  XNOR2HSV1 U56815 ( .A1(n53888), .A2(n53887), .ZN(n53889) );
  XNOR2HSV1 U56816 ( .A1(n53890), .A2(n53889), .ZN(n53892) );
  BUFHSV2 U56817 ( .I(n55018), .Z(n54431) );
  CLKNAND2HSV0 U56818 ( .A1(n54946), .A2(n54716), .ZN(n53891) );
  XOR2HSV0 U56819 ( .A1(n53892), .A2(n53891), .Z(n53893) );
  XOR2HSV0 U56820 ( .A1(n53894), .A2(n53893), .Z(n53895) );
  XNOR2HSV1 U56821 ( .A1(n53896), .A2(n53895), .ZN(n53898) );
  CLKNAND2HSV0 U56822 ( .A1(n55069), .A2(n54724), .ZN(n53897) );
  XNOR2HSV1 U56823 ( .A1(n53898), .A2(n53897), .ZN(n53899) );
  XNOR2HSV1 U56824 ( .A1(n53900), .A2(n53899), .ZN(n53903) );
  INAND2HSV2 U56825 ( .A1(n55529), .B1(\pe1/got [23]), .ZN(n53902) );
  CLKNAND2HSV0 U56826 ( .A1(n55213), .A2(n53520), .ZN(n53901) );
  XOR3HSV2 U56827 ( .A1(n53903), .A2(n53902), .A3(n53901), .Z(n53904) );
  XOR2HSV0 U56828 ( .A1(n53905), .A2(n53904), .Z(n53906) );
  XOR2HSV0 U56829 ( .A1(n53907), .A2(n53906), .Z(n53910) );
  NAND2HSV2 U56830 ( .A1(n25840), .A2(n59374), .ZN(n53909) );
  NAND2HSV0 U56831 ( .A1(n40873), .A2(n55589), .ZN(n53908) );
  XOR3HSV2 U56832 ( .A1(n53910), .A2(n53909), .A3(n53908), .Z(\pe1/poht [4])
         );
  CLKNAND2HSV1 U56833 ( .A1(n55228), .A2(\pe1/got [23]), .ZN(n54025) );
  CLKNAND2HSV0 U56834 ( .A1(n55341), .A2(n40886), .ZN(n54021) );
  NAND2HSV0 U56835 ( .A1(n59422), .A2(n44530), .ZN(n54019) );
  CLKNAND2HSV1 U56836 ( .A1(n54038), .A2(n54716), .ZN(n54015) );
  NOR2HSV1 U56837 ( .A1(n53912), .A2(n53911), .ZN(n54013) );
  CLKNAND2HSV1 U56838 ( .A1(n53522), .A2(n54161), .ZN(n54011) );
  CLKNAND2HSV1 U56839 ( .A1(n54814), .A2(n54241), .ZN(n54009) );
  NOR2HSV1 U56840 ( .A1(n54040), .A2(n54884), .ZN(n54007) );
  NOR2HSV0 U56841 ( .A1(n54731), .A2(n54453), .ZN(n54005) );
  NAND2HSV0 U56842 ( .A1(n53913), .A2(n54970), .ZN(n54002) );
  NAND2HSV0 U56843 ( .A1(n54362), .A2(n55088), .ZN(n54000) );
  NOR2HSV0 U56844 ( .A1(n41566), .A2(n55227), .ZN(n53995) );
  NAND2HSV0 U56845 ( .A1(n54456), .A2(n55448), .ZN(n53991) );
  NAND2HSV0 U56846 ( .A1(n42360), .A2(n55319), .ZN(n53985) );
  NAND2HSV0 U56847 ( .A1(n54904), .A2(n54302), .ZN(n53915) );
  NAND2HSV0 U56848 ( .A1(n59990), .A2(\pe1/bq[17] ), .ZN(n53914) );
  XOR2HSV0 U56849 ( .A1(n53915), .A2(n53914), .Z(n53919) );
  NAND2HSV0 U56850 ( .A1(n41768), .A2(n55379), .ZN(n53917) );
  NAND2HSV0 U56851 ( .A1(\pe1/aot [21]), .A2(\pe1/bq[9] ), .ZN(n53916) );
  XOR2HSV0 U56852 ( .A1(n53917), .A2(n53916), .Z(n53918) );
  XOR2HSV0 U56853 ( .A1(n53919), .A2(n53918), .Z(n53928) );
  NAND2HSV0 U56854 ( .A1(n42132), .A2(n41424), .ZN(n53921) );
  NAND2HSV0 U56855 ( .A1(n54578), .A2(n54048), .ZN(n53920) );
  XOR2HSV0 U56856 ( .A1(n53921), .A2(n53920), .Z(n53926) );
  NAND2HSV0 U56857 ( .A1(\pe1/aot [16]), .A2(n54999), .ZN(n53924) );
  NAND2HSV0 U56858 ( .A1(n59730), .A2(n53922), .ZN(n53923) );
  XOR2HSV0 U56859 ( .A1(n53924), .A2(n53923), .Z(n53925) );
  XOR2HSV0 U56860 ( .A1(n53926), .A2(n53925), .Z(n53927) );
  XOR2HSV0 U56861 ( .A1(n53928), .A2(n53927), .Z(n53946) );
  NAND2HSV0 U56862 ( .A1(n40683), .A2(\pe1/bq[2] ), .ZN(n53930) );
  NAND2HSV0 U56863 ( .A1(\pe1/aot [12]), .A2(\pe1/bq[18] ), .ZN(n53929) );
  XOR2HSV0 U56864 ( .A1(n53930), .A2(n53929), .Z(n53935) );
  NAND2HSV0 U56865 ( .A1(n59389), .A2(n41771), .ZN(n53933) );
  NAND2HSV0 U56866 ( .A1(n53931), .A2(n54371), .ZN(n53932) );
  XOR2HSV0 U56867 ( .A1(n53933), .A2(n53932), .Z(n53934) );
  XOR2HSV0 U56868 ( .A1(n53935), .A2(n53934), .Z(n53944) );
  NAND2HSV0 U56869 ( .A1(n54913), .A2(n42092), .ZN(n53937) );
  XOR2HSV0 U56870 ( .A1(n53938), .A2(n53937), .Z(n53942) );
  NAND2HSV0 U56871 ( .A1(n54307), .A2(n54911), .ZN(n53940) );
  NAND2HSV0 U56872 ( .A1(n41169), .A2(\pe1/bq[8] ), .ZN(n53939) );
  XOR2HSV0 U56873 ( .A1(n53940), .A2(n53939), .Z(n53941) );
  XNOR2HSV1 U56874 ( .A1(n53942), .A2(n53941), .ZN(n53943) );
  XNOR2HSV1 U56875 ( .A1(n53944), .A2(n53943), .ZN(n53945) );
  XNOR2HSV1 U56876 ( .A1(n53946), .A2(n53945), .ZN(n53977) );
  NAND2HSV0 U56877 ( .A1(n54303), .A2(n42366), .ZN(n53948) );
  NAND2HSV0 U56878 ( .A1(\pe1/aot [4]), .A2(\pe1/bq[26] ), .ZN(n53947) );
  XOR2HSV0 U56879 ( .A1(n53948), .A2(n53947), .Z(n53953) );
  NAND2HSV0 U56880 ( .A1(n59992), .A2(n53949), .ZN(n53951) );
  NAND2HSV0 U56881 ( .A1(n55380), .A2(\pe1/bq[21] ), .ZN(n53950) );
  XOR2HSV0 U56882 ( .A1(n53951), .A2(n53950), .Z(n53952) );
  XOR2HSV0 U56883 ( .A1(n53953), .A2(n53952), .Z(n53964) );
  NAND2HSV0 U56884 ( .A1(n53954), .A2(n54274), .ZN(n53956) );
  NAND2HSV0 U56885 ( .A1(n54500), .A2(n42373), .ZN(n53955) );
  XOR2HSV0 U56886 ( .A1(n53956), .A2(n53955), .Z(n53962) );
  NOR2HSV0 U56887 ( .A1(n53957), .A2(n55185), .ZN(n53960) );
  NOR2HSV0 U56888 ( .A1(n54843), .A2(n45814), .ZN(n53959) );
  NAND2HSV2 U56889 ( .A1(\pe1/aot [14]), .A2(n54063), .ZN(n55256) );
  OAI22HSV0 U56890 ( .A1(n53960), .A2(n53959), .B1(n53958), .B2(n55256), .ZN(
        n53961) );
  XNOR2HSV1 U56891 ( .A1(n53962), .A2(n53961), .ZN(n53963) );
  XNOR2HSV1 U56892 ( .A1(n53964), .A2(n53963), .ZN(n53975) );
  NAND2HSV2 U56893 ( .A1(n55397), .A2(n54289), .ZN(n55239) );
  NOR2HSV0 U56894 ( .A1(n53965), .A2(n55239), .ZN(n53967) );
  AOI22HSV0 U56895 ( .A1(\pe1/aot [25]), .A2(n54289), .B1(\pe1/bq[20] ), .B2(
        n55093), .ZN(n53966) );
  NOR2HSV2 U56896 ( .A1(n53967), .A2(n53966), .ZN(n53969) );
  XOR2HSV0 U56897 ( .A1(n53969), .A2(n53968), .Z(n53973) );
  XOR2HSV0 U56898 ( .A1(n53971), .A2(n53970), .Z(n53972) );
  XOR2HSV0 U56899 ( .A1(n53973), .A2(n53972), .Z(n53974) );
  XNOR2HSV1 U56900 ( .A1(n53975), .A2(n53974), .ZN(n53976) );
  XNOR2HSV1 U56901 ( .A1(n53977), .A2(n53976), .ZN(n53981) );
  BUFHSV2 U56902 ( .I(n53978), .Z(n55376) );
  NAND2HSV0 U56903 ( .A1(n53979), .A2(n54455), .ZN(n53980) );
  XNOR2HSV1 U56904 ( .A1(n53981), .A2(n53980), .ZN(n53983) );
  NAND2HSV0 U56905 ( .A1(n59674), .A2(n54104), .ZN(n53982) );
  XNOR2HSV1 U56906 ( .A1(n53983), .A2(n53982), .ZN(n53984) );
  XNOR2HSV1 U56907 ( .A1(n53985), .A2(n53984), .ZN(n53987) );
  NAND2HSV0 U56908 ( .A1(n59686), .A2(n55267), .ZN(n53986) );
  XOR2HSV0 U56909 ( .A1(n53987), .A2(n53986), .Z(n53989) );
  NAND2HSV0 U56910 ( .A1(n59919), .A2(\pe1/got [5]), .ZN(n53988) );
  XOR2HSV0 U56911 ( .A1(n53989), .A2(n53988), .Z(n53990) );
  XNOR2HSV1 U56912 ( .A1(n53991), .A2(n53990), .ZN(n53993) );
  NAND2HSV0 U56913 ( .A1(n41677), .A2(n54894), .ZN(n53992) );
  XOR2HSV0 U56914 ( .A1(n53993), .A2(n53992), .Z(n53994) );
  XNOR2HSV1 U56915 ( .A1(n53995), .A2(n53994), .ZN(n53998) );
  NAND2HSV0 U56916 ( .A1(n53996), .A2(n55145), .ZN(n53997) );
  XOR2HSV0 U56917 ( .A1(n53998), .A2(n53997), .Z(n53999) );
  XNOR2HSV1 U56918 ( .A1(n54000), .A2(n53999), .ZN(n54001) );
  XNOR2HSV1 U56919 ( .A1(n54002), .A2(n54001), .ZN(n54004) );
  NAND2HSV0 U56920 ( .A1(n54521), .A2(\pe1/got [13]), .ZN(n54003) );
  XOR3HSV2 U56921 ( .A1(n54005), .A2(n54004), .A3(n54003), .Z(n54006) );
  XNOR2HSV1 U56922 ( .A1(n54007), .A2(n54006), .ZN(n54008) );
  XNOR2HSV1 U56923 ( .A1(n54009), .A2(n54008), .ZN(n54010) );
  XNOR2HSV1 U56924 ( .A1(n54011), .A2(n54010), .ZN(n54012) );
  XNOR2HSV1 U56925 ( .A1(n54013), .A2(n54012), .ZN(n54014) );
  XNOR2HSV1 U56926 ( .A1(n54015), .A2(n54014), .ZN(n54017) );
  CLKNAND2HSV0 U56927 ( .A1(n54946), .A2(\pe1/got [19]), .ZN(n54016) );
  XOR2HSV0 U56928 ( .A1(n54017), .A2(n54016), .Z(n54018) );
  XNOR2HSV1 U56929 ( .A1(n54019), .A2(n54018), .ZN(n54020) );
  XNOR2HSV1 U56930 ( .A1(n54021), .A2(n54020), .ZN(n54023) );
  CLKNAND2HSV0 U56931 ( .A1(n55069), .A2(n54160), .ZN(n54022) );
  XNOR2HSV1 U56932 ( .A1(n54023), .A2(n54022), .ZN(n54024) );
  XNOR2HSV1 U56933 ( .A1(n54025), .A2(n54024), .ZN(n54028) );
  INAND2HSV2 U56934 ( .A1(n55529), .B1(n53520), .ZN(n54027) );
  CLKNAND2HSV0 U56935 ( .A1(n55213), .A2(\pe1/got [25]), .ZN(n54026) );
  XOR3HSV2 U56936 ( .A1(n54028), .A2(n54027), .A3(n54026), .Z(n54030) );
  CLKNAND2HSV0 U56937 ( .A1(n55289), .A2(n41689), .ZN(n54029) );
  XOR2HSV0 U56938 ( .A1(n54030), .A2(n54029), .Z(n54031) );
  XOR2HSV0 U56939 ( .A1(n54032), .A2(n54031), .Z(n54036) );
  NAND2HSV2 U56940 ( .A1(n55569), .A2(\pe1/got [28]), .ZN(n54035) );
  XOR3HSV2 U56941 ( .A1(n54036), .A2(n54035), .A3(n54034), .Z(\pe1/poht [3])
         );
  CLKNAND2HSV0 U56942 ( .A1(n55488), .A2(\pe1/got [25]), .ZN(n54153) );
  CLKNAND2HSV1 U56943 ( .A1(n55489), .A2(n40913), .ZN(n54151) );
  CLKNAND2HSV1 U56944 ( .A1(n53792), .A2(n54724), .ZN(n54145) );
  NAND2HSV0 U56945 ( .A1(n59995), .A2(n55341), .ZN(n54141) );
  CLKNHSV0 U56946 ( .I(n54037), .ZN(n55375) );
  NAND2HSV0 U56947 ( .A1(n55375), .A2(n54716), .ZN(n54139) );
  CLKNAND2HSV1 U56948 ( .A1(n54038), .A2(n54161), .ZN(n54134) );
  NOR2HSV1 U56949 ( .A1(n53912), .A2(n54039), .ZN(n54132) );
  CLKNAND2HSV0 U56950 ( .A1(n55230), .A2(n54969), .ZN(n54130) );
  CLKNAND2HSV0 U56951 ( .A1(n53392), .A2(\pe1/got [13]), .ZN(n54128) );
  NOR2HSV2 U56952 ( .A1(n54040), .A2(n54453), .ZN(n54126) );
  NOR2HSV0 U56953 ( .A1(n54815), .A2(n54636), .ZN(n54124) );
  CLKNAND2HSV0 U56954 ( .A1(n54557), .A2(\pe1/got [9]), .ZN(n54121) );
  NAND2HSV0 U56955 ( .A1(n54041), .A2(\pe1/got [8]), .ZN(n54119) );
  NOR2HSV0 U56956 ( .A1(n41301), .A2(n55369), .ZN(n54114) );
  NAND2HSV0 U56957 ( .A1(n54456), .A2(n55267), .ZN(n54110) );
  CLKNAND2HSV0 U56958 ( .A1(n41144), .A2(n54455), .ZN(n54103) );
  NAND2HSV0 U56959 ( .A1(n55433), .A2(n54318), .ZN(n54043) );
  NAND2HSV0 U56960 ( .A1(n54913), .A2(n54995), .ZN(n54042) );
  XOR2HSV0 U56961 ( .A1(n54043), .A2(n54042), .Z(n54047) );
  NAND2HSV0 U56962 ( .A1(n54188), .A2(n42092), .ZN(n54045) );
  NAND2HSV0 U56963 ( .A1(\pe1/aot [14]), .A2(n54999), .ZN(n54044) );
  XOR2HSV0 U56964 ( .A1(n54045), .A2(n54044), .Z(n54046) );
  XOR2HSV0 U56965 ( .A1(n54047), .A2(n54046), .Z(n54056) );
  NAND2HSV0 U56966 ( .A1(n59992), .A2(n54302), .ZN(n54050) );
  NAND2HSV0 U56967 ( .A1(n54303), .A2(n54048), .ZN(n54049) );
  XOR2HSV0 U56968 ( .A1(n54050), .A2(n54049), .Z(n54054) );
  NAND2HSV0 U56969 ( .A1(n54364), .A2(\pe1/bq[9] ), .ZN(n54052) );
  NAND2HSV0 U56970 ( .A1(n55186), .A2(n54179), .ZN(n54051) );
  XOR2HSV0 U56971 ( .A1(n54052), .A2(n54051), .Z(n54053) );
  XOR2HSV0 U56972 ( .A1(n54054), .A2(n54053), .Z(n54055) );
  XOR2HSV0 U56973 ( .A1(n54056), .A2(n54055), .Z(n54073) );
  NAND2HSV0 U56974 ( .A1(n42399), .A2(n55379), .ZN(n54058) );
  NAND2HSV0 U56975 ( .A1(n54497), .A2(n55241), .ZN(n54057) );
  XOR2HSV0 U56976 ( .A1(n54058), .A2(n54057), .Z(n54062) );
  NAND2HSV0 U56977 ( .A1(n54578), .A2(\pe1/bq[21] ), .ZN(n54060) );
  NAND2HSV0 U56978 ( .A1(n59730), .A2(n41644), .ZN(n54059) );
  XOR2HSV0 U56979 ( .A1(n54060), .A2(n54059), .Z(n54061) );
  XOR2HSV0 U56980 ( .A1(n54062), .A2(n54061), .Z(n54071) );
  NAND2HSV0 U56981 ( .A1(n59389), .A2(n41173), .ZN(n54065) );
  NAND2HSV2 U56982 ( .A1(n59986), .A2(n54063), .ZN(n54064) );
  XOR2HSV0 U56983 ( .A1(n54065), .A2(n54064), .Z(n54069) );
  NAND2HSV0 U56984 ( .A1(n54904), .A2(n42238), .ZN(n54067) );
  NAND2HSV0 U56985 ( .A1(\pe1/aot [24]), .A2(n54371), .ZN(n54066) );
  XOR2HSV0 U56986 ( .A1(n54067), .A2(n54066), .Z(n54068) );
  XOR2HSV0 U56987 ( .A1(n54069), .A2(n54068), .Z(n54070) );
  XOR2HSV0 U56988 ( .A1(n54071), .A2(n54070), .Z(n54072) );
  XOR2HSV0 U56989 ( .A1(n54073), .A2(n54072), .Z(n54101) );
  NOR2HSV0 U56990 ( .A1(n53672), .A2(n54973), .ZN(n54075) );
  CLKNAND2HSV0 U56991 ( .A1(n44541), .A2(n55110), .ZN(n55255) );
  OAI22HSV0 U56992 ( .A1(n54076), .A2(n54075), .B1(n54074), .B2(n55255), .ZN(
        n54082) );
  CLKNAND2HSV1 U56993 ( .A1(\pe1/aot [12]), .A2(n54911), .ZN(n54976) );
  NOR2HSV0 U56994 ( .A1(n54077), .A2(n54976), .ZN(n54080) );
  AOI22HSV0 U56995 ( .A1(n54078), .A2(n55231), .B1(n54836), .B2(\pe1/aot [12]), 
        .ZN(n54079) );
  NOR2HSV1 U56996 ( .A1(n54080), .A2(n54079), .ZN(n54081) );
  XOR2HSV0 U56997 ( .A1(n54082), .A2(n54081), .Z(n54090) );
  NAND2HSV0 U56998 ( .A1(n54743), .A2(n41771), .ZN(n54086) );
  INHSV2 U56999 ( .I(n55524), .ZN(n54363) );
  NAND2HSV2 U57000 ( .A1(n54363), .A2(n54083), .ZN(n55598) );
  NOR2HSV0 U57001 ( .A1(n54084), .A2(n55598), .ZN(n54085) );
  AOI21HSV2 U57002 ( .A1(n54306), .A2(n54086), .B(n54085), .ZN(n54088) );
  XNOR2HSV1 U57003 ( .A1(n54088), .A2(n54087), .ZN(n54089) );
  XNOR2HSV1 U57004 ( .A1(n54090), .A2(n54089), .ZN(n54099) );
  NAND2HSV0 U57005 ( .A1(n54288), .A2(n54289), .ZN(n54092) );
  NAND2HSV0 U57006 ( .A1(n54669), .A2(n53798), .ZN(n54091) );
  XOR2HSV0 U57007 ( .A1(n54092), .A2(n54091), .Z(n54097) );
  NOR2HSV0 U57008 ( .A1(n41944), .A2(n54093), .ZN(n54095) );
  NAND2HSV0 U57009 ( .A1(n55093), .A2(\pe1/bq[18] ), .ZN(n54094) );
  XOR2HSV0 U57010 ( .A1(n54095), .A2(n54094), .Z(n54096) );
  XOR2HSV0 U57011 ( .A1(n54097), .A2(n54096), .Z(n54098) );
  XOR2HSV0 U57012 ( .A1(n54099), .A2(n54098), .Z(n54100) );
  XNOR2HSV1 U57013 ( .A1(n54101), .A2(n54100), .ZN(n54102) );
  XNOR2HSV1 U57014 ( .A1(n54103), .A2(n54102), .ZN(n54106) );
  NAND2HSV0 U57015 ( .A1(n59686), .A2(n54104), .ZN(n54105) );
  XOR2HSV0 U57016 ( .A1(n54106), .A2(n54105), .Z(n54108) );
  NAND2HSV0 U57017 ( .A1(n59919), .A2(n55319), .ZN(n54107) );
  XOR2HSV0 U57018 ( .A1(n54108), .A2(n54107), .Z(n54109) );
  XNOR2HSV1 U57019 ( .A1(n54110), .A2(n54109), .ZN(n54112) );
  NAND2HSV0 U57020 ( .A1(n29773), .A2(\pe1/got [5]), .ZN(n54111) );
  XOR2HSV0 U57021 ( .A1(n54112), .A2(n54111), .Z(n54113) );
  XNOR2HSV1 U57022 ( .A1(n54114), .A2(n54113), .ZN(n54117) );
  NAND2HSV0 U57023 ( .A1(n54115), .A2(n54894), .ZN(n54116) );
  XOR2HSV0 U57024 ( .A1(n54117), .A2(n54116), .Z(n54118) );
  XNOR2HSV1 U57025 ( .A1(n54119), .A2(n54118), .ZN(n54120) );
  XNOR2HSV1 U57026 ( .A1(n54121), .A2(n54120), .ZN(n54123) );
  NAND2HSV0 U57027 ( .A1(n54521), .A2(\pe1/got [11]), .ZN(n54122) );
  XOR3HSV2 U57028 ( .A1(n54124), .A2(n54123), .A3(n54122), .Z(n54125) );
  XNOR2HSV1 U57029 ( .A1(n54126), .A2(n54125), .ZN(n54127) );
  XNOR2HSV1 U57030 ( .A1(n54128), .A2(n54127), .ZN(n54129) );
  XNOR2HSV1 U57031 ( .A1(n54130), .A2(n54129), .ZN(n54131) );
  XNOR2HSV1 U57032 ( .A1(n54132), .A2(n54131), .ZN(n54133) );
  XNOR2HSV1 U57033 ( .A1(n54134), .A2(n54133), .ZN(n54137) );
  CLKNAND2HSV0 U57034 ( .A1(n54946), .A2(n54135), .ZN(n54136) );
  XOR2HSV0 U57035 ( .A1(n54137), .A2(n54136), .Z(n54138) );
  XNOR2HSV1 U57036 ( .A1(n54139), .A2(n54138), .ZN(n54140) );
  XNOR2HSV1 U57037 ( .A1(n54141), .A2(n54140), .ZN(n54143) );
  NAND2HSV0 U57038 ( .A1(n54541), .A2(n44530), .ZN(n54142) );
  XNOR2HSV1 U57039 ( .A1(n54143), .A2(n54142), .ZN(n54144) );
  XNOR2HSV1 U57040 ( .A1(n54145), .A2(n54144), .ZN(n54149) );
  INHSV2 U57041 ( .I(n54146), .ZN(n55562) );
  INAND2HSV2 U57042 ( .A1(n55562), .B1(n54160), .ZN(n54148) );
  CLKNAND2HSV0 U57043 ( .A1(n55476), .A2(\pe1/got [23]), .ZN(n54147) );
  XOR3HSV2 U57044 ( .A1(n54149), .A2(n54148), .A3(n54147), .Z(n54150) );
  XOR2HSV0 U57045 ( .A1(n54151), .A2(n54150), .Z(n54152) );
  XOR2HSV0 U57046 ( .A1(n54153), .A2(n54152), .Z(n54158) );
  NAND2HSV2 U57047 ( .A1(n25839), .A2(n40605), .ZN(n54157) );
  INHSV2 U57048 ( .I(n54154), .ZN(n54155) );
  XOR3HSV2 U57049 ( .A1(n54158), .A2(n54157), .A3(n54156), .Z(\pe1/poht [5])
         );
  NAND2HSV0 U57050 ( .A1(n55488), .A2(\pe1/got [23]), .ZN(n54259) );
  CLKNAND2HSV1 U57051 ( .A1(n55543), .A2(n54160), .ZN(n54257) );
  INHSV2 U57052 ( .I(n55162), .ZN(n55228) );
  NAND2HSV2 U57053 ( .A1(n55228), .A2(n59995), .ZN(n54252) );
  NAND2HSV0 U57054 ( .A1(n59521), .A2(n54965), .ZN(n54247) );
  NAND2HSV0 U57055 ( .A1(n55375), .A2(n54161), .ZN(n54245) );
  NAND2HSV0 U57056 ( .A1(n53521), .A2(n54969), .ZN(n54240) );
  NOR2HSV2 U57057 ( .A1(n55090), .A2(n54957), .ZN(n54238) );
  CLKNAND2HSV0 U57058 ( .A1(n55230), .A2(\pe1/got [12]), .ZN(n54236) );
  CLKNAND2HSV1 U57059 ( .A1(n53392), .A2(\pe1/got [11]), .ZN(n54234) );
  INHSV2 U57060 ( .I(n53657), .ZN(n54454) );
  NOR2HSV0 U57061 ( .A1(n54454), .A2(n54636), .ZN(n54232) );
  NOR2HSV0 U57062 ( .A1(n54731), .A2(n55227), .ZN(n54230) );
  CLKNAND2HSV0 U57063 ( .A1(n54557), .A2(\pe1/got [7]), .ZN(n54227) );
  NAND2HSV0 U57064 ( .A1(n54162), .A2(\pe1/got [6]), .ZN(n54225) );
  NOR2HSV0 U57065 ( .A1(n42438), .A2(n55444), .ZN(n54221) );
  NAND2HSV0 U57066 ( .A1(n54456), .A2(n59756), .ZN(n54217) );
  NAND2HSV0 U57067 ( .A1(n59919), .A2(n54455), .ZN(n54215) );
  NAND2HSV0 U57068 ( .A1(n54303), .A2(\pe1/bq[21] ), .ZN(n54164) );
  NAND2HSV0 U57069 ( .A1(\pe1/aot [6]), .A2(n54565), .ZN(n54163) );
  XOR2HSV0 U57070 ( .A1(n54164), .A2(n54163), .Z(n54168) );
  NAND2HSV0 U57071 ( .A1(\pe1/aot [21]), .A2(\pe1/bq[5] ), .ZN(n54166) );
  NAND2HSV0 U57072 ( .A1(\pe1/aot [14]), .A2(\pe1/bq[12] ), .ZN(n54165) );
  XOR2HSV0 U57073 ( .A1(n54166), .A2(n54165), .Z(n54167) );
  XOR2HSV0 U57074 ( .A1(n54168), .A2(n54167), .Z(n54176) );
  NAND2HSV0 U57075 ( .A1(n54497), .A2(\pe1/bq[9] ), .ZN(n54170) );
  NAND2HSV0 U57076 ( .A1(n54364), .A2(n54274), .ZN(n54169) );
  XOR2HSV0 U57077 ( .A1(n54170), .A2(n54169), .Z(n54174) );
  NAND2HSV0 U57078 ( .A1(n54913), .A2(n48380), .ZN(n54172) );
  NAND2HSV0 U57079 ( .A1(n59389), .A2(\pe1/bq[23] ), .ZN(n54171) );
  XOR2HSV0 U57080 ( .A1(n54172), .A2(n54171), .Z(n54173) );
  XNOR2HSV1 U57081 ( .A1(n54174), .A2(n54173), .ZN(n54175) );
  XNOR2HSV1 U57082 ( .A1(n54176), .A2(n54175), .ZN(n54197) );
  NAND2HSV0 U57083 ( .A1(n54363), .A2(n41173), .ZN(n54178) );
  NAND2HSV0 U57084 ( .A1(\pe1/aot [16]), .A2(n54847), .ZN(n54177) );
  XOR2HSV0 U57085 ( .A1(n54178), .A2(n54177), .Z(n54183) );
  NAND2HSV0 U57086 ( .A1(n55103), .A2(n54179), .ZN(n54181) );
  NAND2HSV0 U57087 ( .A1(n42093), .A2(n54911), .ZN(n54180) );
  XOR2HSV0 U57088 ( .A1(n54181), .A2(n54180), .Z(n54182) );
  XNOR2HSV1 U57089 ( .A1(n54183), .A2(n54182), .ZN(n54195) );
  NAND2HSV2 U57090 ( .A1(\pe1/aot [2]), .A2(n54988), .ZN(n55607) );
  OAI21HSV0 U57091 ( .A1(n55504), .A2(n54185), .B(n54184), .ZN(n54186) );
  OAI21HSV0 U57092 ( .A1(n54187), .A2(n55607), .B(n54186), .ZN(n54193) );
  NAND2HSV2 U57093 ( .A1(n54371), .A2(n54188), .ZN(n55180) );
  NOR2HSV0 U57094 ( .A1(n54189), .A2(n55180), .ZN(n54191) );
  AOI22HSV0 U57095 ( .A1(n54078), .A2(n55544), .B1(n54995), .B2(n54818), .ZN(
        n54190) );
  NOR2HSV1 U57096 ( .A1(n54191), .A2(n54190), .ZN(n54192) );
  XOR2HSV0 U57097 ( .A1(n54193), .A2(n54192), .Z(n54194) );
  XNOR2HSV1 U57098 ( .A1(n54195), .A2(n54194), .ZN(n54196) );
  XNOR2HSV1 U57099 ( .A1(n54197), .A2(n54196), .ZN(n54213) );
  NAND2HSV0 U57100 ( .A1(n55113), .A2(n54999), .ZN(n54483) );
  NOR2HSV0 U57101 ( .A1(n41974), .A2(n53834), .ZN(n54309) );
  NOR2HSV0 U57102 ( .A1(n55307), .A2(n41963), .ZN(n54199) );
  NAND2HSV2 U57103 ( .A1(n54578), .A2(n55605), .ZN(n55507) );
  OAI22HSV0 U57104 ( .A1(n54309), .A2(n54199), .B1(n54198), .B2(n55507), .ZN(
        n54203) );
  NAND2HSV0 U57105 ( .A1(n54288), .A2(n54668), .ZN(n54201) );
  CLKNAND2HSV0 U57106 ( .A1(n54904), .A2(\pe1/bq[18] ), .ZN(n54200) );
  XOR2HSV0 U57107 ( .A1(n54201), .A2(n54200), .Z(n54202) );
  XOR3HSV1 U57108 ( .A1(n54483), .A2(n54203), .A3(n54202), .Z(n54211) );
  NAND2HSV0 U57109 ( .A1(n55433), .A2(n54465), .ZN(n54205) );
  NAND2HSV0 U57110 ( .A1(n42132), .A2(n55241), .ZN(n54204) );
  XOR2HSV0 U57111 ( .A1(n54205), .A2(n54204), .Z(n54209) );
  NAND2HSV0 U57112 ( .A1(n55397), .A2(\pe1/bq[16] ), .ZN(n54207) );
  NAND2HSV0 U57113 ( .A1(n42399), .A2(n53798), .ZN(n54206) );
  XOR2HSV0 U57114 ( .A1(n54207), .A2(n54206), .Z(n54208) );
  XOR2HSV0 U57115 ( .A1(n54209), .A2(n54208), .Z(n54210) );
  XOR2HSV0 U57116 ( .A1(n54211), .A2(n54210), .Z(n54212) );
  XNOR2HSV1 U57117 ( .A1(n54213), .A2(n54212), .ZN(n54214) );
  XNOR2HSV1 U57118 ( .A1(n54215), .A2(n54214), .ZN(n54216) );
  XNOR2HSV1 U57119 ( .A1(n54217), .A2(n54216), .ZN(n54219) );
  NAND2HSV0 U57120 ( .A1(n29762), .A2(\pe1/got [3]), .ZN(n54218) );
  XOR2HSV0 U57121 ( .A1(n54219), .A2(n54218), .Z(n54220) );
  XNOR2HSV1 U57122 ( .A1(n54221), .A2(n54220), .ZN(n54223) );
  NAND2HSV0 U57123 ( .A1(n54513), .A2(n55475), .ZN(n54222) );
  XOR2HSV0 U57124 ( .A1(n54223), .A2(n54222), .Z(n54224) );
  XNOR2HSV1 U57125 ( .A1(n54225), .A2(n54224), .ZN(n54226) );
  XNOR2HSV1 U57126 ( .A1(n54227), .A2(n54226), .ZN(n54229) );
  NAND2HSV0 U57127 ( .A1(n54521), .A2(\pe1/got [9]), .ZN(n54228) );
  XOR3HSV2 U57128 ( .A1(n54230), .A2(n54229), .A3(n54228), .Z(n54231) );
  XNOR2HSV1 U57129 ( .A1(n54232), .A2(n54231), .ZN(n54233) );
  XNOR2HSV1 U57130 ( .A1(n54234), .A2(n54233), .ZN(n54235) );
  XNOR2HSV1 U57131 ( .A1(n54236), .A2(n54235), .ZN(n54237) );
  XNOR2HSV1 U57132 ( .A1(n54238), .A2(n54237), .ZN(n54239) );
  XNOR2HSV1 U57133 ( .A1(n54240), .A2(n54239), .ZN(n54243) );
  CLKNAND2HSV0 U57134 ( .A1(n54946), .A2(n54241), .ZN(n54242) );
  XOR2HSV0 U57135 ( .A1(n54243), .A2(n54242), .Z(n54244) );
  XNOR2HSV1 U57136 ( .A1(n54245), .A2(n54244), .ZN(n54246) );
  XNOR2HSV1 U57137 ( .A1(n54247), .A2(n54246), .ZN(n54250) );
  NAND2HSV0 U57138 ( .A1(n54541), .A2(n54716), .ZN(n54249) );
  XNOR2HSV1 U57139 ( .A1(n54250), .A2(n54249), .ZN(n54251) );
  XNOR2HSV1 U57140 ( .A1(n54252), .A2(n54251), .ZN(n54255) );
  INAND2HSV2 U57141 ( .A1(n55562), .B1(n44530), .ZN(n54254) );
  INHSV2 U57142 ( .I(n55213), .ZN(n54361) );
  INHSV3 U57143 ( .I(n54361), .ZN(n55427) );
  CLKNAND2HSV1 U57144 ( .A1(n55427), .A2(n54724), .ZN(n54253) );
  XOR3HSV2 U57145 ( .A1(n54255), .A2(n54254), .A3(n54253), .Z(n54256) );
  XOR2HSV0 U57146 ( .A1(n54257), .A2(n54256), .Z(n54258) );
  XOR2HSV0 U57147 ( .A1(n54259), .A2(n54258), .Z(n54262) );
  NAND2HSV2 U57148 ( .A1(n55569), .A2(\pe1/got [24]), .ZN(n54261) );
  XOR3HSV2 U57149 ( .A1(n54262), .A2(n54261), .A3(n54260), .Z(\pe1/poht [7])
         );
  NAND2HSV0 U57150 ( .A1(n59422), .A2(n54965), .ZN(n54360) );
  INHSV4 U57151 ( .I(n54263), .ZN(n55222) );
  NAND2HSV0 U57152 ( .A1(n42085), .A2(n55222), .ZN(n54356) );
  NOR2HSV1 U57153 ( .A1(n55090), .A2(n54884), .ZN(n54354) );
  CLKNAND2HSV0 U57154 ( .A1(n55230), .A2(n42155), .ZN(n54352) );
  CLKNAND2HSV1 U57155 ( .A1(n54814), .A2(\pe1/got [12]), .ZN(n54350) );
  NOR2HSV2 U57156 ( .A1(n54454), .A2(n55082), .ZN(n54348) );
  NOR2HSV0 U57157 ( .A1(n54731), .A2(n55163), .ZN(n54346) );
  NAND2HSV0 U57158 ( .A1(n54557), .A2(\pe1/got [8]), .ZN(n54343) );
  NAND2HSV0 U57159 ( .A1(n54264), .A2(\pe1/got [7]), .ZN(n54341) );
  NOR2HSV0 U57160 ( .A1(n42438), .A2(n55542), .ZN(n54337) );
  NAND2HSV0 U57161 ( .A1(n54265), .A2(n59756), .ZN(n54332) );
  NAND2HSV0 U57162 ( .A1(n59686), .A2(n54455), .ZN(n54330) );
  NAND2HSV0 U57163 ( .A1(n54818), .A2(\pe1/bq[18] ), .ZN(n54267) );
  NAND2HSV0 U57164 ( .A1(n42132), .A2(n42373), .ZN(n54266) );
  XOR2HSV0 U57165 ( .A1(n54267), .A2(n54266), .Z(n54271) );
  NAND2HSV0 U57166 ( .A1(n55093), .A2(n54995), .ZN(n54269) );
  NAND2HSV0 U57167 ( .A1(n54662), .A2(\pe1/bq[16] ), .ZN(n54268) );
  XOR2HSV0 U57168 ( .A1(n54269), .A2(n54268), .Z(n54270) );
  XOR2HSV0 U57169 ( .A1(n54271), .A2(n54270), .Z(n54280) );
  NAND2HSV0 U57170 ( .A1(n53812), .A2(n48380), .ZN(n54273) );
  NAND2HSV0 U57171 ( .A1(n54363), .A2(n41644), .ZN(n54272) );
  XOR2HSV0 U57172 ( .A1(n54273), .A2(n54272), .Z(n54278) );
  NAND2HSV0 U57173 ( .A1(n59737), .A2(n53798), .ZN(n54276) );
  NAND2HSV0 U57174 ( .A1(n42093), .A2(n54274), .ZN(n54275) );
  XOR2HSV0 U57175 ( .A1(n54276), .A2(n54275), .Z(n54277) );
  XOR2HSV0 U57176 ( .A1(n54278), .A2(n54277), .Z(n54279) );
  XOR2HSV0 U57177 ( .A1(n54280), .A2(n54279), .Z(n54301) );
  NAND2HSV0 U57178 ( .A1(n55103), .A2(n41641), .ZN(n54283) );
  NAND2HSV0 U57179 ( .A1(n54497), .A2(n54847), .ZN(n54282) );
  XOR2HSV0 U57180 ( .A1(n54283), .A2(n54282), .Z(n54287) );
  NAND2HSV0 U57181 ( .A1(n59992), .A2(\pe1/bq[21] ), .ZN(n54285) );
  NAND2HSV0 U57182 ( .A1(n54904), .A2(n42092), .ZN(n54284) );
  XOR2HSV0 U57183 ( .A1(n54285), .A2(n54284), .Z(n54286) );
  XNOR2HSV1 U57184 ( .A1(n54287), .A2(n54286), .ZN(n54299) );
  NAND2HSV0 U57185 ( .A1(n54288), .A2(n54371), .ZN(n54291) );
  NAND2HSV0 U57186 ( .A1(n54078), .A2(n54289), .ZN(n54290) );
  XOR2HSV0 U57187 ( .A1(n54291), .A2(n54290), .Z(n54297) );
  NOR2HSV0 U57188 ( .A1(n41944), .A2(n55185), .ZN(n54740) );
  AOI22HSV0 U57189 ( .A1(n54293), .A2(n54292), .B1(n54663), .B2(\pe1/bq[6] ), 
        .ZN(n54294) );
  AOI21HSV0 U57190 ( .A1(n54295), .A2(n54740), .B(n54294), .ZN(n54296) );
  XNOR2HSV1 U57191 ( .A1(n54297), .A2(n54296), .ZN(n54298) );
  XNOR2HSV1 U57192 ( .A1(n54299), .A2(n54298), .ZN(n54300) );
  XNOR2HSV1 U57193 ( .A1(n54301), .A2(n54300), .ZN(n54328) );
  NAND2HSV0 U57194 ( .A1(n55433), .A2(\pe1/bq[23] ), .ZN(n54305) );
  NAND2HSV0 U57195 ( .A1(n54303), .A2(n54302), .ZN(n54304) );
  XOR2HSV0 U57196 ( .A1(n54305), .A2(n54304), .Z(n54326) );
  CLKNHSV0 U57197 ( .I(n54306), .ZN(n54310) );
  AOI22HSV0 U57198 ( .A1(n41743), .A2(n55451), .B1(n54307), .B2(n55518), .ZN(
        n54308) );
  AOI21HSV2 U57199 ( .A1(n54310), .A2(n54309), .B(n54308), .ZN(n54315) );
  NOR2HSV0 U57200 ( .A1(n54843), .A2(n48030), .ZN(n54493) );
  AOI22HSV0 U57201 ( .A1(\pe1/aot [16]), .A2(n54311), .B1(\pe1/aot [14]), .B2(
        n41645), .ZN(n54312) );
  AOI21HSV1 U57202 ( .A1(n54493), .A2(n54313), .B(n54312), .ZN(n54314) );
  XOR2HSV0 U57203 ( .A1(n54315), .A2(n54314), .Z(n54325) );
  NAND2HSV0 U57204 ( .A1(n42399), .A2(\pe1/bq[9] ), .ZN(n54317) );
  NAND2HSV0 U57205 ( .A1(n54578), .A2(n42238), .ZN(n54316) );
  XOR2HSV0 U57206 ( .A1(n54317), .A2(n54316), .Z(n54323) );
  NAND2HSV0 U57207 ( .A1(n59389), .A2(n54318), .ZN(n54321) );
  NAND2HSV0 U57208 ( .A1(n55595), .A2(n54319), .ZN(n54320) );
  XOR2HSV0 U57209 ( .A1(n54321), .A2(n54320), .Z(n54322) );
  XOR2HSV0 U57210 ( .A1(n54323), .A2(n54322), .Z(n54324) );
  XOR3HSV2 U57211 ( .A1(n54326), .A2(n54325), .A3(n54324), .Z(n54327) );
  XNOR2HSV1 U57212 ( .A1(n54328), .A2(n54327), .ZN(n54329) );
  XNOR2HSV1 U57213 ( .A1(n54330), .A2(n54329), .ZN(n54331) );
  XOR2HSV0 U57214 ( .A1(n54332), .A2(n54331), .Z(n54335) );
  NAND2HSV0 U57215 ( .A1(n54456), .A2(\pe1/got [3]), .ZN(n54334) );
  NAND2HSV0 U57216 ( .A1(n29763), .A2(n55410), .ZN(n54333) );
  XOR3HSV2 U57217 ( .A1(n54335), .A2(n54334), .A3(n54333), .Z(n54336) );
  XNOR2HSV1 U57218 ( .A1(n54337), .A2(n54336), .ZN(n54339) );
  NAND2HSV0 U57219 ( .A1(n54513), .A2(\pe1/got [6]), .ZN(n54338) );
  XOR2HSV0 U57220 ( .A1(n54339), .A2(n54338), .Z(n54340) );
  XNOR2HSV1 U57221 ( .A1(n54341), .A2(n54340), .ZN(n54342) );
  XNOR2HSV1 U57222 ( .A1(n54343), .A2(n54342), .ZN(n54345) );
  NOR2HSV0 U57223 ( .A1(n54691), .A2(n54636), .ZN(n54344) );
  XOR3HSV2 U57224 ( .A1(n54346), .A2(n54345), .A3(n54344), .Z(n54347) );
  XNOR2HSV1 U57225 ( .A1(n54348), .A2(n54347), .ZN(n54349) );
  XNOR2HSV1 U57226 ( .A1(n54350), .A2(n54349), .ZN(n54351) );
  XNOR2HSV1 U57227 ( .A1(n54352), .A2(n54351), .ZN(n54353) );
  XOR2HSV0 U57228 ( .A1(n54354), .A2(n54353), .Z(n54355) );
  XNOR2HSV1 U57229 ( .A1(n54356), .A2(n54355), .ZN(n54358) );
  CLKNAND2HSV0 U57230 ( .A1(n54946), .A2(\pe1/got [16]), .ZN(n54357) );
  XOR2HSV0 U57231 ( .A1(n54358), .A2(n54357), .Z(n54359) );
  CLKNAND2HSV0 U57232 ( .A1(n55541), .A2(n54724), .ZN(n54448) );
  CLKNAND2HSV1 U57233 ( .A1(n53792), .A2(n59996), .ZN(n54441) );
  NAND2HSV0 U57234 ( .A1(n59521), .A2(n55222), .ZN(n54437) );
  NAND2HSV0 U57235 ( .A1(n55375), .A2(n54969), .ZN(n54435) );
  NAND2HSV0 U57236 ( .A1(n54813), .A2(\pe1/got [12]), .ZN(n54430) );
  NOR2HSV1 U57237 ( .A1(n53912), .A2(n55082), .ZN(n54428) );
  CLKNAND2HSV0 U57238 ( .A1(n55230), .A2(n55088), .ZN(n54426) );
  NAND2HSV0 U57239 ( .A1(n59592), .A2(n44605), .ZN(n54424) );
  NOR2HSV2 U57240 ( .A1(n54454), .A2(n55227), .ZN(n54422) );
  NOR2HSV1 U57241 ( .A1(n54815), .A2(n55369), .ZN(n54420) );
  NAND2HSV0 U57242 ( .A1(n54557), .A2(\pe1/got [5]), .ZN(n54417) );
  NAND2HSV0 U57243 ( .A1(n54362), .A2(n55410), .ZN(n54415) );
  NOR2HSV0 U57244 ( .A1(n41566), .A2(n55575), .ZN(n54411) );
  NAND2HSV0 U57245 ( .A1(n29763), .A2(n54455), .ZN(n54409) );
  NAND2HSV0 U57246 ( .A1(n54363), .A2(\pe1/bq[23] ), .ZN(n54366) );
  NAND2HSV0 U57247 ( .A1(n54364), .A2(\pe1/bq[5] ), .ZN(n54365) );
  XOR2HSV0 U57248 ( .A1(n54366), .A2(n54365), .Z(n54370) );
  NAND2HSV0 U57249 ( .A1(n59991), .A2(n41641), .ZN(n54368) );
  NAND2HSV0 U57250 ( .A1(n54497), .A2(n55505), .ZN(n54367) );
  XOR2HSV0 U57251 ( .A1(n54368), .A2(n54367), .Z(n54369) );
  XOR2HSV0 U57252 ( .A1(n54370), .A2(n54369), .Z(n54379) );
  NAND2HSV0 U57253 ( .A1(n42093), .A2(n54371), .ZN(n54373) );
  NAND2HSV0 U57254 ( .A1(n42399), .A2(\pe1/bq[6] ), .ZN(n54372) );
  XOR2HSV0 U57255 ( .A1(n54373), .A2(n54372), .Z(n54377) );
  NOR2HSV0 U57256 ( .A1(n54843), .A2(n53723), .ZN(n54375) );
  NAND2HSV0 U57257 ( .A1(n54578), .A2(\pe1/bq[17] ), .ZN(n54374) );
  XOR2HSV0 U57258 ( .A1(n54375), .A2(n54374), .Z(n54376) );
  XOR2HSV0 U57259 ( .A1(n54377), .A2(n54376), .Z(n54378) );
  XOR2HSV0 U57260 ( .A1(n54379), .A2(n54378), .Z(n54390) );
  NOR2HSV0 U57261 ( .A1(n54901), .A2(n41963), .ZN(n54492) );
  NOR2HSV0 U57262 ( .A1(n55430), .A2(n41512), .ZN(n54640) );
  AOI22HSV0 U57263 ( .A1(n55492), .A2(\pe1/bq[18] ), .B1(\pe1/bq[19] ), .B2(
        n59993), .ZN(n54380) );
  AOI21HSV2 U57264 ( .A1(n54492), .A2(n54640), .B(n54380), .ZN(n54388) );
  NAND2HSV0 U57265 ( .A1(n54078), .A2(n55605), .ZN(n54382) );
  NAND2HSV0 U57266 ( .A1(n53954), .A2(n54988), .ZN(n54381) );
  XOR2HSV0 U57267 ( .A1(n54382), .A2(n54381), .Z(n54387) );
  NOR2HSV0 U57268 ( .A1(n55504), .A2(n55385), .ZN(n55342) );
  AOI22HSV0 U57269 ( .A1(n55186), .A2(\pe1/bq[9] ), .B1(n54465), .B2(n59730), 
        .ZN(n54383) );
  AOI21HSV0 U57270 ( .A1(n55342), .A2(n54384), .B(n54383), .ZN(n54385) );
  CLKNAND2HSV1 U57271 ( .A1(n54662), .A2(n54179), .ZN(n54482) );
  XNOR2HSV1 U57272 ( .A1(n54385), .A2(n54482), .ZN(n54386) );
  XOR3HSV2 U57273 ( .A1(n54388), .A2(n54387), .A3(n54386), .Z(n54389) );
  XNOR2HSV1 U57274 ( .A1(n54390), .A2(n54389), .ZN(n54407) );
  NAND2HSV0 U57275 ( .A1(n55433), .A2(n54565), .ZN(n54392) );
  NAND2HSV0 U57276 ( .A1(n55103), .A2(n55241), .ZN(n54391) );
  XOR2HSV0 U57277 ( .A1(n54392), .A2(n54391), .Z(n54396) );
  NAND2HSV0 U57278 ( .A1(\pe1/aot [16]), .A2(n55501), .ZN(n54394) );
  NAND2HSV0 U57279 ( .A1(n55113), .A2(\pe1/bq[12] ), .ZN(n54393) );
  XOR2HSV0 U57280 ( .A1(n54394), .A2(n54393), .Z(n54395) );
  XOR2HSV0 U57281 ( .A1(n54396), .A2(n54395), .Z(n54405) );
  NAND2HSV0 U57282 ( .A1(n54978), .A2(n48380), .ZN(n54398) );
  NAND2HSV0 U57283 ( .A1(n55452), .A2(n55100), .ZN(n54397) );
  XOR2HSV0 U57284 ( .A1(n54398), .A2(n54397), .Z(n54403) );
  NOR2HSV0 U57285 ( .A1(n41944), .A2(n54399), .ZN(n54401) );
  NAND2HSV0 U57286 ( .A1(n55496), .A2(\pe1/bq[21] ), .ZN(n54400) );
  XOR2HSV0 U57287 ( .A1(n54401), .A2(n54400), .Z(n54402) );
  XOR2HSV0 U57288 ( .A1(n54403), .A2(n54402), .Z(n54404) );
  XOR2HSV0 U57289 ( .A1(n54405), .A2(n54404), .Z(n54406) );
  XNOR2HSV1 U57290 ( .A1(n54407), .A2(n54406), .ZN(n54408) );
  XNOR2HSV1 U57291 ( .A1(n54409), .A2(n54408), .ZN(n54410) );
  XNOR2HSV1 U57292 ( .A1(n54411), .A2(n54410), .ZN(n54413) );
  NAND2HSV0 U57293 ( .A1(n54513), .A2(n55319), .ZN(n54412) );
  XOR2HSV0 U57294 ( .A1(n54413), .A2(n54412), .Z(n54414) );
  XNOR2HSV1 U57295 ( .A1(n54415), .A2(n54414), .ZN(n54416) );
  XNOR2HSV1 U57296 ( .A1(n54417), .A2(n54416), .ZN(n54419) );
  NOR2HSV0 U57297 ( .A1(n54691), .A2(n55019), .ZN(n54418) );
  XOR3HSV2 U57298 ( .A1(n54420), .A2(n54419), .A3(n54418), .Z(n54421) );
  XNOR2HSV1 U57299 ( .A1(n54422), .A2(n54421), .ZN(n54423) );
  XNOR2HSV1 U57300 ( .A1(n54424), .A2(n54423), .ZN(n54425) );
  XNOR2HSV1 U57301 ( .A1(n54426), .A2(n54425), .ZN(n54427) );
  XOR2HSV0 U57302 ( .A1(n54428), .A2(n54427), .Z(n54429) );
  XNOR2HSV1 U57303 ( .A1(n54430), .A2(n54429), .ZN(n54433) );
  CLKNAND2HSV0 U57304 ( .A1(n54872), .A2(n55086), .ZN(n54432) );
  XOR2HSV0 U57305 ( .A1(n54433), .A2(n54432), .Z(n54434) );
  XNOR2HSV1 U57306 ( .A1(n54435), .A2(n54434), .ZN(n54436) );
  XNOR2HSV1 U57307 ( .A1(n54437), .A2(n54436), .ZN(n54439) );
  NAND2HSV0 U57308 ( .A1(n54541), .A2(\pe1/got [16]), .ZN(n54438) );
  XNOR2HSV1 U57309 ( .A1(n54439), .A2(n54438), .ZN(n54440) );
  XNOR2HSV1 U57310 ( .A1(n54441), .A2(n54440), .ZN(n54444) );
  INAND2HSV2 U57311 ( .A1(n55562), .B1(n54716), .ZN(n54443) );
  CLKNAND2HSV1 U57312 ( .A1(n55213), .A2(n54728), .ZN(n54442) );
  XOR3HSV2 U57313 ( .A1(n54444), .A2(n54443), .A3(n54442), .Z(n54445) );
  XOR2HSV0 U57314 ( .A1(n54446), .A2(n54445), .Z(n54447) );
  XOR2HSV0 U57315 ( .A1(n54448), .A2(n54447), .Z(n54451) );
  BUFHSV2 U57316 ( .I(n54553), .Z(n55513) );
  XOR3HSV2 U57317 ( .A1(n54451), .A2(n54450), .A3(n54449), .Z(\pe1/poht [9])
         );
  CLKNAND2HSV0 U57318 ( .A1(n55574), .A2(n54452), .ZN(n54552) );
  CLKNAND2HSV1 U57319 ( .A1(n55543), .A2(n54724), .ZN(n54550) );
  CLKNAND2HSV1 U57320 ( .A1(n59736), .A2(n54716), .ZN(n54545) );
  CLKNAND2HSV0 U57321 ( .A1(\pe1/got [16]), .A2(n55341), .ZN(n54540) );
  NAND2HSV0 U57322 ( .A1(n55229), .A2(n55222), .ZN(n54538) );
  NAND2HSV0 U57323 ( .A1(n42085), .A2(n42155), .ZN(n54534) );
  NOR2HSV1 U57324 ( .A1(n42356), .A2(n54453), .ZN(n54532) );
  NAND2HSV0 U57325 ( .A1(n29741), .A2(n55214), .ZN(n54530) );
  CLKNAND2HSV0 U57326 ( .A1(n42358), .A2(n55088), .ZN(n54528) );
  NOR2HSV2 U57327 ( .A1(n54454), .A2(n55163), .ZN(n54526) );
  NOR2HSV1 U57328 ( .A1(n54815), .A2(n55019), .ZN(n54524) );
  NAND2HSV0 U57329 ( .A1(n54557), .A2(\pe1/got [6]), .ZN(n54520) );
  INAND2HSV2 U57330 ( .A1(n55542), .B1(n54362), .ZN(n54518) );
  NAND2HSV0 U57331 ( .A1(n54456), .A2(n54455), .ZN(n54510) );
  NAND2HSV0 U57332 ( .A1(n54912), .A2(n42373), .ZN(n54458) );
  NAND2HSV0 U57333 ( .A1(\pe1/aot [16]), .A2(\pe1/bq[9] ), .ZN(n54457) );
  XOR2HSV0 U57334 ( .A1(n54458), .A2(n54457), .Z(n54462) );
  NAND2HSV0 U57335 ( .A1(\pe1/aot [21]), .A2(n55544), .ZN(n54460) );
  NAND2HSV0 U57336 ( .A1(n53954), .A2(n55605), .ZN(n54459) );
  XOR2HSV0 U57337 ( .A1(n54460), .A2(n54459), .Z(n54461) );
  XOR2HSV0 U57338 ( .A1(n54462), .A2(n54461), .Z(n54471) );
  NAND2HSV0 U57339 ( .A1(n54578), .A2(\pe1/bq[18] ), .ZN(n54464) );
  NAND2HSV0 U57340 ( .A1(n55397), .A2(n48380), .ZN(n54463) );
  XOR2HSV0 U57341 ( .A1(n54464), .A2(n54463), .Z(n54469) );
  NAND2HSV0 U57342 ( .A1(n54669), .A2(n54289), .ZN(n54467) );
  NAND2HSV0 U57343 ( .A1(n55496), .A2(n54465), .ZN(n54466) );
  XOR2HSV0 U57344 ( .A1(n54467), .A2(n54466), .Z(n54468) );
  XOR2HSV0 U57345 ( .A1(n54469), .A2(n54468), .Z(n54470) );
  XOR2HSV0 U57346 ( .A1(n54471), .A2(n54470), .Z(n54491) );
  NAND2HSV0 U57347 ( .A1(n55452), .A2(n54995), .ZN(n54474) );
  NAND2HSV0 U57348 ( .A1(n59495), .A2(n55100), .ZN(n54473) );
  XOR2HSV0 U57349 ( .A1(n54474), .A2(n54473), .Z(n54478) );
  NOR2HSV0 U57350 ( .A1(n41885), .A2(n54399), .ZN(n54476) );
  NAND2HSV0 U57351 ( .A1(n59737), .A2(n55231), .ZN(n54475) );
  XOR2HSV0 U57352 ( .A1(n54476), .A2(n54475), .Z(n54477) );
  XNOR2HSV1 U57353 ( .A1(n54478), .A2(n54477), .ZN(n54489) );
  NAND2HSV0 U57354 ( .A1(n55578), .A2(\pe1/bq[23] ), .ZN(n54481) );
  NAND2HSV0 U57355 ( .A1(n54743), .A2(n54479), .ZN(n54480) );
  XNOR2HSV1 U57356 ( .A1(n54481), .A2(n54480), .ZN(n54487) );
  NOR2HSV0 U57357 ( .A1(n54483), .A2(n54482), .ZN(n54485) );
  AOI22HSV0 U57358 ( .A1(n44533), .A2(n54179), .B1(n54999), .B2(n55393), .ZN(
        n54484) );
  NOR2HSV2 U57359 ( .A1(n54485), .A2(n54484), .ZN(n54486) );
  XNOR2HSV1 U57360 ( .A1(n54487), .A2(n54486), .ZN(n54488) );
  XNOR2HSV1 U57361 ( .A1(n54489), .A2(n54488), .ZN(n54490) );
  XNOR2HSV1 U57362 ( .A1(n54491), .A2(n54490), .ZN(n54508) );
  XOR2HSV0 U57363 ( .A1(n54493), .A2(n54492), .Z(n54496) );
  NAND2HSV0 U57364 ( .A1(n55553), .A2(n42238), .ZN(n54637) );
  NAND2HSV0 U57365 ( .A1(n55433), .A2(\pe1/bq[21] ), .ZN(n54494) );
  XOR2HSV0 U57366 ( .A1(n54637), .A2(n54494), .Z(n54495) );
  XOR2HSV0 U57367 ( .A1(n54496), .A2(n54495), .Z(n54506) );
  NAND2HSV0 U57368 ( .A1(n54497), .A2(n55501), .ZN(n54499) );
  NAND2HSV0 U57369 ( .A1(n42132), .A2(n54847), .ZN(n54498) );
  XOR2HSV0 U57370 ( .A1(n54499), .A2(n54498), .Z(n54504) );
  NOR2HSV0 U57371 ( .A1(n41974), .A2(n55185), .ZN(n54502) );
  NAND2HSV0 U57372 ( .A1(n54500), .A2(n55505), .ZN(n54501) );
  XOR2HSV0 U57373 ( .A1(n54502), .A2(n54501), .Z(n54503) );
  XOR2HSV0 U57374 ( .A1(n54504), .A2(n54503), .Z(n54505) );
  XOR2HSV0 U57375 ( .A1(n54506), .A2(n54505), .Z(n54507) );
  XNOR2HSV1 U57376 ( .A1(n54508), .A2(n54507), .ZN(n54509) );
  XNOR2HSV1 U57377 ( .A1(n54510), .A2(n54509), .ZN(n54512) );
  NAND2HSV0 U57378 ( .A1(n29763), .A2(\pe1/got [2]), .ZN(n54511) );
  XOR2HSV0 U57379 ( .A1(n54512), .A2(n54511), .Z(n54516) );
  NOR2HSV0 U57380 ( .A1(n41301), .A2(n55364), .ZN(n54515) );
  NAND2HSV0 U57381 ( .A1(n54513), .A2(n55410), .ZN(n54514) );
  XOR3HSV1 U57382 ( .A1(n54516), .A2(n54515), .A3(n54514), .Z(n54517) );
  XNOR2HSV1 U57383 ( .A1(n54518), .A2(n54517), .ZN(n54519) );
  XNOR2HSV1 U57384 ( .A1(n54520), .A2(n54519), .ZN(n54523) );
  NAND2HSV0 U57385 ( .A1(n54521), .A2(n55339), .ZN(n54522) );
  XOR3HSV2 U57386 ( .A1(n54524), .A2(n54523), .A3(n54522), .Z(n54525) );
  XNOR2HSV1 U57387 ( .A1(n54526), .A2(n54525), .ZN(n54527) );
  XNOR2HSV1 U57388 ( .A1(n54528), .A2(n54527), .ZN(n54529) );
  XNOR2HSV1 U57389 ( .A1(n54530), .A2(n54529), .ZN(n54531) );
  XNOR2HSV1 U57390 ( .A1(n54532), .A2(n54531), .ZN(n54533) );
  XNOR2HSV1 U57391 ( .A1(n54534), .A2(n54533), .ZN(n54536) );
  CLKNAND2HSV0 U57392 ( .A1(n54872), .A2(n54969), .ZN(n54535) );
  XOR2HSV0 U57393 ( .A1(n54536), .A2(n54535), .Z(n54537) );
  XNOR2HSV1 U57394 ( .A1(n54538), .A2(n54537), .ZN(n54539) );
  XNOR2HSV1 U57395 ( .A1(n54540), .A2(n54539), .ZN(n54543) );
  NAND2HSV0 U57396 ( .A1(n54541), .A2(n54965), .ZN(n54542) );
  XNOR2HSV1 U57397 ( .A1(n54543), .A2(n54542), .ZN(n54544) );
  XNOR2HSV1 U57398 ( .A1(n54545), .A2(n54544), .ZN(n54548) );
  INAND2HSV2 U57399 ( .A1(n55330), .B1(n54728), .ZN(n54547) );
  CLKNAND2HSV1 U57400 ( .A1(n55427), .A2(n44530), .ZN(n54546) );
  XOR3HSV2 U57401 ( .A1(n54548), .A2(n54547), .A3(n54546), .Z(n54549) );
  XOR2HSV0 U57402 ( .A1(n54550), .A2(n54549), .Z(n54551) );
  XOR2HSV0 U57403 ( .A1(n54552), .A2(n54551), .Z(n54556) );
  BUFHSV2 U57404 ( .I(n54553), .Z(n55537) );
  XOR3HSV2 U57405 ( .A1(n54556), .A2(n54555), .A3(n54554), .Z(\pe1/poht [8])
         );
  CLKNAND2HSV0 U57406 ( .A1(n55574), .A2(n54716), .ZN(n54630) );
  CLKNAND2HSV1 U57407 ( .A1(n59736), .A2(n54969), .ZN(n54623) );
  CLKNAND2HSV0 U57408 ( .A1(n55337), .A2(n55341), .ZN(n54619) );
  NAND2HSV0 U57409 ( .A1(n59422), .A2(n55214), .ZN(n54617) );
  BUFHSV2 U57410 ( .I(n59391), .Z(n54813) );
  CLKNAND2HSV1 U57411 ( .A1(n54813), .A2(n55331), .ZN(n54613) );
  NOR2HSV1 U57412 ( .A1(n55090), .A2(n55227), .ZN(n54611) );
  NAND2HSV0 U57413 ( .A1(n54730), .A2(n54894), .ZN(n54609) );
  NAND2HSV0 U57414 ( .A1(n42358), .A2(n55448), .ZN(n54607) );
  CLKNHSV1 U57415 ( .I(n53657), .ZN(n55092) );
  NOR2HSV1 U57416 ( .A1(n55092), .A2(n55542), .ZN(n54605) );
  NOR2HSV0 U57417 ( .A1(n54731), .A2(n55364), .ZN(n54603) );
  CLKNAND2HSV1 U57418 ( .A1(n54557), .A2(n54104), .ZN(n54599) );
  INAND2HSV0 U57419 ( .A1(n55376), .B1(n59534), .ZN(n54597) );
  NAND2HSV0 U57420 ( .A1(n55496), .A2(\pe1/bq[18] ), .ZN(n54638) );
  XOR2HSV0 U57421 ( .A1(n54558), .A2(n54638), .Z(n54562) );
  CLKNAND2HSV0 U57422 ( .A1(\pe1/aot [8]), .A2(n54179), .ZN(n54560) );
  NAND2HSV0 U57423 ( .A1(n59495), .A2(\pe1/bq[12] ), .ZN(n54559) );
  XOR2HSV0 U57424 ( .A1(n54560), .A2(n54559), .Z(n54561) );
  XOR2HSV0 U57425 ( .A1(n54562), .A2(n54561), .Z(n54595) );
  NAND2HSV0 U57426 ( .A1(\pe1/aot [16]), .A2(n54289), .ZN(n54564) );
  NAND2HSV0 U57427 ( .A1(n44541), .A2(n53798), .ZN(n54563) );
  XOR2HSV0 U57428 ( .A1(n54564), .A2(n54563), .Z(n54569) );
  CLKNAND2HSV0 U57429 ( .A1(n55093), .A2(n55166), .ZN(n54567) );
  NAND2HSV0 U57430 ( .A1(n54743), .A2(n54565), .ZN(n54566) );
  XOR2HSV0 U57431 ( .A1(n54567), .A2(n54566), .Z(n54568) );
  XOR2HSV0 U57432 ( .A1(n54569), .A2(n54568), .Z(n54577) );
  NAND2HSV0 U57433 ( .A1(\pe1/aot [14]), .A2(n55045), .ZN(n54571) );
  NAND2HSV0 U57434 ( .A1(n59730), .A2(n42092), .ZN(n54570) );
  XOR2HSV0 U57435 ( .A1(n54571), .A2(n54570), .Z(n54575) );
  NAND2HSV0 U57436 ( .A1(n59737), .A2(n55110), .ZN(n54573) );
  NAND2HSV0 U57437 ( .A1(n54669), .A2(n54988), .ZN(n54572) );
  XOR2HSV0 U57438 ( .A1(n54573), .A2(n54572), .Z(n54574) );
  XNOR2HSV1 U57439 ( .A1(n54575), .A2(n54574), .ZN(n54576) );
  XNOR2HSV1 U57440 ( .A1(n54577), .A2(n54576), .ZN(n54594) );
  NAND2HSV0 U57441 ( .A1(\pe1/aot [4]), .A2(n42098), .ZN(n54580) );
  NAND2HSV0 U57442 ( .A1(n54578), .A2(\pe1/bq[14] ), .ZN(n54579) );
  XOR2HSV0 U57443 ( .A1(n54580), .A2(n54579), .Z(n54584) );
  NAND2HSV0 U57444 ( .A1(n59993), .A2(n54836), .ZN(n54582) );
  CLKNAND2HSV0 U57445 ( .A1(\pe1/aot [6]), .A2(n48380), .ZN(n54581) );
  XOR2HSV0 U57446 ( .A1(n54582), .A2(n54581), .Z(n54583) );
  XOR2HSV0 U57447 ( .A1(n54584), .A2(n54583), .Z(n54592) );
  NAND2HSV0 U57448 ( .A1(n55113), .A2(\pe1/bq[9] ), .ZN(n54586) );
  CLKNAND2HSV0 U57449 ( .A1(n54662), .A2(n54847), .ZN(n54585) );
  XOR2HSV0 U57450 ( .A1(n54586), .A2(n54585), .Z(n54590) );
  NAND2HSV0 U57451 ( .A1(n54900), .A2(n55544), .ZN(n54588) );
  NAND2HSV0 U57452 ( .A1(n59733), .A2(n54668), .ZN(n54587) );
  XOR2HSV0 U57453 ( .A1(n54588), .A2(n54587), .Z(n54589) );
  XOR2HSV0 U57454 ( .A1(n54590), .A2(n54589), .Z(n54591) );
  XOR2HSV0 U57455 ( .A1(n54592), .A2(n54591), .Z(n54593) );
  XOR3HSV2 U57456 ( .A1(n54595), .A2(n54594), .A3(n54593), .Z(n54596) );
  XNOR2HSV1 U57457 ( .A1(n54597), .A2(n54596), .ZN(n54598) );
  XNOR2HSV1 U57458 ( .A1(n54599), .A2(n54598), .ZN(n54602) );
  NAND2HSV0 U57459 ( .A1(n54600), .A2(n55410), .ZN(n54601) );
  XOR3HSV2 U57460 ( .A1(n54603), .A2(n54602), .A3(n54601), .Z(n54604) );
  XNOR2HSV1 U57461 ( .A1(n54605), .A2(n54604), .ZN(n54606) );
  XNOR2HSV1 U57462 ( .A1(n54607), .A2(n54606), .ZN(n54608) );
  XNOR2HSV1 U57463 ( .A1(n54609), .A2(n54608), .ZN(n54610) );
  XNOR2HSV1 U57464 ( .A1(n54611), .A2(n54610), .ZN(n54612) );
  XNOR2HSV1 U57465 ( .A1(n54613), .A2(n54612), .ZN(n54615) );
  CLKNAND2HSV0 U57466 ( .A1(n54872), .A2(n55088), .ZN(n54614) );
  XOR2HSV0 U57467 ( .A1(n54615), .A2(n54614), .Z(n54616) );
  XNOR2HSV1 U57468 ( .A1(n54617), .A2(n54616), .ZN(n54618) );
  XNOR2HSV1 U57469 ( .A1(n54619), .A2(n54618), .ZN(n54621) );
  NAND2HSV0 U57470 ( .A1(n59751), .A2(n42155), .ZN(n54620) );
  XNOR2HSV1 U57471 ( .A1(n54621), .A2(n54620), .ZN(n54622) );
  XNOR2HSV1 U57472 ( .A1(n54623), .A2(n54622), .ZN(n54626) );
  INAND2HSV2 U57473 ( .A1(n55529), .B1(n55222), .ZN(n54625) );
  CLKNAND2HSV1 U57474 ( .A1(n55427), .A2(n42162), .ZN(n54624) );
  XNOR3HSV1 U57475 ( .A1(n54626), .A2(n54625), .A3(n54624), .ZN(n54628) );
  NAND2HSV0 U57476 ( .A1(n55226), .A2(n59996), .ZN(n54627) );
  XNOR2HSV1 U57477 ( .A1(n54628), .A2(n54627), .ZN(n54629) );
  XOR2HSV0 U57478 ( .A1(n54630), .A2(n54629), .Z(n54634) );
  NAND2HSV2 U57479 ( .A1(n25840), .A2(n54728), .ZN(n54633) );
  INHSV2 U57480 ( .I(n54154), .ZN(n54632) );
  INHSV4 U57481 ( .I(n54632), .ZN(n55423) );
  NAND2HSV0 U57482 ( .A1(n55488), .A2(\pe1/got [20]), .ZN(n54723) );
  CLKNAND2HSV1 U57483 ( .A1(n55576), .A2(n54728), .ZN(n54721) );
  CLKNAND2HSV1 U57484 ( .A1(n59736), .A2(n41374), .ZN(n54715) );
  NAND2HSV0 U57485 ( .A1(n54969), .A2(n59521), .ZN(n54710) );
  NAND2HSV0 U57486 ( .A1(n59422), .A2(n54812), .ZN(n54708) );
  CLKNAND2HSV1 U57487 ( .A1(n54813), .A2(n55214), .ZN(n54704) );
  NOR2HSV0 U57488 ( .A1(n53912), .A2(n54636), .ZN(n54702) );
  CLKNAND2HSV0 U57489 ( .A1(n55230), .A2(n44605), .ZN(n54700) );
  CLKNAND2HSV0 U57490 ( .A1(n54814), .A2(n55339), .ZN(n54698) );
  NOR2HSV1 U57491 ( .A1(n55092), .A2(n55019), .ZN(n54696) );
  NOR2HSV0 U57492 ( .A1(n54731), .A2(n55542), .ZN(n54694) );
  NAND2HSV0 U57493 ( .A1(n59725), .A2(n55267), .ZN(n54690) );
  INAND2HSV2 U57494 ( .A1(n55364), .B1(n54162), .ZN(n54688) );
  NOR2HSV0 U57495 ( .A1(n55515), .A2(n48060), .ZN(n54639) );
  OAI22HSV1 U57496 ( .A1(n54640), .A2(n54639), .B1(n54638), .B2(n54637), .ZN(
        n54645) );
  XOR2HSV0 U57497 ( .A1(n54642), .A2(n54641), .Z(n54643) );
  XOR3HSV2 U57498 ( .A1(n54645), .A2(n54644), .A3(n54643), .Z(n54682) );
  NAND2HSV0 U57499 ( .A1(n54578), .A2(n55100), .ZN(n54647) );
  NAND2HSV0 U57500 ( .A1(n54743), .A2(\pe1/bq[22] ), .ZN(n54646) );
  XOR2HSV0 U57501 ( .A1(n54647), .A2(n54646), .Z(n54651) );
  NAND2HSV0 U57502 ( .A1(\pe1/aot [4]), .A2(n42092), .ZN(n54649) );
  NAND2HSV0 U57503 ( .A1(n55234), .A2(n42098), .ZN(n54648) );
  XOR2HSV0 U57504 ( .A1(n54649), .A2(n54648), .Z(n54650) );
  XOR2HSV0 U57505 ( .A1(n54651), .A2(n54650), .Z(n54659) );
  NAND2HSV0 U57506 ( .A1(n54824), .A2(n55544), .ZN(n54653) );
  NAND2HSV0 U57507 ( .A1(n55093), .A2(n54179), .ZN(n54652) );
  XOR2HSV0 U57508 ( .A1(n54653), .A2(n54652), .Z(n54657) );
  NAND2HSV0 U57509 ( .A1(n42132), .A2(n53798), .ZN(n54655) );
  NAND2HSV0 U57510 ( .A1(\pe1/aot [14]), .A2(\pe1/bq[9] ), .ZN(n54654) );
  XOR2HSV0 U57511 ( .A1(n54655), .A2(n54654), .Z(n54656) );
  XNOR2HSV1 U57512 ( .A1(n54657), .A2(n54656), .ZN(n54658) );
  XNOR2HSV1 U57513 ( .A1(n54659), .A2(n54658), .ZN(n54681) );
  NAND2HSV0 U57514 ( .A1(n59733), .A2(n54289), .ZN(n54661) );
  NAND2HSV0 U57515 ( .A1(n54900), .A2(n54911), .ZN(n54660) );
  XOR2HSV0 U57516 ( .A1(n54661), .A2(n54660), .Z(n54667) );
  NAND2HSV0 U57517 ( .A1(n54662), .A2(n42373), .ZN(n54665) );
  NAND2HSV0 U57518 ( .A1(n54663), .A2(n55110), .ZN(n54664) );
  XOR2HSV0 U57519 ( .A1(n54665), .A2(n54664), .Z(n54666) );
  XOR2HSV0 U57520 ( .A1(n54667), .A2(n54666), .Z(n54679) );
  NAND2HSV0 U57521 ( .A1(n54669), .A2(n54668), .ZN(n54671) );
  NAND2HSV0 U57522 ( .A1(n55578), .A2(\pe1/bq[21] ), .ZN(n54670) );
  XOR2HSV0 U57523 ( .A1(n54671), .A2(n54670), .Z(n54677) );
  NOR2HSV0 U57524 ( .A1(n54672), .A2(n48030), .ZN(n54675) );
  NAND2HSV0 U57525 ( .A1(\pe1/aot [16]), .A2(n55045), .ZN(n54674) );
  XOR2HSV0 U57526 ( .A1(n54675), .A2(n54674), .Z(n54676) );
  XOR2HSV0 U57527 ( .A1(n54677), .A2(n54676), .Z(n54678) );
  XOR2HSV0 U57528 ( .A1(n54679), .A2(n54678), .Z(n54680) );
  XOR3HSV2 U57529 ( .A1(n54682), .A2(n54681), .A3(n54680), .Z(n54686) );
  CLKNHSV0 U57530 ( .I(n59755), .ZN(n55594) );
  NOR2HSV0 U57531 ( .A1(n41566), .A2(n55594), .ZN(n54685) );
  NAND2HSV0 U57532 ( .A1(n54683), .A2(\pe1/got [2]), .ZN(n54684) );
  XOR3HSV1 U57533 ( .A1(n54686), .A2(n54685), .A3(n54684), .Z(n54687) );
  XNOR2HSV1 U57534 ( .A1(n54688), .A2(n54687), .ZN(n54689) );
  XNOR2HSV1 U57535 ( .A1(n54690), .A2(n54689), .ZN(n54693) );
  NAND2HSV0 U57536 ( .A1(n54521), .A2(n55448), .ZN(n54692) );
  XOR3HSV2 U57537 ( .A1(n54694), .A2(n54693), .A3(n54692), .Z(n54695) );
  XNOR2HSV1 U57538 ( .A1(n54696), .A2(n54695), .ZN(n54697) );
  XNOR2HSV1 U57539 ( .A1(n54698), .A2(n54697), .ZN(n54699) );
  XNOR2HSV1 U57540 ( .A1(n54700), .A2(n54699), .ZN(n54701) );
  XNOR2HSV1 U57541 ( .A1(n54702), .A2(n54701), .ZN(n54703) );
  XNOR2HSV1 U57542 ( .A1(n54704), .A2(n54703), .ZN(n54706) );
  NAND2HSV0 U57543 ( .A1(n54872), .A2(n55337), .ZN(n54705) );
  XOR2HSV0 U57544 ( .A1(n54706), .A2(n54705), .Z(n54707) );
  XNOR2HSV1 U57545 ( .A1(n54708), .A2(n54707), .ZN(n54709) );
  XNOR2HSV1 U57546 ( .A1(n54710), .A2(n54709), .ZN(n54713) );
  CLKNAND2HSV1 U57547 ( .A1(n55411), .A2(n55222), .ZN(n54712) );
  XNOR2HSV1 U57548 ( .A1(n54713), .A2(n54712), .ZN(n54714) );
  XNOR2HSV1 U57549 ( .A1(n54715), .A2(n54714), .ZN(n54719) );
  INAND2HSV2 U57550 ( .A1(n55512), .B1(n59996), .ZN(n54718) );
  CLKNAND2HSV1 U57551 ( .A1(n55476), .A2(n54716), .ZN(n54717) );
  XOR3HSV2 U57552 ( .A1(n54719), .A2(n54718), .A3(n54717), .Z(n54720) );
  XOR2HSV0 U57553 ( .A1(n54721), .A2(n54720), .Z(n54722) );
  XOR2HSV0 U57554 ( .A1(n54723), .A2(n54722), .Z(n54727) );
  NAND2HSV2 U57555 ( .A1(n55569), .A2(n54724), .ZN(n54726) );
  XOR3HSV2 U57556 ( .A1(n54727), .A2(n54726), .A3(n54725), .Z(\pe1/poht [10])
         );
  NAND2HSV0 U57557 ( .A1(n55541), .A2(n54728), .ZN(n54808) );
  CLKNAND2HSV0 U57558 ( .A1(n59489), .A2(n54716), .ZN(n54806) );
  BUFHSV2 U57559 ( .I(n54729), .Z(n55089) );
  CLKNAND2HSV1 U57560 ( .A1(n55089), .A2(n55222), .ZN(n54801) );
  CLKNAND2HSV0 U57561 ( .A1(n55450), .A2(n54812), .ZN(n54797) );
  NAND2HSV0 U57562 ( .A1(n59422), .A2(n55337), .ZN(n54795) );
  NAND2HSV0 U57563 ( .A1(n54813), .A2(n55088), .ZN(n54791) );
  NOR2HSV1 U57564 ( .A1(n42356), .A2(n55163), .ZN(n54789) );
  NAND2HSV0 U57565 ( .A1(n54730), .A2(n55339), .ZN(n54787) );
  CLKNAND2HSV0 U57566 ( .A1(n42358), .A2(n54894), .ZN(n54785) );
  NOR2HSV1 U57567 ( .A1(n55092), .A2(n55369), .ZN(n54783) );
  NOR2HSV0 U57568 ( .A1(n54731), .A2(n55444), .ZN(n54781) );
  NAND2HSV0 U57569 ( .A1(n59725), .A2(n55319), .ZN(n54778) );
  NAND2HSV0 U57570 ( .A1(n59534), .A2(\pe1/got [2]), .ZN(n54776) );
  NAND2HSV0 U57571 ( .A1(n54732), .A2(\pe1/got [1]), .ZN(n54774) );
  NAND2HSV0 U57572 ( .A1(n55234), .A2(n54836), .ZN(n54733) );
  XNOR2HSV1 U57573 ( .A1(n54734), .A2(n54733), .ZN(n54739) );
  NOR2HSV0 U57574 ( .A1(n54673), .A2(n54735), .ZN(n54737) );
  NAND2HSV0 U57575 ( .A1(\pe1/aot [4]), .A2(\pe1/bq[18] ), .ZN(n54736) );
  XOR2HSV0 U57576 ( .A1(n54737), .A2(n54736), .Z(n54738) );
  XOR3HSV2 U57577 ( .A1(n54740), .A2(n54739), .A3(n54738), .Z(n54772) );
  NAND2HSV0 U57578 ( .A1(n54900), .A2(n54289), .ZN(n54742) );
  NAND2HSV0 U57579 ( .A1(\pe1/aot [14]), .A2(n55501), .ZN(n54741) );
  XOR2HSV0 U57580 ( .A1(n54742), .A2(n54741), .Z(n54747) );
  NAND2HSV0 U57581 ( .A1(n54743), .A2(\pe1/bq[21] ), .ZN(n54745) );
  NAND2HSV0 U57582 ( .A1(n59991), .A2(n42373), .ZN(n54744) );
  XOR2HSV0 U57583 ( .A1(n54745), .A2(n54744), .Z(n54746) );
  XOR2HSV0 U57584 ( .A1(n54747), .A2(n54746), .Z(n54755) );
  NAND2HSV0 U57585 ( .A1(n42132), .A2(n55045), .ZN(n54749) );
  NAND2HSV0 U57586 ( .A1(n55113), .A2(n54847), .ZN(n54748) );
  XOR2HSV0 U57587 ( .A1(n54749), .A2(n54748), .Z(n54753) );
  NAND2HSV0 U57588 ( .A1(n59737), .A2(n55577), .ZN(n54751) );
  NAND2HSV0 U57589 ( .A1(n55547), .A2(\pe1/bq[15] ), .ZN(n54750) );
  XOR2HSV0 U57590 ( .A1(n54751), .A2(n54750), .Z(n54752) );
  XNOR2HSV1 U57591 ( .A1(n54753), .A2(n54752), .ZN(n54754) );
  XNOR2HSV1 U57592 ( .A1(n54755), .A2(n54754), .ZN(n54771) );
  NAND2HSV0 U57593 ( .A1(n55553), .A2(n42098), .ZN(n54757) );
  NAND2HSV0 U57594 ( .A1(n55103), .A2(\pe1/bq[9] ), .ZN(n54756) );
  XOR2HSV0 U57595 ( .A1(n54757), .A2(n54756), .Z(n54761) );
  NAND2HSV0 U57596 ( .A1(\pe1/aot [3]), .A2(n42092), .ZN(n54759) );
  NAND2HSV0 U57597 ( .A1(n42093), .A2(n55110), .ZN(n54758) );
  XOR2HSV0 U57598 ( .A1(n54759), .A2(n54758), .Z(n54760) );
  XOR2HSV0 U57599 ( .A1(n54761), .A2(n54760), .Z(n54769) );
  NAND2HSV0 U57600 ( .A1(n54913), .A2(n55241), .ZN(n54763) );
  NAND2HSV0 U57601 ( .A1(n55380), .A2(n54179), .ZN(n54762) );
  XOR2HSV0 U57602 ( .A1(n54763), .A2(n54762), .Z(n54767) );
  NAND2HSV0 U57603 ( .A1(n59733), .A2(n55544), .ZN(n54765) );
  NAND2HSV0 U57604 ( .A1(n54904), .A2(n41641), .ZN(n54764) );
  XOR2HSV0 U57605 ( .A1(n54765), .A2(n54764), .Z(n54766) );
  XOR2HSV0 U57606 ( .A1(n54767), .A2(n54766), .Z(n54768) );
  XOR2HSV0 U57607 ( .A1(n54769), .A2(n54768), .Z(n54770) );
  XOR3HSV2 U57608 ( .A1(n54772), .A2(n54771), .A3(n54770), .Z(n54773) );
  XNOR2HSV1 U57609 ( .A1(n54774), .A2(n54773), .ZN(n54775) );
  XNOR2HSV1 U57610 ( .A1(n54776), .A2(n54775), .ZN(n54777) );
  XNOR2HSV1 U57611 ( .A1(n54778), .A2(n54777), .ZN(n54780) );
  NAND2HSV0 U57612 ( .A1(n54521), .A2(n55475), .ZN(n54779) );
  XOR3HSV2 U57613 ( .A1(n54781), .A2(n54780), .A3(n54779), .Z(n54782) );
  XNOR2HSV1 U57614 ( .A1(n54783), .A2(n54782), .ZN(n54784) );
  XNOR2HSV1 U57615 ( .A1(n54785), .A2(n54784), .ZN(n54786) );
  XNOR2HSV1 U57616 ( .A1(n54787), .A2(n54786), .ZN(n54788) );
  XNOR2HSV1 U57617 ( .A1(n54789), .A2(n54788), .ZN(n54790) );
  XNOR2HSV1 U57618 ( .A1(n54791), .A2(n54790), .ZN(n54793) );
  CLKNAND2HSV0 U57619 ( .A1(n54872), .A2(n55214), .ZN(n54792) );
  XOR2HSV0 U57620 ( .A1(n54793), .A2(n54792), .Z(n54794) );
  XNOR2HSV1 U57621 ( .A1(n54795), .A2(n54794), .ZN(n54796) );
  XNOR2HSV1 U57622 ( .A1(n54797), .A2(n54796), .ZN(n54799) );
  CLKNAND2HSV1 U57623 ( .A1(n59751), .A2(n54969), .ZN(n54798) );
  XNOR2HSV1 U57624 ( .A1(n54799), .A2(n54798), .ZN(n54800) );
  XNOR2HSV1 U57625 ( .A1(n54801), .A2(n54800), .ZN(n54804) );
  INAND2HSV2 U57626 ( .A1(n55330), .B1(n41374), .ZN(n54803) );
  XOR3HSV2 U57627 ( .A1(n54804), .A2(n54803), .A3(n54802), .Z(n54805) );
  XOR2HSV0 U57628 ( .A1(n54806), .A2(n54805), .Z(n54807) );
  XOR2HSV0 U57629 ( .A1(n54808), .A2(n54807), .Z(n54811) );
  NAND2HSV2 U57630 ( .A1(n55484), .A2(\pe1/got [20]), .ZN(n54810) );
  XOR3HSV2 U57631 ( .A1(n54811), .A2(n54810), .A3(n54809), .Z(\pe1/poht [11])
         );
  CLKNAND2HSV0 U57632 ( .A1(n55593), .A2(n54965), .ZN(n54890) );
  CLKNAND2HSV1 U57633 ( .A1(n55576), .A2(\pe1/got [16]), .ZN(n54888) );
  CLKNAND2HSV1 U57634 ( .A1(n55089), .A2(n54812), .ZN(n54883) );
  NAND2HSV0 U57635 ( .A1(n54970), .A2(n59521), .ZN(n54878) );
  NAND2HSV0 U57636 ( .A1(n55375), .A2(n55088), .ZN(n54876) );
  CLKNAND2HSV1 U57637 ( .A1(n54813), .A2(n55339), .ZN(n54871) );
  CLKNHSV0 U57638 ( .I(n59360), .ZN(n55090) );
  NOR2HSV0 U57639 ( .A1(n55090), .A2(n55019), .ZN(n54869) );
  NAND2HSV0 U57640 ( .A1(n29741), .A2(n55448), .ZN(n54867) );
  NAND2HSV0 U57641 ( .A1(n54814), .A2(n55475), .ZN(n54865) );
  NOR2HSV1 U57642 ( .A1(n55092), .A2(n55444), .ZN(n54863) );
  NOR2HSV1 U57643 ( .A1(n54815), .A2(n55575), .ZN(n54861) );
  NAND2HSV0 U57644 ( .A1(n59725), .A2(\pe1/got [1]), .ZN(n54858) );
  NAND2HSV0 U57645 ( .A1(\pe1/aot [7]), .A2(\pe1/bq[13] ), .ZN(n54817) );
  NAND2HSV0 U57646 ( .A1(n55234), .A2(\pe1/bq[14] ), .ZN(n54816) );
  XOR2HSV0 U57647 ( .A1(n54817), .A2(n54816), .Z(n54822) );
  NAND2HSV0 U57648 ( .A1(n54818), .A2(n55166), .ZN(n54820) );
  CLKNHSV1 U57649 ( .I(n55524), .ZN(n55455) );
  NAND2HSV0 U57650 ( .A1(n55455), .A2(\pe1/bq[19] ), .ZN(n54819) );
  XOR2HSV0 U57651 ( .A1(n54820), .A2(n54819), .Z(n54821) );
  XOR2HSV0 U57652 ( .A1(n54822), .A2(n54821), .Z(n54856) );
  NOR2HSV0 U57653 ( .A1(n54823), .A2(n55607), .ZN(n54826) );
  AOI22HSV0 U57654 ( .A1(n54824), .A2(n55392), .B1(\pe1/bq[18] ), .B2(n55595), 
        .ZN(n54825) );
  NOR2HSV1 U57655 ( .A1(n54826), .A2(n54825), .ZN(n54835) );
  NAND2HSV0 U57656 ( .A1(\pe1/aot [16]), .A2(n55544), .ZN(n54828) );
  NAND2HSV0 U57657 ( .A1(n59993), .A2(\pe1/bq[15] ), .ZN(n54827) );
  XOR2HSV0 U57658 ( .A1(n54828), .A2(n54827), .Z(n54834) );
  NAND2HSV0 U57659 ( .A1(\pe1/aot [12]), .A2(\pe1/bq[8] ), .ZN(n54833) );
  NOR2HSV0 U57660 ( .A1(n54829), .A2(n54399), .ZN(n54831) );
  NAND2HSV0 U57661 ( .A1(n54913), .A2(\pe1/bq[9] ), .ZN(n54830) );
  XOR2HSV0 U57662 ( .A1(n54831), .A2(n54830), .Z(n54832) );
  XOR4HSV1 U57663 ( .A1(n54835), .A2(n54834), .A3(n54833), .A4(n54832), .Z(
        n54855) );
  NAND2HSV0 U57664 ( .A1(\pe1/aot [4]), .A2(n54836), .ZN(n54838) );
  NAND2HSV0 U57665 ( .A1(\pe1/aot [3]), .A2(n42098), .ZN(n54837) );
  XOR2HSV0 U57666 ( .A1(n54838), .A2(n54837), .Z(n54842) );
  NAND2HSV0 U57667 ( .A1(n54904), .A2(n42373), .ZN(n54840) );
  NAND2HSV0 U57668 ( .A1(n42132), .A2(n54289), .ZN(n54839) );
  XOR2HSV0 U57669 ( .A1(n54840), .A2(n54839), .Z(n54841) );
  XOR2HSV0 U57670 ( .A1(n54842), .A2(n54841), .Z(n54853) );
  NAND2HSV0 U57671 ( .A1(n54912), .A2(n55045), .ZN(n54845) );
  NAND2HSV0 U57672 ( .A1(\pe1/aot [14]), .A2(n54911), .ZN(n54844) );
  XOR2HSV0 U57673 ( .A1(n54845), .A2(n54844), .Z(n54851) );
  CLKNHSV0 U57674 ( .I(n54846), .ZN(n55397) );
  NAND2HSV0 U57675 ( .A1(n55397), .A2(n54847), .ZN(n54849) );
  NAND2HSV0 U57676 ( .A1(n59733), .A2(n55605), .ZN(n54848) );
  XOR2HSV0 U57677 ( .A1(n54849), .A2(n54848), .Z(n54850) );
  XOR2HSV0 U57678 ( .A1(n54851), .A2(n54850), .Z(n54852) );
  XOR2HSV0 U57679 ( .A1(n54853), .A2(n54852), .Z(n54854) );
  XOR3HSV2 U57680 ( .A1(n54856), .A2(n54855), .A3(n54854), .Z(n54857) );
  XNOR2HSV1 U57681 ( .A1(n54858), .A2(n54857), .ZN(n54860) );
  NAND2HSV0 U57682 ( .A1(n54521), .A2(n55319), .ZN(n54859) );
  XOR3HSV2 U57683 ( .A1(n54861), .A2(n54860), .A3(n54859), .Z(n54862) );
  XNOR2HSV1 U57684 ( .A1(n54863), .A2(n54862), .ZN(n54864) );
  XNOR2HSV1 U57685 ( .A1(n54865), .A2(n54864), .ZN(n54866) );
  XNOR2HSV1 U57686 ( .A1(n54867), .A2(n54866), .ZN(n54868) );
  XNOR2HSV1 U57687 ( .A1(n54869), .A2(n54868), .ZN(n54870) );
  XNOR2HSV1 U57688 ( .A1(n54871), .A2(n54870), .ZN(n54874) );
  CLKNAND2HSV0 U57689 ( .A1(n54872), .A2(n44605), .ZN(n54873) );
  XOR2HSV0 U57690 ( .A1(n54874), .A2(n54873), .Z(n54875) );
  XNOR2HSV1 U57691 ( .A1(n54876), .A2(n54875), .ZN(n54877) );
  XNOR2HSV1 U57692 ( .A1(n54878), .A2(n54877), .ZN(n54881) );
  CLKNAND2HSV1 U57693 ( .A1(n59751), .A2(n55087), .ZN(n54880) );
  XNOR2HSV1 U57694 ( .A1(n54881), .A2(n54880), .ZN(n54882) );
  XNOR2HSV1 U57695 ( .A1(n54883), .A2(n54882), .ZN(n54887) );
  INAND2HSV2 U57696 ( .A1(n55562), .B1(n54969), .ZN(n54886) );
  CLKNAND2HSV1 U57697 ( .A1(n59931), .A2(n54241), .ZN(n54885) );
  XOR2HSV0 U57698 ( .A1(n54890), .A2(n54889), .Z(n54893) );
  NAND2HSV2 U57699 ( .A1(n59428), .A2(n42359), .ZN(n54892) );
  NAND2HSV2 U57700 ( .A1(n25848), .A2(n59995), .ZN(n54891) );
  XOR3HSV2 U57701 ( .A1(n54893), .A2(n54892), .A3(n54891), .Z(\pe1/poht [13])
         );
  CLKNAND2HSV0 U57702 ( .A1(n55488), .A2(\pe1/got [16]), .ZN(n54964) );
  CLKNAND2HSV1 U57703 ( .A1(n55489), .A2(n54241), .ZN(n54962) );
  CLKNAND2HSV1 U57704 ( .A1(n55089), .A2(n55087), .ZN(n54956) );
  CLKNAND2HSV0 U57705 ( .A1(n55341), .A2(n55088), .ZN(n54952) );
  NAND2HSV0 U57706 ( .A1(n55375), .A2(n55331), .ZN(n54950) );
  CLKNAND2HSV1 U57707 ( .A1(n54813), .A2(n54894), .ZN(n54945) );
  NOR2HSV1 U57708 ( .A1(n55090), .A2(n55369), .ZN(n54943) );
  NAND2HSV0 U57709 ( .A1(n55091), .A2(n55475), .ZN(n54941) );
  NAND2HSV0 U57710 ( .A1(n59592), .A2(n55267), .ZN(n54939) );
  NOR2HSV1 U57711 ( .A1(n55092), .A2(n55364), .ZN(n54937) );
  NAND2HSV0 U57712 ( .A1(n59518), .A2(\pe1/got [1]), .ZN(n54933) );
  NAND2HSV0 U57713 ( .A1(n59495), .A2(n55250), .ZN(n54896) );
  NAND2HSV0 U57714 ( .A1(\pe1/aot [4]), .A2(\pe1/bq[15] ), .ZN(n54895) );
  XOR2HSV0 U57715 ( .A1(n54896), .A2(n54895), .Z(n54899) );
  NAND2HSV0 U57716 ( .A1(n55113), .A2(n55045), .ZN(n55179) );
  CLKNAND2HSV0 U57717 ( .A1(\pe1/aot [7]), .A2(\pe1/bq[12] ), .ZN(n54897) );
  XOR2HSV0 U57718 ( .A1(n55179), .A2(n54897), .Z(n54898) );
  XOR2HSV0 U57719 ( .A1(n54899), .A2(n54898), .Z(n54931) );
  NAND2HSV0 U57720 ( .A1(n54900), .A2(n55605), .ZN(n54903) );
  NAND2HSV0 U57721 ( .A1(n55234), .A2(n54179), .ZN(n54902) );
  XOR2HSV0 U57722 ( .A1(n54903), .A2(n54902), .Z(n54908) );
  NAND2HSV0 U57723 ( .A1(n54904), .A2(n55166), .ZN(n54906) );
  NAND2HSV0 U57724 ( .A1(n59730), .A2(\pe1/bq[17] ), .ZN(n54905) );
  XOR2HSV0 U57725 ( .A1(n54906), .A2(n54905), .Z(n54907) );
  XOR2HSV0 U57726 ( .A1(n54908), .A2(n54907), .Z(n54910) );
  NOR2HSV0 U57727 ( .A1(n55515), .A2(n45814), .ZN(n54975) );
  CLKNAND2HSV0 U57728 ( .A1(n59993), .A2(\pe1/bq[14] ), .ZN(n54998) );
  XOR2HSV0 U57729 ( .A1(n54975), .A2(n54998), .Z(n54909) );
  XNOR2HSV1 U57730 ( .A1(n54910), .A2(n54909), .ZN(n54930) );
  NAND2HSV0 U57731 ( .A1(n54912), .A2(n54911), .ZN(n54915) );
  CLKNAND2HSV0 U57732 ( .A1(n54913), .A2(\pe1/bq[8] ), .ZN(n54914) );
  XOR2HSV0 U57733 ( .A1(n54915), .A2(n54914), .Z(n54920) );
  NAND2HSV0 U57734 ( .A1(n54916), .A2(n54988), .ZN(n54918) );
  NAND2HSV0 U57735 ( .A1(n55455), .A2(\pe1/bq[18] ), .ZN(n54917) );
  XOR2HSV0 U57736 ( .A1(n54918), .A2(n54917), .Z(n54919) );
  XOR2HSV0 U57737 ( .A1(n54920), .A2(n54919), .Z(n54928) );
  NAND2HSV0 U57738 ( .A1(n55186), .A2(n55544), .ZN(n54922) );
  NAND2HSV0 U57739 ( .A1(n55093), .A2(\pe1/bq[9] ), .ZN(n54921) );
  XOR2HSV0 U57740 ( .A1(n54922), .A2(n54921), .Z(n54926) );
  NAND2HSV0 U57741 ( .A1(\pe1/aot [14]), .A2(n54289), .ZN(n54924) );
  NAND2HSV0 U57742 ( .A1(\pe1/aot [16]), .A2(n55577), .ZN(n54923) );
  XOR2HSV0 U57743 ( .A1(n54924), .A2(n54923), .Z(n54925) );
  XOR2HSV0 U57744 ( .A1(n54926), .A2(n54925), .Z(n54927) );
  XOR2HSV0 U57745 ( .A1(n54928), .A2(n54927), .Z(n54929) );
  XOR3HSV2 U57746 ( .A1(n54931), .A2(n54930), .A3(n54929), .Z(n54932) );
  XNOR2HSV1 U57747 ( .A1(n54933), .A2(n54932), .ZN(n54935) );
  CLKNAND2HSV0 U57748 ( .A1(n41850), .A2(n54104), .ZN(n54934) );
  XOR2HSV0 U57749 ( .A1(n54935), .A2(n54934), .Z(n54936) );
  XNOR2HSV1 U57750 ( .A1(n54937), .A2(n54936), .ZN(n54938) );
  XNOR2HSV1 U57751 ( .A1(n54939), .A2(n54938), .ZN(n54940) );
  XNOR2HSV1 U57752 ( .A1(n54941), .A2(n54940), .ZN(n54942) );
  XNOR2HSV1 U57753 ( .A1(n54943), .A2(n54942), .ZN(n54944) );
  XNOR2HSV1 U57754 ( .A1(n54945), .A2(n54944), .ZN(n54948) );
  CLKNAND2HSV0 U57755 ( .A1(n54946), .A2(n55339), .ZN(n54947) );
  XOR2HSV0 U57756 ( .A1(n54948), .A2(n54947), .Z(n54949) );
  XNOR2HSV1 U57757 ( .A1(n54950), .A2(n54949), .ZN(n54951) );
  XNOR2HSV1 U57758 ( .A1(n54952), .A2(n54951), .ZN(n54954) );
  CLKNAND2HSV0 U57759 ( .A1(n55069), .A2(n54970), .ZN(n54953) );
  XNOR2HSV1 U57760 ( .A1(n54954), .A2(n54953), .ZN(n54955) );
  XNOR2HSV1 U57761 ( .A1(n54956), .A2(n54955), .ZN(n54960) );
  INAND2HSV2 U57762 ( .A1(n55330), .B1(n55086), .ZN(n54959) );
  NAND2HSV2 U57763 ( .A1(n55427), .A2(n54969), .ZN(n54958) );
  XOR3HSV2 U57764 ( .A1(n54960), .A2(n54959), .A3(n54958), .Z(n54961) );
  XOR2HSV0 U57765 ( .A1(n54962), .A2(n54961), .Z(n54963) );
  XOR2HSV0 U57766 ( .A1(n54964), .A2(n54963), .Z(n54968) );
  XOR3HSV2 U57767 ( .A1(n54968), .A2(n54967), .A3(n54966), .Z(\pe1/poht [14])
         );
  CLKNAND2HSV0 U57768 ( .A1(n55488), .A2(n54241), .ZN(n55036) );
  CLKNAND2HSV0 U57769 ( .A1(n59489), .A2(n54969), .ZN(n55034) );
  CLKNAND2HSV1 U57770 ( .A1(n55089), .A2(n54970), .ZN(n55029) );
  CLKNAND2HSV0 U57771 ( .A1(n55450), .A2(n55145), .ZN(n55025) );
  NAND2HSV0 U57772 ( .A1(n59422), .A2(n55339), .ZN(n55023) );
  CLKNAND2HSV1 U57773 ( .A1(n54813), .A2(n55448), .ZN(n55017) );
  NOR2HSV1 U57774 ( .A1(n55090), .A2(n55542), .ZN(n55015) );
  NAND2HSV0 U57775 ( .A1(n55091), .A2(n55267), .ZN(n55013) );
  NAND2HSV0 U57776 ( .A1(n59592), .A2(n55319), .ZN(n55011) );
  NOR2HSV1 U57777 ( .A1(n55092), .A2(n55575), .ZN(n55009) );
  CLKNAND2HSV0 U57778 ( .A1(n41850), .A2(\pe1/got [1]), .ZN(n55007) );
  CLKNAND2HSV0 U57779 ( .A1(\pe1/aot [16]), .A2(n55110), .ZN(n54972) );
  NAND2HSV0 U57780 ( .A1(n55103), .A2(n54289), .ZN(n54971) );
  XOR2HSV0 U57781 ( .A1(n54972), .A2(n54971), .Z(n54987) );
  NOR2HSV0 U57782 ( .A1(n55504), .A2(n54973), .ZN(n55119) );
  AOI22HSV0 U57783 ( .A1(n59389), .A2(n48380), .B1(n55100), .B2(n55595), .ZN(
        n54974) );
  AOI21HSV1 U57784 ( .A1(n54975), .A2(n55119), .B(n54974), .ZN(n54977) );
  XOR2HSV0 U57785 ( .A1(n54977), .A2(n54976), .Z(n54986) );
  NAND2HSV0 U57786 ( .A1(n54978), .A2(\pe1/bq[9] ), .ZN(n54980) );
  NAND2HSV0 U57787 ( .A1(n59991), .A2(\pe1/bq[8] ), .ZN(n54979) );
  XOR2HSV0 U57788 ( .A1(n54980), .A2(n54979), .Z(n54984) );
  NAND2HSV0 U57789 ( .A1(\pe1/aot [14]), .A2(n55544), .ZN(n54982) );
  NAND2HSV0 U57790 ( .A1(n54913), .A2(n55394), .ZN(n54981) );
  XOR2HSV0 U57791 ( .A1(n54982), .A2(n54981), .Z(n54983) );
  XNOR2HSV1 U57792 ( .A1(n54984), .A2(n54983), .ZN(n54985) );
  XOR3HSV2 U57793 ( .A1(n54987), .A2(n54986), .A3(n54985), .Z(n55005) );
  NAND2HSV0 U57794 ( .A1(n55186), .A2(n55518), .ZN(n54990) );
  NAND2HSV0 U57795 ( .A1(n54900), .A2(n54988), .ZN(n54989) );
  XOR2HSV0 U57796 ( .A1(n54990), .A2(n54989), .Z(n54994) );
  NOR2HSV0 U57797 ( .A1(n54901), .A2(n53691), .ZN(n54992) );
  NAND2HSV0 U57798 ( .A1(n54904), .A2(n55250), .ZN(n54991) );
  XOR2HSV0 U57799 ( .A1(n54992), .A2(n54991), .Z(n54993) );
  XNOR2HSV1 U57800 ( .A1(n54994), .A2(n54993), .ZN(n55003) );
  CLKNAND2HSV0 U57801 ( .A1(n55455), .A2(n54995), .ZN(n54997) );
  NAND2HSV0 U57802 ( .A1(\pe1/aot [7]), .A2(n55166), .ZN(n54996) );
  XOR2HSV0 U57803 ( .A1(n54997), .A2(n54996), .Z(n55001) );
  CLKNAND2HSV0 U57804 ( .A1(n59619), .A2(n41645), .ZN(n55118) );
  XNOR2HSV1 U57805 ( .A1(n55001), .A2(n55000), .ZN(n55002) );
  XNOR2HSV1 U57806 ( .A1(n55003), .A2(n55002), .ZN(n55004) );
  XNOR2HSV1 U57807 ( .A1(n55005), .A2(n55004), .ZN(n55006) );
  XNOR2HSV1 U57808 ( .A1(n55007), .A2(n55006), .ZN(n55008) );
  XNOR2HSV1 U57809 ( .A1(n55009), .A2(n55008), .ZN(n55010) );
  XNOR2HSV1 U57810 ( .A1(n55011), .A2(n55010), .ZN(n55012) );
  XNOR2HSV1 U57811 ( .A1(n55013), .A2(n55012), .ZN(n55014) );
  XNOR2HSV1 U57812 ( .A1(n55015), .A2(n55014), .ZN(n55016) );
  XNOR2HSV1 U57813 ( .A1(n55017), .A2(n55016), .ZN(n55021) );
  INHSV2 U57814 ( .I(n55019), .ZN(n55570) );
  NAND2HSV0 U57815 ( .A1(n53768), .A2(n55570), .ZN(n55020) );
  XOR2HSV0 U57816 ( .A1(n55021), .A2(n55020), .Z(n55022) );
  XNOR2HSV1 U57817 ( .A1(n55023), .A2(n55022), .ZN(n55024) );
  XNOR2HSV1 U57818 ( .A1(n55025), .A2(n55024), .ZN(n55027) );
  CLKNAND2HSV0 U57819 ( .A1(n55069), .A2(n55088), .ZN(n55026) );
  XNOR2HSV1 U57820 ( .A1(n55027), .A2(n55026), .ZN(n55028) );
  XNOR2HSV1 U57821 ( .A1(n55029), .A2(n55028), .ZN(n55032) );
  INAND2HSV2 U57822 ( .A1(n55562), .B1(n55087), .ZN(n55031) );
  CLKNAND2HSV0 U57823 ( .A1(n55476), .A2(n55086), .ZN(n55030) );
  XOR3HSV2 U57824 ( .A1(n55032), .A2(n55031), .A3(n55030), .Z(n55033) );
  XOR2HSV0 U57825 ( .A1(n55034), .A2(n55033), .Z(n55035) );
  XOR2HSV0 U57826 ( .A1(n55036), .A2(n55035), .Z(n55039) );
  NAND2HSV2 U57827 ( .A1(n25840), .A2(n41374), .ZN(n55038) );
  XOR3HSV2 U57828 ( .A1(n55039), .A2(n55038), .A3(n55037), .Z(\pe1/poht [15])
         );
  CLKNAND2HSV0 U57829 ( .A1(n55541), .A2(n55088), .ZN(n55081) );
  CLKNAND2HSV1 U57830 ( .A1(n55543), .A2(n55145), .ZN(n55079) );
  NAND2HSV0 U57831 ( .A1(n55267), .A2(n55450), .ZN(n55068) );
  NAND2HSV0 U57832 ( .A1(n59422), .A2(n55319), .ZN(n55066) );
  CLKNAND2HSV1 U57833 ( .A1(n55397), .A2(n55518), .ZN(n55041) );
  NAND2HSV0 U57834 ( .A1(n59730), .A2(n55241), .ZN(n55040) );
  XOR2HSV0 U57835 ( .A1(n55041), .A2(n55040), .Z(n55044) );
  CLKNAND2HSV1 U57836 ( .A1(n54913), .A2(n55110), .ZN(n55042) );
  XOR2HSV0 U57837 ( .A1(n55180), .A2(n55042), .Z(n55043) );
  XOR2HSV0 U57838 ( .A1(n55044), .A2(n55043), .Z(n55062) );
  CLKNAND2HSV0 U57839 ( .A1(n59993), .A2(n53708), .ZN(n55047) );
  CLKNAND2HSV1 U57840 ( .A1(n55234), .A2(n55045), .ZN(n55046) );
  XOR2HSV0 U57841 ( .A1(n55047), .A2(n55046), .Z(n55051) );
  CLKNAND2HSV0 U57842 ( .A1(n54904), .A2(\pe1/bq[5] ), .ZN(n55049) );
  NAND2HSV0 U57843 ( .A1(n55113), .A2(n55392), .ZN(n55048) );
  XOR2HSV0 U57844 ( .A1(n55049), .A2(n55048), .Z(n55050) );
  XOR2HSV0 U57845 ( .A1(n55051), .A2(n55050), .Z(n55059) );
  NAND2HSV0 U57846 ( .A1(\pe1/aot [3]), .A2(n54847), .ZN(n55053) );
  CLKNAND2HSV1 U57847 ( .A1(\pe1/aot [4]), .A2(\pe1/bq[9] ), .ZN(n55052) );
  XOR2HSV0 U57848 ( .A1(n55053), .A2(n55052), .Z(n55057) );
  NOR2HSV0 U57849 ( .A1(n55524), .A2(n53691), .ZN(n55055) );
  CLKNAND2HSV1 U57850 ( .A1(n54578), .A2(n55231), .ZN(n55054) );
  XOR2HSV0 U57851 ( .A1(n55055), .A2(n55054), .Z(n55056) );
  XOR2HSV0 U57852 ( .A1(n55057), .A2(n55056), .Z(n55058) );
  XOR2HSV0 U57853 ( .A1(n55059), .A2(n55058), .Z(n55061) );
  CLKNAND2HSV1 U57854 ( .A1(n54038), .A2(\pe1/got [1]), .ZN(n55060) );
  XOR3HSV2 U57855 ( .A1(n55062), .A2(n55061), .A3(n55060), .Z(n55064) );
  NAND2HSV0 U57856 ( .A1(n53768), .A2(n55340), .ZN(n55063) );
  XNOR2HSV1 U57857 ( .A1(n55064), .A2(n55063), .ZN(n55065) );
  XNOR2HSV1 U57858 ( .A1(n55066), .A2(n55065), .ZN(n55067) );
  XNOR2HSV1 U57859 ( .A1(n55068), .A2(n55067), .ZN(n55071) );
  CLKNAND2HSV0 U57860 ( .A1(n55069), .A2(n55475), .ZN(n55070) );
  XNOR2HSV1 U57861 ( .A1(n55071), .A2(n55070), .ZN(n55073) );
  CLKNAND2HSV0 U57862 ( .A1(n55089), .A2(n55448), .ZN(n55072) );
  XOR2HSV0 U57863 ( .A1(n55073), .A2(n55072), .Z(n55075) );
  INAND2HSV2 U57864 ( .A1(n55529), .B1(n55570), .ZN(n55074) );
  XOR2HSV0 U57865 ( .A1(n55075), .A2(n55074), .Z(n55077) );
  CLKNAND2HSV1 U57866 ( .A1(n55427), .A2(n55339), .ZN(n55076) );
  XNOR2HSV1 U57867 ( .A1(n55077), .A2(n55076), .ZN(n55078) );
  XOR2HSV0 U57868 ( .A1(n55079), .A2(n55078), .Z(n55080) );
  XOR2HSV0 U57869 ( .A1(n55081), .A2(n55080), .Z(n55085) );
  NAND2HSV2 U57870 ( .A1(n25839), .A2(n55214), .ZN(n55084) );
  XOR3HSV2 U57871 ( .A1(n55085), .A2(n55084), .A3(n55083), .Z(\pe1/poht [20])
         );
  CLKNAND2HSV0 U57872 ( .A1(n55541), .A2(n54969), .ZN(n55157) );
  CLKNAND2HSV0 U57873 ( .A1(n59489), .A2(n55086), .ZN(n55155) );
  CLKNAND2HSV2 U57874 ( .A1(n55490), .A2(n55087), .ZN(n55151) );
  CLKNAND2HSV1 U57875 ( .A1(n55089), .A2(n55088), .ZN(n55149) );
  NAND2HSV0 U57876 ( .A1(n59521), .A2(n55339), .ZN(n55143) );
  NAND2HSV0 U57877 ( .A1(n55229), .A2(n55570), .ZN(n55141) );
  CLKNAND2HSV1 U57878 ( .A1(n54038), .A2(n55475), .ZN(n55137) );
  NOR2HSV1 U57879 ( .A1(n55090), .A2(n55444), .ZN(n55135) );
  NAND2HSV0 U57880 ( .A1(n55091), .A2(n55319), .ZN(n55133) );
  NAND2HSV0 U57881 ( .A1(n59592), .A2(n55340), .ZN(n55131) );
  NOR2HSV0 U57882 ( .A1(n55092), .A2(n55376), .ZN(n55129) );
  CLKNAND2HSV0 U57883 ( .A1(n55093), .A2(n55394), .ZN(n55095) );
  NAND2HSV0 U57884 ( .A1(\pe1/aot [7]), .A2(n54847), .ZN(n55094) );
  XOR2HSV0 U57885 ( .A1(n55095), .A2(n55094), .Z(n55099) );
  NAND2HSV0 U57886 ( .A1(n59593), .A2(n55231), .ZN(n55097) );
  CLKNAND2HSV0 U57887 ( .A1(\pe1/aot [14]), .A2(n55518), .ZN(n55096) );
  XOR2HSV0 U57888 ( .A1(n55097), .A2(n55096), .Z(n55098) );
  XOR2HSV0 U57889 ( .A1(n55099), .A2(n55098), .Z(n55109) );
  CLKNHSV0 U57890 ( .I(n55524), .ZN(n55290) );
  NAND2HSV0 U57891 ( .A1(n55290), .A2(n55100), .ZN(n55102) );
  CLKNAND2HSV0 U57892 ( .A1(n54303), .A2(n42373), .ZN(n55101) );
  XOR2HSV0 U57893 ( .A1(n55102), .A2(n55101), .Z(n55107) );
  NAND2HSV0 U57894 ( .A1(n55234), .A2(n55241), .ZN(n55105) );
  CLKNAND2HSV0 U57895 ( .A1(n55103), .A2(\pe1/bq[4] ), .ZN(n55104) );
  XOR2HSV0 U57896 ( .A1(n55105), .A2(n55104), .Z(n55106) );
  XOR2HSV0 U57897 ( .A1(n55107), .A2(n55106), .Z(n55108) );
  XOR2HSV0 U57898 ( .A1(n55109), .A2(n55108), .Z(n55127) );
  NAND2HSV0 U57899 ( .A1(\pe1/aot [16]), .A2(n55392), .ZN(n55112) );
  NAND2HSV0 U57900 ( .A1(n55186), .A2(n55110), .ZN(n55111) );
  XOR2HSV0 U57901 ( .A1(n55112), .A2(n55111), .Z(n55117) );
  NAND2HSV0 U57902 ( .A1(n55113), .A2(n54289), .ZN(n55115) );
  NAND2HSV0 U57903 ( .A1(n54904), .A2(\pe1/bq[9] ), .ZN(n55114) );
  XOR2HSV0 U57904 ( .A1(n55115), .A2(n55114), .Z(n55116) );
  XOR2HSV0 U57905 ( .A1(n55117), .A2(n55116), .Z(n55125) );
  XOR2HSV0 U57906 ( .A1(n55119), .A2(n55118), .Z(n55123) );
  NAND2HSV0 U57907 ( .A1(n59495), .A2(n53708), .ZN(n55121) );
  NAND2HSV0 U57908 ( .A1(\pe1/aot [3]), .A2(\pe1/bq[14] ), .ZN(n55120) );
  XOR2HSV0 U57909 ( .A1(n55121), .A2(n55120), .Z(n55122) );
  XOR2HSV0 U57910 ( .A1(n55123), .A2(n55122), .Z(n55124) );
  XOR2HSV0 U57911 ( .A1(n55125), .A2(n55124), .Z(n55126) );
  XOR2HSV0 U57912 ( .A1(n55127), .A2(n55126), .Z(n55128) );
  XNOR2HSV1 U57913 ( .A1(n55129), .A2(n55128), .ZN(n55130) );
  XNOR2HSV1 U57914 ( .A1(n55131), .A2(n55130), .ZN(n55132) );
  XNOR2HSV1 U57915 ( .A1(n55133), .A2(n55132), .ZN(n55134) );
  XNOR2HSV1 U57916 ( .A1(n55135), .A2(n55134), .ZN(n55136) );
  XNOR2HSV1 U57917 ( .A1(n55137), .A2(n55136), .ZN(n55139) );
  NAND2HSV0 U57918 ( .A1(n54946), .A2(n55448), .ZN(n55138) );
  XOR2HSV0 U57919 ( .A1(n55139), .A2(n55138), .Z(n55140) );
  XNOR2HSV1 U57920 ( .A1(n55141), .A2(n55140), .ZN(n55142) );
  XNOR2HSV1 U57921 ( .A1(n55143), .A2(n55142), .ZN(n55147) );
  INHSV1 U57922 ( .I(n55144), .ZN(n55411) );
  CLKNAND2HSV0 U57923 ( .A1(n55411), .A2(n55145), .ZN(n55146) );
  XNOR2HSV1 U57924 ( .A1(n55147), .A2(n55146), .ZN(n55148) );
  XNOR2HSV1 U57925 ( .A1(n55149), .A2(n55148), .ZN(n55150) );
  XNOR2HSV1 U57926 ( .A1(n55151), .A2(n55150), .ZN(n55153) );
  INAND2HSV2 U57927 ( .A1(n55529), .B1(n55214), .ZN(n55152) );
  XNOR2HSV1 U57928 ( .A1(n55153), .A2(n55152), .ZN(n55154) );
  XOR2HSV0 U57929 ( .A1(n55155), .A2(n55154), .Z(n55156) );
  XOR2HSV0 U57930 ( .A1(n55157), .A2(n55156), .Z(n55161) );
  CLKNAND2HSV2 U57931 ( .A1(n55537), .A2(n48339), .ZN(n55160) );
  XOR3HSV2 U57932 ( .A1(n55161), .A2(n55160), .A3(n55159), .Z(\pe1/poht [16])
         );
  CLKNAND2HSV0 U57933 ( .A1(n55541), .A2(n55086), .ZN(n55221) );
  CLKNAND2HSV1 U57934 ( .A1(n55289), .A2(n55087), .ZN(n55219) );
  CLKNAND2HSV1 U57935 ( .A1(n55449), .A2(n55331), .ZN(n55212) );
  NAND2HSV0 U57936 ( .A1(n55450), .A2(n55570), .ZN(n55208) );
  NAND2HSV0 U57937 ( .A1(n55375), .A2(n53523), .ZN(n55206) );
  NAND2HSV0 U57938 ( .A1(n53521), .A2(n55267), .ZN(n55202) );
  NOR2HSV1 U57939 ( .A1(n53391), .A2(n55364), .ZN(n55200) );
  CLKNAND2HSV1 U57940 ( .A1(n29741), .A2(n55340), .ZN(n55198) );
  NAND2HSV0 U57941 ( .A1(n59592), .A2(\pe1/got [1]), .ZN(n55196) );
  NAND2HSV2 U57942 ( .A1(n54578), .A2(\pe1/bq[9] ), .ZN(n55165) );
  CLKNAND2HSV0 U57943 ( .A1(\pe1/aot [4]), .A2(n42373), .ZN(n55164) );
  XOR2HSV0 U57944 ( .A1(n55165), .A2(n55164), .Z(n55170) );
  NAND2HSV0 U57945 ( .A1(n55553), .A2(n55166), .ZN(n55168) );
  NAND2HSV0 U57946 ( .A1(n55234), .A2(n54847), .ZN(n55167) );
  XOR2HSV0 U57947 ( .A1(n55168), .A2(n55167), .Z(n55169) );
  XOR2HSV0 U57948 ( .A1(n55170), .A2(n55169), .Z(n55178) );
  NAND2HSV0 U57949 ( .A1(n54904), .A2(n55501), .ZN(n55172) );
  NAND2HSV0 U57950 ( .A1(\pe1/aot [14]), .A2(n55605), .ZN(n55171) );
  XOR2HSV0 U57951 ( .A1(n55172), .A2(n55171), .Z(n55176) );
  NAND2HSV0 U57952 ( .A1(n59730), .A2(\pe1/bq[14] ), .ZN(n55174) );
  CLKNAND2HSV0 U57953 ( .A1(n55290), .A2(\pe1/bq[15] ), .ZN(n55173) );
  XOR2HSV0 U57954 ( .A1(n55174), .A2(n55173), .Z(n55175) );
  XOR2HSV0 U57955 ( .A1(n55176), .A2(n55175), .Z(n55177) );
  XOR2HSV0 U57956 ( .A1(n55178), .A2(n55177), .Z(n55194) );
  NOR2HSV0 U57957 ( .A1(n55180), .A2(n55179), .ZN(n55182) );
  AOI22HSV0 U57958 ( .A1(n44533), .A2(n55544), .B1(n59495), .B2(n55394), .ZN(
        n55181) );
  NOR2HSV1 U57959 ( .A1(n55182), .A2(n55181), .ZN(n55192) );
  NAND2HSV0 U57960 ( .A1(\pe1/aot [11]), .A2(\pe1/bq[5] ), .ZN(n55184) );
  NAND2HSV0 U57961 ( .A1(n55397), .A2(n55231), .ZN(n55183) );
  XOR2HSV0 U57962 ( .A1(n55184), .A2(n55183), .Z(n55191) );
  NOR2HSV1 U57963 ( .A1(n55515), .A2(n48059), .ZN(n55190) );
  NOR2HSV0 U57964 ( .A1(n53672), .A2(n54399), .ZN(n55188) );
  NAND2HSV0 U57965 ( .A1(n55186), .A2(n55495), .ZN(n55187) );
  XOR2HSV0 U57966 ( .A1(n55188), .A2(n55187), .Z(n55189) );
  XOR4HSV1 U57967 ( .A1(n55192), .A2(n55191), .A3(n55190), .A4(n55189), .Z(
        n55193) );
  XNOR2HSV1 U57968 ( .A1(n55194), .A2(n55193), .ZN(n55195) );
  XNOR2HSV1 U57969 ( .A1(n55196), .A2(n55195), .ZN(n55197) );
  XNOR2HSV1 U57970 ( .A1(n55198), .A2(n55197), .ZN(n55199) );
  XNOR2HSV1 U57971 ( .A1(n55200), .A2(n55199), .ZN(n55201) );
  XNOR2HSV1 U57972 ( .A1(n55202), .A2(n55201), .ZN(n55204) );
  NAND2HSV0 U57973 ( .A1(n54946), .A2(n55475), .ZN(n55203) );
  XOR2HSV0 U57974 ( .A1(n55204), .A2(n55203), .Z(n55205) );
  XNOR2HSV1 U57975 ( .A1(n55206), .A2(n55205), .ZN(n55207) );
  XNOR2HSV1 U57976 ( .A1(n55208), .A2(n55207), .ZN(n55210) );
  CLKNAND2HSV0 U57977 ( .A1(n55411), .A2(n55339), .ZN(n55209) );
  XNOR2HSV1 U57978 ( .A1(n55210), .A2(n55209), .ZN(n55211) );
  XNOR2HSV1 U57979 ( .A1(n55212), .A2(n55211), .ZN(n55217) );
  INAND2HSV2 U57980 ( .A1(n55330), .B1(\pe1/got [10]), .ZN(n55216) );
  NAND2HSV2 U57981 ( .A1(n55332), .A2(n55214), .ZN(n55215) );
  XOR3HSV2 U57982 ( .A1(n55217), .A2(n55216), .A3(n55215), .Z(n55218) );
  XOR2HSV0 U57983 ( .A1(n55219), .A2(n55218), .Z(n55220) );
  XOR2HSV0 U57984 ( .A1(n55221), .A2(n55220), .Z(n55225) );
  XOR3HSV2 U57985 ( .A1(n55225), .A2(n55224), .A3(n55223), .Z(\pe1/poht [17])
         );
  NAND2HSV0 U57986 ( .A1(n55226), .A2(n55214), .ZN(n55283) );
  NAND2HSV2 U57987 ( .A1(n55332), .A2(\pe1/got [10]), .ZN(n55281) );
  INAND2HSV2 U57988 ( .A1(n55529), .B1(n55331), .ZN(n55279) );
  CLKNAND2HSV1 U57989 ( .A1(n55228), .A2(n55339), .ZN(n55277) );
  NAND2HSV0 U57990 ( .A1(n59521), .A2(n55448), .ZN(n55273) );
  NAND2HSV0 U57991 ( .A1(n55229), .A2(\pe1/got [5]), .ZN(n55271) );
  CLKNAND2HSV0 U57992 ( .A1(n53521), .A2(n55319), .ZN(n55266) );
  NOR2HSV1 U57993 ( .A1(n53391), .A2(n55575), .ZN(n55264) );
  CLKNAND2HSV0 U57994 ( .A1(n55230), .A2(\pe1/got [1]), .ZN(n55262) );
  NAND2HSV0 U57995 ( .A1(n54978), .A2(n55231), .ZN(n55233) );
  NAND2HSV0 U57996 ( .A1(n54904), .A2(n55505), .ZN(n55232) );
  XOR2HSV0 U57997 ( .A1(n55233), .A2(n55232), .Z(n55238) );
  NAND2HSV0 U57998 ( .A1(n55234), .A2(\pe1/bq[9] ), .ZN(n55236) );
  NAND2HSV0 U57999 ( .A1(n59593), .A2(\pe1/bq[4] ), .ZN(n55235) );
  XOR2HSV0 U58000 ( .A1(n55236), .A2(n55235), .Z(n55237) );
  XOR2HSV0 U58001 ( .A1(n55238), .A2(n55237), .Z(n55247) );
  XOR2HSV0 U58002 ( .A1(n55240), .A2(n55239), .Z(n55245) );
  NOR2HSV0 U58003 ( .A1(n55515), .A2(n53691), .ZN(n55243) );
  NAND2HSV0 U58004 ( .A1(\pe1/aot [4]), .A2(n55241), .ZN(n55242) );
  XOR2HSV0 U58005 ( .A1(n55243), .A2(n55242), .Z(n55244) );
  XOR2HSV0 U58006 ( .A1(n55245), .A2(n55244), .Z(n55246) );
  XOR2HSV0 U58007 ( .A1(n55247), .A2(n55246), .Z(n55260) );
  NAND2HSV0 U58008 ( .A1(n55595), .A2(\pe1/bq[13] ), .ZN(n55249) );
  CLKNAND2HSV0 U58009 ( .A1(n55290), .A2(n53571), .ZN(n55248) );
  XOR2HSV0 U58010 ( .A1(n55249), .A2(n55248), .Z(n55254) );
  NAND2HSV0 U58011 ( .A1(n55547), .A2(n55501), .ZN(n55252) );
  NAND2HSV0 U58012 ( .A1(\pe1/aot [5]), .A2(n55250), .ZN(n55251) );
  XOR2HSV0 U58013 ( .A1(n55252), .A2(n55251), .Z(n55253) );
  XNOR2HSV1 U58014 ( .A1(n55254), .A2(n55253), .ZN(n55258) );
  XOR2HSV0 U58015 ( .A1(n55256), .A2(n55255), .Z(n55257) );
  XNOR2HSV1 U58016 ( .A1(n55258), .A2(n55257), .ZN(n55259) );
  XNOR2HSV1 U58017 ( .A1(n55260), .A2(n55259), .ZN(n55261) );
  XNOR2HSV1 U58018 ( .A1(n55262), .A2(n55261), .ZN(n55263) );
  XNOR2HSV1 U58019 ( .A1(n55264), .A2(n55263), .ZN(n55265) );
  XNOR2HSV1 U58020 ( .A1(n55266), .A2(n55265), .ZN(n55269) );
  NAND2HSV0 U58021 ( .A1(n54872), .A2(n55267), .ZN(n55268) );
  XOR2HSV0 U58022 ( .A1(n55269), .A2(n55268), .Z(n55270) );
  XNOR2HSV1 U58023 ( .A1(n55271), .A2(n55270), .ZN(n55272) );
  XNOR2HSV1 U58024 ( .A1(n55273), .A2(n55272), .ZN(n55275) );
  NAND2HSV0 U58025 ( .A1(n55411), .A2(n55570), .ZN(n55274) );
  XNOR2HSV1 U58026 ( .A1(n55275), .A2(n55274), .ZN(n55276) );
  XNOR2HSV1 U58027 ( .A1(n55277), .A2(n55276), .ZN(n55278) );
  XOR2HSV0 U58028 ( .A1(n55279), .A2(n55278), .Z(n55280) );
  XNOR2HSV1 U58029 ( .A1(n55281), .A2(n55280), .ZN(n55282) );
  CLKAND2HSV1 U58030 ( .A1(n55593), .A2(n55337), .Z(n55284) );
  XNOR2HSV1 U58031 ( .A1(n55285), .A2(n55284), .ZN(n55288) );
  NAND2HSV2 U58032 ( .A1(n25839), .A2(n55086), .ZN(n55287) );
  NAND2HSV2 U58033 ( .A1(n55423), .A2(\pe1/got [14]), .ZN(n55286) );
  XOR3HSV2 U58034 ( .A1(n55288), .A2(n55287), .A3(n55286), .Z(\pe1/poht [18])
         );
  CLKNAND2HSV0 U58035 ( .A1(n55574), .A2(n55214), .ZN(n55336) );
  CLKNAND2HSV1 U58036 ( .A1(n55449), .A2(n55570), .ZN(n55329) );
  CLKNAND2HSV0 U58037 ( .A1(\pe1/got [5]), .A2(n55450), .ZN(n55325) );
  NAND2HSV0 U58038 ( .A1(n55375), .A2(n55410), .ZN(n55323) );
  NAND2HSV0 U58039 ( .A1(n42085), .A2(n55340), .ZN(n55318) );
  NOR2HSV1 U58040 ( .A1(n42208), .A2(n55376), .ZN(n55316) );
  CLKNAND2HSV1 U58041 ( .A1(n55290), .A2(n54179), .ZN(n55292) );
  NAND2HSV0 U58042 ( .A1(n59991), .A2(\pe1/bq[4] ), .ZN(n55291) );
  XOR2HSV0 U58043 ( .A1(n55292), .A2(n55291), .Z(n55296) );
  CLKNAND2HSV0 U58044 ( .A1(n44533), .A2(n55605), .ZN(n55294) );
  NAND2HSV0 U58045 ( .A1(n55492), .A2(\pe1/bq[8] ), .ZN(n55293) );
  XOR2HSV0 U58046 ( .A1(n55294), .A2(n55293), .Z(n55295) );
  XOR2HSV0 U58047 ( .A1(n55296), .A2(n55295), .Z(n55304) );
  NAND2HSV0 U58048 ( .A1(n55496), .A2(n54311), .ZN(n55298) );
  NAND2HSV0 U58049 ( .A1(\pe1/aot [5]), .A2(\pe1/bq[9] ), .ZN(n55297) );
  XOR2HSV0 U58050 ( .A1(n55298), .A2(n55297), .Z(n55302) );
  CLKNAND2HSV1 U58051 ( .A1(\pe1/aot [4]), .A2(n55352), .ZN(n55300) );
  NAND2HSV0 U58052 ( .A1(n55452), .A2(n55231), .ZN(n55299) );
  XOR2HSV0 U58053 ( .A1(n55300), .A2(n55299), .Z(n55301) );
  XOR2HSV0 U58054 ( .A1(n55302), .A2(n55301), .Z(n55303) );
  XOR2HSV0 U58055 ( .A1(n55304), .A2(n55303), .Z(n55314) );
  NAND2HSV0 U58056 ( .A1(n59593), .A2(n55491), .ZN(n55305) );
  XNOR2HSV1 U58057 ( .A1(n55306), .A2(n55305), .ZN(n55311) );
  NOR2HSV0 U58058 ( .A1(n55307), .A2(n54093), .ZN(n55309) );
  NAND2HSV0 U58059 ( .A1(\pe1/aot [2]), .A2(n42373), .ZN(n55308) );
  XOR2HSV0 U58060 ( .A1(n55309), .A2(n55308), .Z(n55310) );
  XOR3HSV2 U58061 ( .A1(n55312), .A2(n55311), .A3(n55310), .Z(n55313) );
  XNOR2HSV1 U58062 ( .A1(n55314), .A2(n55313), .ZN(n55315) );
  XNOR2HSV1 U58063 ( .A1(n55316), .A2(n55315), .ZN(n55317) );
  XNOR2HSV1 U58064 ( .A1(n55318), .A2(n55317), .ZN(n55321) );
  NAND2HSV0 U58065 ( .A1(n54872), .A2(n55319), .ZN(n55320) );
  XOR2HSV0 U58066 ( .A1(n55321), .A2(n55320), .Z(n55322) );
  XNOR2HSV1 U58067 ( .A1(n55323), .A2(n55322), .ZN(n55324) );
  XNOR2HSV1 U58068 ( .A1(n55325), .A2(n55324), .ZN(n55327) );
  CLKNAND2HSV0 U58069 ( .A1(n55411), .A2(n55448), .ZN(n55326) );
  XNOR2HSV1 U58070 ( .A1(n55327), .A2(n55326), .ZN(n55328) );
  XNOR2HSV1 U58071 ( .A1(n55329), .A2(n55328), .ZN(n55335) );
  INAND2HSV2 U58072 ( .A1(n55330), .B1(n55339), .ZN(n55334) );
  NAND2HSV2 U58073 ( .A1(n55332), .A2(n55331), .ZN(n55333) );
  NAND2HSV2 U58074 ( .A1(n55484), .A2(n55337), .ZN(n55338) );
  CLKNAND2HSV0 U58075 ( .A1(n55574), .A2(n55339), .ZN(n55372) );
  CLKNAND2HSV1 U58076 ( .A1(n55449), .A2(n55410), .ZN(n55368) );
  CLKNAND2HSV0 U58077 ( .A1(n55341), .A2(n55340), .ZN(n55363) );
  NAND2HSV0 U58078 ( .A1(n55375), .A2(n54455), .ZN(n55361) );
  XOR2HSV0 U58079 ( .A1(n55343), .A2(n55342), .Z(n55359) );
  NAND2HSV0 U58080 ( .A1(n59495), .A2(n55605), .ZN(n55345) );
  NAND2HSV0 U58081 ( .A1(n55452), .A2(n55491), .ZN(n55344) );
  XOR2HSV0 U58082 ( .A1(n55345), .A2(n55344), .Z(n55349) );
  NOR2HSV0 U58083 ( .A1(n55430), .A2(n55523), .ZN(n55347) );
  CLKNAND2HSV0 U58084 ( .A1(n55496), .A2(n55501), .ZN(n55346) );
  XOR2HSV0 U58085 ( .A1(n55347), .A2(n55346), .Z(n55348) );
  XNOR2HSV1 U58086 ( .A1(n55349), .A2(n55348), .ZN(n55358) );
  NAND2HSV0 U58087 ( .A1(n55492), .A2(\pe1/bq[5] ), .ZN(n55351) );
  NAND2HSV0 U58088 ( .A1(n55547), .A2(n55544), .ZN(n55350) );
  XOR2HSV0 U58089 ( .A1(n55351), .A2(n55350), .Z(n55356) );
  INHSV2 U58090 ( .I(n55524), .ZN(n55552) );
  NAND2HSV0 U58091 ( .A1(n55552), .A2(n55352), .ZN(n55353) );
  XOR2HSV0 U58092 ( .A1(n55354), .A2(n55353), .Z(n55355) );
  XOR2HSV0 U58093 ( .A1(n55356), .A2(n55355), .Z(n55357) );
  XOR3HSV2 U58094 ( .A1(n55359), .A2(n55358), .A3(n55357), .Z(n55360) );
  XNOR2HSV1 U58095 ( .A1(n55361), .A2(n55360), .ZN(n55362) );
  XNOR2HSV1 U58096 ( .A1(n55363), .A2(n55362), .ZN(n55366) );
  CLKNAND2HSV0 U58097 ( .A1(n55411), .A2(n55514), .ZN(n55365) );
  XNOR2HSV1 U58098 ( .A1(n55366), .A2(n55365), .ZN(n55367) );
  XNOR2HSV1 U58099 ( .A1(n55368), .A2(n55367), .ZN(n55371) );
  INAND2HSV2 U58100 ( .A1(n55562), .B1(n55475), .ZN(n55370) );
  NAND2HSV0 U58101 ( .A1(\pe1/got [10]), .A2(n53513), .ZN(n55373) );
  CLKNAND2HSV0 U58102 ( .A1(n55488), .A2(n55331), .ZN(n55422) );
  CLKNAND2HSV1 U58103 ( .A1(n55489), .A2(n55339), .ZN(n55420) );
  CLKNAND2HSV1 U58104 ( .A1(n55449), .A2(n55475), .ZN(n55415) );
  CLKNAND2HSV0 U58105 ( .A1(n55450), .A2(n55514), .ZN(n55409) );
  NAND2HSV0 U58106 ( .A1(n55375), .A2(n55340), .ZN(n55407) );
  NAND2HSV0 U58107 ( .A1(n59377), .A2(n59755), .ZN(n55405) );
  NAND2HSV0 U58108 ( .A1(n55452), .A2(\pe1/bq[4] ), .ZN(n55378) );
  NAND2HSV0 U58109 ( .A1(n55492), .A2(n55231), .ZN(n55377) );
  XOR2HSV0 U58110 ( .A1(n55378), .A2(n55377), .Z(n55384) );
  CLKNAND2HSV0 U58111 ( .A1(\pe1/aot [2]), .A2(n55379), .ZN(n55382) );
  NAND2HSV0 U58112 ( .A1(n55577), .A2(n55380), .ZN(n55381) );
  XOR2HSV0 U58113 ( .A1(n55382), .A2(n55381), .Z(n55383) );
  XOR2HSV0 U58114 ( .A1(n55384), .A2(n55383), .Z(n55391) );
  NOR2HSV0 U58115 ( .A1(n55515), .A2(n55385), .ZN(n55387) );
  CLKNAND2HSV0 U58116 ( .A1(n55547), .A2(\pe1/bq[5] ), .ZN(n55386) );
  XOR2HSV0 U58117 ( .A1(n55387), .A2(n55386), .Z(n55389) );
  CLKNAND2HSV0 U58118 ( .A1(\pe1/aot [4]), .A2(n55501), .ZN(n55388) );
  XNOR2HSV1 U58119 ( .A1(n55389), .A2(n55388), .ZN(n55390) );
  XNOR2HSV1 U58120 ( .A1(n55391), .A2(n55390), .ZN(n55403) );
  NAND2HSV0 U58121 ( .A1(n55393), .A2(n55392), .ZN(n55396) );
  CLKNAND2HSV0 U58122 ( .A1(n55553), .A2(n55394), .ZN(n55395) );
  XOR2HSV0 U58123 ( .A1(n55396), .A2(n55395), .Z(n55401) );
  NOR2HSV0 U58124 ( .A1(n55524), .A2(n48030), .ZN(n55399) );
  CLKNAND2HSV0 U58125 ( .A1(n55397), .A2(n55451), .ZN(n55398) );
  XOR2HSV0 U58126 ( .A1(n55399), .A2(n55398), .Z(n55400) );
  XOR2HSV0 U58127 ( .A1(n55401), .A2(n55400), .Z(n55402) );
  XNOR2HSV1 U58128 ( .A1(n55403), .A2(n55402), .ZN(n55404) );
  XNOR2HSV1 U58129 ( .A1(n55405), .A2(n55404), .ZN(n55406) );
  XNOR2HSV1 U58130 ( .A1(n55407), .A2(n55406), .ZN(n55408) );
  XNOR2HSV1 U58131 ( .A1(n55409), .A2(n55408), .ZN(n55413) );
  CLKNAND2HSV0 U58132 ( .A1(n55411), .A2(n55410), .ZN(n55412) );
  XNOR2HSV1 U58133 ( .A1(n55413), .A2(n55412), .ZN(n55414) );
  XNOR2HSV1 U58134 ( .A1(n55415), .A2(n55414), .ZN(n55418) );
  INAND2HSV2 U58135 ( .A1(n55562), .B1(n55448), .ZN(n55417) );
  CLKNAND2HSV0 U58136 ( .A1(n55476), .A2(n59750), .ZN(n55416) );
  XOR3HSV2 U58137 ( .A1(n55418), .A2(n55417), .A3(n55416), .Z(n55419) );
  XOR2HSV0 U58138 ( .A1(n55420), .A2(n55419), .Z(n55421) );
  XOR2HSV0 U58139 ( .A1(n55422), .A2(n55421), .Z(n55426) );
  NAND2HSV2 U58140 ( .A1(n59428), .A2(n55088), .ZN(n55425) );
  NAND2HSV2 U58141 ( .A1(n55423), .A2(n55214), .ZN(n55424) );
  XOR3HSV2 U58142 ( .A1(n55426), .A2(n55425), .A3(n55424), .Z(\pe1/poht [21])
         );
  CLKNAND2HSV0 U58143 ( .A1(n55574), .A2(n55514), .ZN(n55443) );
  CLKNAND2HSV1 U58144 ( .A1(n55489), .A2(n59756), .ZN(n55441) );
  NAND2HSV2 U58145 ( .A1(n55427), .A2(n54455), .ZN(n55439) );
  NAND2HSV2 U58146 ( .A1(n55578), .A2(n55544), .ZN(n55429) );
  CLKNAND2HSV0 U58147 ( .A1(n55496), .A2(n55577), .ZN(n55428) );
  XOR2HSV0 U58148 ( .A1(n55429), .A2(n55428), .Z(n55432) );
  NOR2HSV1 U58149 ( .A1(n55430), .A2(n55185), .ZN(n55431) );
  XNOR2HSV1 U58150 ( .A1(n55432), .A2(n55431), .ZN(n55437) );
  CLKNAND2HSV0 U58151 ( .A1(n55552), .A2(\pe1/bq[5] ), .ZN(n55435) );
  CLKNAND2HSV1 U58152 ( .A1(n55433), .A2(n55451), .ZN(n55434) );
  XOR2HSV0 U58153 ( .A1(n55435), .A2(n55434), .Z(n55436) );
  XNOR2HSV1 U58154 ( .A1(n55437), .A2(n55436), .ZN(n55438) );
  XNOR2HSV1 U58155 ( .A1(n55439), .A2(n55438), .ZN(n55440) );
  XOR2HSV0 U58156 ( .A1(n55441), .A2(n55440), .Z(n55442) );
  XOR2HSV0 U58157 ( .A1(n55443), .A2(n55442), .Z(n55447) );
  NAND2HSV2 U58158 ( .A1(n25840), .A2(n53863), .ZN(n55446) );
  NAND2HSV2 U58159 ( .A1(n55608), .A2(n55475), .ZN(n55445) );
  XOR3HSV2 U58160 ( .A1(n55447), .A2(n55446), .A3(n55445), .Z(\pe1/poht [27])
         );
  CLKNAND2HSV0 U58161 ( .A1(n55593), .A2(n59750), .ZN(n55483) );
  CLKNAND2HSV1 U58162 ( .A1(n55489), .A2(n55448), .ZN(n55481) );
  CLKNAND2HSV1 U58163 ( .A1(n55449), .A2(n55514), .ZN(n55474) );
  CLKNAND2HSV0 U58164 ( .A1(n54455), .A2(n55450), .ZN(n55470) );
  CLKNAND2HSV0 U58165 ( .A1(n55452), .A2(n55451), .ZN(n55454) );
  CLKNAND2HSV1 U58166 ( .A1(n55492), .A2(n55544), .ZN(n55453) );
  XOR2HSV0 U58167 ( .A1(n55454), .A2(n55453), .Z(n55468) );
  NAND2HSV2 U58168 ( .A1(n55455), .A2(\pe1/bq[9] ), .ZN(n55457) );
  CLKNAND2HSV0 U58169 ( .A1(\pe1/aot [4]), .A2(\pe1/bq[6] ), .ZN(n55456) );
  XOR2HSV0 U58170 ( .A1(n55457), .A2(n55456), .Z(n55459) );
  CLKNAND2HSV1 U58171 ( .A1(n54978), .A2(n55495), .ZN(n55458) );
  XNOR2HSV1 U58172 ( .A1(n55459), .A2(n55458), .ZN(n55467) );
  CLKNAND2HSV1 U58173 ( .A1(n55595), .A2(n55501), .ZN(n55461) );
  NAND2HSV0 U58174 ( .A1(n55496), .A2(n55505), .ZN(n55460) );
  XOR2HSV0 U58175 ( .A1(n55461), .A2(n55460), .Z(n55465) );
  CLKNAND2HSV0 U58176 ( .A1(n55547), .A2(n55518), .ZN(n55463) );
  NAND2HSV0 U58177 ( .A1(n59993), .A2(\pe1/bq[5] ), .ZN(n55462) );
  XOR2HSV0 U58178 ( .A1(n55463), .A2(n55462), .Z(n55464) );
  XOR2HSV0 U58179 ( .A1(n55465), .A2(n55464), .Z(n55466) );
  XOR3HSV2 U58180 ( .A1(n55468), .A2(n55467), .A3(n55466), .Z(n55469) );
  XNOR2HSV1 U58181 ( .A1(n55470), .A2(n55469), .ZN(n55472) );
  NAND2HSV0 U58182 ( .A1(n59751), .A2(n55340), .ZN(n55471) );
  XNOR2HSV1 U58183 ( .A1(n55472), .A2(n55471), .ZN(n55473) );
  XNOR2HSV1 U58184 ( .A1(n55474), .A2(n55473), .ZN(n55479) );
  INAND2HSV2 U58185 ( .A1(n55512), .B1(\pe1/got [4]), .ZN(n55478) );
  CLKNAND2HSV0 U58186 ( .A1(n55476), .A2(n55475), .ZN(n55477) );
  XOR3HSV2 U58187 ( .A1(n55479), .A2(n55478), .A3(n55477), .Z(n55480) );
  XOR2HSV0 U58188 ( .A1(n55481), .A2(n55480), .Z(n55482) );
  XOR2HSV0 U58189 ( .A1(n55483), .A2(n55482), .Z(n55487) );
  NAND2HSV2 U58190 ( .A1(n55484), .A2(n55339), .ZN(n55486) );
  XOR3HSV2 U58191 ( .A1(n55487), .A2(n55486), .A3(n55485), .Z(\pe1/poht [23])
         );
  CLKNAND2HSV1 U58192 ( .A1(n55492), .A2(n55491), .ZN(n55494) );
  NAND2HSV0 U58193 ( .A1(n55553), .A2(\pe1/bq[4] ), .ZN(n55493) );
  XOR2HSV0 U58194 ( .A1(n55494), .A2(n55493), .Z(n55500) );
  CLKNAND2HSV1 U58195 ( .A1(n54904), .A2(n55495), .ZN(n55498) );
  CLKNAND2HSV0 U58196 ( .A1(n55496), .A2(\pe1/bq[6] ), .ZN(n55497) );
  XOR2HSV0 U58197 ( .A1(n55498), .A2(n55497), .Z(n55499) );
  XOR2HSV0 U58198 ( .A1(n55500), .A2(n55499), .Z(n55511) );
  NAND2HSV0 U58199 ( .A1(\pe1/aot [4]), .A2(\pe1/bq[5] ), .ZN(n55503) );
  NAND2HSV0 U58200 ( .A1(n55552), .A2(n55501), .ZN(n55502) );
  XOR2HSV0 U58201 ( .A1(n55503), .A2(n55502), .Z(n55509) );
  INHSV2 U58202 ( .I(n55504), .ZN(n55578) );
  CLKNAND2HSV0 U58203 ( .A1(n55578), .A2(n55505), .ZN(n55506) );
  XOR2HSV0 U58204 ( .A1(n55507), .A2(n55506), .Z(n55508) );
  XOR2HSV0 U58205 ( .A1(n55509), .A2(n55508), .Z(n55510) );
  CLKNAND2HSV0 U58206 ( .A1(n55541), .A2(n53863), .ZN(n55536) );
  CLKNAND2HSV1 U58207 ( .A1(n55576), .A2(n55514), .ZN(n55534) );
  CLKNAND2HSV0 U58208 ( .A1(\pe1/aot [3]), .A2(n55544), .ZN(n55517) );
  CLKNAND2HSV0 U58209 ( .A1(n59993), .A2(n55605), .ZN(n55516) );
  XOR2HSV0 U58210 ( .A1(n55517), .A2(n55516), .Z(n55522) );
  NOR2HSV2 U58211 ( .A1(n54901), .A2(n55185), .ZN(n55520) );
  CLKNAND2HSV0 U58212 ( .A1(\pe1/aot [4]), .A2(n55518), .ZN(n55519) );
  XOR2HSV0 U58213 ( .A1(n55520), .A2(n55519), .Z(n55521) );
  XNOR2HSV1 U58214 ( .A1(n55522), .A2(n55521), .ZN(n55528) );
  NOR2HSV0 U58215 ( .A1(n55524), .A2(n55523), .ZN(n55526) );
  CLKNAND2HSV0 U58216 ( .A1(n55578), .A2(n54289), .ZN(n55525) );
  XOR2HSV0 U58217 ( .A1(n55526), .A2(n55525), .Z(n55527) );
  XNOR2HSV1 U58218 ( .A1(n55528), .A2(n55527), .ZN(n55532) );
  INAND2HSV2 U58219 ( .A1(n55529), .B1(n54455), .ZN(n55531) );
  NAND2HSV2 U58220 ( .A1(n59931), .A2(n59756), .ZN(n55530) );
  XOR3HSV2 U58221 ( .A1(n55532), .A2(n55531), .A3(n55530), .Z(n55533) );
  XOR2HSV0 U58222 ( .A1(n55534), .A2(n55533), .Z(n55535) );
  XOR2HSV0 U58223 ( .A1(n55536), .A2(n55535), .Z(n55540) );
  CLKNAND2HSV2 U58224 ( .A1(n55537), .A2(n55475), .ZN(n55539) );
  XOR3HSV2 U58225 ( .A1(n55540), .A2(n55539), .A3(n55538), .Z(\pe1/poht [26])
         );
  INAND2HSV0 U58226 ( .A1(n55542), .B1(n55541), .ZN(n55568) );
  CLKNAND2HSV1 U58227 ( .A1(n55543), .A2(n55267), .ZN(n55566) );
  CLKNAND2HSV1 U58228 ( .A1(n59736), .A2(n54455), .ZN(n55561) );
  CLKNAND2HSV1 U58229 ( .A1(n55578), .A2(n55231), .ZN(n55546) );
  NAND2HSV0 U58230 ( .A1(\pe1/aot [4]), .A2(n55544), .ZN(n55545) );
  XOR2HSV0 U58231 ( .A1(n55546), .A2(n55545), .Z(n55551) );
  NAND2HSV0 U58232 ( .A1(n55547), .A2(n55495), .ZN(n55549) );
  CLKNAND2HSV1 U58233 ( .A1(n55496), .A2(\pe1/bq[5] ), .ZN(n55548) );
  XOR2HSV0 U58234 ( .A1(n55549), .A2(n55548), .Z(n55550) );
  XOR2HSV0 U58235 ( .A1(n55551), .A2(n55550), .Z(n55559) );
  NAND2HSV2 U58236 ( .A1(n55552), .A2(n55505), .ZN(n55555) );
  CLKNAND2HSV0 U58237 ( .A1(n55553), .A2(n55577), .ZN(n55554) );
  XOR2HSV0 U58238 ( .A1(n55555), .A2(n55554), .Z(n55557) );
  NOR2HSV1 U58239 ( .A1(n54901), .A2(n53834), .ZN(n55556) );
  XNOR2HSV1 U58240 ( .A1(n55557), .A2(n55556), .ZN(n55558) );
  XNOR2HSV1 U58241 ( .A1(n55559), .A2(n55558), .ZN(n55560) );
  XNOR2HSV1 U58242 ( .A1(n55561), .A2(n55560), .ZN(n55564) );
  INAND2HSV2 U58243 ( .A1(n55562), .B1(n55340), .ZN(n55563) );
  XOR2HSV0 U58244 ( .A1(n55566), .A2(n55565), .Z(n55567) );
  XOR2HSV0 U58245 ( .A1(n55568), .A2(n55567), .Z(n55573) );
  NAND2HSV2 U58246 ( .A1(n55569), .A2(n55448), .ZN(n55572) );
  NAND2HSV0 U58247 ( .A1(n55570), .A2(n53513), .ZN(n55571) );
  XOR3HSV2 U58248 ( .A1(n55573), .A2(n55572), .A3(n55571), .Z(\pe1/poht [25])
         );
  INAND2HSV0 U58249 ( .A1(n55575), .B1(n55574), .ZN(n55588) );
  CLKNAND2HSV1 U58250 ( .A1(n55576), .A2(n59755), .ZN(n55586) );
  NAND2HSV2 U58251 ( .A1(n55578), .A2(n55577), .ZN(n55580) );
  CLKNAND2HSV0 U58252 ( .A1(\pe1/aot [4]), .A2(n55495), .ZN(n55579) );
  XOR2HSV0 U58253 ( .A1(n55580), .A2(n55579), .Z(n55584) );
  CLKNAND2HSV1 U58254 ( .A1(\pe1/aot [3]), .A2(n55605), .ZN(n55582) );
  NAND2HSV0 U58255 ( .A1(n59373), .A2(n55544), .ZN(n55581) );
  XOR2HSV0 U58256 ( .A1(n55582), .A2(n55581), .Z(n55583) );
  XOR2HSV0 U58257 ( .A1(n55584), .A2(n55583), .Z(n55585) );
  XOR2HSV0 U58258 ( .A1(n55586), .A2(n55585), .Z(n55587) );
  XOR2HSV0 U58259 ( .A1(n55588), .A2(n55587), .Z(n55592) );
  NAND2HSV2 U58260 ( .A1(n25839), .A2(n55319), .ZN(n55591) );
  XOR3HSV2 U58261 ( .A1(n55592), .A2(n55591), .A3(n55590), .Z(\pe1/poht [28])
         );
  INAND2HSV2 U58262 ( .A1(n55594), .B1(n55593), .ZN(n55601) );
  CLKNAND2HSV1 U58263 ( .A1(\pe1/aot [3]), .A2(n55495), .ZN(n55597) );
  CLKNAND2HSV1 U58264 ( .A1(n55595), .A2(n55451), .ZN(n55596) );
  XNOR2HSV1 U58265 ( .A1(n55597), .A2(n55596), .ZN(n55599) );
  XNOR2HSV1 U58266 ( .A1(n55599), .A2(n55598), .ZN(n55600) );
  XOR2HSV0 U58267 ( .A1(n55601), .A2(n55600), .Z(n55604) );
  XOR3HSV2 U58268 ( .A1(n55604), .A2(n55603), .A3(n55602), .Z(\pe1/poht [29])
         );
  NAND2HSV0 U58269 ( .A1(n59373), .A2(n55605), .ZN(n55606) );
  XOR2HSV0 U58270 ( .A1(n55607), .A2(n55606), .Z(n55611) );
  NAND2HSV2 U58271 ( .A1(n55608), .A2(n59756), .ZN(n55609) );
  XOR3HSV2 U58272 ( .A1(n55611), .A2(n55610), .A3(n55609), .Z(\pe1/poht [30])
         );
  INHSV2 U58273 ( .I(n55820), .ZN(n56952) );
  INAND2HSV2 U58274 ( .A1(n49314), .B1(n56952), .ZN(n55700) );
  CLKNAND2HSV1 U58275 ( .A1(n56339), .A2(n42999), .ZN(n55698) );
  CLKNAND2HSV0 U58276 ( .A1(n56780), .A2(n55823), .ZN(n55697) );
  CLKNAND2HSV1 U58277 ( .A1(n56340), .A2(n42937), .ZN(n55695) );
  CLKNAND2HSV0 U58278 ( .A1(n55946), .A2(\pe3/got [18]), .ZN(n55693) );
  CLKNHSV0 U58279 ( .I(n55612), .ZN(n55822) );
  CLKNAND2HSV1 U58280 ( .A1(n55822), .A2(\pe3/got [17]), .ZN(n55691) );
  NAND2HSV0 U58281 ( .A1(n59930), .A2(n49252), .ZN(n55689) );
  CLKNAND2HSV0 U58282 ( .A1(n49253), .A2(n56264), .ZN(n55687) );
  BUFHSV2 U58283 ( .I(n55613), .Z(n56497) );
  NAND2HSV2 U58284 ( .A1(n56497), .A2(n56493), .ZN(n55685) );
  CLKNAND2HSV0 U58285 ( .A1(n56562), .A2(n56421), .ZN(n55683) );
  NAND2HSV0 U58286 ( .A1(n55947), .A2(n56557), .ZN(n55679) );
  NAND2HSV0 U58287 ( .A1(n55824), .A2(\pe3/got [10]), .ZN(n55675) );
  CLKNAND2HSV1 U58288 ( .A1(n56067), .A2(n56068), .ZN(n55667) );
  CLKNAND2HSV1 U58289 ( .A1(n56179), .A2(n56069), .ZN(n55665) );
  CLKNAND2HSV0 U58290 ( .A1(n55949), .A2(n59807), .ZN(n55663) );
  NAND2HSV0 U58291 ( .A1(n55895), .A2(\pe3/got [1]), .ZN(n55661) );
  NAND2HSV0 U58292 ( .A1(n56434), .A2(n45807), .ZN(n55615) );
  NAND2HSV0 U58293 ( .A1(n59961), .A2(n56213), .ZN(n55614) );
  XOR2HSV0 U58294 ( .A1(n55615), .A2(n55614), .Z(n55620) );
  NAND2HSV0 U58295 ( .A1(\pe3/aot [8]), .A2(n55616), .ZN(n55618) );
  NAND2HSV0 U58296 ( .A1(n56354), .A2(n56379), .ZN(n55617) );
  XOR2HSV0 U58297 ( .A1(n55618), .A2(n55617), .Z(n55619) );
  XOR2HSV0 U58298 ( .A1(n55620), .A2(n55619), .Z(n55628) );
  NAND2HSV0 U58299 ( .A1(n56370), .A2(n45534), .ZN(n55622) );
  NAND2HSV0 U58300 ( .A1(n55873), .A2(n42971), .ZN(n55621) );
  XOR2HSV0 U58301 ( .A1(n55622), .A2(n55621), .Z(n55626) );
  NAND2HSV0 U58302 ( .A1(n56464), .A2(n55876), .ZN(n55624) );
  NAND2HSV0 U58303 ( .A1(n56508), .A2(\pe3/bq[9] ), .ZN(n55623) );
  XOR2HSV0 U58304 ( .A1(n55624), .A2(n55623), .Z(n55625) );
  XOR2HSV0 U58305 ( .A1(n55626), .A2(n55625), .Z(n55627) );
  XOR2HSV0 U58306 ( .A1(n55628), .A2(n55627), .Z(n55644) );
  NAND2HSV0 U58307 ( .A1(n59646), .A2(n49439), .ZN(n55630) );
  NAND2HSV0 U58308 ( .A1(n42940), .A2(\pe3/bq[4] ), .ZN(n55629) );
  XOR2HSV0 U58309 ( .A1(n55630), .A2(n55629), .Z(n55634) );
  CLKNAND2HSV1 U58310 ( .A1(n42818), .A2(n55828), .ZN(n55632) );
  NAND2HSV0 U58311 ( .A1(n55864), .A2(n56627), .ZN(n55631) );
  XOR2HSV0 U58312 ( .A1(n55632), .A2(n55631), .Z(n55633) );
  XOR2HSV0 U58313 ( .A1(n55634), .A2(n55633), .Z(n55642) );
  NAND2HSV2 U58314 ( .A1(n56188), .A2(n55857), .ZN(n56572) );
  NOR2HSV0 U58315 ( .A1(n55635), .A2(n56572), .ZN(n55637) );
  AOI22HSV0 U58316 ( .A1(n45695), .A2(n56971), .B1(n56188), .B2(\pe3/bq[11] ), 
        .ZN(n55636) );
  NOR2HSV2 U58317 ( .A1(n55637), .A2(n55636), .ZN(n55640) );
  NAND2HSV2 U58318 ( .A1(n55967), .A2(n56529), .ZN(n56837) );
  XOR2HSV0 U58319 ( .A1(n55640), .A2(n55639), .Z(n55641) );
  XNOR2HSV1 U58320 ( .A1(n55642), .A2(n55641), .ZN(n55643) );
  XNOR2HSV1 U58321 ( .A1(n55644), .A2(n55643), .ZN(n55659) );
  NAND2HSV2 U58322 ( .A1(n56221), .A2(n55727), .ZN(n55646) );
  NAND2HSV0 U58323 ( .A1(\pe3/aot [13]), .A2(n56688), .ZN(n55645) );
  XOR2HSV0 U58324 ( .A1(n55646), .A2(n55645), .Z(n55650) );
  CLKNAND2HSV1 U58325 ( .A1(n56113), .A2(n55970), .ZN(n55648) );
  NAND2HSV0 U58326 ( .A1(n56373), .A2(n56640), .ZN(n55647) );
  XOR2HSV0 U58327 ( .A1(n55648), .A2(n55647), .Z(n55649) );
  XOR2HSV0 U58328 ( .A1(n55650), .A2(n55649), .Z(n55657) );
  NAND2HSV0 U58329 ( .A1(n56204), .A2(n56428), .ZN(n56343) );
  XOR2HSV0 U58330 ( .A1(n55651), .A2(n56343), .Z(n55655) );
  NOR2HSV0 U58331 ( .A1(n47447), .A2(n46615), .ZN(n55653) );
  NAND2HSV0 U58332 ( .A1(n42950), .A2(\pe3/bq[7] ), .ZN(n55652) );
  XOR2HSV0 U58333 ( .A1(n55653), .A2(n55652), .Z(n55654) );
  XOR2HSV0 U58334 ( .A1(n55655), .A2(n55654), .Z(n55656) );
  XOR2HSV0 U58335 ( .A1(n55657), .A2(n55656), .Z(n55658) );
  XNOR2HSV1 U58336 ( .A1(n55659), .A2(n55658), .ZN(n55660) );
  XNOR2HSV1 U58337 ( .A1(n55661), .A2(n55660), .ZN(n55662) );
  XNOR2HSV1 U58338 ( .A1(n55663), .A2(n55662), .ZN(n55664) );
  XNOR2HSV1 U58339 ( .A1(n55665), .A2(n55664), .ZN(n55666) );
  XNOR2HSV1 U58340 ( .A1(n55667), .A2(n55666), .ZN(n55670) );
  NOR2HSV2 U58341 ( .A1(n43840), .A2(n56859), .ZN(n55669) );
  NAND2HSV0 U58342 ( .A1(n56683), .A2(n56392), .ZN(n55668) );
  XOR3HSV2 U58343 ( .A1(n55670), .A2(n55669), .A3(n55668), .Z(n55673) );
  NOR2HSV1 U58344 ( .A1(n43844), .A2(n56778), .ZN(n55672) );
  NAND2HSV0 U58345 ( .A1(n56396), .A2(n56855), .ZN(n55671) );
  XOR3HSV2 U58346 ( .A1(n55673), .A2(n55672), .A3(n55671), .Z(n55674) );
  XNOR2HSV1 U58347 ( .A1(n55675), .A2(n55674), .ZN(n55677) );
  CLKNAND2HSV1 U58348 ( .A1(n55912), .A2(\pe3/got [9]), .ZN(n55676) );
  XNOR2HSV1 U58349 ( .A1(n55677), .A2(n55676), .ZN(n55678) );
  XNOR2HSV1 U58350 ( .A1(n55679), .A2(n55678), .ZN(n55681) );
  NOR2HSV1 U58351 ( .A1(n56406), .A2(n50802), .ZN(n55680) );
  XNOR2HSV1 U58352 ( .A1(n55681), .A2(n55680), .ZN(n55682) );
  XNOR2HSV1 U58353 ( .A1(n55683), .A2(n55682), .ZN(n55684) );
  XOR2HSV0 U58354 ( .A1(n55685), .A2(n55684), .Z(n55686) );
  XNOR2HSV1 U58355 ( .A1(n55687), .A2(n55686), .ZN(n55688) );
  XNOR2HSV1 U58356 ( .A1(n55689), .A2(n55688), .ZN(n55690) );
  XNOR2HSV1 U58357 ( .A1(n55691), .A2(n55690), .ZN(n55692) );
  XNOR2HSV1 U58358 ( .A1(n55693), .A2(n55692), .ZN(n55694) );
  XNOR2HSV1 U58359 ( .A1(n55695), .A2(n55694), .ZN(n55696) );
  XNOR2HSV1 U58360 ( .A1(n55700), .A2(n55699), .ZN(n55704) );
  NAND2HSV2 U58361 ( .A1(n56899), .A2(n55701), .ZN(n55703) );
  CLKNAND2HSV1 U58362 ( .A1(n56976), .A2(\pe3/got [23]), .ZN(n55702) );
  XOR3HSV2 U58363 ( .A1(n55704), .A2(n55703), .A3(n55702), .Z(\pe3/poht [8])
         );
  INHSV2 U58364 ( .I(n55820), .ZN(n56905) );
  CLKNAND2HSV1 U58365 ( .A1(n56905), .A2(n56057), .ZN(n55817) );
  CLKNAND2HSV1 U58366 ( .A1(n48480), .A2(n45947), .ZN(n55815) );
  CLKNAND2HSV0 U58367 ( .A1(n55944), .A2(n59384), .ZN(n55813) );
  CLKNAND2HSV1 U58368 ( .A1(n56340), .A2(\pe3/got [24]), .ZN(n55812) );
  CLKNAND2HSV0 U58369 ( .A1(n59527), .A2(n42673), .ZN(n55810) );
  CLKNAND2HSV0 U58370 ( .A1(n55822), .A2(n48485), .ZN(n55808) );
  NAND2HSV0 U58371 ( .A1(n56736), .A2(n43262), .ZN(n55806) );
  CLKNAND2HSV0 U58372 ( .A1(n49253), .A2(n55823), .ZN(n55804) );
  CLKNAND2HSV0 U58373 ( .A1(n59920), .A2(n56489), .ZN(n55802) );
  CLKNAND2HSV0 U58374 ( .A1(n56562), .A2(\pe3/got [18]), .ZN(n55800) );
  NAND2HSV0 U58375 ( .A1(n55947), .A2(n49252), .ZN(n55796) );
  NAND2HSV0 U58376 ( .A1(n55824), .A2(n56264), .ZN(n55792) );
  NAND2HSV0 U58377 ( .A1(n56067), .A2(n59645), .ZN(n55784) );
  NAND2HSV0 U58378 ( .A1(n49255), .A2(n56855), .ZN(n55782) );
  NAND2HSV0 U58379 ( .A1(n55706), .A2(n56241), .ZN(n55780) );
  NAND2HSV0 U58380 ( .A1(n56070), .A2(n56267), .ZN(n55776) );
  NAND2HSV0 U58381 ( .A1(n55707), .A2(n56068), .ZN(n55774) );
  CLKNAND2HSV1 U58382 ( .A1(n37176), .A2(n56069), .ZN(n55772) );
  NAND2HSV0 U58383 ( .A1(n55826), .A2(n59807), .ZN(n55770) );
  NAND2HSV0 U58384 ( .A1(n55873), .A2(n55976), .ZN(n55709) );
  NAND2HSV0 U58385 ( .A1(n59646), .A2(\pe3/bq[26] ), .ZN(n55708) );
  XOR2HSV0 U58386 ( .A1(n55709), .A2(n55708), .Z(n55713) );
  NOR2HSV0 U58387 ( .A1(n45567), .A2(n49272), .ZN(n55711) );
  NAND2HSV0 U58388 ( .A1(n56354), .A2(\pe3/bq[19] ), .ZN(n55710) );
  XOR2HSV0 U58389 ( .A1(n55711), .A2(n55710), .Z(n55712) );
  XNOR2HSV1 U58390 ( .A1(n55713), .A2(n55712), .ZN(n55723) );
  NOR2HSV0 U58391 ( .A1(n55714), .A2(n56914), .ZN(n55716) );
  NAND2HSV0 U58392 ( .A1(\pe3/aot [19]), .A2(\pe3/bq[11] ), .ZN(n55715) );
  XOR2HSV0 U58393 ( .A1(n55716), .A2(n55715), .Z(n55721) );
  NAND2HSV2 U58394 ( .A1(n43030), .A2(n55857), .ZN(n56632) );
  NOR2HSV0 U58395 ( .A1(n55717), .A2(n56632), .ZN(n55719) );
  AOI22HSV0 U58396 ( .A1(n37373), .A2(n56971), .B1(n43030), .B2(n56379), .ZN(
        n55718) );
  NOR2HSV2 U58397 ( .A1(n55719), .A2(n55718), .ZN(n55720) );
  XNOR2HSV1 U58398 ( .A1(n55721), .A2(n55720), .ZN(n55722) );
  XNOR2HSV1 U58399 ( .A1(n55723), .A2(n55722), .ZN(n55732) );
  NAND2HSV0 U58400 ( .A1(n55864), .A2(\pe3/bq[3] ), .ZN(n56650) );
  NAND2HSV0 U58401 ( .A1(n56373), .A2(n56218), .ZN(n55848) );
  XNOR2HSV1 U58402 ( .A1(n55726), .A2(n55848), .ZN(n55730) );
  NAND2HSV0 U58403 ( .A1(n56370), .A2(n55727), .ZN(n55854) );
  NAND2HSV0 U58404 ( .A1(n42940), .A2(n56785), .ZN(n55728) );
  XOR2HSV0 U58405 ( .A1(n55854), .A2(n55728), .Z(n55729) );
  XOR2HSV0 U58406 ( .A1(n55730), .A2(n55729), .Z(n55731) );
  XNOR2HSV1 U58407 ( .A1(n55732), .A2(n55731), .ZN(n55768) );
  NAND2HSV0 U58408 ( .A1(n56434), .A2(n55960), .ZN(n55734) );
  NAND2HSV0 U58409 ( .A1(n56188), .A2(n56640), .ZN(n55733) );
  XOR2HSV0 U58410 ( .A1(n55734), .A2(n55733), .Z(n55739) );
  NAND2HSV0 U58411 ( .A1(n42950), .A2(n56688), .ZN(n55737) );
  NAND2HSV0 U58412 ( .A1(n56970), .A2(n55735), .ZN(n55736) );
  XOR2HSV0 U58413 ( .A1(n55737), .A2(n55736), .Z(n55738) );
  XOR2HSV0 U58414 ( .A1(n55739), .A2(n55738), .Z(n55747) );
  NAND2HSV0 U58415 ( .A1(n59627), .A2(n56213), .ZN(n55741) );
  NAND2HSV0 U58416 ( .A1(\pe3/aot [8]), .A2(n45807), .ZN(n55740) );
  XOR2HSV0 U58417 ( .A1(n55741), .A2(n55740), .Z(n55745) );
  NAND2HSV0 U58418 ( .A1(n55967), .A2(n55872), .ZN(n55743) );
  NAND2HSV0 U58419 ( .A1(n56204), .A2(n56627), .ZN(n55742) );
  XOR2HSV0 U58420 ( .A1(n55743), .A2(n55742), .Z(n55744) );
  XOR2HSV0 U58421 ( .A1(n55745), .A2(n55744), .Z(n55746) );
  XOR2HSV0 U58422 ( .A1(n55747), .A2(n55746), .Z(n55765) );
  NAND2HSV0 U58423 ( .A1(n42743), .A2(\pe3/bq[4] ), .ZN(n55749) );
  NAND2HSV0 U58424 ( .A1(n56087), .A2(n55876), .ZN(n55748) );
  XOR2HSV0 U58425 ( .A1(n55749), .A2(n55748), .Z(n55754) );
  NAND2HSV0 U58426 ( .A1(n42818), .A2(n56832), .ZN(n55752) );
  NAND2HSV0 U58427 ( .A1(n55750), .A2(n55828), .ZN(n55751) );
  XOR2HSV0 U58428 ( .A1(n55752), .A2(n55751), .Z(n55753) );
  XOR2HSV0 U58429 ( .A1(n55754), .A2(n55753), .Z(n55763) );
  NAND2HSV0 U58430 ( .A1(\pe3/aot [13]), .A2(n56433), .ZN(n55757) );
  NAND2HSV0 U58431 ( .A1(n56740), .A2(n42971), .ZN(n55756) );
  XOR2HSV0 U58432 ( .A1(n55757), .A2(n55756), .Z(n55761) );
  NOR2HSV0 U58433 ( .A1(n43527), .A2(n49423), .ZN(n55759) );
  NAND2HSV0 U58434 ( .A1(n59961), .A2(n37280), .ZN(n55758) );
  XOR2HSV0 U58435 ( .A1(n55759), .A2(n55758), .Z(n55760) );
  XOR2HSV0 U58436 ( .A1(n55761), .A2(n55760), .Z(n55762) );
  XOR2HSV0 U58437 ( .A1(n55763), .A2(n55762), .Z(n55764) );
  XOR2HSV0 U58438 ( .A1(n55765), .A2(n55764), .Z(n55767) );
  NAND2HSV0 U58439 ( .A1(n59671), .A2(n56975), .ZN(n55766) );
  XOR3HSV2 U58440 ( .A1(n55768), .A2(n55767), .A3(n55766), .Z(n55769) );
  XNOR2HSV1 U58441 ( .A1(n55770), .A2(n55769), .ZN(n55771) );
  XNOR2HSV1 U58442 ( .A1(n55772), .A2(n55771), .ZN(n55773) );
  XNOR2HSV1 U58443 ( .A1(n55774), .A2(n55773), .ZN(n55775) );
  XNOR2HSV1 U58444 ( .A1(n55776), .A2(n55775), .ZN(n55778) );
  NAND2HSV0 U58445 ( .A1(n56127), .A2(n56683), .ZN(n55777) );
  XNOR2HSV1 U58446 ( .A1(n55778), .A2(n55777), .ZN(n55779) );
  XNOR2HSV1 U58447 ( .A1(n55780), .A2(n55779), .ZN(n55781) );
  XNOR2HSV1 U58448 ( .A1(n55782), .A2(n55781), .ZN(n55783) );
  XNOR2HSV1 U58449 ( .A1(n55784), .A2(n55783), .ZN(n55787) );
  NOR2HSV0 U58450 ( .A1(n56391), .A2(n50756), .ZN(n55786) );
  NAND2HSV0 U58451 ( .A1(n56392), .A2(n56247), .ZN(n55785) );
  XOR3HSV1 U58452 ( .A1(n55787), .A2(n55786), .A3(n55785), .Z(n55790) );
  NOR2HSV1 U58453 ( .A1(n43844), .A2(n50802), .ZN(n55789) );
  NAND2HSV0 U58454 ( .A1(n56396), .A2(n56421), .ZN(n55788) );
  XOR3HSV2 U58455 ( .A1(n55790), .A2(n55789), .A3(n55788), .Z(n55791) );
  XNOR2HSV1 U58456 ( .A1(n55792), .A2(n55791), .ZN(n55794) );
  NAND2HSV0 U58457 ( .A1(n55912), .A2(n56493), .ZN(n55793) );
  XNOR2HSV1 U58458 ( .A1(n55794), .A2(n55793), .ZN(n55795) );
  XNOR2HSV1 U58459 ( .A1(n55796), .A2(n55795), .ZN(n55798) );
  NOR2HSV0 U58460 ( .A1(n56406), .A2(n44693), .ZN(n55797) );
  XNOR2HSV1 U58461 ( .A1(n55798), .A2(n55797), .ZN(n55799) );
  XNOR2HSV1 U58462 ( .A1(n55800), .A2(n55799), .ZN(n55801) );
  XNOR2HSV1 U58463 ( .A1(n55802), .A2(n55801), .ZN(n55803) );
  XNOR2HSV1 U58464 ( .A1(n55804), .A2(n55803), .ZN(n55805) );
  XNOR2HSV1 U58465 ( .A1(n55806), .A2(n55805), .ZN(n55807) );
  XNOR2HSV1 U58466 ( .A1(n55808), .A2(n55807), .ZN(n55809) );
  XNOR2HSV1 U58467 ( .A1(n55810), .A2(n55809), .ZN(n55811) );
  XNOR2HSV1 U58468 ( .A1(n55815), .A2(n55814), .ZN(n55816) );
  CLKNAND2HSV2 U58469 ( .A1(n56676), .A2(n59963), .ZN(n55819) );
  CLKNAND2HSV1 U58470 ( .A1(n56490), .A2(n59964), .ZN(n55818) );
  INHSV2 U58471 ( .I(n55820), .ZN(n56860) );
  CLKNAND2HSV1 U58472 ( .A1(n56860), .A2(n45947), .ZN(n55939) );
  CLKNAND2HSV1 U58473 ( .A1(n56907), .A2(n59384), .ZN(n55937) );
  CLKNAND2HSV0 U58474 ( .A1(n55822), .A2(n56171), .ZN(n55929) );
  NAND2HSV0 U58475 ( .A1(n59930), .A2(n55823), .ZN(n55927) );
  CLKNAND2HSV0 U58476 ( .A1(n56561), .A2(n56489), .ZN(n55925) );
  NAND2HSV0 U58477 ( .A1(n56737), .A2(\pe3/got [18]), .ZN(n55923) );
  NAND2HSV0 U58478 ( .A1(n56685), .A2(n56064), .ZN(n55921) );
  CLKNAND2HSV0 U58479 ( .A1(n56624), .A2(n56174), .ZN(n55916) );
  NAND2HSV0 U58480 ( .A1(n55824), .A2(n56493), .ZN(n55911) );
  NAND2HSV0 U58481 ( .A1(n56067), .A2(n56855), .ZN(n55903) );
  CLKNAND2HSV0 U58482 ( .A1(n56179), .A2(n56241), .ZN(n55901) );
  NAND2HSV0 U58483 ( .A1(n55949), .A2(n56683), .ZN(n55899) );
  NAND2HSV0 U58484 ( .A1(n56070), .A2(n56068), .ZN(n55894) );
  NAND2HSV0 U58485 ( .A1(n55825), .A2(n56069), .ZN(n55892) );
  CLKNAND2HSV1 U58486 ( .A1(n46314), .A2(n55950), .ZN(n55890) );
  NAND2HSV0 U58487 ( .A1(n55826), .A2(\pe3/got [1]), .ZN(n55888) );
  NAND2HSV0 U58488 ( .A1(n55828), .A2(n55827), .ZN(n55985) );
  XOR2HSV0 U58489 ( .A1(n55829), .A2(n55985), .Z(n55833) );
  NOR2HSV0 U58490 ( .A1(n56382), .A2(n46138), .ZN(n55831) );
  NAND2HSV0 U58491 ( .A1(n56464), .A2(n56187), .ZN(n55830) );
  XOR2HSV0 U58492 ( .A1(n55831), .A2(n55830), .Z(n55832) );
  XOR2HSV0 U58493 ( .A1(n55833), .A2(n55832), .Z(n55886) );
  NAND2HSV0 U58494 ( .A1(n56074), .A2(n56071), .ZN(n55835) );
  NAND2HSV0 U58495 ( .A1(n56113), .A2(n56688), .ZN(n55834) );
  XOR2HSV0 U58496 ( .A1(n55835), .A2(n55834), .Z(n55839) );
  NAND2HSV0 U58497 ( .A1(n42950), .A2(\pe3/bq[11] ), .ZN(n55837) );
  NAND2HSV0 U58498 ( .A1(\pe3/aot [14]), .A2(n56094), .ZN(n55836) );
  XOR2HSV0 U58499 ( .A1(n55837), .A2(n55836), .Z(n55838) );
  XOR2HSV0 U58500 ( .A1(n55839), .A2(n55838), .Z(n55847) );
  NAND2HSV0 U58501 ( .A1(\pe3/aot [22]), .A2(n45639), .ZN(n55841) );
  NAND2HSV0 U58502 ( .A1(n56434), .A2(\pe3/bq[26] ), .ZN(n55840) );
  XOR2HSV0 U58503 ( .A1(n55841), .A2(n55840), .Z(n55845) );
  NAND2HSV0 U58504 ( .A1(n43030), .A2(n55975), .ZN(n55843) );
  NAND2HSV0 U58505 ( .A1(n59961), .A2(n55960), .ZN(n55842) );
  XOR2HSV0 U58506 ( .A1(n55843), .A2(n55842), .Z(n55844) );
  XNOR2HSV1 U58507 ( .A1(n55845), .A2(n55844), .ZN(n55846) );
  XNOR2HSV1 U58508 ( .A1(n55847), .A2(n55846), .ZN(n55885) );
  NAND2HSV0 U58509 ( .A1(\pe3/aot [8]), .A2(\pe3/bq[20] ), .ZN(n55991) );
  NOR2HSV0 U58510 ( .A1(n55849), .A2(n56703), .ZN(n55851) );
  AOI22HSV0 U58511 ( .A1(n55988), .A2(n56529), .B1(\pe3/bq[19] ), .B2(n56740), 
        .ZN(n55850) );
  NOR2HSV1 U58512 ( .A1(n55851), .A2(n55850), .ZN(n55852) );
  XOR2HSV0 U58513 ( .A1(n55853), .A2(n55852), .Z(n55863) );
  NAND2HSV0 U58514 ( .A1(\pe3/aot [11]), .A2(n56433), .ZN(n55999) );
  NOR2HSV0 U58515 ( .A1(n55854), .A2(n55999), .ZN(n55856) );
  AOI22HSV0 U58516 ( .A1(n56354), .A2(\pe3/bq[18] ), .B1(n56433), .B2(n56575), 
        .ZN(n55855) );
  NOR2HSV2 U58517 ( .A1(n55856), .A2(n55855), .ZN(n55861) );
  NAND2HSV0 U58518 ( .A1(n55858), .A2(n55857), .ZN(n56097) );
  XNOR2HSV1 U58519 ( .A1(n55861), .A2(n55860), .ZN(n55862) );
  XNOR2HSV1 U58520 ( .A1(n55863), .A2(n55862), .ZN(n55884) );
  NAND2HSV0 U58521 ( .A1(n55864), .A2(n56379), .ZN(n55866) );
  NAND2HSV0 U58522 ( .A1(\pe3/aot [21]), .A2(n55970), .ZN(n55865) );
  XOR2HSV0 U58523 ( .A1(n55866), .A2(n55865), .Z(n55871) );
  NAND2HSV0 U58524 ( .A1(n59511), .A2(n55867), .ZN(n55869) );
  NAND2HSV0 U58525 ( .A1(n56864), .A2(n45807), .ZN(n55868) );
  XOR2HSV0 U58526 ( .A1(n55869), .A2(n55868), .Z(n55870) );
  XOR2HSV0 U58527 ( .A1(n55871), .A2(n55870), .Z(n55882) );
  NAND2HSV0 U58528 ( .A1(n55873), .A2(n55872), .ZN(n55875) );
  NAND2HSV0 U58529 ( .A1(n55967), .A2(n56213), .ZN(n55874) );
  XOR2HSV0 U58530 ( .A1(n55875), .A2(n55874), .Z(n55880) );
  NAND2HSV0 U58531 ( .A1(n42818), .A2(n55876), .ZN(n55878) );
  NAND2HSV0 U58532 ( .A1(n56087), .A2(n56189), .ZN(n55877) );
  XOR2HSV0 U58533 ( .A1(n55878), .A2(n55877), .Z(n55879) );
  XOR2HSV0 U58534 ( .A1(n55880), .A2(n55879), .Z(n55881) );
  XOR2HSV0 U58535 ( .A1(n55882), .A2(n55881), .Z(n55883) );
  XOR4HSV1 U58536 ( .A1(n55886), .A2(n55885), .A3(n55884), .A4(n55883), .Z(
        n55887) );
  XNOR2HSV1 U58537 ( .A1(n55888), .A2(n55887), .ZN(n55889) );
  XNOR2HSV1 U58538 ( .A1(n55890), .A2(n55889), .ZN(n55891) );
  XNOR2HSV1 U58539 ( .A1(n55892), .A2(n55891), .ZN(n55893) );
  XNOR2HSV1 U58540 ( .A1(n55894), .A2(n55893), .ZN(n55897) );
  NAND2HSV0 U58541 ( .A1(n55895), .A2(n56267), .ZN(n55896) );
  XNOR2HSV1 U58542 ( .A1(n55897), .A2(n55896), .ZN(n55898) );
  XNOR2HSV1 U58543 ( .A1(n55899), .A2(n55898), .ZN(n55900) );
  XNOR2HSV1 U58544 ( .A1(n55901), .A2(n55900), .ZN(n55902) );
  XNOR2HSV1 U58545 ( .A1(n55903), .A2(n55902), .ZN(n55906) );
  NOR2HSV1 U58546 ( .A1(n45728), .A2(n56680), .ZN(n55905) );
  NAND2HSV0 U58547 ( .A1(n56422), .A2(n56619), .ZN(n55904) );
  XOR3HSV2 U58548 ( .A1(n55906), .A2(n55905), .A3(n55904), .Z(n55909) );
  NOR2HSV1 U58549 ( .A1(n56475), .A2(n50799), .ZN(n55908) );
  CLKNAND2HSV1 U58550 ( .A1(n56242), .A2(n56494), .ZN(n55907) );
  XOR3HSV2 U58551 ( .A1(n55909), .A2(n55908), .A3(n55907), .Z(n55910) );
  XNOR2HSV1 U58552 ( .A1(n55911), .A2(n55910), .ZN(n55914) );
  CLKNAND2HSV0 U58553 ( .A1(n55912), .A2(n56421), .ZN(n55913) );
  XNOR2HSV1 U58554 ( .A1(n55914), .A2(n55913), .ZN(n55915) );
  XNOR2HSV1 U58555 ( .A1(n55916), .A2(n55915), .ZN(n55919) );
  NOR2HSV0 U58556 ( .A1(n55917), .A2(n45576), .ZN(n55918) );
  XNOR2HSV1 U58557 ( .A1(n55919), .A2(n55918), .ZN(n55920) );
  XNOR2HSV1 U58558 ( .A1(n55921), .A2(n55920), .ZN(n55922) );
  XNOR2HSV1 U58559 ( .A1(n55923), .A2(n55922), .ZN(n55924) );
  XNOR2HSV1 U58560 ( .A1(n55925), .A2(n55924), .ZN(n55926) );
  XNOR2HSV1 U58561 ( .A1(n55927), .A2(n55926), .ZN(n55928) );
  XNOR2HSV1 U58562 ( .A1(n55929), .A2(n55928), .ZN(n55930) );
  XNOR2HSV1 U58563 ( .A1(n55931), .A2(n55930), .ZN(n55932) );
  XNOR2HSV1 U58564 ( .A1(n55933), .A2(n55932), .ZN(n55934) );
  XOR2HSV0 U58565 ( .A1(n55935), .A2(n55934), .Z(n55936) );
  XNOR2HSV1 U58566 ( .A1(n55937), .A2(n55936), .ZN(n55938) );
  CLKNAND2HSV1 U58567 ( .A1(n56490), .A2(n56057), .ZN(n55942) );
  XOR3HSV2 U58568 ( .A1(n55943), .A2(n55942), .A3(n55941), .Z(\pe3/poht [4])
         );
  CLKNAND2HSV1 U58569 ( .A1(n56952), .A2(n37175), .ZN(n56056) );
  CLKNAND2HSV1 U58570 ( .A1(n48480), .A2(n59617), .ZN(n56054) );
  NAND2HSV0 U58571 ( .A1(n55944), .A2(n42673), .ZN(n56052) );
  CLKNAND2HSV1 U58572 ( .A1(n56173), .A2(n48485), .ZN(n56051) );
  CLKNAND2HSV0 U58573 ( .A1(n55946), .A2(n55945), .ZN(n56049) );
  NAND2HSV0 U58574 ( .A1(n56063), .A2(n42996), .ZN(n56047) );
  NAND2HSV0 U58575 ( .A1(n59930), .A2(n56489), .ZN(n56045) );
  CLKNAND2HSV0 U58576 ( .A1(n49253), .A2(\pe3/got [18]), .ZN(n56043) );
  NAND2HSV0 U58577 ( .A1(n56737), .A2(n56335), .ZN(n56041) );
  NAND2HSV0 U58578 ( .A1(n56685), .A2(n49252), .ZN(n56039) );
  NAND2HSV0 U58579 ( .A1(n55947), .A2(n56493), .ZN(n56035) );
  CLKNAND2HSV1 U58580 ( .A1(n56178), .A2(n56421), .ZN(n56031) );
  NAND2HSV0 U58581 ( .A1(n55948), .A2(n56241), .ZN(n56023) );
  NAND2HSV0 U58582 ( .A1(n49255), .A2(n56683), .ZN(n56021) );
  CLKNAND2HSV1 U58583 ( .A1(n55949), .A2(n56623), .ZN(n56019) );
  NAND2HSV0 U58584 ( .A1(n56070), .A2(n56069), .ZN(n56015) );
  NAND2HSV0 U58585 ( .A1(n49405), .A2(n55950), .ZN(n56013) );
  NAND2HSV0 U58586 ( .A1(n55951), .A2(\pe3/got [1]), .ZN(n56011) );
  NAND2HSV0 U58587 ( .A1(n56520), .A2(\pe3/bq[19] ), .ZN(n55953) );
  NAND2HSV0 U58588 ( .A1(\pe3/aot [22]), .A2(n56915), .ZN(n55952) );
  XOR2HSV0 U58589 ( .A1(n55953), .A2(n55952), .Z(n55957) );
  NAND2HSV0 U58590 ( .A1(n59646), .A2(n55872), .ZN(n55955) );
  NAND2HSV0 U58591 ( .A1(\pe3/aot [21]), .A2(n56832), .ZN(n55954) );
  XOR2HSV0 U58592 ( .A1(n55955), .A2(n55954), .Z(n55956) );
  XOR2HSV0 U58593 ( .A1(n55957), .A2(n55956), .Z(n55966) );
  NAND2HSV0 U58594 ( .A1(n56864), .A2(n56106), .ZN(n55959) );
  NAND2HSV0 U58595 ( .A1(\pe3/aot [13]), .A2(n56094), .ZN(n55958) );
  XOR2HSV0 U58596 ( .A1(n55959), .A2(n55958), .Z(n55964) );
  NAND2HSV0 U58597 ( .A1(n42950), .A2(n56187), .ZN(n55962) );
  NAND2HSV0 U58598 ( .A1(n59511), .A2(n55960), .ZN(n55961) );
  XOR2HSV0 U58599 ( .A1(n55962), .A2(n55961), .Z(n55963) );
  XOR2HSV0 U58600 ( .A1(n55964), .A2(n55963), .Z(n55965) );
  XOR2HSV0 U58601 ( .A1(n55966), .A2(n55965), .Z(n55984) );
  NAND2HSV0 U58602 ( .A1(n55967), .A2(n45807), .ZN(n55969) );
  NAND2HSV0 U58603 ( .A1(n56439), .A2(n56213), .ZN(n55968) );
  XOR2HSV0 U58604 ( .A1(n55969), .A2(n55968), .Z(n55974) );
  NAND2HSV0 U58605 ( .A1(n42818), .A2(n56189), .ZN(n55972) );
  NAND2HSV0 U58606 ( .A1(\pe3/aot [20]), .A2(n55970), .ZN(n55971) );
  XOR2HSV0 U58607 ( .A1(n55972), .A2(n55971), .Z(n55973) );
  XOR2HSV0 U58608 ( .A1(n55974), .A2(n55973), .Z(n55982) );
  CLKNAND2HSV0 U58609 ( .A1(n56508), .A2(n56688), .ZN(n56506) );
  CLKNAND2HSV1 U58610 ( .A1(n56378), .A2(n55975), .ZN(n56531) );
  XOR2HSV0 U58611 ( .A1(n56506), .A2(n56531), .Z(n55980) );
  NAND2HSV0 U58612 ( .A1(n56434), .A2(n55976), .ZN(n55978) );
  NAND2HSV0 U58613 ( .A1(n56370), .A2(n56640), .ZN(n55977) );
  XOR2HSV0 U58614 ( .A1(n55978), .A2(n55977), .Z(n55979) );
  XOR2HSV0 U58615 ( .A1(n55980), .A2(n55979), .Z(n55981) );
  XOR2HSV0 U58616 ( .A1(n55982), .A2(n55981), .Z(n55983) );
  XOR2HSV0 U58617 ( .A1(n55984), .A2(n55983), .Z(n56009) );
  NOR2HSV1 U58618 ( .A1(n55986), .A2(n55985), .ZN(n55990) );
  AOI22HSV0 U58619 ( .A1(n55988), .A2(n56892), .B1(n55987), .B2(n56824), .ZN(
        n55989) );
  NOR2HSV2 U58620 ( .A1(n55990), .A2(n55989), .ZN(n55992) );
  XOR2HSV0 U58621 ( .A1(n55992), .A2(n55991), .Z(n56007) );
  NAND2HSV0 U58622 ( .A1(n56464), .A2(\pe3/bq[9] ), .ZN(n55994) );
  NAND2HSV0 U58623 ( .A1(n59961), .A2(\pe3/bq[26] ), .ZN(n55993) );
  XOR2HSV0 U58624 ( .A1(n55994), .A2(n55993), .Z(n55998) );
  NAND2HSV0 U58625 ( .A1(\pe3/aot [10]), .A2(\pe3/bq[18] ), .ZN(n55996) );
  NAND2HSV0 U58626 ( .A1(\pe3/aot [14]), .A2(n56379), .ZN(n55995) );
  XOR2HSV0 U58627 ( .A1(n55996), .A2(n55995), .Z(n55997) );
  XNOR2HSV1 U58628 ( .A1(n55998), .A2(n55997), .ZN(n56006) );
  XOR2HSV0 U58629 ( .A1(n56000), .A2(n55999), .Z(n56004) );
  NOR2HSV0 U58630 ( .A1(n43527), .A2(n56001), .ZN(n56424) );
  XOR2HSV0 U58631 ( .A1(n56424), .A2(n56002), .Z(n56003) );
  XOR2HSV0 U58632 ( .A1(n56004), .A2(n56003), .Z(n56005) );
  XOR3HSV2 U58633 ( .A1(n56007), .A2(n56006), .A3(n56005), .Z(n56008) );
  XNOR2HSV1 U58634 ( .A1(n56009), .A2(n56008), .ZN(n56010) );
  XNOR2HSV1 U58635 ( .A1(n56011), .A2(n56010), .ZN(n56012) );
  XNOR2HSV1 U58636 ( .A1(n56013), .A2(n56012), .ZN(n56014) );
  XNOR2HSV1 U58637 ( .A1(n56015), .A2(n56014), .ZN(n56017) );
  NAND2HSV0 U58638 ( .A1(n56127), .A2(n56068), .ZN(n56016) );
  XNOR2HSV1 U58639 ( .A1(n56017), .A2(n56016), .ZN(n56018) );
  XNOR2HSV1 U58640 ( .A1(n56019), .A2(n56018), .ZN(n56020) );
  XNOR2HSV1 U58641 ( .A1(n56021), .A2(n56020), .ZN(n56022) );
  XNOR2HSV1 U58642 ( .A1(n56023), .A2(n56022), .ZN(n56026) );
  NOR2HSV0 U58643 ( .A1(n43840), .A2(n56496), .ZN(n56025) );
  NAND2HSV0 U58644 ( .A1(n56620), .A2(n56392), .ZN(n56024) );
  XOR3HSV1 U58645 ( .A1(n56026), .A2(n56025), .A3(n56024), .Z(n56029) );
  NOR2HSV1 U58646 ( .A1(n56475), .A2(n50756), .ZN(n56028) );
  CLKNAND2HSV0 U58647 ( .A1(n56242), .A2(n56247), .ZN(n56027) );
  XOR3HSV2 U58648 ( .A1(n56029), .A2(n56028), .A3(n56027), .Z(n56030) );
  XNOR2HSV1 U58649 ( .A1(n56031), .A2(n56030), .ZN(n56033) );
  CLKNAND2HSV0 U58650 ( .A1(n46052), .A2(n56494), .ZN(n56032) );
  XNOR2HSV1 U58651 ( .A1(n56033), .A2(n56032), .ZN(n56034) );
  XNOR2HSV1 U58652 ( .A1(n56035), .A2(n56034), .ZN(n56037) );
  NAND2HSV0 U58653 ( .A1(n43463), .A2(n56174), .ZN(n56036) );
  XNOR2HSV1 U58654 ( .A1(n56037), .A2(n56036), .ZN(n56038) );
  XNOR2HSV1 U58655 ( .A1(n56039), .A2(n56038), .ZN(n56040) );
  XNOR2HSV1 U58656 ( .A1(n56041), .A2(n56040), .ZN(n56042) );
  XNOR2HSV1 U58657 ( .A1(n56043), .A2(n56042), .ZN(n56044) );
  XNOR2HSV1 U58658 ( .A1(n56045), .A2(n56044), .ZN(n56046) );
  XNOR2HSV1 U58659 ( .A1(n56047), .A2(n56046), .ZN(n56048) );
  XNOR2HSV1 U58660 ( .A1(n56049), .A2(n56048), .ZN(n56050) );
  XOR2HSV0 U58661 ( .A1(n56054), .A2(n56053), .Z(n56055) );
  XNOR2HSV1 U58662 ( .A1(n56056), .A2(n56055), .ZN(n56062) );
  NAND2HSV2 U58663 ( .A1(n56899), .A2(n56057), .ZN(n56061) );
  CLKNAND2HSV1 U58664 ( .A1(n56900), .A2(n45947), .ZN(n56060) );
  XOR3HSV2 U58665 ( .A1(n56062), .A2(n56061), .A3(n56060), .Z(\pe3/poht [5])
         );
  CLKNAND2HSV0 U58666 ( .A1(n56905), .A2(n42673), .ZN(n56167) );
  CLKNAND2HSV1 U58667 ( .A1(n59527), .A2(n59965), .ZN(n56162) );
  NAND2HSV0 U58668 ( .A1(n56063), .A2(\pe3/got [18]), .ZN(n56160) );
  CLKNAND2HSV0 U58669 ( .A1(n56783), .A2(n56064), .ZN(n56158) );
  CLKNAND2HSV1 U58670 ( .A1(n56561), .A2(n56065), .ZN(n56156) );
  CLKNAND2HSV1 U58671 ( .A1(n56497), .A2(n56174), .ZN(n56154) );
  NAND2HSV0 U58672 ( .A1(n56066), .A2(n56493), .ZN(n56152) );
  CLKNAND2HSV1 U58673 ( .A1(n53228), .A2(n56176), .ZN(n56148) );
  CLKNAND2HSV1 U58674 ( .A1(n45636), .A2(n56247), .ZN(n56144) );
  NAND2HSV0 U58675 ( .A1(n56067), .A2(n56822), .ZN(n56135) );
  CLKNAND2HSV1 U58676 ( .A1(n43373), .A2(n56068), .ZN(n56133) );
  NAND2HSV0 U58677 ( .A1(n56180), .A2(n56069), .ZN(n56131) );
  NAND2HSV0 U58678 ( .A1(n56070), .A2(\pe3/got [1]), .ZN(n56126) );
  NAND2HSV0 U58679 ( .A1(n59511), .A2(n56071), .ZN(n56073) );
  NAND2HSV0 U58680 ( .A1(n56740), .A2(n56640), .ZN(n56072) );
  XOR2HSV0 U58681 ( .A1(n56073), .A2(n56072), .Z(n56078) );
  NAND2HSV0 U58682 ( .A1(n59961), .A2(n43052), .ZN(n56076) );
  NAND2HSV0 U58683 ( .A1(n56074), .A2(n56222), .ZN(n56075) );
  XOR2HSV0 U58684 ( .A1(n56076), .A2(n56075), .Z(n56077) );
  XOR2HSV0 U58685 ( .A1(n56078), .A2(n56077), .Z(n56086) );
  CLKNAND2HSV0 U58686 ( .A1(n56434), .A2(n56213), .ZN(n56080) );
  CLKNAND2HSV0 U58687 ( .A1(n56221), .A2(\pe3/bq[19] ), .ZN(n56079) );
  XOR2HSV0 U58688 ( .A1(n56080), .A2(n56079), .Z(n56084) );
  NAND2HSV0 U58689 ( .A1(\pe3/aot [8]), .A2(\pe3/bq[18] ), .ZN(n56082) );
  NAND2HSV0 U58690 ( .A1(n56911), .A2(n42971), .ZN(n56081) );
  XOR2HSV0 U58691 ( .A1(n56082), .A2(n56081), .Z(n56083) );
  XOR2HSV0 U58692 ( .A1(n56084), .A2(n56083), .Z(n56085) );
  XOR2HSV0 U58693 ( .A1(n56086), .A2(n56085), .Z(n56105) );
  NAND2HSV0 U58694 ( .A1(n42940), .A2(n56189), .ZN(n56089) );
  NAND2HSV0 U58695 ( .A1(n56087), .A2(n56348), .ZN(n56088) );
  XOR2HSV0 U58696 ( .A1(n56089), .A2(n56088), .Z(n56093) );
  NOR2HSV0 U58697 ( .A1(n56295), .A2(n49272), .ZN(n56091) );
  NAND2HSV0 U58698 ( .A1(\pe3/aot [22]), .A2(\pe3/bq[4] ), .ZN(n56090) );
  XOR2HSV0 U58699 ( .A1(n56091), .A2(n56090), .Z(n56092) );
  XNOR2HSV1 U58700 ( .A1(n56093), .A2(n56092), .ZN(n56103) );
  NAND2HSV0 U58701 ( .A1(n56204), .A2(n56915), .ZN(n56096) );
  NAND2HSV0 U58702 ( .A1(n56197), .A2(n56094), .ZN(n56095) );
  XOR2HSV0 U58703 ( .A1(n56096), .A2(n56095), .Z(n56101) );
  NAND2HSV2 U58704 ( .A1(n56520), .A2(n55857), .ZN(n56791) );
  OAI21HSV0 U58705 ( .A1(n56567), .A2(n55755), .B(n56097), .ZN(n56098) );
  OAI21HSV0 U58706 ( .A1(n56791), .A2(n56099), .B(n56098), .ZN(n56100) );
  XNOR2HSV1 U58707 ( .A1(n56101), .A2(n56100), .ZN(n56102) );
  XNOR2HSV1 U58708 ( .A1(n56103), .A2(n56102), .ZN(n56104) );
  XNOR2HSV1 U58709 ( .A1(n56105), .A2(n56104), .ZN(n56124) );
  NAND2HSV0 U58710 ( .A1(n55873), .A2(n56106), .ZN(n56108) );
  NAND2HSV0 U58711 ( .A1(n56508), .A2(n56187), .ZN(n56107) );
  XOR2HSV0 U58712 ( .A1(n56108), .A2(n56107), .Z(n56112) );
  NAND2HSV0 U58713 ( .A1(\pe3/aot [14]), .A2(n56688), .ZN(n56110) );
  NAND2HSV0 U58714 ( .A1(n56378), .A2(\pe3/bq[11] ), .ZN(n56109) );
  XOR2HSV0 U58715 ( .A1(n56110), .A2(n56109), .Z(n56111) );
  XOR2HSV0 U58716 ( .A1(n56112), .A2(n56111), .Z(n56122) );
  NAND2HSV0 U58717 ( .A1(n56113), .A2(n56529), .ZN(n56426) );
  NAND2HSV0 U58718 ( .A1(n42728), .A2(n56832), .ZN(n56118) );
  NAND2HSV0 U58719 ( .A1(n56455), .A2(n48499), .ZN(n56117) );
  XOR2HSV0 U58720 ( .A1(n56118), .A2(n56117), .Z(n56119) );
  XOR2HSV0 U58721 ( .A1(n56120), .A2(n56119), .Z(n56121) );
  XOR2HSV0 U58722 ( .A1(n56122), .A2(n56121), .Z(n56123) );
  XNOR2HSV1 U58723 ( .A1(n56124), .A2(n56123), .ZN(n56125) );
  XNOR2HSV1 U58724 ( .A1(n56126), .A2(n56125), .ZN(n56129) );
  NAND2HSV0 U58725 ( .A1(n56127), .A2(n56541), .ZN(n56128) );
  XOR2HSV0 U58726 ( .A1(n56129), .A2(n56128), .Z(n56130) );
  XNOR2HSV1 U58727 ( .A1(n56131), .A2(n56130), .ZN(n56132) );
  XNOR2HSV1 U58728 ( .A1(n56133), .A2(n56132), .ZN(n56134) );
  XNOR2HSV1 U58729 ( .A1(n56135), .A2(n56134), .ZN(n56139) );
  NOR2HSV0 U58730 ( .A1(n43840), .A2(n56821), .ZN(n56138) );
  NAND2HSV0 U58731 ( .A1(n56136), .A2(n56266), .ZN(n56137) );
  XOR3HSV1 U58732 ( .A1(n56139), .A2(n56138), .A3(n56137), .Z(n56142) );
  NOR2HSV1 U58733 ( .A1(n43844), .A2(n56496), .ZN(n56141) );
  CLKNAND2HSV1 U58734 ( .A1(n56242), .A2(\pe3/got [9]), .ZN(n56140) );
  XOR3HSV2 U58735 ( .A1(n56142), .A2(n56141), .A3(n56140), .Z(n56143) );
  XNOR2HSV1 U58736 ( .A1(n56144), .A2(n56143), .ZN(n56146) );
  NAND2HSV0 U58737 ( .A1(n55912), .A2(n56619), .ZN(n56145) );
  XNOR2HSV1 U58738 ( .A1(n56146), .A2(n56145), .ZN(n56147) );
  XNOR2HSV1 U58739 ( .A1(n56148), .A2(n56147), .ZN(n56150) );
  NOR2HSV0 U58740 ( .A1(n56406), .A2(n46406), .ZN(n56149) );
  XNOR2HSV1 U58741 ( .A1(n56150), .A2(n56149), .ZN(n56151) );
  XNOR2HSV1 U58742 ( .A1(n56152), .A2(n56151), .ZN(n56153) );
  XOR2HSV0 U58743 ( .A1(n56154), .A2(n56153), .Z(n56155) );
  XNOR2HSV1 U58744 ( .A1(n56156), .A2(n56155), .ZN(n56157) );
  XNOR2HSV1 U58745 ( .A1(n56158), .A2(n56157), .ZN(n56159) );
  XNOR2HSV1 U58746 ( .A1(n56160), .A2(n56159), .ZN(n56161) );
  XNOR2HSV1 U58747 ( .A1(n56162), .A2(n56161), .ZN(n56163) );
  CLKNAND2HSV1 U58748 ( .A1(n56953), .A2(\pe3/got [22]), .ZN(n56164) );
  XNOR2HSV1 U58749 ( .A1(n56165), .A2(n56164), .ZN(n56166) );
  XNOR2HSV1 U58750 ( .A1(n56167), .A2(n56166), .ZN(n56170) );
  CLKNAND2HSV1 U58751 ( .A1(n59823), .A2(n59617), .ZN(n56168) );
  XOR3HSV2 U58752 ( .A1(n56170), .A2(n56169), .A3(n56168), .Z(\pe3/poht [7])
         );
  CLKNAND2HSV1 U58753 ( .A1(n56339), .A2(n45581), .ZN(n56257) );
  NAND2HSV2 U58754 ( .A1(n25989), .A2(n59965), .ZN(n56255) );
  CLKNAND2HSV1 U58755 ( .A1(n56341), .A2(n56335), .ZN(n56251) );
  INHSV2 U58756 ( .I(n45576), .ZN(n56675) );
  CLKNAND2HSV0 U58757 ( .A1(n56621), .A2(n56675), .ZN(n56249) );
  NAND2HSV0 U58758 ( .A1(n56178), .A2(n56177), .ZN(n56246) );
  INAND2HSV0 U58759 ( .A1(n56906), .B1(n59620), .ZN(n56237) );
  NAND2HSV0 U58760 ( .A1(n56179), .A2(n56541), .ZN(n56235) );
  NAND2HSV0 U58761 ( .A1(n56180), .A2(\pe3/got [1]), .ZN(n56233) );
  NAND2HSV2 U58762 ( .A1(n56373), .A2(n56529), .ZN(n56754) );
  NOR2HSV0 U58763 ( .A1(n56181), .A2(n56754), .ZN(n56184) );
  AOI22HSV0 U58764 ( .A1(n56182), .A2(n56529), .B1(n56641), .B2(n59808), .ZN(
        n56183) );
  NOR2HSV1 U58765 ( .A1(n56184), .A2(n56183), .ZN(n56194) );
  NAND2HSV0 U58766 ( .A1(n42818), .A2(n55857), .ZN(n56186) );
  NAND2HSV0 U58767 ( .A1(\pe3/aot [8]), .A2(n43544), .ZN(n56185) );
  XNOR2HSV1 U58768 ( .A1(n56186), .A2(n56185), .ZN(n56193) );
  NAND2HSV0 U58769 ( .A1(n56188), .A2(n56187), .ZN(n56353) );
  NAND2HSV0 U58770 ( .A1(n56464), .A2(n56189), .ZN(n56191) );
  NAND2HSV0 U58771 ( .A1(n56508), .A2(n56827), .ZN(n56190) );
  XOR2HSV0 U58772 ( .A1(n56191), .A2(n56190), .Z(n56192) );
  XOR4HSV1 U58773 ( .A1(n56194), .A2(n56193), .A3(n56353), .A4(n56192), .Z(
        n56231) );
  NAND2HSV0 U58774 ( .A1(n55967), .A2(\pe3/bq[18] ), .ZN(n56196) );
  NAND2HSV0 U58775 ( .A1(n56740), .A2(n48499), .ZN(n56195) );
  XOR2HSV0 U58776 ( .A1(n56196), .A2(n56195), .Z(n56201) );
  NAND2HSV0 U58777 ( .A1(\pe3/aot [13]), .A2(\pe3/bq[11] ), .ZN(n56199) );
  NAND2HSV0 U58778 ( .A1(n56197), .A2(n45534), .ZN(n56198) );
  XOR2HSV0 U58779 ( .A1(n56199), .A2(n56198), .Z(n56200) );
  XOR2HSV0 U58780 ( .A1(n56201), .A2(n56200), .Z(n56210) );
  NAND2HSV0 U58781 ( .A1(n59344), .A2(\pe3/bq[7] ), .ZN(n56203) );
  NAND2HSV0 U58782 ( .A1(n56455), .A2(n56688), .ZN(n56202) );
  XOR2HSV0 U58783 ( .A1(n56203), .A2(n56202), .Z(n56208) );
  NAND2HSV0 U58784 ( .A1(n56378), .A2(n56785), .ZN(n56206) );
  NAND2HSV0 U58785 ( .A1(n56204), .A2(\pe3/bq[4] ), .ZN(n56205) );
  XOR2HSV0 U58786 ( .A1(n56206), .A2(n56205), .Z(n56207) );
  XOR2HSV0 U58787 ( .A1(n56208), .A2(n56207), .Z(n56209) );
  XOR2HSV0 U58788 ( .A1(n56210), .A2(n56209), .Z(n56230) );
  NAND2HSV0 U58789 ( .A1(\pe3/aot [4]), .A2(n42971), .ZN(n56212) );
  NAND2HSV0 U58790 ( .A1(n56439), .A2(\pe3/bq[19] ), .ZN(n56211) );
  XOR2HSV0 U58791 ( .A1(n56212), .A2(n56211), .Z(n56217) );
  NAND2HSV0 U58792 ( .A1(n59511), .A2(n56213), .ZN(n56215) );
  NAND2HSV0 U58793 ( .A1(\pe3/aot [22]), .A2(n56348), .ZN(n56214) );
  XOR2HSV0 U58794 ( .A1(n56215), .A2(n56214), .Z(n56216) );
  XOR2HSV0 U58795 ( .A1(n56217), .A2(n56216), .Z(n56228) );
  NAND2HSV0 U58796 ( .A1(n53250), .A2(n56218), .ZN(n56220) );
  NAND2HSV0 U58797 ( .A1(n42950), .A2(n56915), .ZN(n56219) );
  XOR2HSV0 U58798 ( .A1(n56220), .A2(n56219), .Z(n56226) );
  CLKNAND2HSV0 U58799 ( .A1(n56221), .A2(n56433), .ZN(n56224) );
  NAND2HSV0 U58800 ( .A1(n59961), .A2(n56222), .ZN(n56223) );
  XOR2HSV0 U58801 ( .A1(n56224), .A2(n56223), .Z(n56225) );
  XOR2HSV0 U58802 ( .A1(n56226), .A2(n56225), .Z(n56227) );
  XOR2HSV0 U58803 ( .A1(n56228), .A2(n56227), .Z(n56229) );
  XOR3HSV2 U58804 ( .A1(n56231), .A2(n56230), .A3(n56229), .Z(n56232) );
  XNOR2HSV1 U58805 ( .A1(n56233), .A2(n56232), .ZN(n56234) );
  XNOR2HSV1 U58806 ( .A1(n56235), .A2(n56234), .ZN(n56236) );
  XNOR2HSV1 U58807 ( .A1(n56237), .A2(n56236), .ZN(n56240) );
  NOR2HSV0 U58808 ( .A1(n56391), .A2(n56904), .ZN(n56239) );
  NAND2HSV0 U58809 ( .A1(n56734), .A2(n56422), .ZN(n56238) );
  XOR3HSV1 U58810 ( .A1(n56240), .A2(n56239), .A3(n56238), .Z(n56245) );
  NOR2HSV1 U58811 ( .A1(n56475), .A2(n56821), .ZN(n56244) );
  CLKNAND2HSV1 U58812 ( .A1(n56242), .A2(n56241), .ZN(n56243) );
  XNOR2HSV1 U58813 ( .A1(n56249), .A2(n56248), .ZN(n56250) );
  XNOR2HSV1 U58814 ( .A1(n56251), .A2(n56250), .ZN(n56252) );
  XNOR2HSV1 U58815 ( .A1(n56259), .A2(n56258), .ZN(n56263) );
  NAND2HSV2 U58816 ( .A1(n56490), .A2(n42770), .ZN(n56262) );
  CLKNAND2HSV1 U58817 ( .A1(n56676), .A2(n42673), .ZN(n56261) );
  XOR3HSV2 U58818 ( .A1(n56263), .A2(n56262), .A3(n56261), .Z(\pe3/poht [9])
         );
  CLKAND2HSV2 U58819 ( .A1(n56907), .A2(n56264), .Z(n56332) );
  CLKNAND2HSV1 U58820 ( .A1(n56340), .A2(n56421), .ZN(n56328) );
  CLKNAND2HSV0 U58821 ( .A1(n55946), .A2(n56618), .ZN(n56326) );
  CLKNAND2HSV0 U58822 ( .A1(n59359), .A2(n56342), .ZN(n56324) );
  CLKNAND2HSV0 U58823 ( .A1(n56783), .A2(n56495), .ZN(n56322) );
  CLKNAND2HSV1 U58824 ( .A1(n56561), .A2(n56559), .ZN(n56320) );
  NAND2HSV0 U58825 ( .A1(n59920), .A2(\pe3/got [8]), .ZN(n56318) );
  CLKNAND2HSV0 U58826 ( .A1(n59500), .A2(n56266), .ZN(n56316) );
  NAND2HSV0 U58827 ( .A1(n43754), .A2(n56267), .ZN(n56312) );
  NAND2HSV0 U58828 ( .A1(n55824), .A2(n56781), .ZN(n56308) );
  NAND2HSV0 U58829 ( .A1(\pe3/aot [14]), .A2(n56937), .ZN(n56573) );
  NAND2HSV0 U58830 ( .A1(n59961), .A2(n56433), .ZN(n56268) );
  XOR2HSV0 U58831 ( .A1(n56573), .A2(n56268), .Z(n56286) );
  NOR2HSV2 U58832 ( .A1(n45662), .A2(n56269), .ZN(n56564) );
  AOI22HSV0 U58833 ( .A1(n59808), .A2(n56627), .B1(\pe3/bq[14] ), .B2(n59816), 
        .ZN(n56270) );
  AOI21HSV1 U58834 ( .A1(n56564), .A2(n56271), .B(n56270), .ZN(n56276) );
  AOI22HSV0 U58835 ( .A1(n56508), .A2(n56529), .B1(n53249), .B2(n56272), .ZN(
        n56273) );
  AOI21HSV0 U58836 ( .A1(n56578), .A2(n56274), .B(n56273), .ZN(n56275) );
  XOR2HSV0 U58837 ( .A1(n56276), .A2(n56275), .Z(n56285) );
  NAND2HSV0 U58838 ( .A1(n56695), .A2(n45639), .ZN(n56279) );
  NAND2HSV0 U58839 ( .A1(n56740), .A2(n56785), .ZN(n56278) );
  XOR2HSV0 U58840 ( .A1(n56279), .A2(n56278), .Z(n56283) );
  NAND2HSV0 U58841 ( .A1(n59344), .A2(n56348), .ZN(n56281) );
  NAND2HSV0 U58842 ( .A1(n59511), .A2(\pe3/bq[18] ), .ZN(n56280) );
  XOR2HSV0 U58843 ( .A1(n56281), .A2(n56280), .Z(n56282) );
  XOR2HSV0 U58844 ( .A1(n56283), .A2(n56282), .Z(n56284) );
  XOR3HSV2 U58845 ( .A1(n56286), .A2(n56285), .A3(n56284), .Z(n56303) );
  NAND2HSV0 U58846 ( .A1(n56795), .A2(n56460), .ZN(n56288) );
  NAND2HSV0 U58847 ( .A1(\pe3/aot [8]), .A2(\pe3/bq[11] ), .ZN(n56287) );
  XOR2HSV0 U58848 ( .A1(n56288), .A2(n56287), .Z(n56292) );
  NAND2HSV0 U58849 ( .A1(n56378), .A2(\pe3/bq[4] ), .ZN(n56290) );
  NAND2HSV0 U58850 ( .A1(n56197), .A2(n56454), .ZN(n56289) );
  XOR2HSV0 U58851 ( .A1(n56290), .A2(n56289), .Z(n56291) );
  XOR2HSV0 U58852 ( .A1(n56292), .A2(n56291), .Z(n56301) );
  NAND2HSV0 U58853 ( .A1(n53250), .A2(n43544), .ZN(n56294) );
  NAND2HSV0 U58854 ( .A1(n56788), .A2(n56641), .ZN(n56293) );
  XOR2HSV0 U58855 ( .A1(n56294), .A2(n56293), .Z(n56299) );
  NOR2HSV0 U58856 ( .A1(n56295), .A2(n49275), .ZN(n56297) );
  NAND2HSV0 U58857 ( .A1(\pe3/aot [7]), .A2(n56507), .ZN(n56296) );
  XOR2HSV0 U58858 ( .A1(n56297), .A2(n56296), .Z(n56298) );
  XOR2HSV0 U58859 ( .A1(n56299), .A2(n56298), .Z(n56300) );
  XOR2HSV0 U58860 ( .A1(n56301), .A2(n56300), .Z(n56302) );
  XOR2HSV0 U58861 ( .A1(n56303), .A2(n56302), .Z(n56306) );
  NOR2HSV0 U58862 ( .A1(n56475), .A2(n47431), .ZN(n56305) );
  CLKNAND2HSV0 U58863 ( .A1(n56396), .A2(n56541), .ZN(n56304) );
  XOR3HSV1 U58864 ( .A1(n56306), .A2(n56305), .A3(n56304), .Z(n56307) );
  XNOR2HSV1 U58865 ( .A1(n56308), .A2(n56307), .ZN(n56310) );
  NAND2HSV0 U58866 ( .A1(n59811), .A2(n59356), .ZN(n56309) );
  XNOR2HSV1 U58867 ( .A1(n56310), .A2(n56309), .ZN(n56311) );
  XNOR2HSV1 U58868 ( .A1(n56312), .A2(n56311), .ZN(n56314) );
  NOR2HSV0 U58869 ( .A1(n56406), .A2(n56821), .ZN(n56313) );
  XNOR2HSV1 U58870 ( .A1(n56314), .A2(n56313), .ZN(n56315) );
  XNOR2HSV1 U58871 ( .A1(n56316), .A2(n56315), .ZN(n56317) );
  XNOR2HSV1 U58872 ( .A1(n56318), .A2(n56317), .ZN(n56319) );
  XNOR2HSV1 U58873 ( .A1(n56320), .A2(n56319), .ZN(n56321) );
  XNOR2HSV1 U58874 ( .A1(n56322), .A2(n56321), .ZN(n56323) );
  XNOR2HSV1 U58875 ( .A1(n56324), .A2(n56323), .ZN(n56325) );
  XNOR2HSV1 U58876 ( .A1(n56326), .A2(n56325), .ZN(n56327) );
  XNOR2HSV1 U58877 ( .A1(n56328), .A2(n56327), .ZN(n56329) );
  XNOR2HSV1 U58878 ( .A1(n56330), .A2(n56329), .ZN(n56331) );
  XNOR2HSV1 U58879 ( .A1(n56332), .A2(n56331), .ZN(n56334) );
  XNOR2HSV1 U58880 ( .A1(n56334), .A2(n56333), .ZN(n56338) );
  NAND2HSV2 U58881 ( .A1(n56490), .A2(n56335), .ZN(n56337) );
  XOR3HSV2 U58882 ( .A1(n56338), .A2(n56337), .A3(n56336), .Z(\pe3/poht [14])
         );
  CLKNAND2HSV0 U58883 ( .A1(n56736), .A2(n56618), .ZN(n56416) );
  CLKNAND2HSV1 U58884 ( .A1(n56622), .A2(n56342), .ZN(n56414) );
  NAND2HSV2 U58885 ( .A1(n56497), .A2(n56495), .ZN(n56412) );
  NAND2HSV0 U58886 ( .A1(n56685), .A2(n56559), .ZN(n56410) );
  CLKNAND2HSV1 U58887 ( .A1(n55947), .A2(n56888), .ZN(n56405) );
  CLKNAND2HSV0 U58888 ( .A1(n56178), .A2(n56683), .ZN(n56401) );
  NOR2HSV1 U58889 ( .A1(n56343), .A2(n56632), .ZN(n56345) );
  AOI22HSV0 U58890 ( .A1(n56204), .A2(n56971), .B1(n45645), .B2(n56867), .ZN(
        n56344) );
  NOR2HSV2 U58891 ( .A1(n56345), .A2(n56344), .ZN(n56361) );
  NAND2HSV0 U58892 ( .A1(n56434), .A2(\pe3/bq[18] ), .ZN(n56347) );
  NAND2HSV0 U58893 ( .A1(\pe3/aot [8]), .A2(n56460), .ZN(n56346) );
  XOR2HSV0 U58894 ( .A1(n56347), .A2(n56346), .Z(n56360) );
  NAND2HSV0 U58895 ( .A1(n56349), .A2(n56348), .ZN(n56438) );
  CLKNHSV0 U58896 ( .I(n56438), .ZN(n56352) );
  AOI22HSV0 U58897 ( .A1(n56464), .A2(n56348), .B1(n56349), .B2(n56529), .ZN(
        n56350) );
  AOI21HSV2 U58898 ( .A1(n56352), .A2(n56351), .B(n56350), .ZN(n56358) );
  CLKNAND2HSV0 U58899 ( .A1(n56354), .A2(n56832), .ZN(n56511) );
  NOR2HSV0 U58900 ( .A1(n56353), .A2(n56511), .ZN(n56356) );
  AOI22HSV0 U58901 ( .A1(n56188), .A2(n56832), .B1(n56354), .B2(n56627), .ZN(
        n56355) );
  NOR2HSV1 U58902 ( .A1(n56356), .A2(n56355), .ZN(n56357) );
  XOR2HSV0 U58903 ( .A1(n56358), .A2(n56357), .Z(n56359) );
  XOR3HSV2 U58904 ( .A1(n56361), .A2(n56360), .A3(n56359), .Z(n56369) );
  NAND2HSV0 U58905 ( .A1(n56439), .A2(n56498), .ZN(n56363) );
  NAND2HSV0 U58906 ( .A1(n59960), .A2(\pe3/bq[11] ), .ZN(n56362) );
  XOR2HSV0 U58907 ( .A1(n56363), .A2(n56362), .Z(n56367) );
  NOR2HSV0 U58908 ( .A1(n56784), .A2(n45810), .ZN(n56365) );
  CLKNAND2HSV0 U58909 ( .A1(n56788), .A2(n56433), .ZN(n56364) );
  XOR2HSV0 U58910 ( .A1(n56365), .A2(n56364), .Z(n56366) );
  XOR2HSV0 U58911 ( .A1(n56367), .A2(n56366), .Z(n56368) );
  XNOR2HSV1 U58912 ( .A1(n56369), .A2(n56368), .ZN(n56390) );
  NAND2HSV0 U58913 ( .A1(n59961), .A2(\pe3/bq[19] ), .ZN(n56372) );
  NAND2HSV0 U58914 ( .A1(n56370), .A2(n56785), .ZN(n56371) );
  XOR2HSV0 U58915 ( .A1(n56372), .A2(n56371), .Z(n56377) );
  NAND2HSV0 U58916 ( .A1(n56373), .A2(n45982), .ZN(n56375) );
  NAND2HSV0 U58917 ( .A1(n56795), .A2(n56641), .ZN(n56374) );
  XOR2HSV0 U58918 ( .A1(n56375), .A2(n56374), .Z(n56376) );
  XOR2HSV0 U58919 ( .A1(n56377), .A2(n56376), .Z(n56388) );
  NAND2HSV0 U58920 ( .A1(n56378), .A2(n56835), .ZN(n56381) );
  NAND2HSV0 U58921 ( .A1(\pe3/aot [7]), .A2(n56379), .ZN(n56380) );
  XOR2HSV0 U58922 ( .A1(n56381), .A2(n56380), .Z(n56386) );
  NOR2HSV0 U58923 ( .A1(n56382), .A2(n49272), .ZN(n56384) );
  NAND2HSV0 U58924 ( .A1(n59344), .A2(\pe3/bq[4] ), .ZN(n56383) );
  XOR2HSV0 U58925 ( .A1(n56384), .A2(n56383), .Z(n56385) );
  XOR2HSV0 U58926 ( .A1(n56386), .A2(n56385), .Z(n56387) );
  XOR2HSV0 U58927 ( .A1(n56388), .A2(n56387), .Z(n56389) );
  XNOR2HSV1 U58928 ( .A1(n56390), .A2(n56389), .ZN(n56395) );
  NOR2HSV0 U58929 ( .A1(n56391), .A2(n47431), .ZN(n56394) );
  NAND2HSV0 U58930 ( .A1(n56392), .A2(n56541), .ZN(n56393) );
  XOR3HSV1 U58931 ( .A1(n56395), .A2(n56394), .A3(n56393), .Z(n56399) );
  NOR2HSV0 U58932 ( .A1(n56475), .A2(n56906), .ZN(n56398) );
  NAND2HSV0 U58933 ( .A1(n56396), .A2(n56781), .ZN(n56397) );
  XOR3HSV2 U58934 ( .A1(n56399), .A2(n56398), .A3(n56397), .Z(n56400) );
  XNOR2HSV1 U58935 ( .A1(n56401), .A2(n56400), .ZN(n56403) );
  NAND2HSV0 U58936 ( .A1(n59811), .A2(n56734), .ZN(n56402) );
  XNOR2HSV1 U58937 ( .A1(n56403), .A2(n56402), .ZN(n56404) );
  XNOR2HSV1 U58938 ( .A1(n56405), .A2(n56404), .ZN(n56408) );
  NOR2HSV0 U58939 ( .A1(n56406), .A2(n56496), .ZN(n56407) );
  XNOR2HSV1 U58940 ( .A1(n56408), .A2(n56407), .ZN(n56409) );
  XNOR2HSV1 U58941 ( .A1(n56410), .A2(n56409), .ZN(n56411) );
  XNOR2HSV1 U58942 ( .A1(n56412), .A2(n56411), .ZN(n56413) );
  XNOR2HSV1 U58943 ( .A1(n56414), .A2(n56413), .ZN(n56415) );
  CLKNAND2HSV1 U58944 ( .A1(n48480), .A2(n56675), .ZN(n56486) );
  NAND2HSV2 U58945 ( .A1(n25989), .A2(n56419), .ZN(n56484) );
  CLKNAND2HSV1 U58946 ( .A1(n48481), .A2(n56493), .ZN(n56482) );
  CLKNAND2HSV0 U58947 ( .A1(n59527), .A2(n56421), .ZN(n56480) );
  NAND2HSV0 U58948 ( .A1(n59359), .A2(n56618), .ZN(n56478) );
  NAND2HSV0 U58949 ( .A1(n56422), .A2(\pe3/got [1]), .ZN(n56474) );
  NAND2HSV0 U58950 ( .A1(n56423), .A2(\pe3/bq[11] ), .ZN(n56655) );
  CLKNHSV0 U58951 ( .I(n56754), .ZN(n56425) );
  AOI22HSV2 U58952 ( .A1(n56426), .A2(n56655), .B1(n56425), .B2(n56424), .ZN(
        n56432) );
  NAND2HSV0 U58953 ( .A1(\pe3/aot [8]), .A2(n56937), .ZN(n56702) );
  NOR2HSV0 U58954 ( .A1(n56427), .A2(n56702), .ZN(n56430) );
  AOI22HSV0 U58955 ( .A1(n56651), .A2(n56428), .B1(n45982), .B2(\pe3/aot [8]), 
        .ZN(n56429) );
  NOR2HSV2 U58956 ( .A1(n56430), .A2(n56429), .ZN(n56431) );
  XNOR2HSV1 U58957 ( .A1(n56432), .A2(n56431), .ZN(n56443) );
  NAND2HSV0 U58958 ( .A1(n56434), .A2(n56433), .ZN(n56437) );
  CLKNAND2HSV1 U58959 ( .A1(n56434), .A2(n56969), .ZN(n56954) );
  NOR2HSV0 U58960 ( .A1(n56435), .A2(n56954), .ZN(n56436) );
  AOI21HSV2 U58961 ( .A1(n56438), .A2(n56437), .B(n56436), .ZN(n56441) );
  NAND2HSV0 U58962 ( .A1(n56439), .A2(n56641), .ZN(n56440) );
  XNOR2HSV1 U58963 ( .A1(n56441), .A2(n56440), .ZN(n56442) );
  XNOR2HSV1 U58964 ( .A1(n56443), .A2(n56442), .ZN(n56451) );
  NAND2HSV0 U58965 ( .A1(n45973), .A2(\pe3/bq[14] ), .ZN(n56445) );
  NAND2HSV0 U58966 ( .A1(n45645), .A2(\pe3/bq[4] ), .ZN(n56444) );
  XOR2HSV0 U58967 ( .A1(n56445), .A2(n56444), .Z(n56449) );
  NOR2HSV1 U58968 ( .A1(n47447), .A2(n56269), .ZN(n56447) );
  NAND2HSV0 U58969 ( .A1(n59511), .A2(\pe3/bq[19] ), .ZN(n56446) );
  XOR2HSV0 U58970 ( .A1(n56447), .A2(n56446), .Z(n56448) );
  XOR2HSV0 U58971 ( .A1(n56449), .A2(n56448), .Z(n56450) );
  XOR2HSV0 U58972 ( .A1(n56451), .A2(n56450), .Z(n56472) );
  NAND2HSV0 U58973 ( .A1(n43280), .A2(n56832), .ZN(n56453) );
  NAND2HSV0 U58974 ( .A1(n56188), .A2(n56915), .ZN(n56452) );
  XOR2HSV0 U58975 ( .A1(n56453), .A2(n56452), .Z(n56459) );
  CLKNAND2HSV1 U58976 ( .A1(n56455), .A2(n56454), .ZN(n56457) );
  NAND2HSV0 U58977 ( .A1(n56197), .A2(n56785), .ZN(n56456) );
  XOR2HSV0 U58978 ( .A1(n56457), .A2(n56456), .Z(n56458) );
  XNOR2HSV1 U58979 ( .A1(n56459), .A2(n56458), .ZN(n56470) );
  NAND2HSV0 U58980 ( .A1(\pe3/aot [2]), .A2(\pe3/bq[18] ), .ZN(n56462) );
  NAND2HSV0 U58981 ( .A1(\pe3/aot [7]), .A2(n56460), .ZN(n56461) );
  XOR2HSV0 U58982 ( .A1(n56462), .A2(n56461), .Z(n56468) );
  NAND2HSV2 U58983 ( .A1(n56788), .A2(n56824), .ZN(n56955) );
  NOR2HSV0 U58984 ( .A1(n56463), .A2(n56955), .ZN(n56466) );
  AOI22HSV0 U58985 ( .A1(n56464), .A2(n56824), .B1(n56498), .B2(n56788), .ZN(
        n56465) );
  NOR2HSV2 U58986 ( .A1(n56466), .A2(n56465), .ZN(n56467) );
  XNOR2HSV1 U58987 ( .A1(n56468), .A2(n56467), .ZN(n56469) );
  XNOR2HSV1 U58988 ( .A1(n56470), .A2(n56469), .ZN(n56471) );
  XNOR2HSV1 U58989 ( .A1(n56472), .A2(n56471), .ZN(n56473) );
  NOR2HSV0 U58990 ( .A1(n56475), .A2(n56936), .ZN(n56476) );
  XNOR2HSV1 U58991 ( .A1(n56478), .A2(n56477), .ZN(n56479) );
  XNOR2HSV1 U58992 ( .A1(n56480), .A2(n56479), .ZN(n56481) );
  XNOR2HSV1 U58993 ( .A1(n56482), .A2(n56481), .ZN(n56483) );
  XOR2HSV0 U58994 ( .A1(n56484), .A2(n56483), .Z(n56485) );
  XOR2HSV0 U58995 ( .A1(n56486), .A2(n56485), .Z(n56487) );
  CLKNAND2HSV2 U58996 ( .A1(n56965), .A2(n56489), .ZN(n56492) );
  CLKNAND2HSV1 U58997 ( .A1(n56490), .A2(\pe3/got [18]), .ZN(n56491) );
  CLKNAND2HSV1 U58998 ( .A1(n56952), .A2(n56419), .ZN(n56553) );
  CLKNAND2HSV0 U58999 ( .A1(n56953), .A2(n56493), .ZN(n56551) );
  CLKNAND2HSV1 U59000 ( .A1(n48481), .A2(n56494), .ZN(n56547) );
  CLKNAND2HSV1 U59001 ( .A1(n56621), .A2(n56495), .ZN(n56543) );
  NAND2HSV0 U59002 ( .A1(n59821), .A2(n56823), .ZN(n56540) );
  NAND2HSV0 U59003 ( .A1(n59810), .A2(\pe3/got [1]), .ZN(n56539) );
  NAND2HSV0 U59004 ( .A1(\pe3/aot [8]), .A2(n56627), .ZN(n56500) );
  NAND2HSV0 U59005 ( .A1(\pe3/aot [2]), .A2(n56498), .ZN(n56499) );
  XOR2HSV0 U59006 ( .A1(n56500), .A2(n56499), .Z(n56504) );
  NAND2HSV0 U59007 ( .A1(n56695), .A2(n56835), .ZN(n56502) );
  NAND2HSV0 U59008 ( .A1(n43280), .A2(n56867), .ZN(n56501) );
  XOR2HSV0 U59009 ( .A1(n56502), .A2(n56501), .Z(n56503) );
  XOR2HSV0 U59010 ( .A1(n56504), .A2(n56503), .Z(n56518) );
  CLKNAND2HSV1 U59011 ( .A1(n45973), .A2(n56505), .ZN(n56869) );
  NOR2HSV0 U59012 ( .A1(n56506), .A2(n56869), .ZN(n56510) );
  AOI22HSV0 U59013 ( .A1(n56508), .A2(n56348), .B1(n56507), .B2(n56795), .ZN(
        n56509) );
  NOR2HSV2 U59014 ( .A1(n56510), .A2(n56509), .ZN(n56512) );
  XNOR2HSV1 U59015 ( .A1(n56512), .A2(n56511), .ZN(n56516) );
  NAND2HSV0 U59016 ( .A1(n56740), .A2(n55970), .ZN(n56513) );
  XOR2HSV0 U59017 ( .A1(n56514), .A2(n56513), .Z(n56515) );
  XOR2HSV0 U59018 ( .A1(n56516), .A2(n56515), .Z(n56517) );
  XOR2HSV0 U59019 ( .A1(n56518), .A2(n56517), .Z(n56537) );
  NAND2HSV0 U59020 ( .A1(n59511), .A2(n56519), .ZN(n56522) );
  NAND2HSV0 U59021 ( .A1(n56520), .A2(n53232), .ZN(n56521) );
  XOR2HSV0 U59022 ( .A1(n56522), .A2(n56521), .Z(n56526) );
  CLKNAND2HSV1 U59023 ( .A1(n53250), .A2(n56641), .ZN(n56524) );
  NAND2HSV0 U59024 ( .A1(n56188), .A2(\pe3/bq[4] ), .ZN(n56523) );
  XOR2HSV0 U59025 ( .A1(n56524), .A2(n56523), .Z(n56525) );
  XOR2HSV0 U59026 ( .A1(n56526), .A2(n56525), .Z(n56535) );
  NAND2HSV0 U59027 ( .A1(n56074), .A2(\pe3/bq[14] ), .ZN(n56528) );
  NAND2HSV0 U59028 ( .A1(n59627), .A2(\pe3/bq[11] ), .ZN(n56527) );
  XOR2HSV0 U59029 ( .A1(n56528), .A2(n56527), .Z(n56533) );
  CLKNAND2HSV1 U59030 ( .A1(\pe3/aot [5]), .A2(n56529), .ZN(n56874) );
  OAI21HSV0 U59031 ( .A1(n45662), .A2(n49423), .B(n56650), .ZN(n56530) );
  OAI21HSV0 U59032 ( .A1(n56874), .A2(n56531), .B(n56530), .ZN(n56532) );
  XNOR2HSV1 U59033 ( .A1(n56533), .A2(n56532), .ZN(n56534) );
  XNOR2HSV1 U59034 ( .A1(n56535), .A2(n56534), .ZN(n56536) );
  XNOR2HSV1 U59035 ( .A1(n56537), .A2(n56536), .ZN(n56538) );
  XNOR2HSV1 U59036 ( .A1(n56543), .A2(n56542), .ZN(n56544) );
  XNOR2HSV1 U59037 ( .A1(n56545), .A2(n56544), .ZN(n56546) );
  XNOR2HSV1 U59038 ( .A1(n56547), .A2(n56546), .ZN(n56548) );
  XOR2HSV0 U59039 ( .A1(n56549), .A2(n56548), .Z(n56550) );
  XOR2HSV0 U59040 ( .A1(n56551), .A2(n56550), .Z(n56552) );
  XNOR2HSV1 U59041 ( .A1(n56553), .A2(n56552), .ZN(n56556) );
  INHSV2 U59042 ( .I(n56854), .ZN(n56817) );
  CLKNAND2HSV1 U59043 ( .A1(n59823), .A2(n56675), .ZN(n56554) );
  XOR3HSV2 U59044 ( .A1(n56556), .A2(n56555), .A3(n56554), .Z(\pe3/poht [15])
         );
  CLKNAND2HSV1 U59045 ( .A1(n56905), .A2(n56618), .ZN(n56614) );
  CLKNAND2HSV1 U59046 ( .A1(n48480), .A2(n56557), .ZN(n56612) );
  NAND2HSV2 U59047 ( .A1(n56909), .A2(n56558), .ZN(n56610) );
  CLKNAND2HSV1 U59048 ( .A1(n48481), .A2(n56559), .ZN(n56608) );
  CLKNAND2HSV0 U59049 ( .A1(n55946), .A2(n56855), .ZN(n56606) );
  CLKNAND2HSV1 U59050 ( .A1(n56621), .A2(n56266), .ZN(n56604) );
  CLKNAND2HSV0 U59051 ( .A1(n56736), .A2(n56560), .ZN(n56602) );
  CLKNAND2HSV1 U59052 ( .A1(n56561), .A2(n56623), .ZN(n56600) );
  NAND2HSV0 U59053 ( .A1(n56737), .A2(n56684), .ZN(n56598) );
  CLKNAND2HSV0 U59054 ( .A1(n56562), .A2(n56823), .ZN(n56596) );
  NAND2HSV0 U59055 ( .A1(n55947), .A2(\pe3/got [1]), .ZN(n56592) );
  XOR2HSV0 U59056 ( .A1(n56564), .A2(n56563), .Z(n56590) );
  NAND2HSV2 U59057 ( .A1(\pe3/aot [8]), .A2(\pe3/bq[7] ), .ZN(n56566) );
  NAND2HSV0 U59058 ( .A1(n53250), .A2(n56507), .ZN(n56565) );
  XOR2HSV0 U59059 ( .A1(n56566), .A2(n56565), .Z(n56571) );
  NOR2HSV0 U59060 ( .A1(n56567), .A2(n49258), .ZN(n56569) );
  NAND2HSV0 U59061 ( .A1(\pe3/aot [11]), .A2(\pe3/bq[4] ), .ZN(n56568) );
  XOR2HSV0 U59062 ( .A1(n56569), .A2(n56568), .Z(n56570) );
  XNOR2HSV1 U59063 ( .A1(n56571), .A2(n56570), .ZN(n56589) );
  AOI22HSV0 U59064 ( .A1(n56575), .A2(n56529), .B1(\pe3/aot [13]), .B2(n56348), 
        .ZN(n56576) );
  AOI21HSV0 U59065 ( .A1(n56578), .A2(n56577), .B(n56576), .ZN(n56579) );
  XOR2HSV0 U59066 ( .A1(n56580), .A2(n56579), .Z(n56588) );
  NAND2HSV0 U59067 ( .A1(n45973), .A2(n53232), .ZN(n56582) );
  NAND2HSV0 U59068 ( .A1(n59961), .A2(n56644), .ZN(n56581) );
  XOR2HSV0 U59069 ( .A1(n56582), .A2(n56581), .Z(n56586) );
  NAND2HSV0 U59070 ( .A1(n59511), .A2(n48499), .ZN(n56584) );
  NAND2HSV0 U59071 ( .A1(n56221), .A2(n56454), .ZN(n56583) );
  XOR2HSV0 U59072 ( .A1(n56584), .A2(n56583), .Z(n56585) );
  XOR2HSV0 U59073 ( .A1(n56586), .A2(n56585), .Z(n56587) );
  XOR4HSV1 U59074 ( .A1(n56590), .A2(n56589), .A3(n56588), .A4(n56587), .Z(
        n56591) );
  XNOR2HSV1 U59075 ( .A1(n56592), .A2(n56591), .ZN(n56594) );
  INHSV2 U59076 ( .I(n56936), .ZN(n56862) );
  NAND2HSV0 U59077 ( .A1(n56662), .A2(n56862), .ZN(n56593) );
  XNOR2HSV1 U59078 ( .A1(n56594), .A2(n56593), .ZN(n56595) );
  XNOR2HSV1 U59079 ( .A1(n56596), .A2(n56595), .ZN(n56597) );
  XNOR2HSV1 U59080 ( .A1(n56598), .A2(n56597), .ZN(n56599) );
  XNOR2HSV1 U59081 ( .A1(n56600), .A2(n56599), .ZN(n56601) );
  XNOR2HSV1 U59082 ( .A1(n56602), .A2(n56601), .ZN(n56603) );
  XNOR2HSV1 U59083 ( .A1(n56604), .A2(n56603), .ZN(n56605) );
  XNOR2HSV1 U59084 ( .A1(n56606), .A2(n56605), .ZN(n56607) );
  XNOR2HSV1 U59085 ( .A1(n56608), .A2(n56607), .ZN(n56609) );
  CLKNAND2HSV2 U59086 ( .A1(n56817), .A2(n56493), .ZN(n56616) );
  CLKNAND2HSV1 U59087 ( .A1(n59823), .A2(n43829), .ZN(n56615) );
  XOR3HSV2 U59088 ( .A1(n56617), .A2(n56616), .A3(n56615), .Z(\pe3/poht [18])
         );
  CLKNAND2HSV0 U59089 ( .A1(n56860), .A2(\pe3/got [14]), .ZN(n56674) );
  CLKNAND2HSV1 U59090 ( .A1(n48480), .A2(n56421), .ZN(n56672) );
  CLKNAND2HSV1 U59091 ( .A1(n48481), .A2(n56342), .ZN(n56668) );
  CLKNAND2HSV1 U59092 ( .A1(n56341), .A2(n56619), .ZN(n56666) );
  CLKNAND2HSV1 U59093 ( .A1(n56621), .A2(n56620), .ZN(n56664) );
  NAND2HSV0 U59094 ( .A1(n56197), .A2(n56915), .ZN(n56626) );
  NAND2HSV0 U59095 ( .A1(n53249), .A2(\pe3/bq[4] ), .ZN(n56625) );
  XOR2HSV0 U59096 ( .A1(n56626), .A2(n56625), .Z(n56631) );
  NAND2HSV0 U59097 ( .A1(n56740), .A2(n56832), .ZN(n56629) );
  NAND2HSV0 U59098 ( .A1(n56221), .A2(n56627), .ZN(n56628) );
  XOR2HSV0 U59099 ( .A1(n56629), .A2(n56628), .Z(n56630) );
  XOR2HSV0 U59100 ( .A1(n56631), .A2(n56630), .Z(n56639) );
  XOR2HSV0 U59101 ( .A1(n56633), .A2(n56632), .Z(n56637) );
  NAND2HSV0 U59102 ( .A1(\pe3/aot [8]), .A2(n53232), .ZN(n56634) );
  XOR2HSV0 U59103 ( .A1(n56635), .A2(n56634), .Z(n56636) );
  XOR2HSV0 U59104 ( .A1(n56637), .A2(n56636), .Z(n56638) );
  NAND2HSV0 U59105 ( .A1(n59511), .A2(n56640), .ZN(n56643) );
  NAND2HSV0 U59106 ( .A1(\pe3/aot [2]), .A2(n56641), .ZN(n56642) );
  XOR2HSV0 U59107 ( .A1(n56643), .A2(n56642), .Z(n56648) );
  NAND2HSV0 U59108 ( .A1(n53250), .A2(\pe3/bq[14] ), .ZN(n56646) );
  NAND2HSV0 U59109 ( .A1(n56074), .A2(n56644), .ZN(n56645) );
  XOR2HSV0 U59110 ( .A1(n56646), .A2(n56645), .Z(n56647) );
  XNOR2HSV1 U59111 ( .A1(n56648), .A2(n56647), .ZN(n56661) );
  NOR2HSV0 U59112 ( .A1(n56650), .A2(n56649), .ZN(n56653) );
  AOI22HSV0 U59113 ( .A1(n56188), .A2(n56529), .B1(n56651), .B2(n56892), .ZN(
        n56652) );
  NOR2HSV2 U59114 ( .A1(n56653), .A2(n56652), .ZN(n56659) );
  NOR2HSV1 U59115 ( .A1(n56655), .A2(n56654), .ZN(n56657) );
  AOI22HSV0 U59116 ( .A1(n59808), .A2(n56454), .B1(\pe3/bq[11] ), .B2(n56911), 
        .ZN(n56656) );
  NOR2HSV2 U59117 ( .A1(n56657), .A2(n56656), .ZN(n56658) );
  XOR2HSV0 U59118 ( .A1(n56659), .A2(n56658), .Z(n56660) );
  XNOR2HSV1 U59119 ( .A1(n56664), .A2(n56663), .ZN(n56665) );
  XNOR2HSV1 U59120 ( .A1(n56666), .A2(n56665), .ZN(n56667) );
  XNOR2HSV1 U59121 ( .A1(n56668), .A2(n56667), .ZN(n56669) );
  XOR2HSV0 U59122 ( .A1(n56670), .A2(n56669), .Z(n56671) );
  XOR2HSV0 U59123 ( .A1(n56672), .A2(n56671), .Z(n56673) );
  XNOR2HSV1 U59124 ( .A1(n56674), .A2(n56673), .ZN(n56679) );
  CLKNAND2HSV2 U59125 ( .A1(n56948), .A2(n56675), .ZN(n56678) );
  CLKNAND2HSV1 U59126 ( .A1(n56900), .A2(n56419), .ZN(n56677) );
  XOR3HSV2 U59127 ( .A1(n56679), .A2(n56678), .A3(n56677), .Z(\pe3/poht [16])
         );
  CLKNAND2HSV1 U59128 ( .A1(n56860), .A2(n56619), .ZN(n56730) );
  CLKNAND2HSV1 U59129 ( .A1(n48480), .A2(n56559), .ZN(n56728) );
  CLKNHSV0 U59130 ( .I(n56855), .ZN(n56681) );
  NOR2HSV2 U59131 ( .A1(n56682), .A2(n56681), .ZN(n56726) );
  CLKNAND2HSV1 U59132 ( .A1(n48481), .A2(n56771), .ZN(n56724) );
  CLKNAND2HSV0 U59133 ( .A1(n59527), .A2(n56683), .ZN(n56722) );
  CLKNAND2HSV0 U59134 ( .A1(n59359), .A2(n56822), .ZN(n56720) );
  CLKNAND2HSV0 U59135 ( .A1(n56783), .A2(n56684), .ZN(n56718) );
  CLKNAND2HSV0 U59136 ( .A1(n49253), .A2(n56735), .ZN(n56716) );
  CLKNAND2HSV0 U59137 ( .A1(n59920), .A2(n56782), .ZN(n56714) );
  NAND2HSV0 U59138 ( .A1(n56685), .A2(\pe3/got [1]), .ZN(n56712) );
  NAND2HSV0 U59139 ( .A1(n59808), .A2(\pe3/bq[4] ), .ZN(n56687) );
  NAND2HSV0 U59140 ( .A1(n55873), .A2(n56827), .ZN(n56686) );
  XOR2HSV0 U59141 ( .A1(n56687), .A2(n56686), .Z(n56692) );
  CLKNAND2HSV0 U59142 ( .A1(n59511), .A2(n56688), .ZN(n56690) );
  NAND2HSV0 U59143 ( .A1(n59961), .A2(\pe3/bq[11] ), .ZN(n56689) );
  XOR2HSV0 U59144 ( .A1(n56690), .A2(n56689), .Z(n56691) );
  XOR2HSV0 U59145 ( .A1(n56692), .A2(n56691), .Z(n56701) );
  NAND2HSV0 U59146 ( .A1(n56911), .A2(\pe3/bq[7] ), .ZN(n56694) );
  NAND2HSV0 U59147 ( .A1(n56788), .A2(n56785), .ZN(n56693) );
  XOR2HSV0 U59148 ( .A1(n56694), .A2(n56693), .Z(n56699) );
  CLKNAND2HSV1 U59149 ( .A1(n56695), .A2(\pe3/bq[1] ), .ZN(n56697) );
  NAND2HSV0 U59150 ( .A1(\pe3/aot [11]), .A2(n56892), .ZN(n56696) );
  XOR2HSV0 U59151 ( .A1(n56697), .A2(n56696), .Z(n56698) );
  XOR2HSV0 U59152 ( .A1(n56699), .A2(n56698), .Z(n56700) );
  XOR2HSV0 U59153 ( .A1(n56701), .A2(n56700), .Z(n56710) );
  XOR2HSV0 U59154 ( .A1(n56703), .A2(n56702), .Z(n56708) );
  NOR2HSV0 U59155 ( .A1(n56704), .A2(n56269), .ZN(n56706) );
  NAND2HSV0 U59156 ( .A1(n56221), .A2(n56272), .ZN(n56705) );
  XOR2HSV0 U59157 ( .A1(n56706), .A2(n56705), .Z(n56707) );
  XOR2HSV0 U59158 ( .A1(n56708), .A2(n56707), .Z(n56709) );
  XNOR2HSV1 U59159 ( .A1(n56710), .A2(n56709), .ZN(n56711) );
  XNOR2HSV1 U59160 ( .A1(n56712), .A2(n56711), .ZN(n56713) );
  XNOR2HSV1 U59161 ( .A1(n56714), .A2(n56713), .ZN(n56715) );
  XNOR2HSV1 U59162 ( .A1(n56716), .A2(n56715), .ZN(n56717) );
  XNOR2HSV1 U59163 ( .A1(n56718), .A2(n56717), .ZN(n56719) );
  XNOR2HSV1 U59164 ( .A1(n56720), .A2(n56719), .ZN(n56721) );
  XNOR2HSV1 U59165 ( .A1(n56722), .A2(n56721), .ZN(n56723) );
  XNOR2HSV1 U59166 ( .A1(n56724), .A2(n56723), .ZN(n56725) );
  XNOR2HSV1 U59167 ( .A1(n56730), .A2(n56729), .ZN(n56733) );
  CLKNAND2HSV1 U59168 ( .A1(n56976), .A2(n59967), .ZN(n56731) );
  XOR3HSV2 U59169 ( .A1(n56733), .A2(n56732), .A3(n56731), .Z(\pe3/poht [20])
         );
  CLKNAND2HSV1 U59170 ( .A1(n56935), .A2(n56177), .ZN(n56774) );
  CLKNAND2HSV0 U59171 ( .A1(n55946), .A2(n56734), .ZN(n56768) );
  NAND2HSV0 U59172 ( .A1(n59359), .A2(n56861), .ZN(n56766) );
  CLKNAND2HSV0 U59173 ( .A1(n56736), .A2(n56735), .ZN(n56764) );
  NAND2HSV0 U59174 ( .A1(n56622), .A2(n56782), .ZN(n56762) );
  NAND2HSV0 U59175 ( .A1(n56737), .A2(\pe3/got [1]), .ZN(n56760) );
  NAND2HSV0 U59176 ( .A1(n45973), .A2(n56915), .ZN(n56739) );
  NAND2HSV0 U59177 ( .A1(\pe3/aot [8]), .A2(\pe3/bq[4] ), .ZN(n56738) );
  XOR2HSV0 U59178 ( .A1(n56739), .A2(n56738), .Z(n56744) );
  NAND2HSV0 U59179 ( .A1(n56740), .A2(n56892), .ZN(n56742) );
  NAND2HSV0 U59180 ( .A1(n53250), .A2(n56785), .ZN(n56741) );
  XOR2HSV0 U59181 ( .A1(n56742), .A2(n56741), .Z(n56743) );
  XOR2HSV0 U59182 ( .A1(n56744), .A2(n56743), .Z(n56750) );
  NAND2HSV2 U59183 ( .A1(n56972), .A2(n56627), .ZN(n56746) );
  CLKNAND2HSV0 U59184 ( .A1(n56788), .A2(n56827), .ZN(n56745) );
  XOR2HSV0 U59185 ( .A1(n56746), .A2(n56745), .Z(n56748) );
  XNOR2HSV1 U59186 ( .A1(n56748), .A2(n56747), .ZN(n56749) );
  XNOR2HSV1 U59187 ( .A1(n56750), .A2(n56749), .ZN(n56758) );
  CLKNAND2HSV0 U59188 ( .A1(n59816), .A2(n56832), .ZN(n56752) );
  CLKNAND2HSV1 U59189 ( .A1(n59511), .A2(\pe3/bq[11] ), .ZN(n56751) );
  XOR2HSV0 U59190 ( .A1(n56752), .A2(n56751), .Z(n56756) );
  NAND2HSV0 U59191 ( .A1(n56221), .A2(n56937), .ZN(n56753) );
  XOR2HSV0 U59192 ( .A1(n56754), .A2(n56753), .Z(n56755) );
  XOR2HSV0 U59193 ( .A1(n56756), .A2(n56755), .Z(n56757) );
  XNOR2HSV1 U59194 ( .A1(n56758), .A2(n56757), .ZN(n56759) );
  XNOR2HSV1 U59195 ( .A1(n56760), .A2(n56759), .ZN(n56761) );
  XNOR2HSV1 U59196 ( .A1(n56762), .A2(n56761), .ZN(n56763) );
  XNOR2HSV1 U59197 ( .A1(n56764), .A2(n56763), .ZN(n56765) );
  XNOR2HSV1 U59198 ( .A1(n56766), .A2(n56765), .ZN(n56767) );
  XNOR2HSV1 U59199 ( .A1(n56768), .A2(n56767), .ZN(n56770) );
  CLKNAND2HSV0 U59200 ( .A1(n48481), .A2(n56779), .ZN(n56769) );
  NAND2HSV2 U59201 ( .A1(n26151), .A2(n56771), .ZN(n56773) );
  CLKNAND2HSV0 U59202 ( .A1(n56953), .A2(n56855), .ZN(n56772) );
  CLKNAND2HSV2 U59203 ( .A1(n56817), .A2(n59967), .ZN(n56776) );
  CLKNAND2HSV1 U59204 ( .A1(n56490), .A2(n56619), .ZN(n56775) );
  XOR3HSV2 U59205 ( .A1(n56777), .A2(n56775), .A3(n56776), .Z(\pe3/poht [21])
         );
  CLKNAND2HSV1 U59206 ( .A1(n56905), .A2(n56888), .ZN(n56816) );
  CLKNAND2HSV0 U59207 ( .A1(n56953), .A2(n56779), .ZN(n56814) );
  CLKNAND2HSV0 U59208 ( .A1(n56780), .A2(n56822), .ZN(n56812) );
  INAND2HSV2 U59209 ( .A1(n56910), .B1(n56781), .ZN(n56810) );
  NAND2HSV0 U59210 ( .A1(n59527), .A2(n59356), .ZN(n56808) );
  CLKNAND2HSV0 U59211 ( .A1(n59359), .A2(n56782), .ZN(n56806) );
  CLKNAND2HSV0 U59212 ( .A1(n56783), .A2(\pe3/got [1]), .ZN(n56804) );
  NAND2HSV2 U59213 ( .A1(n59961), .A2(n56827), .ZN(n56787) );
  NAND2HSV0 U59214 ( .A1(n59511), .A2(n56785), .ZN(n56786) );
  XOR2HSV0 U59215 ( .A1(n56787), .A2(n56786), .Z(n56802) );
  CLKNAND2HSV0 U59216 ( .A1(n56788), .A2(n56272), .ZN(n56790) );
  NAND2HSV0 U59217 ( .A1(\pe3/aot [5]), .A2(n56937), .ZN(n56789) );
  XOR2HSV0 U59218 ( .A1(n56790), .A2(n56789), .Z(n56792) );
  XNOR2HSV1 U59219 ( .A1(n56792), .A2(n56791), .ZN(n56801) );
  NAND2HSV0 U59220 ( .A1(n53250), .A2(n56832), .ZN(n56794) );
  NAND2HSV0 U59221 ( .A1(\pe3/aot [8]), .A2(n56892), .ZN(n56793) );
  XOR2HSV0 U59222 ( .A1(n56794), .A2(n56793), .Z(n56799) );
  NAND2HSV0 U59223 ( .A1(n56864), .A2(n56529), .ZN(n56797) );
  NAND2HSV0 U59224 ( .A1(n56795), .A2(\pe3/bq[4] ), .ZN(n56796) );
  XOR2HSV0 U59225 ( .A1(n56797), .A2(n56796), .Z(n56798) );
  XOR2HSV0 U59226 ( .A1(n56799), .A2(n56798), .Z(n56800) );
  XOR3HSV2 U59227 ( .A1(n56802), .A2(n56801), .A3(n56800), .Z(n56803) );
  XNOR2HSV1 U59228 ( .A1(n56804), .A2(n56803), .ZN(n56805) );
  XNOR2HSV1 U59229 ( .A1(n56806), .A2(n56805), .ZN(n56807) );
  XNOR2HSV1 U59230 ( .A1(n56808), .A2(n56807), .ZN(n56809) );
  XNOR2HSV1 U59231 ( .A1(n56810), .A2(n56809), .ZN(n56811) );
  XOR2HSV0 U59232 ( .A1(n56812), .A2(n56811), .Z(n56813) );
  XOR2HSV0 U59233 ( .A1(n56814), .A2(n56813), .Z(n56815) );
  XNOR2HSV1 U59234 ( .A1(n56816), .A2(n56815), .ZN(n56820) );
  CLKNAND2HSV2 U59235 ( .A1(n59441), .A2(n56177), .ZN(n56819) );
  CLKNAND2HSV1 U59236 ( .A1(n56976), .A2(n56855), .ZN(n56818) );
  XOR3HSV2 U59237 ( .A1(n56820), .A2(n56819), .A3(n56818), .Z(\pe3/poht [23])
         );
  CLKNAND2HSV1 U59238 ( .A1(n56860), .A2(n56779), .ZN(n56853) );
  CLKNAND2HSV1 U59239 ( .A1(n48480), .A2(n56822), .ZN(n56851) );
  NAND2HSV2 U59240 ( .A1(n56909), .A2(n56861), .ZN(n56849) );
  INAND2HSV2 U59241 ( .A1(n56910), .B1(n56823), .ZN(n56847) );
  CLKNAND2HSV0 U59242 ( .A1(n59527), .A2(n56908), .ZN(n56845) );
  NAND2HSV0 U59243 ( .A1(n59359), .A2(\pe3/got [1]), .ZN(n56843) );
  CLKNAND2HSV0 U59244 ( .A1(n59816), .A2(\pe3/bq[4] ), .ZN(n56826) );
  NAND2HSV0 U59245 ( .A1(\pe3/aot [8]), .A2(n56824), .ZN(n56825) );
  XOR2HSV0 U59246 ( .A1(n56826), .A2(n56825), .Z(n56831) );
  CLKNAND2HSV0 U59247 ( .A1(n56864), .A2(n56969), .ZN(n56829) );
  NAND2HSV0 U59248 ( .A1(\pe3/aot [1]), .A2(n56827), .ZN(n56828) );
  XOR2HSV0 U59249 ( .A1(n56829), .A2(n56828), .Z(n56830) );
  XOR2HSV0 U59250 ( .A1(n56831), .A2(n56830), .Z(n56841) );
  NAND2HSV2 U59251 ( .A1(n59961), .A2(n56832), .ZN(n56834) );
  NAND2HSV0 U59252 ( .A1(n56788), .A2(n56867), .ZN(n56833) );
  XOR2HSV0 U59253 ( .A1(n56834), .A2(n56833), .Z(n56839) );
  NAND2HSV0 U59254 ( .A1(n53250), .A2(n56835), .ZN(n56836) );
  XOR2HSV0 U59255 ( .A1(n56837), .A2(n56836), .Z(n56838) );
  XOR2HSV0 U59256 ( .A1(n56839), .A2(n56838), .Z(n56840) );
  XOR2HSV0 U59257 ( .A1(n56841), .A2(n56840), .Z(n56842) );
  XNOR2HSV1 U59258 ( .A1(n56843), .A2(n56842), .ZN(n56844) );
  XNOR2HSV1 U59259 ( .A1(n56845), .A2(n56844), .ZN(n56846) );
  XNOR2HSV1 U59260 ( .A1(n56847), .A2(n56846), .ZN(n56848) );
  NAND2HSV2 U59261 ( .A1(n56899), .A2(n56855), .ZN(n56857) );
  CLKNAND2HSV1 U59262 ( .A1(n56900), .A2(n56888), .ZN(n56856) );
  XOR3HSV2 U59263 ( .A1(n56858), .A2(n56857), .A3(n56856), .Z(\pe3/poht [24])
         );
  CLKNAND2HSV1 U59264 ( .A1(n56860), .A2(n56822), .ZN(n56887) );
  CLKNAND2HSV1 U59265 ( .A1(n48480), .A2(n56861), .ZN(n56885) );
  INAND2HSV2 U59266 ( .A1(n56910), .B1(n56862), .ZN(n56881) );
  NAND2HSV2 U59267 ( .A1(n59511), .A2(n56832), .ZN(n56866) );
  NAND2HSV0 U59268 ( .A1(n56864), .A2(n56971), .ZN(n56865) );
  XOR2HSV0 U59269 ( .A1(n56866), .A2(n56865), .Z(n56871) );
  NAND2HSV0 U59270 ( .A1(n53250), .A2(n56867), .ZN(n56868) );
  XOR2HSV0 U59271 ( .A1(n56869), .A2(n56868), .Z(n56870) );
  XOR2HSV0 U59272 ( .A1(n56871), .A2(n56870), .Z(n56877) );
  NOR2HSV2 U59273 ( .A1(n56956), .A2(n49258), .ZN(n56873) );
  CLKNAND2HSV0 U59274 ( .A1(n56788), .A2(\pe3/bq[4] ), .ZN(n56872) );
  XOR2HSV0 U59275 ( .A1(n56873), .A2(n56872), .Z(n56875) );
  XNOR2HSV1 U59276 ( .A1(n56875), .A2(n56874), .ZN(n56876) );
  XNOR2HSV1 U59277 ( .A1(n56877), .A2(n56876), .ZN(n56878) );
  XNOR2HSV1 U59278 ( .A1(n56879), .A2(n56878), .ZN(n56880) );
  XNOR2HSV1 U59279 ( .A1(n56881), .A2(n56880), .ZN(n56882) );
  XNOR2HSV1 U59280 ( .A1(n56887), .A2(n56886), .ZN(n56891) );
  CLKNAND2HSV1 U59281 ( .A1(n59823), .A2(n56560), .ZN(n56889) );
  XOR3HSV2 U59282 ( .A1(n56891), .A2(n56890), .A3(n56889), .Z(\pe3/poht [25])
         );
  CLKNAND2HSV1 U59283 ( .A1(n56905), .A2(\pe3/got [1]), .ZN(n56898) );
  NAND2HSV2 U59284 ( .A1(n59511), .A2(n56529), .ZN(n56894) );
  CLKNAND2HSV1 U59285 ( .A1(n56972), .A2(n56892), .ZN(n56893) );
  XOR2HSV0 U59286 ( .A1(n56894), .A2(n56893), .Z(n56896) );
  NAND2HSV0 U59287 ( .A1(n56434), .A2(n56971), .ZN(n56895) );
  XNOR2HSV1 U59288 ( .A1(n56896), .A2(n56895), .ZN(n56897) );
  XNOR2HSV1 U59289 ( .A1(n56898), .A2(n56897), .ZN(n56903) );
  CLKNAND2HSV2 U59290 ( .A1(n56948), .A2(n59356), .ZN(n56902) );
  CLKNAND2HSV1 U59291 ( .A1(n56900), .A2(n56908), .ZN(n56901) );
  XOR3HSV2 U59292 ( .A1(n56903), .A2(n56902), .A3(n56901), .Z(\pe3/poht [29])
         );
  CLKNAND2HSV1 U59293 ( .A1(n56905), .A2(n56861), .ZN(n56931) );
  CLKNAND2HSV1 U59294 ( .A1(n56907), .A2(n56735), .ZN(n56929) );
  NAND2HSV2 U59295 ( .A1(n56909), .A2(n56908), .ZN(n56927) );
  INAND2HSV2 U59296 ( .A1(n56910), .B1(\pe3/got [1]), .ZN(n56925) );
  CLKNAND2HSV0 U59297 ( .A1(n53250), .A2(\pe3/bq[4] ), .ZN(n56913) );
  CLKNAND2HSV0 U59298 ( .A1(n56911), .A2(n56971), .ZN(n56912) );
  XOR2HSV0 U59299 ( .A1(n56913), .A2(n56912), .Z(n56919) );
  NOR2HSV0 U59300 ( .A1(n56956), .A2(n56914), .ZN(n56917) );
  CLKNAND2HSV0 U59301 ( .A1(\pe3/aot [1]), .A2(n56915), .ZN(n56916) );
  XOR2HSV0 U59302 ( .A1(n56917), .A2(n56916), .Z(n56918) );
  XNOR2HSV1 U59303 ( .A1(n56919), .A2(n56918), .ZN(n56923) );
  NOR2HSV2 U59304 ( .A1(n45662), .A2(n48495), .ZN(n56921) );
  CLKNAND2HSV1 U59305 ( .A1(n59646), .A2(n56529), .ZN(n56920) );
  XOR2HSV0 U59306 ( .A1(n56921), .A2(n56920), .Z(n56922) );
  XNOR2HSV1 U59307 ( .A1(n56923), .A2(n56922), .ZN(n56924) );
  XNOR2HSV1 U59308 ( .A1(n56925), .A2(n56924), .ZN(n56926) );
  NAND2HSV2 U59309 ( .A1(n56490), .A2(n56822), .ZN(n56933) );
  XOR3HSV2 U59310 ( .A1(n56934), .A2(n56933), .A3(n56932), .Z(\pe3/poht [26])
         );
  CLKNAND2HSV1 U59311 ( .A1(n56935), .A2(n56823), .ZN(n56947) );
  CLKNAND2HSV1 U59312 ( .A1(\pe3/aot [4]), .A2(n56892), .ZN(n56939) );
  CLKNAND2HSV0 U59313 ( .A1(n56970), .A2(n56937), .ZN(n56938) );
  XOR2HSV0 U59314 ( .A1(n56939), .A2(n56938), .Z(n56941) );
  XNOR2HSV1 U59315 ( .A1(n56941), .A2(n56940), .ZN(n56945) );
  CLKNAND2HSV1 U59316 ( .A1(n56972), .A2(\pe3/bq[4] ), .ZN(n56943) );
  CLKNAND2HSV0 U59317 ( .A1(n59816), .A2(n56971), .ZN(n56942) );
  XOR2HSV0 U59318 ( .A1(n56943), .A2(n56942), .Z(n56944) );
  XNOR2HSV1 U59319 ( .A1(n56945), .A2(n56944), .ZN(n56946) );
  NAND2HSV2 U59320 ( .A1(n56490), .A2(n56861), .ZN(n56950) );
  CLKNAND2HSV1 U59321 ( .A1(n56948), .A2(n56822), .ZN(n56949) );
  XOR3HSV2 U59322 ( .A1(n56951), .A2(n56950), .A3(n56949), .Z(\pe3/poht [27])
         );
  CLKNAND2HSV1 U59323 ( .A1(n56952), .A2(n56908), .ZN(n56964) );
  CLKNAND2HSV1 U59324 ( .A1(n56907), .A2(n56975), .ZN(n56962) );
  XOR2HSV0 U59325 ( .A1(n56955), .A2(n56954), .Z(n56960) );
  NOR2HSV1 U59326 ( .A1(n56956), .A2(n50722), .ZN(n56958) );
  CLKNAND2HSV0 U59327 ( .A1(n56970), .A2(\pe3/bq[4] ), .ZN(n56957) );
  XOR2HSV0 U59328 ( .A1(n56958), .A2(n56957), .Z(n56959) );
  XOR2HSV0 U59329 ( .A1(n56960), .A2(n56959), .Z(n56961) );
  XOR2HSV0 U59330 ( .A1(n56962), .A2(n56961), .Z(n56963) );
  XNOR2HSV1 U59331 ( .A1(n56964), .A2(n56963), .ZN(n56968) );
  NAND2HSV2 U59332 ( .A1(n56058), .A2(n56861), .ZN(n56967) );
  CLKNAND2HSV1 U59333 ( .A1(n59823), .A2(n56823), .ZN(n56966) );
  XOR3HSV2 U59334 ( .A1(n56968), .A2(n56967), .A3(n56966), .Z(\pe3/poht [28])
         );
  NAND2HSV2 U59335 ( .A1(n56970), .A2(n56969), .ZN(n56974) );
  NAND2HSV0 U59336 ( .A1(n56972), .A2(n56971), .ZN(n56973) );
  XOR2HSV0 U59337 ( .A1(n56974), .A2(n56973), .Z(n56979) );
  CLKNAND2HSV1 U59338 ( .A1(n56976), .A2(n56975), .ZN(n56977) );
  XOR3HSV2 U59339 ( .A1(n56979), .A2(n56978), .A3(n56977), .Z(\pe3/poht [30])
         );
  CLKNAND2HSV1 U59340 ( .A1(n58217), .A2(n57574), .ZN(n57079) );
  CLKNAND2HSV1 U59341 ( .A1(n58193), .A2(n59369), .ZN(n57077) );
  CLKNAND2HSV1 U59342 ( .A1(n58112), .A2(n34042), .ZN(n57068) );
  NAND2HSV0 U59343 ( .A1(n57675), .A2(n50189), .ZN(n57058) );
  NAND2HSV0 U59344 ( .A1(n57324), .A2(n57646), .ZN(n57056) );
  NAND2HSV0 U59345 ( .A1(n57209), .A2(n57180), .ZN(n57053) );
  NAND2HSV0 U59346 ( .A1(n57458), .A2(\pe4/got [7]), .ZN(n57049) );
  NAND2HSV0 U59347 ( .A1(n57140), .A2(\pe4/bq[11] ), .ZN(n56981) );
  NAND2HSV0 U59348 ( .A1(n33947), .A2(n58156), .ZN(n56980) );
  XOR2HSV0 U59349 ( .A1(n56981), .A2(n56980), .Z(n56985) );
  NAND2HSV0 U59350 ( .A1(n59632), .A2(n57476), .ZN(n56983) );
  NAND2HSV0 U59351 ( .A1(n57506), .A2(n33711), .ZN(n56982) );
  XOR2HSV0 U59352 ( .A1(n56983), .A2(n56982), .Z(n56984) );
  XOR2HSV0 U59353 ( .A1(n56985), .A2(n56984), .Z(n56993) );
  NAND2HSV0 U59354 ( .A1(n57210), .A2(\pe4/bq[2] ), .ZN(n56987) );
  NAND2HSV0 U59355 ( .A1(n59831), .A2(n57691), .ZN(n56986) );
  XOR2HSV0 U59356 ( .A1(n56987), .A2(n56986), .Z(n56991) );
  NAND2HSV0 U59357 ( .A1(n57138), .A2(n57911), .ZN(n56989) );
  NAND2HSV0 U59358 ( .A1(n59954), .A2(\pe4/bq[27] ), .ZN(n56988) );
  XOR2HSV0 U59359 ( .A1(n56989), .A2(n56988), .Z(n56990) );
  XOR2HSV0 U59360 ( .A1(n56991), .A2(n56990), .Z(n56992) );
  XOR2HSV0 U59361 ( .A1(n56993), .A2(n56992), .Z(n57009) );
  NAND2HSV0 U59362 ( .A1(n33965), .A2(\pe4/bq[8] ), .ZN(n56995) );
  NAND2HSV0 U59363 ( .A1(\pe4/aot [23]), .A2(n57684), .ZN(n56994) );
  XOR2HSV0 U59364 ( .A1(n56995), .A2(n56994), .Z(n56999) );
  NAND2HSV0 U59365 ( .A1(n34743), .A2(\pe4/bq[10] ), .ZN(n56997) );
  NAND2HSV0 U59366 ( .A1(\pe4/aot [2]), .A2(\pe4/bq[28] ), .ZN(n56996) );
  XOR2HSV0 U59367 ( .A1(n56997), .A2(n56996), .Z(n56998) );
  XOR2HSV0 U59368 ( .A1(n56999), .A2(n56998), .Z(n57007) );
  NAND2HSV0 U59369 ( .A1(\pe4/aot [1]), .A2(n33533), .ZN(n57001) );
  NAND2HSV0 U59370 ( .A1(n47718), .A2(n57785), .ZN(n57000) );
  XOR2HSV0 U59371 ( .A1(n57001), .A2(n57000), .Z(n57005) );
  NOR2HSV0 U59372 ( .A1(n44338), .A2(n47809), .ZN(n57003) );
  NAND2HSV0 U59373 ( .A1(n59951), .A2(n58113), .ZN(n57002) );
  XOR2HSV0 U59374 ( .A1(n57003), .A2(n57002), .Z(n57004) );
  XOR2HSV0 U59375 ( .A1(n57005), .A2(n57004), .Z(n57006) );
  XOR2HSV0 U59376 ( .A1(n57007), .A2(n57006), .Z(n57008) );
  XOR2HSV0 U59377 ( .A1(n57009), .A2(n57008), .Z(n57037) );
  NOR2HSV0 U59378 ( .A1(n33250), .A2(n57010), .ZN(n57224) );
  NOR2HSV0 U59379 ( .A1(n57011), .A2(n33350), .ZN(n57013) );
  NAND2HSV2 U59380 ( .A1(n57230), .A2(n58196), .ZN(n58267) );
  OAI22HSV0 U59381 ( .A1(n57224), .A2(n57013), .B1(n57012), .B2(n58267), .ZN(
        n57018) );
  NOR2HSV0 U59382 ( .A1(n35175), .A2(n47818), .ZN(n57245) );
  AOI22HSV0 U59383 ( .A1(n57014), .A2(n58127), .B1(n59953), .B2(n57348), .ZN(
        n57015) );
  AOI21HSV0 U59384 ( .A1(n57016), .A2(n57245), .B(n57015), .ZN(n57017) );
  XOR2HSV0 U59385 ( .A1(n57018), .A2(n57017), .Z(n57035) );
  NAND2HSV0 U59386 ( .A1(n57338), .A2(n33712), .ZN(n57020) );
  NAND2HSV0 U59387 ( .A1(\pe4/aot [11]), .A2(n57929), .ZN(n57019) );
  XOR2HSV0 U59388 ( .A1(n57020), .A2(n57019), .Z(n57024) );
  NOR2HSV0 U59389 ( .A1(n34470), .A2(n48024), .ZN(n57022) );
  NAND2HSV0 U59390 ( .A1(n59343), .A2(n57089), .ZN(n57021) );
  XOR2HSV0 U59391 ( .A1(n57022), .A2(n57021), .Z(n57023) );
  XOR2HSV0 U59392 ( .A1(n57024), .A2(n57023), .Z(n57034) );
  NAND2HSV0 U59393 ( .A1(n57504), .A2(n34254), .ZN(n57125) );
  NOR2HSV0 U59394 ( .A1(n57025), .A2(n57841), .ZN(n57220) );
  NOR2HSV0 U59395 ( .A1(n57026), .A2(n48032), .ZN(n57029) );
  OAI22HSV0 U59396 ( .A1(n57220), .A2(n57029), .B1(n57028), .B2(n57027), .ZN(
        n57032) );
  NOR2HSV0 U59397 ( .A1(n57030), .A2(n57387), .ZN(n57839) );
  NAND2HSV0 U59398 ( .A1(n57727), .A2(n57851), .ZN(n57494) );
  XOR2HSV0 U59399 ( .A1(n57839), .A2(n57494), .Z(n57031) );
  XOR3HSV2 U59400 ( .A1(n57125), .A2(n57032), .A3(n57031), .Z(n57033) );
  XOR3HSV2 U59401 ( .A1(n57035), .A2(n57034), .A3(n57033), .Z(n57036) );
  XNOR2HSV1 U59402 ( .A1(n57037), .A2(n57036), .ZN(n57039) );
  NAND2HSV0 U59403 ( .A1(n59501), .A2(n58282), .ZN(n57038) );
  XNOR2HSV1 U59404 ( .A1(n57039), .A2(n57038), .ZN(n57042) );
  NAND2HSV0 U59405 ( .A1(n59524), .A2(n58314), .ZN(n57041) );
  NAND2HSV0 U59406 ( .A1(n29738), .A2(n57584), .ZN(n57040) );
  XOR3HSV2 U59407 ( .A1(n57042), .A2(n57041), .A3(n57040), .Z(n57045) );
  NAND2HSV0 U59408 ( .A1(n59667), .A2(n59832), .ZN(n57044) );
  NAND2HSV0 U59409 ( .A1(n57405), .A2(n57677), .ZN(n57043) );
  XOR3HSV2 U59410 ( .A1(n57045), .A2(n57044), .A3(n57043), .Z(n57047) );
  NAND2HSV0 U59411 ( .A1(n33608), .A2(n58184), .ZN(n57046) );
  XOR2HSV0 U59412 ( .A1(n57047), .A2(n57046), .Z(n57048) );
  XNOR2HSV1 U59413 ( .A1(n57049), .A2(n57048), .ZN(n57051) );
  NAND2HSV0 U59414 ( .A1(n57183), .A2(n57177), .ZN(n57050) );
  XNOR2HSV1 U59415 ( .A1(n57051), .A2(n57050), .ZN(n57052) );
  XNOR2HSV1 U59416 ( .A1(n57053), .A2(n57052), .ZN(n57055) );
  NAND2HSV0 U59417 ( .A1(n59845), .A2(n58153), .ZN(n57054) );
  XOR3HSV2 U59418 ( .A1(n57056), .A2(n57055), .A3(n57054), .Z(n57057) );
  XNOR2HSV1 U59419 ( .A1(n57058), .A2(n57057), .ZN(n57060) );
  NAND2HSV0 U59420 ( .A1(n59932), .A2(n57820), .ZN(n57059) );
  XNOR2HSV1 U59421 ( .A1(n57060), .A2(n57059), .ZN(n57063) );
  NAND2HSV0 U59422 ( .A1(n34409), .A2(n57424), .ZN(n57062) );
  NAND2HSV0 U59423 ( .A1(n57817), .A2(n59664), .ZN(n57061) );
  XOR3HSV2 U59424 ( .A1(n57063), .A2(n57062), .A3(n57061), .Z(n57066) );
  CLKNAND2HSV1 U59425 ( .A1(n35577), .A2(n57753), .ZN(n57065) );
  CLKNAND2HSV0 U59426 ( .A1(n57554), .A2(n57189), .ZN(n57064) );
  XOR3HSV2 U59427 ( .A1(n57066), .A2(n57065), .A3(n57064), .Z(n57067) );
  XNOR2HSV1 U59428 ( .A1(n57068), .A2(n57067), .ZN(n57071) );
  CLKNAND2HSV0 U59429 ( .A1(n47841), .A2(n59386), .ZN(n57070) );
  NAND2HSV0 U59430 ( .A1(n57560), .A2(n35321), .ZN(n57069) );
  XOR3HSV2 U59431 ( .A1(n57071), .A2(n57070), .A3(n57069), .Z(n57073) );
  NAND2HSV0 U59432 ( .A1(n57889), .A2(n57760), .ZN(n57072) );
  XNOR2HSV1 U59433 ( .A1(n57073), .A2(n57072), .ZN(n57075) );
  NAND2HSV0 U59434 ( .A1(n57310), .A2(n59601), .ZN(n57074) );
  XNOR2HSV1 U59435 ( .A1(n57075), .A2(n57074), .ZN(n57076) );
  XNOR2HSV1 U59436 ( .A1(n57077), .A2(n57076), .ZN(n57078) );
  XOR2HSV0 U59437 ( .A1(n57079), .A2(n57078), .Z(n57081) );
  CLKNAND2HSV0 U59438 ( .A1(n59348), .A2(\pe4/got [25]), .ZN(n57080) );
  XNOR2HSV1 U59439 ( .A1(n57081), .A2(n57080), .ZN(n57083) );
  INAND2HSV0 U59440 ( .A1(n35587), .B1(n26692), .ZN(n57082) );
  XNOR2HSV1 U59441 ( .A1(n57083), .A2(n57082), .ZN(n57084) );
  INHSV2 U59442 ( .I(n26413), .ZN(n57900) );
  NAND2HSV2 U59443 ( .A1(n57900), .A2(n59956), .ZN(n57086) );
  XOR3HSV2 U59444 ( .A1(n57088), .A2(n57087), .A3(n57086), .Z(\pe4/poht [3])
         );
  NAND2HSV2 U59445 ( .A1(n50318), .A2(n35445), .ZN(n57203) );
  NAND2HSV0 U59446 ( .A1(n59837), .A2(n34020), .ZN(n57194) );
  NAND2HSV0 U59447 ( .A1(n59667), .A2(n58036), .ZN(n57176) );
  NAND2HSV0 U59448 ( .A1(n59524), .A2(n57677), .ZN(n57172) );
  NAND2HSV0 U59449 ( .A1(\pe4/aot [15]), .A2(n57089), .ZN(n57091) );
  NAND2HSV0 U59450 ( .A1(n57506), .A2(n57337), .ZN(n57090) );
  XOR2HSV0 U59451 ( .A1(n57091), .A2(n57090), .Z(n57095) );
  NAND2HSV0 U59452 ( .A1(n59632), .A2(n57460), .ZN(n57093) );
  NAND2HSV0 U59453 ( .A1(n33965), .A2(\pe4/bq[11] ), .ZN(n57092) );
  XOR2HSV0 U59454 ( .A1(n57093), .A2(n57092), .Z(n57094) );
  XOR2HSV0 U59455 ( .A1(n57095), .A2(n57094), .Z(n57104) );
  NAND2HSV0 U59456 ( .A1(n33716), .A2(n58116), .ZN(n57097) );
  NAND2HSV0 U59457 ( .A1(n57338), .A2(n33427), .ZN(n57096) );
  XOR2HSV0 U59458 ( .A1(n57097), .A2(n57096), .Z(n57102) );
  NAND2HSV0 U59459 ( .A1(n57692), .A2(n57098), .ZN(n57100) );
  NAND2HSV0 U59460 ( .A1(n57510), .A2(n57851), .ZN(n57099) );
  XOR2HSV0 U59461 ( .A1(n57100), .A2(n57099), .Z(n57101) );
  XOR2HSV0 U59462 ( .A1(n57102), .A2(n57101), .Z(n57103) );
  XOR2HSV0 U59463 ( .A1(n57104), .A2(n57103), .Z(n57122) );
  NAND2HSV0 U59464 ( .A1(n57106), .A2(n57911), .ZN(n57347) );
  NOR2HSV0 U59465 ( .A1(n57105), .A2(n57347), .ZN(n57108) );
  AOI22HSV0 U59466 ( .A1(n33727), .A2(n57241), .B1(n57106), .B2(n58301), .ZN(
        n57107) );
  NOR2HSV1 U59467 ( .A1(n57108), .A2(n57107), .ZN(n57120) );
  NAND2HSV0 U59468 ( .A1(\pe4/pq ), .A2(n34054), .ZN(n57110) );
  NAND2HSV0 U59469 ( .A1(\pe4/aot [14]), .A2(n57368), .ZN(n57109) );
  XOR2HSV0 U59470 ( .A1(n57110), .A2(n57109), .Z(n57119) );
  AOI22HSV0 U59471 ( .A1(n57114), .A2(n57113), .B1(n57112), .B2(n57111), .ZN(
        n57118) );
  NOR2HSV0 U59472 ( .A1(n44338), .A2(n48023), .ZN(n57116) );
  NAND2HSV0 U59473 ( .A1(n33867), .A2(n57348), .ZN(n57115) );
  XOR2HSV0 U59474 ( .A1(n57116), .A2(n57115), .Z(n57117) );
  XOR4HSV1 U59475 ( .A1(n57120), .A2(n57119), .A3(n57118), .A4(n57117), .Z(
        n57121) );
  XNOR2HSV1 U59476 ( .A1(n57122), .A2(n57121), .ZN(n57170) );
  NAND2HSV0 U59477 ( .A1(n57251), .A2(n57584), .ZN(n57148) );
  NOR2HSV0 U59478 ( .A1(n57509), .A2(n50114), .ZN(n57329) );
  NOR2HSV0 U59479 ( .A1(n57026), .A2(n48028), .ZN(n57124) );
  NAND2HSV0 U59480 ( .A1(n59838), .A2(n57684), .ZN(n57497) );
  OAI22HSV0 U59481 ( .A1(n57329), .A2(n57124), .B1(n57123), .B2(n57497), .ZN(
        n57130) );
  NOR2HSV0 U59482 ( .A1(n57126), .A2(n57125), .ZN(n57128) );
  AOI22HSV0 U59483 ( .A1(n59343), .A2(n57505), .B1(n33712), .B2(\pe4/aot [9]), 
        .ZN(n57127) );
  NOR2HSV2 U59484 ( .A1(n57128), .A2(n57127), .ZN(n57129) );
  XNOR2HSV1 U59485 ( .A1(n57130), .A2(n57129), .ZN(n57133) );
  NAND2HSV0 U59486 ( .A1(n59523), .A2(\pe4/bq[2] ), .ZN(n57240) );
  XOR2HSV0 U59487 ( .A1(n57131), .A2(n57240), .Z(n57132) );
  XNOR2HSV1 U59488 ( .A1(n57133), .A2(n57132), .ZN(n57146) );
  NAND2HSV0 U59489 ( .A1(\pe4/aot [3]), .A2(n57134), .ZN(n57137) );
  NAND2HSV0 U59490 ( .A1(n57727), .A2(n57135), .ZN(n57136) );
  XOR2HSV0 U59491 ( .A1(n57137), .A2(n57136), .Z(n57144) );
  NAND2HSV0 U59492 ( .A1(n57138), .A2(n58156), .ZN(n57142) );
  NAND2HSV0 U59493 ( .A1(n57140), .A2(n57139), .ZN(n57141) );
  XOR2HSV0 U59494 ( .A1(n57142), .A2(n57141), .Z(n57143) );
  XOR2HSV0 U59495 ( .A1(n57144), .A2(n57143), .Z(n57145) );
  XOR2HSV0 U59496 ( .A1(n57146), .A2(n57145), .Z(n57147) );
  XOR2HSV0 U59497 ( .A1(n57148), .A2(n57147), .Z(n57169) );
  NAND2HSV0 U59498 ( .A1(n59951), .A2(n57986), .ZN(n57150) );
  NAND2HSV0 U59499 ( .A1(n47718), .A2(\pe4/bq[23] ), .ZN(n57149) );
  XOR2HSV0 U59500 ( .A1(n57150), .A2(n57149), .Z(n57154) );
  NAND2HSV0 U59501 ( .A1(\pe4/aot [11]), .A2(n34044), .ZN(n57152) );
  NAND2HSV0 U59502 ( .A1(n57234), .A2(n57926), .ZN(n57151) );
  XOR2HSV0 U59503 ( .A1(n57152), .A2(n57151), .Z(n57153) );
  XOR2HSV0 U59504 ( .A1(n57154), .A2(n57153), .Z(n57163) );
  NAND2HSV0 U59505 ( .A1(n59831), .A2(\pe4/bq[28] ), .ZN(n57156) );
  NAND2HSV0 U59506 ( .A1(n57230), .A2(n57254), .ZN(n57155) );
  XOR2HSV0 U59507 ( .A1(n57156), .A2(n57155), .Z(n57161) );
  NAND2HSV0 U59508 ( .A1(n59958), .A2(n57157), .ZN(n57159) );
  NAND2HSV0 U59509 ( .A1(\pe4/aot [2]), .A2(n33103), .ZN(n57158) );
  XOR2HSV0 U59510 ( .A1(n57159), .A2(n57158), .Z(n57160) );
  XOR2HSV0 U59511 ( .A1(n57161), .A2(n57160), .Z(n57162) );
  XOR2HSV0 U59512 ( .A1(n57163), .A2(n57162), .Z(n57165) );
  NAND2HSV0 U59513 ( .A1(n34127), .A2(n58314), .ZN(n57164) );
  XNOR2HSV1 U59514 ( .A1(n57165), .A2(n57164), .ZN(n57168) );
  NAND2HSV0 U59515 ( .A1(n57166), .A2(n59832), .ZN(n57167) );
  XOR4HSV1 U59516 ( .A1(n57170), .A2(n57169), .A3(n57168), .A4(n57167), .Z(
        n57171) );
  XNOR2HSV1 U59517 ( .A1(n57172), .A2(n57171), .ZN(n57174) );
  NAND2HSV0 U59518 ( .A1(n34396), .A2(n58184), .ZN(n57173) );
  XNOR2HSV1 U59519 ( .A1(n57174), .A2(n57173), .ZN(n57175) );
  XNOR2HSV1 U59520 ( .A1(n57176), .A2(n57175), .ZN(n57179) );
  NAND2HSV0 U59521 ( .A1(n57405), .A2(n57177), .ZN(n57178) );
  XNOR2HSV1 U59522 ( .A1(n57179), .A2(n57178), .ZN(n57182) );
  NAND2HSV0 U59523 ( .A1(n35401), .A2(n57180), .ZN(n57181) );
  XOR2HSV0 U59524 ( .A1(n57182), .A2(n57181), .Z(n57186) );
  NAND2HSV0 U59525 ( .A1(n57458), .A2(n57646), .ZN(n57185) );
  NAND2HSV0 U59526 ( .A1(n57183), .A2(n58153), .ZN(n57184) );
  XOR3HSV1 U59527 ( .A1(n57186), .A2(n57185), .A3(n57184), .Z(n57187) );
  CLKNAND2HSV0 U59528 ( .A1(n35033), .A2(n57190), .ZN(n57191) );
  XNOR2HSV1 U59529 ( .A1(n57192), .A2(n57191), .ZN(n57193) );
  XNOR2HSV1 U59530 ( .A1(n57194), .A2(n57193), .ZN(n57198) );
  CLKNAND2HSV1 U59531 ( .A1(n58217), .A2(n59350), .ZN(n57197) );
  CLKNAND2HSV0 U59532 ( .A1(n57970), .A2(n57195), .ZN(n57196) );
  XOR3HSV2 U59533 ( .A1(n57198), .A2(n57197), .A3(n57196), .Z(n57201) );
  INAND2HSV0 U59534 ( .A1(n57199), .B1(n26692), .ZN(n57200) );
  XNOR2HSV1 U59535 ( .A1(n57201), .A2(n57200), .ZN(n57202) );
  XNOR2HSV1 U59536 ( .A1(n57203), .A2(n57202), .ZN(n57207) );
  NOR2HSV2 U59537 ( .A1(n29774), .A2(n57204), .ZN(n57206) );
  XOR3HSV2 U59538 ( .A1(n57207), .A2(n57206), .A3(n57205), .Z(po4) );
  CLKNAND2HSV1 U59539 ( .A1(n50318), .A2(n57208), .ZN(n57320) );
  CLKNAND2HSV1 U59540 ( .A1(n58104), .A2(n34020), .ZN(n57314) );
  CLKNAND2HSV0 U59541 ( .A1(n58218), .A2(n35318), .ZN(n57312) );
  NAND2HSV0 U59542 ( .A1(n57324), .A2(n57888), .ZN(n57306) );
  NAND2HSV0 U59543 ( .A1(n57209), .A2(n58153), .ZN(n57304) );
  NAND2HSV0 U59544 ( .A1(n57404), .A2(n58184), .ZN(n57295) );
  NAND2HSV0 U59545 ( .A1(n59524), .A2(n59832), .ZN(n57291) );
  NAND2HSV0 U59546 ( .A1(n57210), .A2(n58156), .ZN(n57212) );
  NAND2HSV0 U59547 ( .A1(n33965), .A2(n58116), .ZN(n57211) );
  XOR2HSV0 U59548 ( .A1(n57212), .A2(n57211), .Z(n57216) );
  NOR2HSV0 U59549 ( .A1(n58174), .A2(n33350), .ZN(n57214) );
  NAND2HSV0 U59550 ( .A1(n57506), .A2(n33712), .ZN(n57213) );
  XOR2HSV0 U59551 ( .A1(n57214), .A2(n57213), .Z(n57215) );
  XNOR2HSV1 U59552 ( .A1(n57216), .A2(n57215), .ZN(n57229) );
  CLKNHSV0 U59553 ( .I(n57217), .ZN(n57221) );
  AOI22HSV0 U59554 ( .A1(n34743), .A2(n57986), .B1(n57218), .B2(n58069), .ZN(
        n57219) );
  AOI21HSV2 U59555 ( .A1(n57221), .A2(n57220), .B(n57219), .ZN(n57227) );
  CLKNHSV0 U59556 ( .I(n57222), .ZN(n57225) );
  AOI22HSV0 U59557 ( .A1(n59834), .A2(n58301), .B1(n57510), .B2(n57837), .ZN(
        n57223) );
  AOI21HSV2 U59558 ( .A1(n57225), .A2(n57224), .B(n57223), .ZN(n57226) );
  XOR2HSV0 U59559 ( .A1(n57227), .A2(n57226), .Z(n57228) );
  XNOR2HSV1 U59560 ( .A1(n57229), .A2(n57228), .ZN(n57250) );
  NAND2HSV0 U59561 ( .A1(n57230), .A2(\pe4/bq[28] ), .ZN(n57233) );
  AOI22HSV0 U59562 ( .A1(n57497), .A2(n57233), .B1(n57232), .B2(n57231), .ZN(
        n57239) );
  NAND2HSV0 U59563 ( .A1(n57234), .A2(n34480), .ZN(n57516) );
  NOR2HSV0 U59564 ( .A1(n57235), .A2(n57516), .ZN(n57237) );
  AOI22HSV0 U59565 ( .A1(n57140), .A2(n58127), .B1(n49943), .B2(n59952), .ZN(
        n57236) );
  NOR2HSV1 U59566 ( .A1(n57237), .A2(n57236), .ZN(n57238) );
  XOR2HSV0 U59567 ( .A1(n57239), .A2(n57238), .Z(n57248) );
  NOR2HSV0 U59568 ( .A1(n57240), .A2(n57347), .ZN(n57244) );
  AOI22HSV0 U59569 ( .A1(n35377), .A2(n57241), .B1(n59383), .B2(\pe4/bq[2] ), 
        .ZN(n57243) );
  NOR2HSV2 U59570 ( .A1(n57244), .A2(n57243), .ZN(n57246) );
  XOR2HSV0 U59571 ( .A1(n57246), .A2(n57245), .Z(n57247) );
  XOR2HSV0 U59572 ( .A1(n57248), .A2(n57247), .Z(n57249) );
  XNOR2HSV1 U59573 ( .A1(n57250), .A2(n57249), .ZN(n57289) );
  NAND2HSV0 U59574 ( .A1(n57251), .A2(n58314), .ZN(n57268) );
  NAND2HSV0 U59575 ( .A1(n59951), .A2(\pe4/bq[11] ), .ZN(n57253) );
  NAND2HSV0 U59576 ( .A1(n57504), .A2(n57476), .ZN(n57252) );
  XOR2HSV0 U59577 ( .A1(n57253), .A2(n57252), .Z(n57258) );
  NAND2HSV0 U59578 ( .A1(\pe4/aot [11]), .A2(n34254), .ZN(n57256) );
  NAND2HSV0 U59579 ( .A1(n59954), .A2(n57254), .ZN(n57255) );
  XOR2HSV0 U59580 ( .A1(n57256), .A2(n57255), .Z(n57257) );
  XOR2HSV0 U59581 ( .A1(n57258), .A2(n57257), .Z(n57266) );
  NAND2HSV0 U59582 ( .A1(n59661), .A2(n57851), .ZN(n57259) );
  XOR2HSV0 U59583 ( .A1(n57849), .A2(n57259), .Z(n57264) );
  NOR2HSV0 U59584 ( .A1(n49929), .A2(n57260), .ZN(n57262) );
  NAND2HSV0 U59585 ( .A1(n57727), .A2(n58130), .ZN(n57261) );
  XOR2HSV0 U59586 ( .A1(n57262), .A2(n57261), .Z(n57263) );
  XOR2HSV0 U59587 ( .A1(n57264), .A2(n57263), .Z(n57265) );
  XOR2HSV0 U59588 ( .A1(n57266), .A2(n57265), .Z(n57267) );
  XOR2HSV0 U59589 ( .A1(n57268), .A2(n57267), .Z(n57288) );
  NAND2HSV0 U59590 ( .A1(\pe4/aot [2]), .A2(n46617), .ZN(n57270) );
  NAND2HSV0 U59591 ( .A1(n57463), .A2(n57368), .ZN(n57269) );
  XOR2HSV0 U59592 ( .A1(n57270), .A2(n57269), .Z(n57274) );
  NAND2HSV0 U59593 ( .A1(\pe4/aot [1]), .A2(n33423), .ZN(n57272) );
  NAND2HSV0 U59594 ( .A1(n47718), .A2(n34044), .ZN(n57271) );
  XOR2HSV0 U59595 ( .A1(n57272), .A2(n57271), .Z(n57273) );
  XOR2HSV0 U59596 ( .A1(n57274), .A2(n57273), .Z(n57282) );
  NAND2HSV0 U59597 ( .A1(n59632), .A2(n57337), .ZN(n57276) );
  NAND2HSV0 U59598 ( .A1(n59343), .A2(\pe4/bq[20] ), .ZN(n57275) );
  XOR2HSV0 U59599 ( .A1(n57276), .A2(n57275), .Z(n57280) );
  NAND2HSV0 U59600 ( .A1(\pe4/aot [14]), .A2(n57906), .ZN(n57278) );
  NAND2HSV0 U59601 ( .A1(n33716), .A2(n58113), .ZN(n57277) );
  XOR2HSV0 U59602 ( .A1(n57278), .A2(n57277), .Z(n57279) );
  XOR2HSV0 U59603 ( .A1(n57280), .A2(n57279), .Z(n57281) );
  XOR2HSV0 U59604 ( .A1(n57282), .A2(n57281), .Z(n57284) );
  NAND2HSV0 U59605 ( .A1(n34127), .A2(n57680), .ZN(n57283) );
  XNOR2HSV1 U59606 ( .A1(n57284), .A2(n57283), .ZN(n57287) );
  NAND2HSV0 U59607 ( .A1(n57285), .A2(n57584), .ZN(n57286) );
  XOR4HSV1 U59608 ( .A1(n57289), .A2(n57288), .A3(n57287), .A4(n57286), .Z(
        n57290) );
  XNOR2HSV1 U59609 ( .A1(n57291), .A2(n57290), .ZN(n57293) );
  NAND2HSV0 U59610 ( .A1(n59662), .A2(n57951), .ZN(n57292) );
  XNOR2HSV1 U59611 ( .A1(n57293), .A2(n57292), .ZN(n57294) );
  XNOR2HSV1 U59612 ( .A1(n57295), .A2(n57294), .ZN(n57297) );
  NAND2HSV0 U59613 ( .A1(n57405), .A2(n58036), .ZN(n57296) );
  XNOR2HSV1 U59614 ( .A1(n57297), .A2(n57296), .ZN(n57299) );
  NAND2HSV0 U59615 ( .A1(n57679), .A2(\pe4/got [8]), .ZN(n57298) );
  XOR2HSV0 U59616 ( .A1(n57299), .A2(n57298), .Z(n57302) );
  NAND2HSV0 U59617 ( .A1(n57458), .A2(n58041), .ZN(n57301) );
  CLKNAND2HSV0 U59618 ( .A1(n57183), .A2(n59663), .ZN(n57300) );
  XOR3HSV1 U59619 ( .A1(n57302), .A2(n57301), .A3(n57300), .Z(n57303) );
  XNOR2HSV1 U59620 ( .A1(n57304), .A2(n57303), .ZN(n57305) );
  XOR2HSV0 U59621 ( .A1(n57312), .A2(n57311), .Z(n57313) );
  XOR2HSV0 U59622 ( .A1(n57314), .A2(n57313), .Z(n57316) );
  CLKNAND2HSV0 U59623 ( .A1(n57970), .A2(n59350), .ZN(n57315) );
  XNOR2HSV1 U59624 ( .A1(n57316), .A2(n57315), .ZN(n57318) );
  INAND2HSV0 U59625 ( .A1(n35034), .B1(n26692), .ZN(n57317) );
  XOR2HSV0 U59626 ( .A1(n57318), .A2(n57317), .Z(n57319) );
  XNOR2HSV1 U59627 ( .A1(n57320), .A2(n57319), .ZN(n57323) );
  OR2HSV1 U59628 ( .A1(n26413), .A2(n34718), .Z(n57321) );
  XOR3HSV2 U59629 ( .A1(n57323), .A2(n57322), .A3(n57321), .Z(\pe4/poht [1])
         );
  NAND2HSV2 U59630 ( .A1(n58299), .A2(\pe4/got [28]), .ZN(n57452) );
  CLKNAND2HSV1 U59631 ( .A1(n58141), .A2(\pe4/got [25]), .ZN(n57446) );
  CLKNAND2HSV1 U59632 ( .A1(n58218), .A2(n57574), .ZN(n57444) );
  CLKNAND2HSV0 U59633 ( .A1(n58112), .A2(n50404), .ZN(n57435) );
  NAND2HSV0 U59634 ( .A1(n57675), .A2(n57820), .ZN(n57423) );
  NAND2HSV0 U59635 ( .A1(n57324), .A2(n58153), .ZN(n57421) );
  CLKNAND2HSV0 U59636 ( .A1(n57678), .A2(n57646), .ZN(n57418) );
  NAND2HSV0 U59637 ( .A1(n57458), .A2(\pe4/got [8]), .ZN(n57412) );
  NAND2HSV0 U59638 ( .A1(n57325), .A2(n57584), .ZN(n57401) );
  NOR2HSV0 U59639 ( .A1(n57326), .A2(n48032), .ZN(n57496) );
  AOI22HSV0 U59640 ( .A1(n57327), .A2(\pe4/bq[5] ), .B1(n57727), .B2(n57684), 
        .ZN(n57328) );
  AOI21HSV1 U59641 ( .A1(n57329), .A2(n57496), .B(n57328), .ZN(n57334) );
  NAND2HSV0 U59642 ( .A1(n59951), .A2(n58196), .ZN(n57604) );
  NOR2HSV0 U59643 ( .A1(n57330), .A2(n57604), .ZN(n57332) );
  AOI22HSV0 U59644 ( .A1(n35533), .A2(n58301), .B1(n59951), .B2(n58116), .ZN(
        n57331) );
  NOR2HSV1 U59645 ( .A1(n57332), .A2(n57331), .ZN(n57333) );
  XOR2HSV0 U59646 ( .A1(n57334), .A2(n57333), .Z(n57358) );
  NAND2HSV0 U59647 ( .A1(n47718), .A2(n57505), .ZN(n57336) );
  NAND2HSV0 U59648 ( .A1(n57504), .A2(n34044), .ZN(n57335) );
  XOR2HSV0 U59649 ( .A1(n57336), .A2(n57335), .Z(n57342) );
  NAND2HSV0 U59650 ( .A1(n57506), .A2(n57476), .ZN(n57340) );
  NAND2HSV0 U59651 ( .A1(n57338), .A2(n57337), .ZN(n57339) );
  XOR2HSV0 U59652 ( .A1(n57340), .A2(n57339), .Z(n57341) );
  XNOR2HSV1 U59653 ( .A1(n57342), .A2(n57341), .ZN(n57357) );
  NAND2HSV0 U59654 ( .A1(n59954), .A2(n35194), .ZN(n57346) );
  CLKNHSV0 U59655 ( .I(n57343), .ZN(n57345) );
  AOI22HSV0 U59656 ( .A1(n57347), .A2(n57346), .B1(n57345), .B2(n57344), .ZN(
        n57351) );
  NAND2HSV0 U59657 ( .A1(\pe4/aot [11]), .A2(n57348), .ZN(n57731) );
  XOR2HSV0 U59658 ( .A1(n57351), .A2(n57350), .Z(n57355) );
  NAND2HSV0 U59659 ( .A1(n33867), .A2(n58127), .ZN(n57352) );
  XOR2HSV0 U59660 ( .A1(n57353), .A2(n57352), .Z(n57354) );
  XNOR2HSV1 U59661 ( .A1(n57355), .A2(n57354), .ZN(n57356) );
  XOR3HSV2 U59662 ( .A1(n57358), .A2(n57357), .A3(n57356), .Z(n57361) );
  NAND2HSV0 U59663 ( .A1(n57359), .A2(n57680), .ZN(n57360) );
  XNOR2HSV1 U59664 ( .A1(n57361), .A2(n57360), .ZN(n57397) );
  NAND2HSV0 U59665 ( .A1(n59838), .A2(n57851), .ZN(n57363) );
  NAND2HSV0 U59666 ( .A1(n58198), .A2(n33712), .ZN(n57362) );
  XOR2HSV0 U59667 ( .A1(n57363), .A2(n57362), .Z(n57367) );
  NAND2HSV0 U59668 ( .A1(n59953), .A2(\pe4/bq[16] ), .ZN(n57365) );
  NAND2HSV0 U59669 ( .A1(n57463), .A2(n57906), .ZN(n57364) );
  XOR2HSV0 U59670 ( .A1(n57365), .A2(n57364), .Z(n57366) );
  XOR2HSV0 U59671 ( .A1(n57367), .A2(n57366), .Z(n57376) );
  NAND2HSV0 U59672 ( .A1(n58307), .A2(n33427), .ZN(n57370) );
  NAND2HSV0 U59673 ( .A1(\pe4/aot [12]), .A2(n57368), .ZN(n57369) );
  XOR2HSV0 U59674 ( .A1(n57370), .A2(n57369), .Z(n57374) );
  NAND2HSV0 U59675 ( .A1(\pe4/aot [14]), .A2(\pe4/bq[17] ), .ZN(n57372) );
  NAND2HSV0 U59676 ( .A1(n58223), .A2(n57460), .ZN(n57371) );
  XOR2HSV0 U59677 ( .A1(n57372), .A2(n57371), .Z(n57373) );
  XOR2HSV0 U59678 ( .A1(n57374), .A2(n57373), .Z(n57375) );
  XOR2HSV0 U59679 ( .A1(n57376), .A2(n57375), .Z(n57395) );
  NAND2HSV0 U59680 ( .A1(n59834), .A2(\pe4/bq[2] ), .ZN(n57379) );
  NAND2HSV0 U59681 ( .A1(\pe4/aot [2]), .A2(n57377), .ZN(n57378) );
  XOR2HSV0 U59682 ( .A1(n57379), .A2(n57378), .Z(n57383) );
  NAND2HSV0 U59683 ( .A1(n57140), .A2(n57986), .ZN(n57381) );
  NAND2HSV0 U59684 ( .A1(n58230), .A2(n46617), .ZN(n57380) );
  XOR2HSV0 U59685 ( .A1(n57381), .A2(n57380), .Z(n57382) );
  XOR2HSV0 U59686 ( .A1(n57383), .A2(n57382), .Z(n57393) );
  NAND2HSV0 U59687 ( .A1(n57384), .A2(n58130), .ZN(n57386) );
  NAND2HSV0 U59688 ( .A1(n57510), .A2(n58156), .ZN(n57385) );
  XOR2HSV0 U59689 ( .A1(n57386), .A2(n57385), .Z(n57391) );
  NOR2HSV0 U59690 ( .A1(n35175), .A2(n57387), .ZN(n57389) );
  NAND2HSV0 U59691 ( .A1(n34743), .A2(\pe4/bq[11] ), .ZN(n57388) );
  XOR2HSV0 U59692 ( .A1(n57389), .A2(n57388), .Z(n57390) );
  XOR2HSV0 U59693 ( .A1(n57391), .A2(n57390), .Z(n57392) );
  XOR2HSV0 U59694 ( .A1(n57393), .A2(n57392), .Z(n57394) );
  XOR2HSV0 U59695 ( .A1(n57395), .A2(n57394), .Z(n57396) );
  XNOR2HSV1 U59696 ( .A1(n57397), .A2(n57396), .ZN(n57399) );
  NOR2HSV0 U59697 ( .A1(n33437), .A2(n58325), .ZN(n57398) );
  XNOR2HSV1 U59698 ( .A1(n57399), .A2(n57398), .ZN(n57400) );
  XNOR2HSV1 U59699 ( .A1(n57401), .A2(n57400), .ZN(n57403) );
  NAND2HSV0 U59700 ( .A1(n29780), .A2(n57744), .ZN(n57402) );
  XNOR2HSV1 U59701 ( .A1(n57403), .A2(n57402), .ZN(n57408) );
  NAND2HSV0 U59702 ( .A1(n57404), .A2(n57677), .ZN(n57407) );
  NAND2HSV0 U59703 ( .A1(n57405), .A2(n58184), .ZN(n57406) );
  XOR3HSV2 U59704 ( .A1(n57408), .A2(n57407), .A3(n57406), .Z(n57410) );
  NAND2HSV0 U59705 ( .A1(n35401), .A2(\pe4/got [7]), .ZN(n57409) );
  XOR2HSV0 U59706 ( .A1(n57410), .A2(n57409), .Z(n57411) );
  XNOR2HSV1 U59707 ( .A1(n57412), .A2(n57411), .ZN(n57416) );
  NAND2HSV0 U59708 ( .A1(n57414), .A2(n57413), .ZN(n57415) );
  XNOR2HSV1 U59709 ( .A1(n57416), .A2(n57415), .ZN(n57417) );
  XNOR2HSV1 U59710 ( .A1(n57418), .A2(n57417), .ZN(n57420) );
  NAND2HSV0 U59711 ( .A1(n25409), .A2(n57888), .ZN(n57419) );
  XOR3HSV2 U59712 ( .A1(n57421), .A2(n57420), .A3(n57419), .Z(n57422) );
  XNOR2HSV1 U59713 ( .A1(n57423), .A2(n57422), .ZN(n57426) );
  NAND2HSV0 U59714 ( .A1(n57985), .A2(n57424), .ZN(n57425) );
  XNOR2HSV1 U59715 ( .A1(n57426), .A2(n57425), .ZN(n57430) );
  NAND2HSV0 U59716 ( .A1(n57550), .A2(n57752), .ZN(n57429) );
  CLKNAND2HSV0 U59717 ( .A1(n57427), .A2(n47656), .ZN(n57428) );
  XOR3HSV1 U59718 ( .A1(n57430), .A2(n57429), .A3(n57428), .Z(n57433) );
  CLKNAND2HSV1 U59719 ( .A1(n58029), .A2(n57834), .ZN(n57432) );
  CLKNAND2HSV0 U59720 ( .A1(n57554), .A2(n57457), .ZN(n57431) );
  XOR3HSV2 U59721 ( .A1(n57433), .A2(n57432), .A3(n57431), .Z(n57434) );
  XNOR2HSV1 U59722 ( .A1(n57435), .A2(n57434), .ZN(n57438) );
  NAND2HSV2 U59723 ( .A1(n47841), .A2(n57760), .ZN(n57437) );
  NAND2HSV0 U59724 ( .A1(n57560), .A2(n57564), .ZN(n57436) );
  XOR3HSV2 U59725 ( .A1(n57438), .A2(n57437), .A3(n57436), .Z(n57440) );
  CLKNAND2HSV0 U59726 ( .A1(n25427), .A2(n59601), .ZN(n57439) );
  XNOR2HSV1 U59727 ( .A1(n57440), .A2(n57439), .ZN(n57442) );
  CLKNAND2HSV0 U59728 ( .A1(n35033), .A2(\pe4/got [23]), .ZN(n57441) );
  XNOR2HSV1 U59729 ( .A1(n57442), .A2(n57441), .ZN(n57443) );
  XNOR2HSV1 U59730 ( .A1(n57444), .A2(n57443), .ZN(n57445) );
  XOR2HSV0 U59731 ( .A1(n57446), .A2(n57445), .Z(n57448) );
  CLKNAND2HSV0 U59732 ( .A1(n57970), .A2(n33708), .ZN(n57447) );
  XNOR2HSV1 U59733 ( .A1(n57452), .A2(n57451), .ZN(n57456) );
  NOR2HSV2 U59734 ( .A1(n29774), .A2(n57453), .ZN(n57455) );
  NAND2HSV2 U59735 ( .A1(n57900), .A2(n35445), .ZN(n57454) );
  XOR3HSV2 U59736 ( .A1(n57456), .A2(n57455), .A3(n57454), .Z(\pe4/poht [2])
         );
  NAND2HSV2 U59737 ( .A1(n26417), .A2(n33708), .ZN(n57580) );
  CLKNAND2HSV1 U59738 ( .A1(n58141), .A2(n34239), .ZN(n57573) );
  CLKNAND2HSV1 U59739 ( .A1(n58218), .A2(n59601), .ZN(n57571) );
  CLKNAND2HSV1 U59740 ( .A1(n50065), .A2(n57457), .ZN(n57559) );
  CLKNAND2HSV1 U59741 ( .A1(n59378), .A2(n58153), .ZN(n57546) );
  NAND2HSV0 U59742 ( .A1(n59835), .A2(n58140), .ZN(n57544) );
  NAND2HSV0 U59743 ( .A1(n57678), .A2(\pe4/got [8]), .ZN(n57541) );
  NAND2HSV0 U59744 ( .A1(n57458), .A2(n58137), .ZN(n57537) );
  NAND2HSV0 U59745 ( .A1(n58307), .A2(n57459), .ZN(n57462) );
  NAND2HSV0 U59746 ( .A1(\pe4/aot [3]), .A2(n57460), .ZN(n57461) );
  XOR2HSV0 U59747 ( .A1(n57462), .A2(n57461), .Z(n57467) );
  NAND2HSV0 U59748 ( .A1(n47718), .A2(n50250), .ZN(n57465) );
  NAND2HSV0 U59749 ( .A1(n57463), .A2(\pe4/bq[16] ), .ZN(n57464) );
  XOR2HSV0 U59750 ( .A1(n57465), .A2(n57464), .Z(n57466) );
  XOR2HSV0 U59751 ( .A1(n57467), .A2(n57466), .Z(n57475) );
  CLKNAND2HSV0 U59752 ( .A1(\pe4/aot [2]), .A2(n34598), .ZN(n57469) );
  NAND2HSV0 U59753 ( .A1(n58230), .A2(n33966), .ZN(n57468) );
  XOR2HSV0 U59754 ( .A1(n57469), .A2(n57468), .Z(n57473) );
  NAND2HSV0 U59755 ( .A1(n59951), .A2(n58130), .ZN(n57471) );
  NAND2HSV0 U59756 ( .A1(n34743), .A2(n57798), .ZN(n57470) );
  XOR2HSV0 U59757 ( .A1(n57471), .A2(n57470), .Z(n57472) );
  XOR2HSV0 U59758 ( .A1(n57473), .A2(n57472), .Z(n57474) );
  XOR2HSV0 U59759 ( .A1(n57475), .A2(n57474), .Z(n57492) );
  NAND2HSV0 U59760 ( .A1(n58223), .A2(n34120), .ZN(n57478) );
  NAND2HSV0 U59761 ( .A1(n59352), .A2(n57476), .ZN(n57477) );
  XOR2HSV0 U59762 ( .A1(n57478), .A2(n57477), .Z(n57482) );
  NAND2HSV0 U59763 ( .A1(n57140), .A2(n58116), .ZN(n57480) );
  NAND2HSV0 U59764 ( .A1(n35533), .A2(n57241), .ZN(n57479) );
  XOR2HSV0 U59765 ( .A1(n57480), .A2(n57479), .Z(n57481) );
  XOR2HSV0 U59766 ( .A1(n57482), .A2(n57481), .Z(n57490) );
  NAND2HSV0 U59767 ( .A1(n58198), .A2(\pe4/bq[22] ), .ZN(n57484) );
  NAND2HSV0 U59768 ( .A1(n33867), .A2(\pe4/bq[11] ), .ZN(n57483) );
  XOR2HSV0 U59769 ( .A1(n57484), .A2(n57483), .Z(n57488) );
  NAND2HSV0 U59770 ( .A1(\pe4/aot [17]), .A2(n58077), .ZN(n57486) );
  NAND2HSV0 U59771 ( .A1(n34873), .A2(\pe4/bq[17] ), .ZN(n57485) );
  XOR2HSV0 U59772 ( .A1(n57486), .A2(n57485), .Z(n57487) );
  XOR2HSV0 U59773 ( .A1(n57488), .A2(n57487), .Z(n57489) );
  XOR2HSV0 U59774 ( .A1(n57490), .A2(n57489), .Z(n57491) );
  XOR2HSV0 U59775 ( .A1(n57492), .A2(n57491), .Z(n57525) );
  NOR2HSV0 U59776 ( .A1(n46143), .A2(n50351), .ZN(n57495) );
  OAI22HSV2 U59777 ( .A1(n57496), .A2(n57495), .B1(n57494), .B2(n57493), .ZN(
        n57503) );
  NAND2HSV0 U59778 ( .A1(\pe4/aot [22]), .A2(n58156), .ZN(n57722) );
  NOR2HSV0 U59779 ( .A1(n57497), .A2(n57722), .ZN(n57501) );
  AOI22HSV0 U59780 ( .A1(n57499), .A2(n57498), .B1(\pe4/aot [22]), .B2(n58197), 
        .ZN(n57500) );
  NOR2HSV1 U59781 ( .A1(n57501), .A2(n57500), .ZN(n57502) );
  XOR2HSV0 U59782 ( .A1(n57503), .A2(n57502), .Z(n57523) );
  NAND2HSV0 U59783 ( .A1(n57504), .A2(n57785), .ZN(n57508) );
  NAND2HSV0 U59784 ( .A1(n57506), .A2(n57505), .ZN(n57507) );
  XOR2HSV0 U59785 ( .A1(n57508), .A2(n57507), .Z(n57514) );
  NOR2HSV0 U59786 ( .A1(n57509), .A2(n57010), .ZN(n57512) );
  NAND2HSV0 U59787 ( .A1(n57510), .A2(\pe4/bq[2] ), .ZN(n57511) );
  XOR2HSV0 U59788 ( .A1(n57512), .A2(n57511), .Z(n57513) );
  XNOR2HSV1 U59789 ( .A1(n57514), .A2(n57513), .ZN(n57522) );
  NAND2HSV0 U59790 ( .A1(\pe4/aot [15]), .A2(n58126), .ZN(n57515) );
  XOR2HSV0 U59791 ( .A1(n57516), .A2(n57515), .Z(n57520) );
  NOR2HSV0 U59792 ( .A1(n34470), .A2(n47818), .ZN(n57518) );
  NAND2HSV0 U59793 ( .A1(\pe4/aot [11]), .A2(\pe4/bq[18] ), .ZN(n57517) );
  XOR2HSV0 U59794 ( .A1(n57518), .A2(n57517), .Z(n57519) );
  XOR2HSV0 U59795 ( .A1(n57520), .A2(n57519), .Z(n57521) );
  XOR3HSV2 U59796 ( .A1(n57523), .A2(n57522), .A3(n57521), .Z(n57524) );
  XNOR2HSV1 U59797 ( .A1(n57525), .A2(n57524), .ZN(n57529) );
  NAND2HSV0 U59798 ( .A1(n59524), .A2(n59958), .ZN(n57528) );
  NAND2HSV0 U59799 ( .A1(n34396), .A2(n59346), .ZN(n57527) );
  XOR3HSV2 U59800 ( .A1(n57529), .A2(n57528), .A3(n57527), .Z(n57533) );
  NAND2HSV0 U59801 ( .A1(n57530), .A2(n57584), .ZN(n57532) );
  NAND2HSV0 U59802 ( .A1(n59681), .A2(n57744), .ZN(n57531) );
  XOR3HSV2 U59803 ( .A1(n57533), .A2(n57532), .A3(n57531), .Z(n57535) );
  NAND2HSV0 U59804 ( .A1(n47742), .A2(n58246), .ZN(n57534) );
  XOR2HSV0 U59805 ( .A1(n57535), .A2(n57534), .Z(n57536) );
  XNOR2HSV1 U59806 ( .A1(n57537), .A2(n57536), .ZN(n57539) );
  CLKNAND2HSV1 U59807 ( .A1(n59928), .A2(\pe4/got [7]), .ZN(n57538) );
  XNOR2HSV1 U59808 ( .A1(n57539), .A2(n57538), .ZN(n57540) );
  XNOR2HSV1 U59809 ( .A1(n57541), .A2(n57540), .ZN(n57543) );
  NAND2HSV2 U59810 ( .A1(n59845), .A2(n57646), .ZN(n57542) );
  XOR3HSV2 U59811 ( .A1(n57544), .A2(n57543), .A3(n57542), .Z(n57545) );
  XNOR2HSV1 U59812 ( .A1(n57546), .A2(n57545), .ZN(n57549) );
  NAND2HSV0 U59813 ( .A1(n25284), .A2(n57888), .ZN(n57548) );
  XNOR2HSV1 U59814 ( .A1(n57549), .A2(n57548), .ZN(n57553) );
  NAND2HSV0 U59815 ( .A1(n57550), .A2(n57820), .ZN(n57552) );
  CLKNAND2HSV1 U59816 ( .A1(n49951), .A2(n57674), .ZN(n57551) );
  XOR3HSV1 U59817 ( .A1(n57553), .A2(n57552), .A3(n57551), .Z(n57557) );
  NAND2HSV2 U59818 ( .A1(n57189), .A2(n57308), .ZN(n57556) );
  CLKNAND2HSV1 U59819 ( .A1(n57554), .A2(n57752), .ZN(n57555) );
  XOR3HSV2 U59820 ( .A1(n57557), .A2(n57556), .A3(n57555), .Z(n57558) );
  XNOR2HSV1 U59821 ( .A1(n57559), .A2(n57558), .ZN(n57563) );
  NAND2HSV2 U59822 ( .A1(n47841), .A2(n35321), .ZN(n57562) );
  NAND2HSV0 U59823 ( .A1(n57560), .A2(n57754), .ZN(n57561) );
  XOR3HSV2 U59824 ( .A1(n57563), .A2(n57562), .A3(n57561), .Z(n57566) );
  CLKNAND2HSV1 U59825 ( .A1(n47904), .A2(n57564), .ZN(n57565) );
  XNOR2HSV1 U59826 ( .A1(n57566), .A2(n57565), .ZN(n57569) );
  CLKNAND2HSV0 U59827 ( .A1(n35033), .A2(n57567), .ZN(n57568) );
  XNOR2HSV1 U59828 ( .A1(n57569), .A2(n57568), .ZN(n57570) );
  XOR2HSV0 U59829 ( .A1(n57571), .A2(n57570), .Z(n57572) );
  XOR2HSV0 U59830 ( .A1(n57573), .A2(n57572), .Z(n57576) );
  CLKNAND2HSV0 U59831 ( .A1(n57970), .A2(n57574), .ZN(n57575) );
  XNOR2HSV1 U59832 ( .A1(n57576), .A2(n57575), .ZN(n57578) );
  XOR2HSV0 U59833 ( .A1(n57578), .A2(n57577), .Z(n57579) );
  XNOR2HSV1 U59834 ( .A1(n57580), .A2(n57579), .ZN(n57583) );
  INAND2HSV2 U59835 ( .A1(n26413), .B1(n34966), .ZN(n57581) );
  XOR3HSV2 U59836 ( .A1(n57583), .A2(n57582), .A3(n57581), .Z(\pe4/poht [4])
         );
  NAND2HSV2 U59837 ( .A1(n50318), .A2(n57760), .ZN(n57668) );
  CLKNAND2HSV1 U59838 ( .A1(n58141), .A2(n57754), .ZN(n57662) );
  CLKNAND2HSV1 U59839 ( .A1(n57673), .A2(n34797), .ZN(n57660) );
  CLKNAND2HSV0 U59840 ( .A1(n50065), .A2(n59631), .ZN(n57651) );
  NAND2HSV0 U59841 ( .A1(n57675), .A2(n58184), .ZN(n57640) );
  CLKNAND2HSV0 U59842 ( .A1(n57676), .A2(n57744), .ZN(n57638) );
  CLKNAND2HSV0 U59843 ( .A1(n57678), .A2(n57584), .ZN(n57635) );
  NAND2HSV0 U59844 ( .A1(n59682), .A2(n57680), .ZN(n57631) );
  NAND2HSV0 U59845 ( .A1(n57585), .A2(\pe4/bq[11] ), .ZN(n57587) );
  NAND2HSV0 U59846 ( .A1(n57234), .A2(\pe4/bq[8] ), .ZN(n57586) );
  XOR2HSV0 U59847 ( .A1(n57587), .A2(n57586), .Z(n57591) );
  NAND2HSV0 U59848 ( .A1(\pe4/aot [22]), .A2(\pe4/bq[2] ), .ZN(n57589) );
  NAND2HSV0 U59849 ( .A1(\pe4/aot [17]), .A2(n57684), .ZN(n57588) );
  XOR2HSV0 U59850 ( .A1(n57589), .A2(n57588), .Z(n57590) );
  XOR2HSV0 U59851 ( .A1(n57591), .A2(n57590), .Z(n57601) );
  NAND2HSV0 U59852 ( .A1(\pe4/aot [7]), .A2(n57926), .ZN(n57594) );
  NAND2HSV0 U59853 ( .A1(n58230), .A2(n57592), .ZN(n57593) );
  XOR2HSV0 U59854 ( .A1(n57594), .A2(n57593), .Z(n57599) );
  NAND2HSV0 U59855 ( .A1(n34743), .A2(n57595), .ZN(n57597) );
  NAND2HSV0 U59856 ( .A1(n57852), .A2(n57798), .ZN(n57596) );
  XOR2HSV0 U59857 ( .A1(n57597), .A2(n57596), .Z(n57598) );
  XNOR2HSV1 U59858 ( .A1(n57599), .A2(n57598), .ZN(n57600) );
  XNOR2HSV1 U59859 ( .A1(n57601), .A2(n57600), .ZN(n57613) );
  NOR2HSV0 U59860 ( .A1(n58174), .A2(n48026), .ZN(n57720) );
  NAND2HSV0 U59861 ( .A1(\pe4/aot [18]), .A2(n57784), .ZN(n57603) );
  NAND2HSV0 U59862 ( .A1(n34873), .A2(\pe4/bq[12] ), .ZN(n57602) );
  XOR2HSV0 U59863 ( .A1(n57603), .A2(n57602), .Z(n57611) );
  CLKNHSV1 U59864 ( .I(n57604), .ZN(n57606) );
  NOR2HSV0 U59865 ( .A1(n57605), .A2(n48032), .ZN(n57781) );
  NAND2HSV0 U59866 ( .A1(\pe4/aot [21]), .A2(n58010), .ZN(n57726) );
  CLKNAND2HSV1 U59867 ( .A1(n50215), .A2(\pe4/bq[3] ), .ZN(n57782) );
  OAI22HSV1 U59868 ( .A1(n57606), .A2(n57781), .B1(n57726), .B2(n57782), .ZN(
        n57610) );
  NAND2HSV0 U59869 ( .A1(\pe4/aot [9]), .A2(n57348), .ZN(n57608) );
  NAND2HSV0 U59870 ( .A1(n34022), .A2(n57911), .ZN(n57607) );
  XOR2HSV0 U59871 ( .A1(n57608), .A2(n57607), .Z(n57609) );
  XOR4HSV1 U59872 ( .A1(n57720), .A2(n57611), .A3(n57610), .A4(n57609), .Z(
        n57612) );
  XNOR2HSV1 U59873 ( .A1(n57613), .A2(n57612), .ZN(n57629) );
  CLKNAND2HSV0 U59874 ( .A1(\pe4/aot [14]), .A2(n58116), .ZN(n57615) );
  NAND2HSV0 U59875 ( .A1(\pe4/aot [3]), .A2(n57505), .ZN(n57614) );
  XOR2HSV0 U59876 ( .A1(n57615), .A2(n57614), .Z(n57619) );
  CLKNAND2HSV1 U59877 ( .A1(\pe4/aot [2]), .A2(n33711), .ZN(n57617) );
  NAND2HSV0 U59878 ( .A1(n57683), .A2(n58126), .ZN(n57616) );
  XOR2HSV0 U59879 ( .A1(n57617), .A2(n57616), .Z(n57618) );
  XOR2HSV0 U59880 ( .A1(n57619), .A2(n57618), .Z(n57627) );
  NAND2HSV0 U59881 ( .A1(\pe4/aot [11]), .A2(n58127), .ZN(n57621) );
  NAND2HSV0 U59882 ( .A1(n58199), .A2(n57785), .ZN(n57620) );
  XOR2HSV0 U59883 ( .A1(n57621), .A2(n57620), .Z(n57625) );
  NOR2HSV0 U59884 ( .A1(n57775), .A2(n48024), .ZN(n57623) );
  NAND2HSV0 U59885 ( .A1(\pe4/aot [5]), .A2(n50250), .ZN(n57622) );
  XOR2HSV0 U59886 ( .A1(n57623), .A2(n57622), .Z(n57624) );
  XOR2HSV0 U59887 ( .A1(n57625), .A2(n57624), .Z(n57626) );
  XOR2HSV0 U59888 ( .A1(n57627), .A2(n57626), .Z(n57628) );
  XNOR2HSV1 U59889 ( .A1(n57629), .A2(n57628), .ZN(n57630) );
  XNOR2HSV1 U59890 ( .A1(n57631), .A2(n57630), .ZN(n57633) );
  CLKNAND2HSV0 U59891 ( .A1(n59928), .A2(n59346), .ZN(n57632) );
  XNOR2HSV1 U59892 ( .A1(n57633), .A2(n57632), .ZN(n57634) );
  XNOR2HSV1 U59893 ( .A1(n57635), .A2(n57634), .ZN(n57637) );
  NAND2HSV0 U59894 ( .A1(n25243), .A2(\pe4/got [5]), .ZN(n57636) );
  XOR3HSV2 U59895 ( .A1(n57638), .A2(n57637), .A3(n57636), .Z(n57639) );
  XNOR2HSV1 U59896 ( .A1(n57640), .A2(n57639), .ZN(n57642) );
  NOR2HSV0 U59897 ( .A1(n57816), .A2(n50064), .ZN(n57641) );
  XNOR2HSV1 U59898 ( .A1(n57642), .A2(n57641), .ZN(n57645) );
  NAND2HSV0 U59899 ( .A1(n34409), .A2(n58111), .ZN(n57644) );
  CLKNAND2HSV0 U59900 ( .A1(n49951), .A2(n57818), .ZN(n57643) );
  XOR3HSV1 U59901 ( .A1(n57645), .A2(n57644), .A3(n57643), .Z(n57649) );
  CLKNAND2HSV1 U59902 ( .A1(n58096), .A2(n58153), .ZN(n57648) );
  NAND2HSV0 U59903 ( .A1(n59935), .A2(n57646), .ZN(n57647) );
  XOR3HSV2 U59904 ( .A1(n57649), .A2(n57648), .A3(n57647), .Z(n57650) );
  XNOR2HSV1 U59905 ( .A1(n57651), .A2(n57650), .ZN(n57654) );
  CLKNAND2HSV0 U59906 ( .A1(n58183), .A2(n57674), .ZN(n57653) );
  CLKNAND2HSV0 U59907 ( .A1(n57960), .A2(\pe4/got [13]), .ZN(n57652) );
  XOR3HSV2 U59908 ( .A1(n57654), .A2(n57653), .A3(n57652), .Z(n57656) );
  CLKNAND2HSV1 U59909 ( .A1(n57889), .A2(n57752), .ZN(n57655) );
  XNOR2HSV1 U59910 ( .A1(n57656), .A2(n57655), .ZN(n57658) );
  CLKNAND2HSV0 U59911 ( .A1(n57755), .A2(n59604), .ZN(n57657) );
  XNOR2HSV1 U59912 ( .A1(n57658), .A2(n57657), .ZN(n57659) );
  XNOR2HSV1 U59913 ( .A1(n57660), .A2(n57659), .ZN(n57661) );
  XOR2HSV0 U59914 ( .A1(n57662), .A2(n57661), .Z(n57664) );
  CLKNAND2HSV0 U59915 ( .A1(n59348), .A2(n57770), .ZN(n57663) );
  CLKNAND2HSV1 U59916 ( .A1(n26516), .A2(n33831), .ZN(n57665) );
  XNOR2HSV1 U59917 ( .A1(n57668), .A2(n57667), .ZN(n57671) );
  NOR2HSV2 U59918 ( .A1(n29774), .A2(n49965), .ZN(n57670) );
  XOR3HSV2 U59919 ( .A1(n57671), .A2(n57670), .A3(n57669), .Z(\pe4/poht [9])
         );
  NAND2HSV2 U59920 ( .A1(n26417), .A2(n57672), .ZN(n57766) );
  CLKNAND2HSV1 U59921 ( .A1(n58141), .A2(n33831), .ZN(n57759) );
  CLKNAND2HSV1 U59922 ( .A1(n57673), .A2(n57770), .ZN(n57757) );
  CLKNAND2HSV0 U59923 ( .A1(n57676), .A2(n58137), .ZN(n57751) );
  CLKNAND2HSV0 U59924 ( .A1(n57678), .A2(n57677), .ZN(n57748) );
  NAND2HSV0 U59925 ( .A1(n59682), .A2(n58298), .ZN(n57743) );
  NAND2HSV0 U59926 ( .A1(n57679), .A2(n59346), .ZN(n57741) );
  NAND2HSV0 U59927 ( .A1(n59681), .A2(n57680), .ZN(n57739) );
  NAND2HSV0 U59928 ( .A1(\pe4/aot [14]), .A2(\pe4/bq[12] ), .ZN(n57682) );
  NAND2HSV0 U59929 ( .A1(n59632), .A2(n50250), .ZN(n57681) );
  XOR2HSV0 U59930 ( .A1(n57682), .A2(n57681), .Z(n57688) );
  NAND2HSV0 U59931 ( .A1(n57683), .A2(n49943), .ZN(n57686) );
  NAND2HSV0 U59932 ( .A1(n57859), .A2(n57684), .ZN(n57685) );
  XOR2HSV0 U59933 ( .A1(n57686), .A2(n57685), .Z(n57687) );
  XOR2HSV0 U59934 ( .A1(n57688), .A2(n57687), .Z(n57698) );
  NAND2HSV0 U59935 ( .A1(n57234), .A2(n58116), .ZN(n57690) );
  NAND2HSV0 U59936 ( .A1(n57230), .A2(\pe4/bq[22] ), .ZN(n57689) );
  XOR2HSV0 U59937 ( .A1(n57690), .A2(n57689), .Z(n57696) );
  NAND2HSV0 U59938 ( .A1(n57692), .A2(n57691), .ZN(n57694) );
  NAND2HSV0 U59939 ( .A1(n59839), .A2(n57784), .ZN(n57693) );
  XOR2HSV0 U59940 ( .A1(n57694), .A2(n57693), .Z(n57695) );
  XOR2HSV0 U59941 ( .A1(n57696), .A2(n57695), .Z(n57697) );
  XOR2HSV0 U59942 ( .A1(n57698), .A2(n57697), .Z(n57716) );
  NAND2HSV0 U59943 ( .A1(n34873), .A2(n58126), .ZN(n57700) );
  NAND2HSV0 U59944 ( .A1(\pe4/aot [5]), .A2(n34636), .ZN(n57699) );
  XOR2HSV0 U59945 ( .A1(n57700), .A2(n57699), .Z(n57704) );
  NOR2HSV0 U59946 ( .A1(n44338), .A2(n53219), .ZN(n57702) );
  NAND2HSV0 U59947 ( .A1(\pe4/aot [15]), .A2(\pe4/bq[11] ), .ZN(n57701) );
  XOR2HSV0 U59948 ( .A1(n57702), .A2(n57701), .Z(n57703) );
  XNOR2HSV1 U59949 ( .A1(n57704), .A2(n57703), .ZN(n57714) );
  NAND2HSV0 U59950 ( .A1(n57384), .A2(\pe4/bq[3] ), .ZN(n57706) );
  NAND2HSV0 U59951 ( .A1(\pe4/aot [2]), .A2(n34120), .ZN(n57705) );
  XOR2HSV0 U59952 ( .A1(n57706), .A2(n57705), .Z(n57712) );
  NOR2HSV0 U59953 ( .A1(n57026), .A2(n58013), .ZN(n57710) );
  NOR2HSV0 U59954 ( .A1(n57707), .A2(n47809), .ZN(n57709) );
  NAND2HSV2 U59955 ( .A1(\pe4/aot [9]), .A2(n57911), .ZN(n58222) );
  OAI22HSV0 U59956 ( .A1(n57710), .A2(n57709), .B1(n57708), .B2(n58222), .ZN(
        n57711) );
  XNOR2HSV1 U59957 ( .A1(n57712), .A2(n57711), .ZN(n57713) );
  XNOR2HSV1 U59958 ( .A1(n57714), .A2(n57713), .ZN(n57715) );
  XNOR2HSV1 U59959 ( .A1(n57716), .A2(n57715), .ZN(n57737) );
  CLKNHSV0 U59960 ( .I(n57717), .ZN(n57721) );
  AOI21HSV0 U59961 ( .A1(n59352), .A2(n57785), .B(n57718), .ZN(n57719) );
  AOI21HSV2 U59962 ( .A1(n57721), .A2(n57720), .B(n57719), .ZN(n57725) );
  XOR2HSV0 U59963 ( .A1(n57723), .A2(n57722), .Z(n57724) );
  XOR3HSV2 U59964 ( .A1(n57726), .A2(n57725), .A3(n57724), .Z(n57735) );
  NAND2HSV0 U59965 ( .A1(n57727), .A2(\pe4/bq[2] ), .ZN(n57729) );
  NAND2HSV0 U59966 ( .A1(n57014), .A2(n57135), .ZN(n57728) );
  XOR2HSV0 U59967 ( .A1(n57729), .A2(n57728), .Z(n57733) );
  NAND2HSV0 U59968 ( .A1(n59605), .A2(\pe4/bq[8] ), .ZN(n57730) );
  XOR2HSV0 U59969 ( .A1(n57731), .A2(n57730), .Z(n57732) );
  XOR2HSV0 U59970 ( .A1(n57733), .A2(n57732), .Z(n57734) );
  XOR2HSV0 U59971 ( .A1(n57735), .A2(n57734), .Z(n57736) );
  XNOR2HSV1 U59972 ( .A1(n57737), .A2(n57736), .ZN(n57738) );
  XNOR2HSV1 U59973 ( .A1(n57739), .A2(n57738), .ZN(n57740) );
  XNOR2HSV1 U59974 ( .A1(n57741), .A2(n57740), .ZN(n57742) );
  XNOR2HSV1 U59975 ( .A1(n57743), .A2(n57742), .ZN(n57746) );
  CLKNAND2HSV0 U59976 ( .A1(n34405), .A2(n57744), .ZN(n57745) );
  XNOR2HSV1 U59977 ( .A1(n57746), .A2(n57745), .ZN(n57747) );
  XNOR2HSV1 U59978 ( .A1(n57748), .A2(n57747), .ZN(n57750) );
  XNOR2HSV1 U59979 ( .A1(n57757), .A2(n57756), .ZN(n57758) );
  XOR2HSV0 U59980 ( .A1(n57759), .A2(n57758), .Z(n57762) );
  NAND2HSV0 U59981 ( .A1(n57760), .A2(n59348), .ZN(n57761) );
  XNOR2HSV1 U59982 ( .A1(n57762), .A2(n57761), .ZN(n57764) );
  CLKNAND2HSV1 U59983 ( .A1(n26516), .A2(n59601), .ZN(n57763) );
  XOR2HSV0 U59984 ( .A1(n57764), .A2(n57763), .Z(n57765) );
  XNOR2HSV1 U59985 ( .A1(n57766), .A2(n57765), .ZN(n57769) );
  NOR2HSV2 U59986 ( .A1(n29752), .A2(n35319), .ZN(n57768) );
  NAND2HSV2 U59987 ( .A1(n57900), .A2(n35318), .ZN(n57767) );
  XOR3HSV2 U59988 ( .A1(n57769), .A2(n57768), .A3(n57767), .Z(\pe4/poht [7])
         );
  NAND2HSV2 U59989 ( .A1(n50318), .A2(n57770), .ZN(n57829) );
  CLKNAND2HSV1 U59990 ( .A1(n57983), .A2(n57982), .ZN(n57822) );
  NAND2HSV0 U59991 ( .A1(n59835), .A2(n58314), .ZN(n57815) );
  NAND2HSV0 U59992 ( .A1(n59833), .A2(n58219), .ZN(n57814) );
  NAND2HSV0 U59993 ( .A1(n58230), .A2(n57505), .ZN(n57772) );
  NAND2HSV0 U59994 ( .A1(\pe4/aot [7]), .A2(n58084), .ZN(n57771) );
  XOR2HSV0 U59995 ( .A1(n57772), .A2(n57771), .Z(n57795) );
  NAND2HSV0 U59996 ( .A1(n35347), .A2(n58003), .ZN(n57774) );
  NAND2HSV0 U59997 ( .A1(\pe4/aot [11]), .A2(\pe4/bq[11] ), .ZN(n57773) );
  XOR2HSV0 U59998 ( .A1(n57774), .A2(n57773), .Z(n57780) );
  NOR2HSV0 U59999 ( .A1(n57775), .A2(n53217), .ZN(n57778) );
  NAND2HSV0 U60000 ( .A1(n59954), .A2(n50250), .ZN(n57777) );
  XOR2HSV0 U60001 ( .A1(n57778), .A2(n57777), .Z(n57779) );
  XNOR2HSV1 U60002 ( .A1(n57780), .A2(n57779), .ZN(n57794) );
  NAND2HSV0 U60003 ( .A1(n57014), .A2(n58010), .ZN(n57919) );
  NOR2HSV0 U60004 ( .A1(n35175), .A2(n57010), .ZN(n57921) );
  AOI22HSV2 U60005 ( .A1(n57782), .A2(n57919), .B1(n57921), .B2(n57781), .ZN(
        n57783) );
  NOR2HSV0 U60006 ( .A1(n58174), .A2(n48024), .ZN(n57848) );
  XOR2HSV0 U60007 ( .A1(n57783), .A2(n57848), .Z(n57793) );
  NAND2HSV0 U60008 ( .A1(n59952), .A2(n57784), .ZN(n57787) );
  NAND2HSV0 U60009 ( .A1(\pe4/aot [2]), .A2(n57785), .ZN(n57786) );
  XOR2HSV0 U60010 ( .A1(n57787), .A2(n57786), .Z(n57791) );
  NAND2HSV0 U60011 ( .A1(n59343), .A2(n58116), .ZN(n57789) );
  NAND2HSV0 U60012 ( .A1(\pe4/aot [21]), .A2(n57911), .ZN(n57788) );
  XOR2HSV0 U60013 ( .A1(n57789), .A2(n57788), .Z(n57790) );
  XOR2HSV0 U60014 ( .A1(n57791), .A2(n57790), .Z(n57792) );
  XOR4HSV1 U60015 ( .A1(n57795), .A2(n57794), .A3(n57793), .A4(n57792), .Z(
        n57812) );
  CLKNAND2HSV1 U60016 ( .A1(\pe4/aot [10]), .A2(n57986), .ZN(n57797) );
  NAND2HSV0 U60017 ( .A1(\pe4/aot [18]), .A2(n57595), .ZN(n57796) );
  XOR2HSV0 U60018 ( .A1(n57797), .A2(n57796), .Z(n57802) );
  NAND2HSV0 U60019 ( .A1(n59839), .A2(\pe4/bq[2] ), .ZN(n57800) );
  NAND2HSV0 U60020 ( .A1(n58163), .A2(n57798), .ZN(n57799) );
  XOR2HSV0 U60021 ( .A1(n57800), .A2(n57799), .Z(n57801) );
  XOR2HSV0 U60022 ( .A1(n57802), .A2(n57801), .Z(n57810) );
  NAND2HSV0 U60023 ( .A1(\pe4/aot [14]), .A2(n35184), .ZN(n57804) );
  NAND2HSV0 U60024 ( .A1(\pe4/aot [9]), .A2(n58127), .ZN(n57803) );
  XOR2HSV0 U60025 ( .A1(n57804), .A2(n57803), .Z(n57808) );
  NOR2HSV0 U60026 ( .A1(n49929), .A2(n47809), .ZN(n57806) );
  NAND2HSV0 U60027 ( .A1(\pe4/aot [4]), .A2(\pe4/bq[18] ), .ZN(n57805) );
  XOR2HSV0 U60028 ( .A1(n57806), .A2(n57805), .Z(n57807) );
  XOR2HSV0 U60029 ( .A1(n57808), .A2(n57807), .Z(n57809) );
  XOR2HSV0 U60030 ( .A1(n57810), .A2(n57809), .Z(n57811) );
  XNOR2HSV1 U60031 ( .A1(n57812), .A2(n57811), .ZN(n57813) );
  XNOR2HSV1 U60032 ( .A1(n57822), .A2(n57821), .ZN(n57825) );
  CLKNAND2HSV1 U60033 ( .A1(n58048), .A2(n57974), .ZN(n57824) );
  CLKNAND2HSV0 U60034 ( .A1(n34797), .A2(n59348), .ZN(n57823) );
  XOR3HSV2 U60035 ( .A1(n57825), .A2(n57824), .A3(n57823), .Z(n57827) );
  CLKNAND2HSV0 U60036 ( .A1(n58207), .A2(n57834), .ZN(n57826) );
  XNOR2HSV1 U60037 ( .A1(n57827), .A2(n57826), .ZN(n57828) );
  XNOR2HSV1 U60038 ( .A1(n57829), .A2(n57828), .ZN(n57833) );
  NOR2HSV2 U60039 ( .A1(n29752), .A2(n57830), .ZN(n57832) );
  NOR2HSV2 U60040 ( .A1(n26761), .A2(n50207), .ZN(n57831) );
  XOR3HSV2 U60041 ( .A1(n57833), .A2(n57832), .A3(n57831), .Z(\pe4/poht [11])
         );
  NAND2HSV2 U60042 ( .A1(n26417), .A2(n57834), .ZN(n57899) );
  NAND2HSV0 U60043 ( .A1(n57835), .A2(n57982), .ZN(n57893) );
  CLKNAND2HSV1 U60044 ( .A1(n58218), .A2(n58052), .ZN(n57891) );
  NAND2HSV0 U60045 ( .A1(n59835), .A2(n58219), .ZN(n57885) );
  AOI22HSV0 U60046 ( .A1(n59952), .A2(n57837), .B1(n58069), .B2(n58198), .ZN(
        n57838) );
  AOI21HSV0 U60047 ( .A1(n57840), .A2(n57839), .B(n57838), .ZN(n57845) );
  NOR2HSV0 U60048 ( .A1(n58194), .A2(n57841), .ZN(n58136) );
  AOI22HSV0 U60049 ( .A1(\pe4/aot [9]), .A2(n57986), .B1(n57906), .B2(n58283), 
        .ZN(n57842) );
  AOI21HSV0 U60050 ( .A1(n57843), .A2(n58136), .B(n57842), .ZN(n57844) );
  XOR2HSV0 U60051 ( .A1(n57845), .A2(n57844), .Z(n57858) );
  NOR2HSV0 U60052 ( .A1(n49929), .A2(n47818), .ZN(n57922) );
  AOI22HSV0 U60053 ( .A1(n59352), .A2(n57846), .B1(n49943), .B2(n58306), .ZN(
        n57847) );
  AOI21HSV1 U60054 ( .A1(n57848), .A2(n57922), .B(n57847), .ZN(n57856) );
  NAND2HSV2 U60055 ( .A1(\pe4/aot [4]), .A2(n58014), .ZN(n58226) );
  NOR2HSV0 U60056 ( .A1(n57849), .A2(n58226), .ZN(n57854) );
  AOI22HSV0 U60057 ( .A1(n57852), .A2(n57851), .B1(n57850), .B2(n58199), .ZN(
        n57853) );
  NOR2HSV1 U60058 ( .A1(n57854), .A2(n57853), .ZN(n57855) );
  XOR2HSV0 U60059 ( .A1(n57856), .A2(n57855), .Z(n57857) );
  XOR2HSV0 U60060 ( .A1(n57858), .A2(n57857), .Z(n57867) );
  NAND2HSV0 U60061 ( .A1(n57859), .A2(\pe4/bq[2] ), .ZN(n57861) );
  NAND2HSV0 U60062 ( .A1(\pe4/aot [17]), .A2(\pe4/bq[4] ), .ZN(n57860) );
  XOR2HSV0 U60063 ( .A1(n57861), .A2(n57860), .Z(n57865) );
  NAND2HSV0 U60064 ( .A1(\pe4/aot [11]), .A2(n58116), .ZN(n57863) );
  NAND2HSV0 U60065 ( .A1(n59343), .A2(\pe4/bq[9] ), .ZN(n57862) );
  XOR2HSV0 U60066 ( .A1(n57863), .A2(n57862), .Z(n57864) );
  XOR2HSV0 U60067 ( .A1(n57865), .A2(n57864), .Z(n57866) );
  XOR2HSV0 U60068 ( .A1(n57867), .A2(n57866), .Z(n57883) );
  NAND2HSV0 U60069 ( .A1(n57218), .A2(n58301), .ZN(n57869) );
  CLKNAND2HSV0 U60070 ( .A1(n47718), .A2(\pe4/bq[11] ), .ZN(n57868) );
  XOR2HSV0 U60071 ( .A1(n57869), .A2(n57868), .Z(n57873) );
  NAND2HSV0 U60072 ( .A1(n58230), .A2(n57785), .ZN(n57871) );
  NAND2HSV0 U60073 ( .A1(\pe4/aot [2]), .A2(n50250), .ZN(n57870) );
  XOR2HSV0 U60074 ( .A1(n57871), .A2(n57870), .Z(n57872) );
  XOR2HSV0 U60075 ( .A1(n57873), .A2(n57872), .Z(n57881) );
  NAND2HSV0 U60076 ( .A1(n58163), .A2(n35184), .ZN(n57875) );
  NAND2HSV0 U60077 ( .A1(n59839), .A2(n57911), .ZN(n57874) );
  XOR2HSV0 U60078 ( .A1(n57875), .A2(n57874), .Z(n57879) );
  NAND2HSV0 U60079 ( .A1(\pe4/aot [14]), .A2(n58003), .ZN(n57877) );
  NAND2HSV0 U60080 ( .A1(n58087), .A2(\pe4/bq[13] ), .ZN(n57876) );
  XOR2HSV0 U60081 ( .A1(n57877), .A2(n57876), .Z(n57878) );
  XOR2HSV0 U60082 ( .A1(n57879), .A2(n57878), .Z(n57880) );
  XOR2HSV0 U60083 ( .A1(n57881), .A2(n57880), .Z(n57882) );
  XNOR2HSV1 U60084 ( .A1(n57883), .A2(n57882), .ZN(n57884) );
  XNOR2HSV1 U60085 ( .A1(n57885), .A2(n57884), .ZN(n57886) );
  XNOR2HSV1 U60086 ( .A1(n57891), .A2(n57890), .ZN(n57892) );
  XOR2HSV0 U60087 ( .A1(n57893), .A2(n57892), .Z(n57895) );
  NAND2HSV0 U60088 ( .A1(n58272), .A2(n57974), .ZN(n57894) );
  XNOR2HSV1 U60089 ( .A1(n57895), .A2(n57894), .ZN(n57897) );
  CLKNAND2HSV0 U60090 ( .A1(n58207), .A2(n34797), .ZN(n57896) );
  XNOR2HSV1 U60091 ( .A1(n57897), .A2(n57896), .ZN(n57898) );
  XNOR2HSV1 U60092 ( .A1(n57899), .A2(n57898), .ZN(n57903) );
  NOR2HSV2 U60093 ( .A1(n29774), .A2(n50052), .ZN(n57902) );
  NAND2HSV2 U60094 ( .A1(n57900), .A2(n57564), .ZN(n57901) );
  XOR3HSV2 U60095 ( .A1(n57903), .A2(n57902), .A3(n57901), .Z(\pe4/poht [12])
         );
  CLKNAND2HSV1 U60096 ( .A1(n57983), .A2(n35400), .ZN(n57969) );
  CLKNAND2HSV0 U60097 ( .A1(n58112), .A2(n58111), .ZN(n57959) );
  NAND2HSV0 U60098 ( .A1(n59378), .A2(\pe4/got [2]), .ZN(n57948) );
  NAND2HSV0 U60099 ( .A1(n25243), .A2(n58219), .ZN(n57946) );
  CLKNAND2HSV0 U60100 ( .A1(n57993), .A2(n57986), .ZN(n57905) );
  CLKNAND2HSV0 U60101 ( .A1(\pe4/aot [6]), .A2(n58126), .ZN(n57904) );
  XOR2HSV0 U60102 ( .A1(n57905), .A2(n57904), .Z(n57910) );
  NAND2HSV0 U60103 ( .A1(n57218), .A2(\pe4/bq[2] ), .ZN(n57908) );
  NAND2HSV0 U60104 ( .A1(\pe4/aot [2]), .A2(n57906), .ZN(n57907) );
  XOR2HSV0 U60105 ( .A1(n57908), .A2(n57907), .Z(n57909) );
  XOR2HSV0 U60106 ( .A1(n57910), .A2(n57909), .Z(n57944) );
  CLKNAND2HSV0 U60107 ( .A1(n50215), .A2(n57911), .ZN(n57913) );
  NAND2HSV0 U60108 ( .A1(n59952), .A2(n58156), .ZN(n57912) );
  XOR2HSV0 U60109 ( .A1(n57913), .A2(n57912), .Z(n57917) );
  NOR2HSV0 U60110 ( .A1(n44338), .A2(n50114), .ZN(n57915) );
  NAND2HSV0 U60111 ( .A1(n57683), .A2(n58116), .ZN(n57914) );
  XOR2HSV0 U60112 ( .A1(n57915), .A2(n57914), .Z(n57916) );
  XNOR2HSV1 U60113 ( .A1(n57917), .A2(n57916), .ZN(n57925) );
  NOR2HSV0 U60114 ( .A1(n57918), .A2(n48032), .ZN(n57920) );
  NAND2HSV0 U60115 ( .A1(n35347), .A2(n58301), .ZN(n57991) );
  OAI22HSV1 U60116 ( .A1(n57921), .A2(n57920), .B1(n57991), .B2(n57919), .ZN(
        n57923) );
  XOR2HSV0 U60117 ( .A1(n57923), .A2(n57922), .Z(n57924) );
  XNOR2HSV1 U60118 ( .A1(n57925), .A2(n57924), .ZN(n57943) );
  NAND2HSV0 U60119 ( .A1(\pe4/aot [4]), .A2(\pe4/bq[16] ), .ZN(n57928) );
  NAND2HSV0 U60120 ( .A1(n59954), .A2(n57926), .ZN(n57927) );
  XOR2HSV0 U60121 ( .A1(n57928), .A2(n57927), .Z(n57933) );
  NAND2HSV0 U60122 ( .A1(\pe4/aot [9]), .A2(\pe4/bq[11] ), .ZN(n57931) );
  NAND2HSV0 U60123 ( .A1(n58230), .A2(n57929), .ZN(n57930) );
  XOR2HSV0 U60124 ( .A1(n57931), .A2(n57930), .Z(n57932) );
  XOR2HSV0 U60125 ( .A1(n57933), .A2(n57932), .Z(n57941) );
  NAND2HSV0 U60126 ( .A1(n59343), .A2(n35184), .ZN(n57935) );
  NAND2HSV0 U60127 ( .A1(\pe4/aot [11]), .A2(n57135), .ZN(n57934) );
  XOR2HSV0 U60128 ( .A1(n57935), .A2(n57934), .Z(n57939) );
  NAND2HSV0 U60129 ( .A1(\pe4/aot [7]), .A2(\pe4/bq[13] ), .ZN(n57937) );
  NAND2HSV0 U60130 ( .A1(\pe4/aot [14]), .A2(n58014), .ZN(n57936) );
  XOR2HSV0 U60131 ( .A1(n57937), .A2(n57936), .Z(n57938) );
  XOR2HSV0 U60132 ( .A1(n57939), .A2(n57938), .Z(n57940) );
  XOR2HSV0 U60133 ( .A1(n57941), .A2(n57940), .Z(n57942) );
  XOR3HSV2 U60134 ( .A1(n57944), .A2(n57943), .A3(n57942), .Z(n57945) );
  XNOR2HSV1 U60135 ( .A1(n57946), .A2(n57945), .ZN(n57947) );
  XNOR2HSV1 U60136 ( .A1(n57948), .A2(n57947), .ZN(n57950) );
  NAND2HSV0 U60137 ( .A1(n57985), .A2(n58298), .ZN(n57949) );
  XNOR2HSV1 U60138 ( .A1(n57950), .A2(n57949), .ZN(n57954) );
  NAND2HSV0 U60139 ( .A1(n57984), .A2(n58030), .ZN(n57953) );
  CLKNAND2HSV0 U60140 ( .A1(n58060), .A2(n57951), .ZN(n57952) );
  XOR3HSV2 U60141 ( .A1(n57954), .A2(n57953), .A3(n57952), .Z(n57957) );
  CLKNAND2HSV1 U60142 ( .A1(n58096), .A2(n58036), .ZN(n57956) );
  NAND2HSV0 U60143 ( .A1(n59935), .A2(\pe4/got [6]), .ZN(n57955) );
  XOR3HSV2 U60144 ( .A1(n57957), .A2(n57956), .A3(n57955), .Z(n57958) );
  XNOR2HSV1 U60145 ( .A1(n57959), .A2(n57958), .ZN(n57963) );
  CLKNAND2HSV0 U60146 ( .A1(n47841), .A2(\pe4/got [10]), .ZN(n57962) );
  CLKNAND2HSV1 U60147 ( .A1(n57960), .A2(n58041), .ZN(n57961) );
  XOR3HSV2 U60148 ( .A1(n57963), .A2(n57962), .A3(n57961), .Z(n57965) );
  CLKNAND2HSV1 U60149 ( .A1(n58103), .A2(n58153), .ZN(n57964) );
  XNOR2HSV1 U60150 ( .A1(n57965), .A2(n57964), .ZN(n57967) );
  CLKNAND2HSV0 U60151 ( .A1(n58185), .A2(n58110), .ZN(n57966) );
  XNOR2HSV1 U60152 ( .A1(n57967), .A2(n57966), .ZN(n57968) );
  XNOR2HSV1 U60153 ( .A1(n57969), .A2(n57968), .ZN(n57973) );
  CLKNAND2HSV1 U60154 ( .A1(n58048), .A2(n58052), .ZN(n57972) );
  CLKNAND2HSV0 U60155 ( .A1(n57970), .A2(n57982), .ZN(n57971) );
  XOR3HSV2 U60156 ( .A1(n57973), .A2(n57972), .A3(n57971), .Z(n57976) );
  CLKNAND2HSV1 U60157 ( .A1(n58207), .A2(n57974), .ZN(n57975) );
  XNOR2HSV1 U60158 ( .A1(n57976), .A2(n57975), .ZN(n57977) );
  XNOR2HSV1 U60159 ( .A1(n57978), .A2(n57977), .ZN(n57981) );
  XOR3HSV2 U60160 ( .A1(n57981), .A2(n57980), .A3(n57979), .Z(\pe4/poht [13])
         );
  NAND2HSV2 U60161 ( .A1(n50318), .A2(n57982), .ZN(n58056) );
  CLKNAND2HSV0 U60162 ( .A1(n57983), .A2(\pe4/got [11]), .ZN(n58047) );
  CLKNAND2HSV0 U60163 ( .A1(n58154), .A2(n58184), .ZN(n58035) );
  NAND2HSV0 U60164 ( .A1(n57984), .A2(n58314), .ZN(n58026) );
  NAND2HSV0 U60165 ( .A1(n57547), .A2(n58282), .ZN(n58024) );
  NAND2HSV0 U60166 ( .A1(n58070), .A2(n57986), .ZN(n57987) );
  XOR2HSV0 U60167 ( .A1(n57988), .A2(n57987), .Z(n58002) );
  NAND2HSV0 U60168 ( .A1(n57234), .A2(\pe4/bq[2] ), .ZN(n57990) );
  NAND2HSV0 U60169 ( .A1(n58198), .A2(\pe4/bq[11] ), .ZN(n57989) );
  XOR2HSV0 U60170 ( .A1(n57990), .A2(n57989), .Z(n57992) );
  XNOR2HSV1 U60171 ( .A1(n57992), .A2(n57991), .ZN(n58001) );
  NAND2HSV0 U60172 ( .A1(n57993), .A2(n58116), .ZN(n57995) );
  NAND2HSV0 U60173 ( .A1(n57230), .A2(n58069), .ZN(n57994) );
  XOR2HSV0 U60174 ( .A1(n57995), .A2(n57994), .Z(n57999) );
  NAND2HSV0 U60175 ( .A1(n59831), .A2(n58127), .ZN(n57997) );
  NAND2HSV0 U60176 ( .A1(\pe4/aot [10]), .A2(n35184), .ZN(n57996) );
  XOR2HSV0 U60177 ( .A1(n57997), .A2(n57996), .Z(n57998) );
  XOR2HSV0 U60178 ( .A1(n57999), .A2(n57998), .Z(n58000) );
  XOR3HSV2 U60179 ( .A1(n58002), .A2(n58001), .A3(n58000), .Z(n58022) );
  NAND2HSV0 U60180 ( .A1(\pe4/aot [14]), .A2(n58156), .ZN(n58005) );
  NAND2HSV0 U60181 ( .A1(n59683), .A2(n58003), .ZN(n58004) );
  XOR2HSV0 U60182 ( .A1(n58005), .A2(n58004), .Z(n58009) );
  NAND2HSV0 U60183 ( .A1(\pe4/aot [2]), .A2(n49943), .ZN(n58007) );
  NAND2HSV0 U60184 ( .A1(n58283), .A2(n57348), .ZN(n58006) );
  XOR2HSV0 U60185 ( .A1(n58007), .A2(n58006), .Z(n58008) );
  XOR2HSV0 U60186 ( .A1(n58009), .A2(n58008), .Z(n58020) );
  NAND2HSV0 U60187 ( .A1(\pe4/aot [9]), .A2(n57798), .ZN(n58012) );
  NAND2HSV0 U60188 ( .A1(n59857), .A2(n58010), .ZN(n58011) );
  XOR2HSV0 U60189 ( .A1(n58012), .A2(n58011), .Z(n58018) );
  NOR2HSV0 U60190 ( .A1(n35175), .A2(n58013), .ZN(n58016) );
  NAND2HSV0 U60191 ( .A1(n59343), .A2(n58014), .ZN(n58015) );
  XOR2HSV0 U60192 ( .A1(n58016), .A2(n58015), .Z(n58017) );
  XOR2HSV0 U60193 ( .A1(n58018), .A2(n58017), .Z(n58019) );
  XOR2HSV0 U60194 ( .A1(n58020), .A2(n58019), .Z(n58021) );
  XNOR2HSV1 U60195 ( .A1(n58022), .A2(n58021), .ZN(n58023) );
  XNOR2HSV1 U60196 ( .A1(n58024), .A2(n58023), .ZN(n58025) );
  XNOR2HSV1 U60197 ( .A1(n58026), .A2(n58025), .ZN(n58028) );
  CLKNAND2HSV0 U60198 ( .A1(n58060), .A2(n58298), .ZN(n58027) );
  XNOR2HSV1 U60199 ( .A1(n58028), .A2(n58027), .ZN(n58033) );
  NAND2HSV2 U60200 ( .A1(n58029), .A2(n57951), .ZN(n58032) );
  CLKNAND2HSV0 U60201 ( .A1(n58097), .A2(n58030), .ZN(n58031) );
  XOR3HSV2 U60202 ( .A1(n58033), .A2(n58032), .A3(n58031), .Z(n58034) );
  XNOR2HSV1 U60203 ( .A1(n58035), .A2(n58034), .ZN(n58040) );
  NAND2HSV2 U60204 ( .A1(n58183), .A2(n58111), .ZN(n58039) );
  NAND2HSV0 U60205 ( .A1(n58037), .A2(n58036), .ZN(n58038) );
  XOR3HSV2 U60206 ( .A1(n58040), .A2(n58039), .A3(n58038), .Z(n58043) );
  CLKNAND2HSV1 U60207 ( .A1(n57889), .A2(n58041), .ZN(n58042) );
  XNOR2HSV1 U60208 ( .A1(n58043), .A2(n58042), .ZN(n58045) );
  CLKNAND2HSV0 U60209 ( .A1(n57310), .A2(n59663), .ZN(n58044) );
  XNOR2HSV1 U60210 ( .A1(n58045), .A2(n58044), .ZN(n58046) );
  XNOR2HSV1 U60211 ( .A1(n58047), .A2(n58046), .ZN(n58051) );
  CLKNAND2HSV1 U60212 ( .A1(n58048), .A2(n58110), .ZN(n58050) );
  NAND2HSV0 U60213 ( .A1(n58272), .A2(n35400), .ZN(n58049) );
  XOR3HSV2 U60214 ( .A1(n58051), .A2(n58050), .A3(n58049), .Z(n58054) );
  CLKNAND2HSV1 U60215 ( .A1(n58207), .A2(n58052), .ZN(n58053) );
  XNOR2HSV1 U60216 ( .A1(n58054), .A2(n58053), .ZN(n58055) );
  XNOR2HSV1 U60217 ( .A1(n58056), .A2(n58055), .ZN(n58059) );
  NOR2HSV3 U60218 ( .A1(n29752), .A2(n50294), .ZN(n58058) );
  NOR2HSV2 U60219 ( .A1(n26761), .A2(n47861), .ZN(n58057) );
  XOR3HSV2 U60220 ( .A1(n58059), .A2(n58058), .A3(n58057), .Z(\pe4/poht [15])
         );
  NAND2HSV0 U60221 ( .A1(n58060), .A2(n58282), .ZN(n58095) );
  NAND2HSV0 U60222 ( .A1(\pe4/aot [14]), .A2(\pe4/bq[2] ), .ZN(n58062) );
  NAND2HSV0 U60223 ( .A1(n58198), .A2(n58113), .ZN(n58061) );
  XOR2HSV0 U60224 ( .A1(n58062), .A2(n58061), .Z(n58066) );
  NAND2HSV0 U60225 ( .A1(n59857), .A2(n58301), .ZN(n58064) );
  NAND2HSV0 U60226 ( .A1(n57683), .A2(n58265), .ZN(n58063) );
  XOR2HSV0 U60227 ( .A1(n58064), .A2(n58063), .Z(n58065) );
  XOR2HSV0 U60228 ( .A1(n58066), .A2(n58065), .Z(n58076) );
  NAND2HSV0 U60229 ( .A1(n58283), .A2(n58127), .ZN(n58068) );
  NAND2HSV0 U60230 ( .A1(n59953), .A2(n58322), .ZN(n58067) );
  XOR2HSV0 U60231 ( .A1(n58068), .A2(n58067), .Z(n58074) );
  CLKNAND2HSV1 U60232 ( .A1(\pe4/aot [2]), .A2(n58069), .ZN(n58072) );
  CLKNAND2HSV0 U60233 ( .A1(n58070), .A2(\pe4/bq[10] ), .ZN(n58071) );
  XOR2HSV0 U60234 ( .A1(n58072), .A2(n58071), .Z(n58073) );
  XOR2HSV0 U60235 ( .A1(n58074), .A2(n58073), .Z(n58075) );
  XOR2HSV0 U60236 ( .A1(n58076), .A2(n58075), .Z(n58093) );
  CLKNAND2HSV0 U60237 ( .A1(\pe4/aot [12]), .A2(n57595), .ZN(n58079) );
  NAND2HSV0 U60238 ( .A1(n57230), .A2(n58077), .ZN(n58078) );
  XOR2HSV0 U60239 ( .A1(n58079), .A2(n58078), .Z(n58083) );
  NAND2HSV0 U60240 ( .A1(n59831), .A2(\pe4/bq[11] ), .ZN(n58081) );
  NAND2HSV0 U60241 ( .A1(n59683), .A2(n58155), .ZN(n58080) );
  XOR2HSV0 U60242 ( .A1(n58081), .A2(n58080), .Z(n58082) );
  XOR2HSV0 U60243 ( .A1(n58083), .A2(n58082), .Z(n58091) );
  NAND2HSV0 U60244 ( .A1(n57692), .A2(n58084), .ZN(n58086) );
  NAND2HSV0 U60245 ( .A1(\pe4/aot [9]), .A2(n58197), .ZN(n58085) );
  XOR2HSV0 U60246 ( .A1(n58086), .A2(n58085), .Z(n58089) );
  CLKNAND2HSV1 U60247 ( .A1(n58087), .A2(n58130), .ZN(n58088) );
  XNOR2HSV1 U60248 ( .A1(n58089), .A2(n58088), .ZN(n58090) );
  XNOR2HSV1 U60249 ( .A1(n58091), .A2(n58090), .ZN(n58092) );
  XNOR2HSV1 U60250 ( .A1(n58093), .A2(n58092), .ZN(n58094) );
  XNOR2HSV1 U60251 ( .A1(n58095), .A2(n58094), .ZN(n58100) );
  NAND2HSV2 U60252 ( .A1(n58096), .A2(n58298), .ZN(n58099) );
  CLKNAND2HSV1 U60253 ( .A1(n58097), .A2(n58314), .ZN(n58098) );
  XOR3HSV2 U60254 ( .A1(n58100), .A2(n58099), .A3(n58098), .Z(n58101) );
  XNOR2HSV1 U60255 ( .A1(n58106), .A2(n58105), .ZN(n58109) );
  NOR2HSV2 U60256 ( .A1(n29774), .A2(n50042), .ZN(n58108) );
  NOR2HSV2 U60257 ( .A1(n26761), .A2(n50212), .ZN(n58107) );
  XOR3HSV2 U60258 ( .A1(n58109), .A2(n58108), .A3(n58107), .Z(\pe4/poht [17])
         );
  CLKNAND2HSV1 U60259 ( .A1(n26417), .A2(n58110), .ZN(n58149) );
  NAND2HSV0 U60260 ( .A1(n59837), .A2(n58111), .ZN(n58139) );
  NAND2HSV0 U60261 ( .A1(n58070), .A2(n58113), .ZN(n58115) );
  NAND2HSV0 U60262 ( .A1(n59683), .A2(n58156), .ZN(n58114) );
  XOR2HSV0 U60263 ( .A1(n58115), .A2(n58114), .Z(n58120) );
  NAND2HSV0 U60264 ( .A1(n58306), .A2(n58116), .ZN(n58118) );
  NAND2HSV0 U60265 ( .A1(n57993), .A2(n58197), .ZN(n58117) );
  XOR2HSV0 U60266 ( .A1(n58118), .A2(n58117), .Z(n58119) );
  CLKNAND2HSV0 U60267 ( .A1(\pe4/aot [10]), .A2(n58155), .ZN(n58122) );
  NAND2HSV0 U60268 ( .A1(\pe4/aot [9]), .A2(n58195), .ZN(n58121) );
  NAND2HSV0 U60269 ( .A1(n59857), .A2(\pe4/bq[2] ), .ZN(n58124) );
  NAND2HSV0 U60270 ( .A1(\pe4/aot [14]), .A2(n58322), .ZN(n58123) );
  XOR2HSV0 U60271 ( .A1(n58124), .A2(n58123), .Z(n58125) );
  CLKNAND2HSV0 U60272 ( .A1(n57692), .A2(n58126), .ZN(n58129) );
  NAND2HSV0 U60273 ( .A1(\pe4/aot [2]), .A2(n58127), .ZN(n58128) );
  XOR2HSV0 U60274 ( .A1(n58129), .A2(n58128), .Z(n58134) );
  CLKNAND2HSV1 U60275 ( .A1(n59632), .A2(n58130), .ZN(n58132) );
  NAND2HSV0 U60276 ( .A1(\pe4/aot [12]), .A2(n58301), .ZN(n58131) );
  XOR2HSV0 U60277 ( .A1(n58132), .A2(n58131), .Z(n58133) );
  NAND2HSV0 U60278 ( .A1(n58199), .A2(\pe4/bq[11] ), .ZN(n58135) );
  XNOR2HSV1 U60279 ( .A1(n58139), .A2(n58138), .ZN(n58144) );
  CLKNAND2HSV1 U60280 ( .A1(n58141), .A2(n58140), .ZN(n58143) );
  CLKNAND2HSV0 U60281 ( .A1(n59663), .A2(n59348), .ZN(n58142) );
  XOR3HSV2 U60282 ( .A1(n58144), .A2(n58143), .A3(n58142), .Z(n58147) );
  CLKNAND2HSV0 U60283 ( .A1(n26692), .A2(n58153), .ZN(n58146) );
  XNOR2HSV1 U60284 ( .A1(n58147), .A2(n58146), .ZN(n58148) );
  XNOR2HSV1 U60285 ( .A1(n58149), .A2(n58148), .ZN(n58152) );
  NOR2HSV2 U60286 ( .A1(n29774), .A2(n58189), .ZN(n58151) );
  NOR2HSV2 U60287 ( .A1(n26761), .A2(n50042), .ZN(n58150) );
  XOR3HSV2 U60288 ( .A1(n58152), .A2(n58151), .A3(n58150), .Z(\pe4/poht [18])
         );
  NAND2HSV0 U60289 ( .A1(n59665), .A2(n58300), .ZN(n58182) );
  NAND2HSV0 U60290 ( .A1(\pe4/aot [9]), .A2(n58155), .ZN(n58158) );
  NAND2HSV0 U60291 ( .A1(\pe4/aot [10]), .A2(n58156), .ZN(n58157) );
  XOR2HSV0 U60292 ( .A1(n58158), .A2(n58157), .Z(n58162) );
  CLKNAND2HSV0 U60293 ( .A1(n58230), .A2(n58127), .ZN(n58160) );
  NAND2HSV0 U60294 ( .A1(n58223), .A2(n58113), .ZN(n58159) );
  XOR2HSV0 U60295 ( .A1(n58160), .A2(n58159), .Z(n58161) );
  XOR2HSV0 U60296 ( .A1(n58162), .A2(n58161), .Z(n58171) );
  NAND2HSV0 U60297 ( .A1(n58163), .A2(n57241), .ZN(n58165) );
  NAND2HSV0 U60298 ( .A1(n59683), .A2(n58196), .ZN(n58164) );
  XOR2HSV0 U60299 ( .A1(n58165), .A2(n58164), .Z(n58169) );
  NAND2HSV0 U60300 ( .A1(n59954), .A2(\pe4/bq[11] ), .ZN(n58167) );
  NAND2HSV0 U60301 ( .A1(n59343), .A2(\pe4/bq[2] ), .ZN(n58166) );
  XOR2HSV0 U60302 ( .A1(n58167), .A2(n58166), .Z(n58168) );
  XOR2HSV0 U60303 ( .A1(n58169), .A2(n58168), .Z(n58170) );
  XOR2HSV0 U60304 ( .A1(n58171), .A2(n58170), .Z(n58181) );
  CLKNAND2HSV1 U60305 ( .A1(\pe4/aot [2]), .A2(n58077), .ZN(n58173) );
  NAND2HSV0 U60306 ( .A1(n57993), .A2(n58265), .ZN(n58172) );
  XOR2HSV0 U60307 ( .A1(n58173), .A2(n58172), .Z(n58178) );
  NOR2HSV0 U60308 ( .A1(n58174), .A2(n48028), .ZN(n58176) );
  NAND2HSV0 U60309 ( .A1(n59632), .A2(n58197), .ZN(n58175) );
  XOR2HSV0 U60310 ( .A1(n58176), .A2(n58175), .Z(n58177) );
  XOR3HSV2 U60311 ( .A1(n58179), .A2(n58178), .A3(n58177), .Z(n58180) );
  XNOR2HSV1 U60312 ( .A1(n58188), .A2(n58187), .ZN(n58192) );
  NOR2HSV2 U60313 ( .A1(n26761), .A2(n58189), .ZN(n58190) );
  XOR3HSV2 U60314 ( .A1(n58192), .A2(n58191), .A3(n58190), .Z(\pe4/poht [19])
         );
  CLKNAND2HSV1 U60315 ( .A1(n58217), .A2(n58314), .ZN(n58203) );
  CLKNAND2HSV1 U60316 ( .A1(n58193), .A2(n58300), .ZN(n58201) );
  XNOR2HSV1 U60317 ( .A1(n58201), .A2(n58200), .ZN(n58202) );
  NAND2HSV0 U60318 ( .A1(n58272), .A2(n58298), .ZN(n58204) );
  XNOR2HSV1 U60319 ( .A1(n58205), .A2(n58204), .ZN(n58209) );
  CLKNAND2HSV0 U60320 ( .A1(n58207), .A2(n58206), .ZN(n58208) );
  XOR2HSV0 U60321 ( .A1(n58209), .A2(n58208), .Z(n58210) );
  XNOR2HSV1 U60322 ( .A1(n58211), .A2(n58210), .ZN(n58215) );
  XOR3HSV2 U60323 ( .A1(n58215), .A2(n58214), .A3(n58213), .Z(\pe4/poht [25])
         );
  CLKNAND2HSV1 U60324 ( .A1(n58217), .A2(n58258), .ZN(n58245) );
  CLKNAND2HSV1 U60325 ( .A1(n58218), .A2(\pe4/got [3]), .ZN(n58243) );
  CLKNAND2HSV0 U60326 ( .A1(n35033), .A2(n58314), .ZN(n58241) );
  CLKNAND2HSV1 U60327 ( .A1(n58220), .A2(n58219), .ZN(n58239) );
  NAND2HSV0 U60328 ( .A1(\pe4/aot [2]), .A2(n58130), .ZN(n58221) );
  XOR2HSV0 U60329 ( .A1(n58222), .A2(n58221), .Z(n58237) );
  NAND2HSV0 U60330 ( .A1(n57993), .A2(\pe4/bq[2] ), .ZN(n58225) );
  CLKNAND2HSV0 U60331 ( .A1(n58223), .A2(n58155), .ZN(n58224) );
  XOR2HSV0 U60332 ( .A1(n58225), .A2(n58224), .Z(n58227) );
  XNOR2HSV1 U60333 ( .A1(n58227), .A2(n58226), .ZN(n58236) );
  NAND2HSV0 U60334 ( .A1(n58070), .A2(n58156), .ZN(n58229) );
  NAND2HSV0 U60335 ( .A1(n59954), .A2(n58003), .ZN(n58228) );
  XOR2HSV0 U60336 ( .A1(n58229), .A2(n58228), .Z(n58234) );
  NOR2HSV1 U60337 ( .A1(n35042), .A2(n57010), .ZN(n58232) );
  CLKNAND2HSV0 U60338 ( .A1(n58230), .A2(n58113), .ZN(n58231) );
  XOR2HSV0 U60339 ( .A1(n58232), .A2(n58231), .Z(n58233) );
  XOR2HSV0 U60340 ( .A1(n58234), .A2(n58233), .Z(n58235) );
  XOR3HSV2 U60341 ( .A1(n58237), .A2(n58236), .A3(n58235), .Z(n58238) );
  XNOR2HSV1 U60342 ( .A1(n58239), .A2(n58238), .ZN(n58240) );
  XNOR2HSV1 U60343 ( .A1(n58241), .A2(n58240), .ZN(n58242) );
  XNOR2HSV1 U60344 ( .A1(n58243), .A2(n58242), .ZN(n58244) );
  NAND2HSV0 U60345 ( .A1(n58246), .A2(n50199), .ZN(n58247) );
  XNOR2HSV1 U60346 ( .A1(n58248), .A2(n58247), .ZN(n58250) );
  XOR2HSV0 U60347 ( .A1(n58250), .A2(n58249), .Z(n58251) );
  XNOR2HSV1 U60348 ( .A1(n58252), .A2(n58251), .ZN(n58257) );
  NOR2HSV2 U60349 ( .A1(n29774), .A2(n58253), .ZN(n58256) );
  CLKNAND2HSV1 U60350 ( .A1(n58254), .A2(n58140), .ZN(n58255) );
  XOR3HSV2 U60351 ( .A1(n58257), .A2(n58256), .A3(n58255), .Z(\pe4/poht [23])
         );
  CLKNAND2HSV1 U60352 ( .A1(n58141), .A2(n58282), .ZN(n58271) );
  NAND2HSV0 U60353 ( .A1(\pe4/aot [2]), .A2(n58010), .ZN(n58260) );
  CLKNAND2HSV0 U60354 ( .A1(\pe4/aot [5]), .A2(\pe4/bq[2] ), .ZN(n58259) );
  XOR2HSV0 U60355 ( .A1(n58260), .A2(n58259), .Z(n58264) );
  CLKNAND2HSV0 U60356 ( .A1(n58283), .A2(n57498), .ZN(n58262) );
  NAND2HSV0 U60357 ( .A1(n59352), .A2(n57241), .ZN(n58261) );
  XOR2HSV0 U60358 ( .A1(n58262), .A2(n58261), .Z(n58263) );
  XOR2HSV0 U60359 ( .A1(n58264), .A2(n58263), .Z(n58269) );
  NAND2HSV0 U60360 ( .A1(\pe4/aot [1]), .A2(n58265), .ZN(n58266) );
  XOR2HSV0 U60361 ( .A1(n58267), .A2(n58266), .Z(n58268) );
  XNOR2HSV1 U60362 ( .A1(n58269), .A2(n58268), .ZN(n58270) );
  XOR2HSV0 U60363 ( .A1(n58271), .A2(n58270), .Z(n58274) );
  NAND2HSV0 U60364 ( .A1(n58272), .A2(n58314), .ZN(n58273) );
  NAND2HSV0 U60365 ( .A1(n58207), .A2(n58298), .ZN(n58275) );
  XNOR2HSV1 U60366 ( .A1(n58278), .A2(n58277), .ZN(n58281) );
  NOR2HSV2 U60367 ( .A1(n58212), .A2(n50095), .ZN(n58280) );
  NOR2HSV2 U60368 ( .A1(n26761), .A2(n50214), .ZN(n58279) );
  XOR3HSV2 U60369 ( .A1(n58281), .A2(n58280), .A3(n58279), .Z(\pe4/poht [26])
         );
  NAND2HSV0 U60370 ( .A1(n58207), .A2(n58282), .ZN(n58291) );
  CLKNAND2HSV1 U60371 ( .A1(n58283), .A2(\pe4/bq[2] ), .ZN(n58285) );
  NAND2HSV0 U60372 ( .A1(\pe4/aot [1]), .A2(n57498), .ZN(n58284) );
  XOR2HSV0 U60373 ( .A1(n58285), .A2(n58284), .Z(n58289) );
  CLKNAND2HSV0 U60374 ( .A1(\pe4/aot [2]), .A2(n58301), .ZN(n58286) );
  XOR2HSV0 U60375 ( .A1(n58287), .A2(n58286), .Z(n58288) );
  XOR2HSV0 U60376 ( .A1(n58289), .A2(n58288), .Z(n58290) );
  XNOR2HSV1 U60377 ( .A1(n58291), .A2(n58290), .ZN(n58292) );
  XNOR2HSV1 U60378 ( .A1(n58293), .A2(n58292), .ZN(n58297) );
  XOR3HSV2 U60379 ( .A1(n58297), .A2(n58296), .A3(n58295), .Z(\pe4/poht [28])
         );
  CLKNAND2HSV1 U60380 ( .A1(n58299), .A2(n58298), .ZN(n58318) );
  CLKNAND2HSV1 U60381 ( .A1(n59348), .A2(n58300), .ZN(n58313) );
  CLKNAND2HSV0 U60382 ( .A1(\pe4/aot [2]), .A2(n57595), .ZN(n58303) );
  CLKNAND2HSV0 U60383 ( .A1(n58283), .A2(n58301), .ZN(n58302) );
  XOR2HSV0 U60384 ( .A1(n58303), .A2(n58302), .Z(n58305) );
  XNOR2HSV1 U60385 ( .A1(n58305), .A2(n58304), .ZN(n58311) );
  CLKNAND2HSV1 U60386 ( .A1(n58306), .A2(n58322), .ZN(n58309) );
  CLKNAND2HSV0 U60387 ( .A1(n58307), .A2(\pe4/bq[2] ), .ZN(n58308) );
  XOR2HSV0 U60388 ( .A1(n58309), .A2(n58308), .Z(n58310) );
  XNOR2HSV1 U60389 ( .A1(n58311), .A2(n58310), .ZN(n58312) );
  XNOR2HSV1 U60390 ( .A1(n58313), .A2(n58312), .ZN(n58316) );
  CLKNAND2HSV1 U60391 ( .A1(n26516), .A2(n58314), .ZN(n58315) );
  XOR2HSV0 U60392 ( .A1(n58316), .A2(n58315), .Z(n58317) );
  XNOR2HSV1 U60393 ( .A1(n58318), .A2(n58317), .ZN(n58321) );
  XOR3HSV2 U60394 ( .A1(n58321), .A2(n58320), .A3(n58319), .Z(\pe4/poht [27])
         );
  NAND2HSV2 U60395 ( .A1(n58230), .A2(\pe4/bq[2] ), .ZN(n58324) );
  CLKNAND2HSV1 U60396 ( .A1(\pe4/aot [2]), .A2(n58322), .ZN(n58323) );
  XOR2HSV0 U60397 ( .A1(n58324), .A2(n58323), .Z(n58328) );
  NOR2HSV2 U60398 ( .A1(n29774), .A2(n49967), .ZN(n58327) );
  NOR2HSV2 U60399 ( .A1(n26761), .A2(n58325), .ZN(n58326) );
  XOR3HSV2 U60400 ( .A1(n58328), .A2(n58327), .A3(n58326), .Z(\pe4/poht [30])
         );
  NAND2HSV2 U60401 ( .A1(n58360), .A2(\pe6/aot [1]), .ZN(n58330) );
  NAND2HSV0 U60402 ( .A1(n58336), .A2(n58579), .ZN(n58329) );
  XOR2HSV0 U60403 ( .A1(n58330), .A2(n58329), .Z(n58334) );
  CLKNAND2HSV1 U60404 ( .A1(n25849), .A2(\pe6/got [1]), .ZN(n58333) );
  NAND2HSV2 U60405 ( .A1(n59023), .A2(n58331), .ZN(n58332) );
  XOR3HSV2 U60406 ( .A1(n58334), .A2(n58333), .A3(n58332), .Z(\pe6/poht [30])
         );
  CLKNAND2HSV1 U60407 ( .A1(n58724), .A2(n59169), .ZN(n58347) );
  CLKNHSV0 U60408 ( .I(n58817), .ZN(n58335) );
  INAND2HSV2 U60409 ( .A1(n58335), .B1(n49181), .ZN(n58345) );
  NAND2HSV0 U60410 ( .A1(n58336), .A2(n58459), .ZN(n58338) );
  CLKNAND2HSV0 U60411 ( .A1(n58360), .A2(n58353), .ZN(n58337) );
  XOR2HSV0 U60412 ( .A1(n58338), .A2(n58337), .Z(n58343) );
  CLKNAND2HSV0 U60413 ( .A1(n58339), .A2(n58579), .ZN(n58340) );
  XOR2HSV0 U60414 ( .A1(n58341), .A2(n58340), .Z(n58342) );
  XOR2HSV0 U60415 ( .A1(n58343), .A2(n58342), .Z(n58344) );
  XNOR2HSV1 U60416 ( .A1(n58345), .A2(n58344), .ZN(n58346) );
  XNOR2HSV1 U60417 ( .A1(n58347), .A2(n58346), .ZN(n58351) );
  CLKNHSV0 U60418 ( .I(n58724), .ZN(n58352) );
  INAND2HSV0 U60419 ( .A1(n58352), .B1(n58656), .ZN(n58368) );
  INHSV2 U60420 ( .I(n58447), .ZN(n58809) );
  CLKNAND2HSV1 U60421 ( .A1(n58809), .A2(\pe6/got [1]), .ZN(n58366) );
  INHSV2 U60422 ( .I(n49327), .ZN(n58408) );
  CLKNAND2HSV1 U60423 ( .A1(n58408), .A2(n58353), .ZN(n58355) );
  CLKNAND2HSV0 U60424 ( .A1(n59062), .A2(n58579), .ZN(n58354) );
  XOR2HSV0 U60425 ( .A1(n58355), .A2(n58354), .Z(n58358) );
  CLKNAND2HSV0 U60426 ( .A1(n58356), .A2(\pe6/aot [1]), .ZN(n58357) );
  XNOR2HSV1 U60427 ( .A1(n58358), .A2(n58357), .ZN(n58364) );
  NOR2HSV2 U60428 ( .A1(n48887), .A2(n58359), .ZN(n58362) );
  CLKNAND2HSV0 U60429 ( .A1(n58360), .A2(n58459), .ZN(n58361) );
  XOR2HSV0 U60430 ( .A1(n58362), .A2(n58361), .Z(n58363) );
  XNOR2HSV1 U60431 ( .A1(n58364), .A2(n58363), .ZN(n58365) );
  XNOR2HSV1 U60432 ( .A1(n58366), .A2(n58365), .ZN(n58367) );
  XOR2HSV0 U60433 ( .A1(n58368), .A2(n58367), .Z(n58371) );
  NAND2HSV0 U60434 ( .A1(n58369), .A2(n58423), .ZN(n58370) );
  XOR2HSV0 U60435 ( .A1(n58371), .A2(n58370), .Z(n58375) );
  XOR3HSV2 U60436 ( .A1(n58375), .A2(n58374), .A3(n58373), .Z(\pe6/poht [27])
         );
  CLKNAND2HSV1 U60437 ( .A1(n58405), .A2(\pe6/aot [1]), .ZN(n58377) );
  CLKNAND2HSV0 U60438 ( .A1(n58408), .A2(n58459), .ZN(n58376) );
  NAND2HSV2 U60439 ( .A1(n59041), .A2(n58378), .ZN(n58380) );
  CLKNAND2HSV1 U60440 ( .A1(n59277), .A2(\pe6/aot [6]), .ZN(n58379) );
  CLKNAND2HSV1 U60441 ( .A1(n58460), .A2(\pe6/aot [1]), .ZN(n58387) );
  CLKNAND2HSV0 U60442 ( .A1(n58408), .A2(n49847), .ZN(n58386) );
  XOR2HSV0 U60443 ( .A1(n58387), .A2(n58386), .Z(n58391) );
  CLKNAND2HSV1 U60444 ( .A1(n58452), .A2(n58404), .ZN(n58389) );
  NAND2HSV0 U60445 ( .A1(n58405), .A2(n58579), .ZN(n58388) );
  XOR2HSV0 U60446 ( .A1(n58389), .A2(n58388), .Z(n58390) );
  XOR2HSV0 U60447 ( .A1(n58391), .A2(n58390), .Z(n58397) );
  NOR2HSV1 U60448 ( .A1(n48887), .A2(n58392), .ZN(n58394) );
  CLKNAND2HSV1 U60449 ( .A1(n58360), .A2(n59266), .ZN(n58393) );
  XOR2HSV0 U60450 ( .A1(n58394), .A2(n58393), .Z(n58396) );
  CLKNAND2HSV0 U60451 ( .A1(n58399), .A2(n58575), .ZN(n58432) );
  CLKNAND2HSV1 U60452 ( .A1(n58576), .A2(n58400), .ZN(n58430) );
  CLKNAND2HSV0 U60453 ( .A1(n58385), .A2(n58401), .ZN(n58428) );
  NAND2HSV0 U60454 ( .A1(n58402), .A2(n58816), .ZN(n58426) );
  NAND2HSV0 U60455 ( .A1(n58480), .A2(n58403), .ZN(n58422) );
  CLKNAND2HSV1 U60456 ( .A1(n58452), .A2(n58459), .ZN(n58407) );
  CLKNAND2HSV0 U60457 ( .A1(n58405), .A2(n58404), .ZN(n58406) );
  XOR2HSV0 U60458 ( .A1(n58407), .A2(n58406), .Z(n58412) );
  CLKNAND2HSV1 U60459 ( .A1(\pe6/bq[4] ), .A2(n49847), .ZN(n58410) );
  CLKNAND2HSV0 U60460 ( .A1(n58408), .A2(\pe6/aot [6]), .ZN(n58409) );
  XOR2HSV0 U60461 ( .A1(n58410), .A2(n58409), .Z(n58411) );
  XOR2HSV0 U60462 ( .A1(n58412), .A2(n58411), .Z(n58420) );
  CLKNAND2HSV1 U60463 ( .A1(n58619), .A2(\pe6/aot [1]), .ZN(n58414) );
  NAND2HSV0 U60464 ( .A1(n58460), .A2(n58579), .ZN(n58413) );
  XOR2HSV0 U60465 ( .A1(n58414), .A2(n58413), .Z(n58418) );
  NOR2HSV1 U60466 ( .A1(n48887), .A2(n58483), .ZN(n58416) );
  CLKNAND2HSV0 U60467 ( .A1(n58360), .A2(\pe6/aot [7]), .ZN(n58415) );
  XOR2HSV0 U60468 ( .A1(n58416), .A2(n58415), .Z(n58417) );
  XOR2HSV0 U60469 ( .A1(n58418), .A2(n58417), .Z(n58419) );
  XOR2HSV0 U60470 ( .A1(n58420), .A2(n58419), .Z(n58421) );
  XNOR2HSV1 U60471 ( .A1(n58422), .A2(n58421), .ZN(n58425) );
  NAND2HSV0 U60472 ( .A1(n59528), .A2(n58423), .ZN(n58424) );
  XOR3HSV2 U60473 ( .A1(n58426), .A2(n58425), .A3(n58424), .Z(n58427) );
  XNOR2HSV1 U60474 ( .A1(n58428), .A2(n58427), .ZN(n58429) );
  XOR2HSV0 U60475 ( .A1(n58430), .A2(n58429), .Z(n58431) );
  XOR2HSV0 U60476 ( .A1(n58432), .A2(n58431), .Z(n58446) );
  CLKNAND2HSV2 U60477 ( .A1(n59021), .A2(n36109), .ZN(n58445) );
  NOR3HSV2 U60478 ( .A1(n58435), .A2(n58434), .A3(n58433), .ZN(n58436) );
  INAND2HSV2 U60479 ( .A1(n58437), .B1(n58436), .ZN(n58443) );
  NAND3HSV0 U60480 ( .A1(n58439), .A2(n58438), .A3(n59182), .ZN(n58440) );
  OAI22HSV1 U60481 ( .A1(n58443), .A2(n25886), .B1(n58441), .B2(n58440), .ZN(
        n58444) );
  XOR3HSV2 U60482 ( .A1(n58446), .A2(n58445), .A3(n58444), .Z(\pe6/poht [24])
         );
  NAND2HSV0 U60483 ( .A1(n58448), .A2(n58817), .ZN(n58473) );
  CLKNAND2HSV1 U60484 ( .A1(n58496), .A2(n58449), .ZN(n58450) );
  XOR2HSV0 U60485 ( .A1(n58451), .A2(n58450), .Z(n58471) );
  CLKNAND2HSV0 U60486 ( .A1(n58452), .A2(\pe6/aot [6]), .ZN(n58454) );
  CLKNAND2HSV1 U60487 ( .A1(n58360), .A2(n58495), .ZN(n58453) );
  XOR2HSV0 U60488 ( .A1(n58454), .A2(n58453), .Z(n58458) );
  NOR2HSV2 U60489 ( .A1(n46147), .A2(n58359), .ZN(n58456) );
  CLKNAND2HSV0 U60490 ( .A1(n58962), .A2(\pe6/aot [1]), .ZN(n58455) );
  XOR2HSV0 U60491 ( .A1(n58456), .A2(n58455), .Z(n58457) );
  XNOR2HSV1 U60492 ( .A1(n58458), .A2(n58457), .ZN(n58470) );
  CLKNAND2HSV0 U60493 ( .A1(n58460), .A2(n58459), .ZN(n58462) );
  CLKNAND2HSV0 U60494 ( .A1(n58619), .A2(\pe6/aot [3]), .ZN(n58461) );
  XOR2HSV0 U60495 ( .A1(n58462), .A2(n58461), .Z(n58468) );
  NOR2HSV0 U60496 ( .A1(n48887), .A2(n58463), .ZN(n58466) );
  CLKNAND2HSV1 U60497 ( .A1(\pe6/bq[9] ), .A2(n58464), .ZN(n58465) );
  XOR2HSV0 U60498 ( .A1(n58466), .A2(n58465), .Z(n58467) );
  XOR2HSV0 U60499 ( .A1(n58468), .A2(n58467), .Z(n58469) );
  XOR3HSV2 U60500 ( .A1(n58471), .A2(n58470), .A3(n58469), .Z(n58472) );
  XNOR2HSV1 U60501 ( .A1(n58473), .A2(n58472), .ZN(n58475) );
  CLKNAND2HSV0 U60502 ( .A1(n58805), .A2(n59231), .ZN(n58474) );
  CLKNAND2HSV0 U60503 ( .A1(n58477), .A2(n59169), .ZN(n58522) );
  CLKNAND2HSV0 U60504 ( .A1(n59514), .A2(n58526), .ZN(n58520) );
  CLKNAND2HSV1 U60505 ( .A1(n58562), .A2(n59026), .ZN(n58518) );
  CLKNAND2HSV0 U60506 ( .A1(n58934), .A2(n58478), .ZN(n58516) );
  NAND2HSV0 U60507 ( .A1(n58480), .A2(n58479), .ZN(n58512) );
  CLKNAND2HSV1 U60508 ( .A1(n58660), .A2(n59039), .ZN(n58508) );
  CLKNAND2HSV1 U60509 ( .A1(n46825), .A2(n58817), .ZN(n58506) );
  NAND2HSV0 U60510 ( .A1(n58962), .A2(n58579), .ZN(n58482) );
  CLKNAND2HSV1 U60511 ( .A1(n58356), .A2(\pe6/aot [7]), .ZN(n58481) );
  XOR2HSV0 U60512 ( .A1(n58482), .A2(n58481), .Z(n58487) );
  NOR2HSV1 U60513 ( .A1(n48042), .A2(n58530), .ZN(n58485) );
  CLKNAND2HSV1 U60514 ( .A1(n59062), .A2(n35632), .ZN(n58484) );
  XOR2HSV0 U60515 ( .A1(n58485), .A2(n58484), .Z(n58486) );
  XOR2HSV0 U60516 ( .A1(n58487), .A2(n58486), .Z(n58494) );
  CLKNAND2HSV0 U60517 ( .A1(n59277), .A2(\pe6/aot [11]), .ZN(n58490) );
  NAND2HSV0 U60518 ( .A1(n58360), .A2(n58488), .ZN(n58489) );
  XOR2HSV0 U60519 ( .A1(n58490), .A2(n58489), .Z(n58492) );
  XNOR2HSV1 U60520 ( .A1(n58492), .A2(n58491), .ZN(n58493) );
  XNOR2HSV1 U60521 ( .A1(n58494), .A2(n58493), .ZN(n58504) );
  CLKNAND2HSV1 U60522 ( .A1(n58496), .A2(n58495), .ZN(n58498) );
  CLKNAND2HSV0 U60523 ( .A1(n35750), .A2(\pe6/aot [1]), .ZN(n58497) );
  XOR2HSV0 U60524 ( .A1(n58498), .A2(n58497), .Z(n58502) );
  CLKNAND2HSV0 U60525 ( .A1(n58628), .A2(\pe6/aot [3]), .ZN(n58500) );
  INHSV1 U60526 ( .I(n48041), .ZN(n58675) );
  CLKNAND2HSV1 U60527 ( .A1(n58675), .A2(n59250), .ZN(n58499) );
  XOR2HSV0 U60528 ( .A1(n58500), .A2(n58499), .Z(n58501) );
  XOR2HSV0 U60529 ( .A1(n58502), .A2(n58501), .Z(n58503) );
  XNOR2HSV1 U60530 ( .A1(n58504), .A2(n58503), .ZN(n58505) );
  XNOR2HSV1 U60531 ( .A1(n58506), .A2(n58505), .ZN(n58507) );
  XNOR2HSV1 U60532 ( .A1(n58508), .A2(n58507), .ZN(n58510) );
  CLKNAND2HSV0 U60533 ( .A1(n59161), .A2(n58527), .ZN(n58509) );
  XOR2HSV0 U60534 ( .A1(n58510), .A2(n58509), .Z(n58511) );
  XNOR2HSV1 U60535 ( .A1(n58512), .A2(n58511), .ZN(n58515) );
  NAND2HSV0 U60536 ( .A1(n59528), .A2(n58513), .ZN(n58514) );
  XOR3HSV2 U60537 ( .A1(n58516), .A2(n58515), .A3(n58514), .Z(n58517) );
  XNOR2HSV1 U60538 ( .A1(n58518), .A2(n58517), .ZN(n58519) );
  XOR2HSV0 U60539 ( .A1(n58520), .A2(n58519), .Z(n58521) );
  XOR2HSV0 U60540 ( .A1(n58522), .A2(n58521), .Z(n58524) );
  CLKNAND2HSV1 U60541 ( .A1(n25849), .A2(n58812), .ZN(n58523) );
  CLKNAND2HSV1 U60542 ( .A1(\pe6/got [10]), .A2(n58575), .ZN(n58571) );
  NAND2HSV2 U60543 ( .A1(n58656), .A2(n58525), .ZN(n58569) );
  CLKNAND2HSV1 U60544 ( .A1(n58809), .A2(n58526), .ZN(n58567) );
  CLKNAND2HSV0 U60545 ( .A1(n58934), .A2(n58659), .ZN(n58565) );
  NAND2HSV0 U60546 ( .A1(n58611), .A2(n58661), .ZN(n58561) );
  CLKNAND2HSV1 U60547 ( .A1(n58660), .A2(n58527), .ZN(n58557) );
  CLKNAND2HSV1 U60548 ( .A1(n46769), .A2(n58816), .ZN(n58555) );
  NAND2HSV0 U60549 ( .A1(n58601), .A2(n58817), .ZN(n58553) );
  CLKNAND2HSV1 U60550 ( .A1(\pe6/bq[12] ), .A2(\pe6/aot [1]), .ZN(n58529) );
  BUFHSV2 U60551 ( .I(\pe6/aot [6]), .Z(n58665) );
  CLKNAND2HSV0 U60552 ( .A1(n58675), .A2(n58665), .ZN(n58528) );
  XOR2HSV0 U60553 ( .A1(n58529), .A2(n58528), .Z(n58534) );
  CLKNAND2HSV1 U60554 ( .A1(n58356), .A2(n35632), .ZN(n58532) );
  NAND2HSV0 U60555 ( .A1(n58628), .A2(\pe6/aot [4]), .ZN(n58531) );
  XOR2HSV0 U60556 ( .A1(n58532), .A2(n58531), .Z(n58533) );
  XOR2HSV0 U60557 ( .A1(n58534), .A2(n58533), .Z(n58543) );
  NAND2HSV0 U60558 ( .A1(n35750), .A2(n58579), .ZN(n58536) );
  NAND2HSV0 U60559 ( .A1(n58360), .A2(\pe6/aot [11]), .ZN(n58535) );
  XOR2HSV0 U60560 ( .A1(n58536), .A2(n58535), .Z(n58541) );
  CLKNAND2HSV1 U60561 ( .A1(n58618), .A2(\pe6/aot [7]), .ZN(n58539) );
  CLKNAND2HSV1 U60562 ( .A1(n49106), .A2(n58999), .ZN(n58538) );
  XOR2HSV0 U60563 ( .A1(n58539), .A2(n58538), .Z(n58540) );
  XOR2HSV0 U60564 ( .A1(n58541), .A2(n58540), .Z(n58542) );
  XOR2HSV0 U60565 ( .A1(n58543), .A2(n58542), .Z(n58551) );
  XOR2HSV0 U60566 ( .A1(n58545), .A2(n58544), .Z(n58549) );
  CLKNAND2HSV0 U60567 ( .A1(n59277), .A2(n58631), .ZN(n58547) );
  CLKNAND2HSV0 U60568 ( .A1(n58619), .A2(\pe6/aot [5]), .ZN(n58546) );
  XOR2HSV0 U60569 ( .A1(n58547), .A2(n58546), .Z(n58548) );
  XOR2HSV0 U60570 ( .A1(n58549), .A2(n58548), .Z(n58550) );
  XNOR2HSV1 U60571 ( .A1(n58551), .A2(n58550), .ZN(n58552) );
  XNOR2HSV1 U60572 ( .A1(n58553), .A2(n58552), .ZN(n58554) );
  XNOR2HSV1 U60573 ( .A1(n58555), .A2(n58554), .ZN(n58556) );
  XNOR2HSV1 U60574 ( .A1(n58557), .A2(n58556), .ZN(n58559) );
  CLKNAND2HSV0 U60575 ( .A1(n58805), .A2(n46173), .ZN(n58558) );
  XOR2HSV0 U60576 ( .A1(n58559), .A2(n58558), .Z(n58560) );
  XNOR2HSV1 U60577 ( .A1(n58561), .A2(n58560), .ZN(n58564) );
  CLKNAND2HSV0 U60578 ( .A1(n29753), .A2(n58562), .ZN(n58563) );
  XOR3HSV2 U60579 ( .A1(n58565), .A2(n58564), .A3(n58563), .Z(n58566) );
  XNOR2HSV1 U60580 ( .A1(n58567), .A2(n58566), .ZN(n58568) );
  XNOR2HSV1 U60581 ( .A1(n58569), .A2(n58568), .ZN(n58570) );
  XNOR2HSV1 U60582 ( .A1(n58571), .A2(n58570), .ZN(n58574) );
  NAND2HSV2 U60583 ( .A1(n25849), .A2(n58572), .ZN(n58573) );
  CLKNAND2HSV1 U60584 ( .A1(n58660), .A2(n46173), .ZN(n58608) );
  CLKNAND2HSV1 U60585 ( .A1(n46769), .A2(n48891), .ZN(n58606) );
  CLKNAND2HSV0 U60586 ( .A1(n58962), .A2(\pe6/aot [4]), .ZN(n58578) );
  CLKNHSV0 U60587 ( .I(n49327), .ZN(n59216) );
  CLKNAND2HSV0 U60588 ( .A1(n59216), .A2(\pe6/aot [11]), .ZN(n58577) );
  XOR2HSV0 U60589 ( .A1(n58578), .A2(n58577), .Z(n58583) );
  CLKNAND2HSV1 U60590 ( .A1(n36143), .A2(\pe6/aot [1]), .ZN(n58581) );
  NAND2HSV0 U60591 ( .A1(\pe6/bq[12] ), .A2(n58579), .ZN(n58580) );
  XOR2HSV0 U60592 ( .A1(n58581), .A2(n58580), .Z(n58582) );
  XOR2HSV0 U60593 ( .A1(n58583), .A2(n58582), .Z(n58591) );
  NAND2HSV0 U60594 ( .A1(n35750), .A2(n58404), .ZN(n58585) );
  CLKNAND2HSV0 U60595 ( .A1(n49106), .A2(\pe6/aot [10]), .ZN(n58584) );
  XOR2HSV0 U60596 ( .A1(n58585), .A2(n58584), .Z(n58589) );
  CLKNAND2HSV0 U60597 ( .A1(n58619), .A2(n58665), .ZN(n58587) );
  CLKNAND2HSV0 U60598 ( .A1(n58452), .A2(n58999), .ZN(n58586) );
  XOR2HSV0 U60599 ( .A1(n58587), .A2(n58586), .Z(n58588) );
  XOR2HSV0 U60600 ( .A1(n58589), .A2(n58588), .Z(n58590) );
  XOR2HSV0 U60601 ( .A1(n58591), .A2(n58590), .Z(n58600) );
  CLKNAND2HSV0 U60602 ( .A1(n58618), .A2(n58449), .ZN(n58593) );
  NAND2HSV0 U60603 ( .A1(n59277), .A2(\pe6/aot [13]), .ZN(n58592) );
  XOR2HSV0 U60604 ( .A1(n58593), .A2(n58592), .Z(n58597) );
  XOR2HSV0 U60605 ( .A1(n58595), .A2(n58594), .Z(n58596) );
  XOR3HSV2 U60606 ( .A1(n58598), .A2(n58597), .A3(n58596), .Z(n58599) );
  XNOR2HSV1 U60607 ( .A1(n58600), .A2(n58599), .ZN(n58604) );
  NAND2HSV0 U60608 ( .A1(n58662), .A2(n58403), .ZN(n58603) );
  NAND2HSV0 U60609 ( .A1(n58601), .A2(n59231), .ZN(n58602) );
  XOR3HSV2 U60610 ( .A1(n58604), .A2(n58603), .A3(n58602), .Z(n58605) );
  XNOR2HSV1 U60611 ( .A1(n58606), .A2(n58605), .ZN(n58607) );
  XNOR2HSV1 U60612 ( .A1(n58608), .A2(n58607), .ZN(n58610) );
  CLKNAND2HSV0 U60613 ( .A1(n59335), .A2(n58661), .ZN(n58609) );
  CLKNAND2HSV1 U60614 ( .A1(n58660), .A2(n58661), .ZN(n58651) );
  CLKNAND2HSV0 U60615 ( .A1(n58718), .A2(n46173), .ZN(n58649) );
  NAND2HSV0 U60616 ( .A1(n58662), .A2(n59231), .ZN(n58645) );
  NAND2HSV0 U60617 ( .A1(n58663), .A2(n58403), .ZN(n58643) );
  NAND2HSV0 U60618 ( .A1(n58668), .A2(\pe6/aot [1]), .ZN(n58613) );
  NAND2HSV0 U60619 ( .A1(n58990), .A2(n58943), .ZN(n58612) );
  XOR2HSV0 U60620 ( .A1(n58613), .A2(n58612), .Z(n58617) );
  CLKNAND2HSV0 U60621 ( .A1(n58675), .A2(n58449), .ZN(n58615) );
  NAND2HSV0 U60622 ( .A1(n36143), .A2(n59260), .ZN(n58614) );
  XOR2HSV0 U60623 ( .A1(n58615), .A2(n58614), .Z(n58616) );
  XOR2HSV0 U60624 ( .A1(n58617), .A2(n58616), .Z(n58627) );
  NAND2HSV0 U60625 ( .A1(n58618), .A2(n58999), .ZN(n58621) );
  NAND2HSV0 U60626 ( .A1(n58619), .A2(\pe6/aot [7]), .ZN(n58620) );
  XOR2HSV0 U60627 ( .A1(n58621), .A2(n58620), .Z(n58625) );
  CLKNAND2HSV0 U60628 ( .A1(n58452), .A2(\pe6/aot [10]), .ZN(n58623) );
  NAND2HSV0 U60629 ( .A1(\pe6/bq[12] ), .A2(n58404), .ZN(n58622) );
  XOR2HSV0 U60630 ( .A1(n58623), .A2(n58622), .Z(n58624) );
  XOR2HSV0 U60631 ( .A1(n58625), .A2(n58624), .Z(n58626) );
  XOR2HSV0 U60632 ( .A1(n58627), .A2(n58626), .Z(n58641) );
  NAND2HSV0 U60633 ( .A1(n58628), .A2(n58665), .ZN(n58630) );
  CLKNAND2HSV0 U60634 ( .A1(n49106), .A2(\pe6/aot [11]), .ZN(n58629) );
  XOR2HSV0 U60635 ( .A1(n58630), .A2(n58629), .Z(n58635) );
  CLKNAND2HSV0 U60636 ( .A1(n59216), .A2(n58631), .ZN(n58633) );
  CLKNAND2HSV1 U60637 ( .A1(n58360), .A2(\pe6/aot [13]), .ZN(n58632) );
  XOR2HSV0 U60638 ( .A1(n58633), .A2(n58632), .Z(n58634) );
  XNOR2HSV1 U60639 ( .A1(n58635), .A2(n58634), .ZN(n58639) );
  NAND2HSV0 U60640 ( .A1(n35750), .A2(\pe6/aot [4]), .ZN(n58636) );
  XOR2HSV0 U60641 ( .A1(n58637), .A2(n58636), .Z(n58638) );
  XNOR2HSV1 U60642 ( .A1(n58639), .A2(n58638), .ZN(n58640) );
  XNOR2HSV1 U60643 ( .A1(n58641), .A2(n58640), .ZN(n58642) );
  XNOR2HSV1 U60644 ( .A1(n58643), .A2(n58642), .ZN(n58644) );
  XNOR2HSV1 U60645 ( .A1(n58645), .A2(n58644), .ZN(n58647) );
  CLKNAND2HSV1 U60646 ( .A1(n58702), .A2(n48891), .ZN(n58646) );
  XNOR2HSV1 U60647 ( .A1(n58647), .A2(n58646), .ZN(n58648) );
  XNOR2HSV1 U60648 ( .A1(n58649), .A2(n58648), .ZN(n58650) );
  XNOR2HSV1 U60649 ( .A1(n58651), .A2(n58650), .ZN(n58653) );
  CLKNAND2HSV0 U60650 ( .A1(n59335), .A2(n58659), .ZN(n58652) );
  CLKNAND2HSV0 U60651 ( .A1(n58660), .A2(n58659), .ZN(n58708) );
  CLKNAND2HSV0 U60652 ( .A1(n58936), .A2(n58661), .ZN(n58706) );
  NAND2HSV0 U60653 ( .A1(n58662), .A2(n58527), .ZN(n58701) );
  NAND2HSV0 U60654 ( .A1(n58663), .A2(n59231), .ZN(n58699) );
  NAND2HSV0 U60655 ( .A1(n58664), .A2(n58403), .ZN(n58697) );
  CLKNAND2HSV1 U60656 ( .A1(n59240), .A2(n58459), .ZN(n58667) );
  NAND2HSV0 U60657 ( .A1(n58962), .A2(n58665), .ZN(n58666) );
  XOR2HSV0 U60658 ( .A1(n58667), .A2(n58666), .Z(n58672) );
  NAND2HSV0 U60659 ( .A1(n35750), .A2(n58378), .ZN(n58670) );
  NAND2HSV0 U60660 ( .A1(n58668), .A2(n58464), .ZN(n58669) );
  XOR2HSV0 U60661 ( .A1(n58670), .A2(n58669), .Z(n58671) );
  XOR2HSV0 U60662 ( .A1(n58672), .A2(n58671), .Z(n58681) );
  CLKNAND2HSV1 U60663 ( .A1(n59265), .A2(n59252), .ZN(n58674) );
  CLKNAND2HSV0 U60664 ( .A1(n48038), .A2(\pe6/aot [10]), .ZN(n58673) );
  XOR2HSV0 U60665 ( .A1(n58674), .A2(n58673), .Z(n58679) );
  NAND2HSV0 U60666 ( .A1(n58675), .A2(n58999), .ZN(n58676) );
  XOR2HSV0 U60667 ( .A1(n58677), .A2(n58676), .Z(n58678) );
  XOR2HSV0 U60668 ( .A1(n58679), .A2(n58678), .Z(n58680) );
  XOR2HSV0 U60669 ( .A1(n58681), .A2(n58680), .Z(n58695) );
  CLKNAND2HSV0 U60670 ( .A1(n58682), .A2(\pe6/aot [1]), .ZN(n58684) );
  CLKNAND2HSV0 U60671 ( .A1(n59216), .A2(\pe6/aot [13]), .ZN(n58683) );
  XOR2HSV0 U60672 ( .A1(n58684), .A2(n58683), .Z(n58688) );
  NAND2HSV2 U60673 ( .A1(n58731), .A2(\pe6/aot [11]), .ZN(n58686) );
  NAND2HSV0 U60674 ( .A1(n59041), .A2(\pe6/aot [14]), .ZN(n58685) );
  XOR2HSV0 U60675 ( .A1(n58686), .A2(n58685), .Z(n58687) );
  XOR2HSV0 U60676 ( .A1(n58688), .A2(n58687), .Z(n58693) );
  CLKNAND2HSV1 U60677 ( .A1(n59084), .A2(\pe6/aot [7]), .ZN(n58690) );
  CLKNAND2HSV0 U60678 ( .A1(n58990), .A2(n33024), .ZN(n58689) );
  XOR2HSV0 U60679 ( .A1(n58690), .A2(n58689), .Z(n58691) );
  NOR2HSV0 U60680 ( .A1(n48042), .A2(n58483), .ZN(n58860) );
  XNOR2HSV1 U60681 ( .A1(n58691), .A2(n58860), .ZN(n58692) );
  XNOR2HSV1 U60682 ( .A1(n58693), .A2(n58692), .ZN(n58694) );
  XNOR2HSV1 U60683 ( .A1(n58695), .A2(n58694), .ZN(n58696) );
  XNOR2HSV1 U60684 ( .A1(n58697), .A2(n58696), .ZN(n58698) );
  XNOR2HSV1 U60685 ( .A1(n58699), .A2(n58698), .ZN(n58700) );
  XNOR2HSV1 U60686 ( .A1(n58701), .A2(n58700), .ZN(n58704) );
  CLKNAND2HSV0 U60687 ( .A1(n58702), .A2(\pe6/got [4]), .ZN(n58703) );
  XNOR2HSV1 U60688 ( .A1(n58704), .A2(n58703), .ZN(n58705) );
  XNOR2HSV1 U60689 ( .A1(n58706), .A2(n58705), .ZN(n58707) );
  CLKNAND2HSV0 U60690 ( .A1(n59335), .A2(n58709), .ZN(n58710) );
  CLKNAND2HSV1 U60691 ( .A1(n58935), .A2(\pe6/got [15]), .ZN(n58804) );
  CLKNAND2HSV0 U60692 ( .A1(n58718), .A2(n58810), .ZN(n58802) );
  NAND2HSV0 U60693 ( .A1(n59177), .A2(n58719), .ZN(n58798) );
  CLKNAND2HSV1 U60694 ( .A1(n53112), .A2(n58720), .ZN(n58796) );
  CLKNAND2HSV1 U60695 ( .A1(n58938), .A2(\pe6/got [10]), .ZN(n58794) );
  CLKNAND2HSV1 U60696 ( .A1(n53114), .A2(n58721), .ZN(n58792) );
  NAND2HSV0 U60697 ( .A1(n58722), .A2(\pe6/got [7]), .ZN(n58788) );
  CLKNAND2HSV1 U60698 ( .A1(n59033), .A2(n58723), .ZN(n58786) );
  NAND2HSV0 U60699 ( .A1(n58813), .A2(n58478), .ZN(n58784) );
  NAND2HSV0 U60700 ( .A1(n59036), .A2(n58479), .ZN(n58782) );
  NAND2HSV0 U60701 ( .A1(n32165), .A2(n58527), .ZN(n58780) );
  NAND2HSV0 U60702 ( .A1(n58886), .A2(n58403), .ZN(n58776) );
  NAND2HSV0 U60703 ( .A1(n59066), .A2(n49831), .ZN(n58726) );
  NAND2HSV0 U60704 ( .A1(n48038), .A2(\pe6/aot [19]), .ZN(n58725) );
  XOR2HSV0 U60705 ( .A1(n58726), .A2(n58725), .Z(n58730) );
  NAND2HSV0 U60706 ( .A1(n59084), .A2(n59044), .ZN(n58728) );
  CLKNAND2HSV0 U60707 ( .A1(\pe6/bq[2] ), .A2(\pe6/aot [23]), .ZN(n58727) );
  XOR2HSV0 U60708 ( .A1(n58728), .A2(n58727), .Z(n58729) );
  XOR2HSV0 U60709 ( .A1(n58730), .A2(n58729), .Z(n58740) );
  NAND2HSV0 U60710 ( .A1(n58731), .A2(n59264), .ZN(n58733) );
  NAND2HSV0 U60711 ( .A1(\pe6/bq[21] ), .A2(\pe6/aot [4]), .ZN(n58732) );
  XOR2HSV0 U60712 ( .A1(n58733), .A2(n58732), .Z(n58738) );
  NAND2HSV0 U60713 ( .A1(n32886), .A2(n58734), .ZN(n58736) );
  NAND2HSV0 U60714 ( .A1(n58962), .A2(n58842), .ZN(n58735) );
  XOR2HSV0 U60715 ( .A1(n58736), .A2(n58735), .Z(n58737) );
  XOR2HSV0 U60716 ( .A1(n58738), .A2(n58737), .Z(n58739) );
  XOR2HSV0 U60717 ( .A1(n58740), .A2(n58739), .Z(n58757) );
  NAND2HSV0 U60718 ( .A1(n59050), .A2(\pe6/aot [1]), .ZN(n58742) );
  NAND2HSV0 U60719 ( .A1(n44702), .A2(n59260), .ZN(n58741) );
  XOR2HSV0 U60720 ( .A1(n58742), .A2(n58741), .Z(n58746) );
  NAND2HSV0 U60721 ( .A1(n59224), .A2(n59266), .ZN(n58744) );
  NAND2HSV0 U60722 ( .A1(n58976), .A2(\pe6/aot [13]), .ZN(n58743) );
  XOR2HSV0 U60723 ( .A1(n58744), .A2(n58743), .Z(n58745) );
  XOR2HSV0 U60724 ( .A1(n58746), .A2(n58745), .Z(n58755) );
  NOR2HSV0 U60725 ( .A1(n46853), .A2(n49188), .ZN(n58748) );
  NAND2HSV0 U60726 ( .A1(n58668), .A2(\pe6/aot [11]), .ZN(n58747) );
  XOR2HSV0 U60727 ( .A1(n58748), .A2(n58747), .Z(n58753) );
  AOI22HSV0 U60728 ( .A1(n59062), .A2(\pe6/aot [21]), .B1(n58749), .B2(n58990), 
        .ZN(n58750) );
  AOI21HSV1 U60729 ( .A1(n58751), .A2(n58855), .B(n58750), .ZN(n58752) );
  XNOR2HSV1 U60730 ( .A1(n58753), .A2(n58752), .ZN(n58754) );
  XNOR2HSV1 U60731 ( .A1(n58755), .A2(n58754), .ZN(n58756) );
  XNOR2HSV1 U60732 ( .A1(n58757), .A2(n58756), .ZN(n58774) );
  NAND2HSV0 U60733 ( .A1(n46210), .A2(n49208), .ZN(n58759) );
  NAND2HSV0 U60734 ( .A1(n59246), .A2(\pe6/aot [17]), .ZN(n58758) );
  XOR2HSV0 U60735 ( .A1(n58759), .A2(n58758), .Z(n58764) );
  NAND2HSV0 U60736 ( .A1(n59273), .A2(n58760), .ZN(n58762) );
  NAND2HSV0 U60737 ( .A1(\pe6/bq[18] ), .A2(\pe6/aot [7]), .ZN(n58761) );
  XOR2HSV0 U60738 ( .A1(n58762), .A2(n58761), .Z(n58763) );
  XOR2HSV0 U60739 ( .A1(n58764), .A2(n58763), .Z(n58772) );
  NAND2HSV0 U60740 ( .A1(n58833), .A2(n59099), .ZN(n58765) );
  XOR2HSV0 U60741 ( .A1(n58766), .A2(n58765), .Z(n58770) );
  NOR2HSV0 U60742 ( .A1(n46688), .A2(n58483), .ZN(n58768) );
  NAND2HSV0 U60743 ( .A1(n59045), .A2(\pe6/aot [10]), .ZN(n58767) );
  XOR2HSV0 U60744 ( .A1(n58768), .A2(n58767), .Z(n58769) );
  XOR2HSV0 U60745 ( .A1(n58770), .A2(n58769), .Z(n58771) );
  XOR2HSV0 U60746 ( .A1(n58772), .A2(n58771), .Z(n58773) );
  XNOR2HSV1 U60747 ( .A1(n58774), .A2(n58773), .ZN(n58775) );
  XNOR2HSV1 U60748 ( .A1(n58776), .A2(n58775), .ZN(n58777) );
  XNOR2HSV1 U60749 ( .A1(n58778), .A2(n58777), .ZN(n58779) );
  XNOR2HSV1 U60750 ( .A1(n58780), .A2(n58779), .ZN(n58781) );
  XNOR2HSV1 U60751 ( .A1(n58782), .A2(n58781), .ZN(n58783) );
  XNOR2HSV1 U60752 ( .A1(n58784), .A2(n58783), .ZN(n58785) );
  XNOR2HSV1 U60753 ( .A1(n58786), .A2(n58785), .ZN(n58787) );
  XNOR2HSV1 U60754 ( .A1(n58788), .A2(n58787), .ZN(n58790) );
  CLKNAND2HSV0 U60755 ( .A1(n59144), .A2(n58526), .ZN(n58789) );
  XNOR2HSV1 U60756 ( .A1(n58790), .A2(n58789), .ZN(n58791) );
  XNOR2HSV1 U60757 ( .A1(n58792), .A2(n58791), .ZN(n58793) );
  XNOR2HSV1 U60758 ( .A1(n58794), .A2(n58793), .ZN(n58795) );
  XNOR2HSV1 U60759 ( .A1(n58796), .A2(n58795), .ZN(n58797) );
  XNOR2HSV1 U60760 ( .A1(n58798), .A2(n58797), .ZN(n58800) );
  CLKNAND2HSV1 U60761 ( .A1(n59915), .A2(\pe6/got [13]), .ZN(n58799) );
  XNOR2HSV1 U60762 ( .A1(n58800), .A2(n58799), .ZN(n58801) );
  XNOR2HSV1 U60763 ( .A1(n58802), .A2(n58801), .ZN(n58803) );
  CLKNAND2HSV0 U60764 ( .A1(n58805), .A2(n58937), .ZN(n58806) );
  CLKNAND2HSV1 U60765 ( .A1(n59173), .A2(n59169), .ZN(n58930) );
  CLKNAND2HSV1 U60766 ( .A1(n59514), .A2(n59165), .ZN(n58928) );
  CLKNAND2HSV1 U60767 ( .A1(n58809), .A2(n59027), .ZN(n58926) );
  CLKNAND2HSV0 U60768 ( .A1(n58934), .A2(n59328), .ZN(n58924) );
  CLKNAND2HSV1 U60769 ( .A1(n59028), .A2(n59029), .ZN(n58921) );
  CLKNAND2HSV1 U60770 ( .A1(n58935), .A2(n53101), .ZN(n58917) );
  CLKNAND2HSV1 U60771 ( .A1(n58718), .A2(n32971), .ZN(n58915) );
  NAND2HSV0 U60772 ( .A1(n59177), .A2(\pe6/got [15]), .ZN(n58911) );
  NAND2HSV0 U60773 ( .A1(n59916), .A2(n58810), .ZN(n58909) );
  CLKNAND2HSV0 U60774 ( .A1(n58938), .A2(n58811), .ZN(n58907) );
  NAND2HSV0 U60775 ( .A1(n53114), .A2(\pe6/got [12]), .ZN(n58905) );
  NAND2HSV0 U60776 ( .A1(n46632), .A2(n58812), .ZN(n58900) );
  NAND2HSV0 U60777 ( .A1(n46172), .A2(n59037), .ZN(n58898) );
  NAND2HSV0 U60778 ( .A1(n58813), .A2(n58526), .ZN(n58896) );
  NAND2HSV0 U60779 ( .A1(n59036), .A2(n58814), .ZN(n58894) );
  NAND2HSV0 U60780 ( .A1(n58815), .A2(n58659), .ZN(n58892) );
  NAND2HSV0 U60781 ( .A1(n32218), .A2(n48891), .ZN(n58885) );
  NAND2HSV0 U60782 ( .A1(n59183), .A2(n58816), .ZN(n58883) );
  NAND2HSV0 U60783 ( .A1(n25218), .A2(n58817), .ZN(n58881) );
  NAND2HSV0 U60784 ( .A1(n32172), .A2(\pe6/aot [7]), .ZN(n58819) );
  NAND2HSV0 U60785 ( .A1(\pe6/bq[25] ), .A2(n58404), .ZN(n58818) );
  XOR2HSV0 U60786 ( .A1(n58819), .A2(n58818), .Z(n58823) );
  NAND2HSV0 U60787 ( .A1(n32886), .A2(n58665), .ZN(n58821) );
  NAND2HSV0 U60788 ( .A1(n44702), .A2(n59250), .ZN(n58820) );
  XOR2HSV0 U60789 ( .A1(n58821), .A2(n58820), .Z(n58822) );
  XOR2HSV0 U60790 ( .A1(n58823), .A2(n58822), .Z(n58832) );
  NAND2HSV0 U60791 ( .A1(n59066), .A2(n58824), .ZN(n58826) );
  NAND2HSV0 U60792 ( .A1(n58965), .A2(\pe6/aot [1]), .ZN(n58825) );
  XOR2HSV0 U60793 ( .A1(n58826), .A2(n58825), .Z(n58830) );
  NAND2HSV0 U60794 ( .A1(\pe6/bq[17] ), .A2(\pe6/aot [11]), .ZN(n58828) );
  NAND2HSV0 U60795 ( .A1(n58975), .A2(n49831), .ZN(n58827) );
  XOR2HSV0 U60796 ( .A1(n58828), .A2(n58827), .Z(n58829) );
  XOR2HSV0 U60797 ( .A1(n58830), .A2(n58829), .Z(n58831) );
  XOR2HSV0 U60798 ( .A1(n58832), .A2(n58831), .Z(n58850) );
  NAND2HSV0 U60799 ( .A1(n58833), .A2(n58631), .ZN(n58835) );
  NAND2HSV0 U60800 ( .A1(n59050), .A2(n58459), .ZN(n58834) );
  XOR2HSV0 U60801 ( .A1(n58835), .A2(n58834), .Z(n58839) );
  NAND2HSV0 U60802 ( .A1(n58336), .A2(n32588), .ZN(n58837) );
  NAND2HSV0 U60803 ( .A1(n36150), .A2(\pe6/aot [10]), .ZN(n58836) );
  XOR2HSV0 U60804 ( .A1(n58837), .A2(n58836), .Z(n58838) );
  XOR2HSV0 U60805 ( .A1(n58839), .A2(n58838), .Z(n58848) );
  NAND2HSV0 U60806 ( .A1(\pe6/bq[5] ), .A2(\pe6/aot [23]), .ZN(n58841) );
  NAND2HSV0 U60807 ( .A1(n59075), .A2(\pe6/aot [21]), .ZN(n58840) );
  XOR2HSV0 U60808 ( .A1(n58841), .A2(n58840), .Z(n58846) );
  NAND2HSV0 U60809 ( .A1(n35751), .A2(\pe6/aot [13]), .ZN(n58844) );
  NAND2HSV0 U60810 ( .A1(n59089), .A2(n58842), .ZN(n58843) );
  XOR2HSV0 U60811 ( .A1(n58844), .A2(n58843), .Z(n58845) );
  XOR2HSV0 U60812 ( .A1(n58846), .A2(n58845), .Z(n58847) );
  XOR2HSV0 U60813 ( .A1(n58848), .A2(n58847), .Z(n58849) );
  XOR2HSV0 U60814 ( .A1(n58850), .A2(n58849), .Z(n58879) );
  NOR2HSV0 U60815 ( .A1(n46850), .A2(n58851), .ZN(n58854) );
  OAI22HSV0 U60816 ( .A1(n58855), .A2(n58854), .B1(n58853), .B2(n58852), .ZN(
        n58862) );
  AOI22HSV0 U60817 ( .A1(n59098), .A2(n58857), .B1(n58856), .B2(\pe6/bq[8] ), 
        .ZN(n58858) );
  AOI21HSV0 U60818 ( .A1(n58860), .A2(n58859), .B(n58858), .ZN(n58861) );
  XOR2HSV0 U60819 ( .A1(n58862), .A2(n58861), .Z(n58869) );
  NAND2HSV0 U60820 ( .A1(n58668), .A2(n58943), .ZN(n58865) );
  NOR2HSV0 U60821 ( .A1(n58863), .A2(n59188), .ZN(n58864) );
  AOI21HSV0 U60822 ( .A1(n58866), .A2(n58865), .B(n58864), .ZN(n58867) );
  XOR2HSV0 U60823 ( .A1(n58867), .A2(n59108), .Z(n58868) );
  XNOR2HSV1 U60824 ( .A1(n58869), .A2(n58868), .ZN(n58877) );
  NAND2HSV0 U60825 ( .A1(n58962), .A2(n59088), .ZN(n58870) );
  XOR2HSV0 U60826 ( .A1(n58871), .A2(n58870), .Z(n58875) );
  NAND2HSV0 U60827 ( .A1(n59084), .A2(\pe6/aot [19]), .ZN(n58873) );
  NAND2HSV0 U60828 ( .A1(\pe6/bq[2] ), .A2(n32876), .ZN(n58872) );
  XOR2HSV0 U60829 ( .A1(n58873), .A2(n58872), .Z(n58874) );
  XOR2HSV0 U60830 ( .A1(n58875), .A2(n58874), .Z(n58876) );
  XNOR2HSV1 U60831 ( .A1(n58877), .A2(n58876), .ZN(n58878) );
  XNOR2HSV1 U60832 ( .A1(n58879), .A2(n58878), .ZN(n58880) );
  XNOR2HSV1 U60833 ( .A1(n58881), .A2(n58880), .ZN(n58882) );
  XNOR2HSV1 U60834 ( .A1(n58883), .A2(n58882), .ZN(n58884) );
  XNOR2HSV1 U60835 ( .A1(n58885), .A2(n58884), .ZN(n58888) );
  NAND2HSV0 U60836 ( .A1(n58886), .A2(n58479), .ZN(n58887) );
  XNOR2HSV1 U60837 ( .A1(n58888), .A2(n58887), .ZN(n58889) );
  XNOR2HSV1 U60838 ( .A1(n58890), .A2(n58889), .ZN(n58891) );
  XNOR2HSV1 U60839 ( .A1(n58892), .A2(n58891), .ZN(n58893) );
  XNOR2HSV1 U60840 ( .A1(n58894), .A2(n58893), .ZN(n58895) );
  XNOR2HSV1 U60841 ( .A1(n58896), .A2(n58895), .ZN(n58897) );
  XNOR2HSV1 U60842 ( .A1(n58898), .A2(n58897), .ZN(n58899) );
  XNOR2HSV1 U60843 ( .A1(n58900), .A2(n58899), .ZN(n58903) );
  CLKNAND2HSV0 U60844 ( .A1(n58901), .A2(n59181), .ZN(n58902) );
  XNOR2HSV1 U60845 ( .A1(n58903), .A2(n58902), .ZN(n58904) );
  XOR2HSV0 U60846 ( .A1(n58905), .A2(n58904), .Z(n58906) );
  XOR2HSV0 U60847 ( .A1(n58907), .A2(n58906), .Z(n58908) );
  XNOR2HSV1 U60848 ( .A1(n58909), .A2(n58908), .ZN(n58910) );
  XNOR2HSV1 U60849 ( .A1(n58911), .A2(n58910), .ZN(n58913) );
  CLKNAND2HSV1 U60850 ( .A1(n49726), .A2(n58937), .ZN(n58912) );
  XNOR2HSV1 U60851 ( .A1(n58913), .A2(n58912), .ZN(n58914) );
  XNOR2HSV1 U60852 ( .A1(n58915), .A2(n58914), .ZN(n58916) );
  XOR2HSV0 U60853 ( .A1(n58917), .A2(n58916), .Z(n58919) );
  CLKNAND2HSV0 U60854 ( .A1(n59161), .A2(\pe6/got [19]), .ZN(n58918) );
  XOR2HSV0 U60855 ( .A1(n58919), .A2(n58918), .Z(n58920) );
  XNOR2HSV1 U60856 ( .A1(n58921), .A2(n58920), .ZN(n58923) );
  XOR3HSV2 U60857 ( .A1(n58924), .A2(n58923), .A3(n58922), .Z(n58925) );
  XNOR2HSV1 U60858 ( .A1(n58926), .A2(n58925), .ZN(n58927) );
  XNOR2HSV1 U60859 ( .A1(n58928), .A2(n58927), .ZN(n58929) );
  XNOR2HSV1 U60860 ( .A1(n58930), .A2(n58929), .ZN(n58933) );
  NAND2HSV2 U60861 ( .A1(n59021), .A2(n59025), .ZN(n58932) );
  XOR3HSV2 U60862 ( .A1(n58933), .A2(n58932), .A3(n58931), .Z(\pe6/poht [5])
         );
  CLKNAND2HSV1 U60863 ( .A1(n58935), .A2(n35922), .ZN(n59019) );
  NAND2HSV0 U60864 ( .A1(n59678), .A2(n58479), .ZN(n59017) );
  NAND2HSV0 U60865 ( .A1(n59183), .A2(n58527), .ZN(n59015) );
  NAND2HSV0 U60866 ( .A1(n58940), .A2(n59235), .ZN(n59010) );
  NAND2HSV0 U60867 ( .A1(n59041), .A2(n32588), .ZN(n58942) );
  NAND2HSV0 U60868 ( .A1(n59066), .A2(n32876), .ZN(n58941) );
  XOR2HSV0 U60869 ( .A1(n58942), .A2(n58941), .Z(n58947) );
  NAND2HSV0 U60870 ( .A1(n58682), .A2(n58943), .ZN(n58945) );
  NAND2HSV0 U60871 ( .A1(n58668), .A2(n58842), .ZN(n58944) );
  XOR2HSV0 U60872 ( .A1(n58945), .A2(n58944), .Z(n58946) );
  XOR2HSV0 U60873 ( .A1(n58947), .A2(n58946), .Z(n58955) );
  NAND2HSV0 U60874 ( .A1(n32172), .A2(n35632), .ZN(n58949) );
  NAND2HSV0 U60875 ( .A1(\pe6/bq[25] ), .A2(n58459), .ZN(n58948) );
  XOR2HSV0 U60876 ( .A1(n58949), .A2(n58948), .Z(n58953) );
  NAND2HSV0 U60877 ( .A1(n48035), .A2(n58353), .ZN(n58951) );
  NAND2HSV0 U60878 ( .A1(\pe6/bq[11] ), .A2(n59088), .ZN(n58950) );
  XOR2HSV0 U60879 ( .A1(n58951), .A2(n58950), .Z(n58952) );
  XOR2HSV0 U60880 ( .A1(n58953), .A2(n58952), .Z(n58954) );
  XOR2HSV0 U60881 ( .A1(n58955), .A2(n58954), .Z(n58973) );
  NAND2HSV0 U60882 ( .A1(n59054), .A2(n58665), .ZN(n58957) );
  NAND2HSV0 U60883 ( .A1(n59050), .A2(n59250), .ZN(n58956) );
  XOR2HSV0 U60884 ( .A1(n58957), .A2(n58956), .Z(n58961) );
  NAND2HSV0 U60885 ( .A1(n59084), .A2(n59264), .ZN(n58959) );
  NAND2HSV0 U60886 ( .A1(n33023), .A2(\pe6/aot [11]), .ZN(n58958) );
  XOR2HSV0 U60887 ( .A1(n58959), .A2(n58958), .Z(n58960) );
  XOR2HSV0 U60888 ( .A1(n58961), .A2(n58960), .Z(n58971) );
  NAND2HSV0 U60889 ( .A1(n59273), .A2(n33004), .ZN(n58964) );
  NAND2HSV0 U60890 ( .A1(n58962), .A2(\pe6/aot [19]), .ZN(n58963) );
  XOR2HSV0 U60891 ( .A1(n58964), .A2(n58963), .Z(n58969) );
  NAND2HSV0 U60892 ( .A1(n58965), .A2(\pe6/aot [2]), .ZN(n58967) );
  NAND2HSV0 U60893 ( .A1(n59251), .A2(\pe6/aot [1]), .ZN(n58966) );
  XOR2HSV0 U60894 ( .A1(n58967), .A2(n58966), .Z(n58968) );
  XOR2HSV0 U60895 ( .A1(n58969), .A2(n58968), .Z(n58970) );
  XOR2HSV0 U60896 ( .A1(n58971), .A2(n58970), .Z(n58972) );
  XOR2HSV0 U60897 ( .A1(n58973), .A2(n58972), .Z(n59008) );
  CLKNHSV0 U60898 ( .I(n58974), .ZN(n58979) );
  AOI22HSV0 U60899 ( .A1(n58976), .A2(\pe6/aot [17]), .B1(\pe6/aot [23]), .B2(
        n58975), .ZN(n58977) );
  AOI21HSV0 U60900 ( .A1(n58979), .A2(n58978), .B(n58977), .ZN(n58998) );
  NAND2HSV0 U60901 ( .A1(\pe6/bq[17] ), .A2(n58631), .ZN(n58981) );
  NAND2HSV0 U60902 ( .A1(\pe6/bq[5] ), .A2(n59239), .ZN(n58980) );
  XOR2HSV0 U60903 ( .A1(n58981), .A2(n58980), .Z(n58997) );
  CLKNHSV0 U60904 ( .I(n58982), .ZN(n58987) );
  NOR2HSV0 U60905 ( .A1(n58984), .A2(n58983), .ZN(n59107) );
  OAI22HSV0 U60906 ( .A1(n58987), .A2(n59107), .B1(n58986), .B2(n58985), .ZN(
        n58995) );
  NOR2HSV0 U60907 ( .A1(n58989), .A2(n58988), .ZN(n58993) );
  AOI22HSV0 U60908 ( .A1(n59062), .A2(n59087), .B1(n58991), .B2(n58990), .ZN(
        n58992) );
  NOR2HSV2 U60909 ( .A1(n58993), .A2(n58992), .ZN(n58994) );
  XNOR2HSV1 U60910 ( .A1(n58995), .A2(n58994), .ZN(n58996) );
  XOR3HSV2 U60911 ( .A1(n58998), .A2(n58997), .A3(n58996), .Z(n59006) );
  NAND2HSV0 U60912 ( .A1(n59098), .A2(n58999), .ZN(n59097) );
  XOR2HSV0 U60913 ( .A1(n59000), .A2(n59097), .Z(n59004) );
  NAND2HSV0 U60914 ( .A1(n59100), .A2(\pe6/aot [7]), .ZN(n59002) );
  NAND2HSV0 U60915 ( .A1(n59224), .A2(\pe6/aot [10]), .ZN(n59001) );
  XOR2HSV0 U60916 ( .A1(n59002), .A2(n59001), .Z(n59003) );
  XOR2HSV0 U60917 ( .A1(n59004), .A2(n59003), .Z(n59005) );
  XNOR2HSV1 U60918 ( .A1(n59006), .A2(n59005), .ZN(n59007) );
  XNOR2HSV1 U60919 ( .A1(n59008), .A2(n59007), .ZN(n59009) );
  XNOR2HSV1 U60920 ( .A1(n59010), .A2(n59009), .ZN(n59013) );
  NAND2HSV0 U60921 ( .A1(n25218), .A2(n59039), .ZN(n59012) );
  XOR2HSV0 U60922 ( .A1(n59013), .A2(n59012), .Z(n59014) );
  XNOR2HSV1 U60923 ( .A1(n59015), .A2(n59014), .ZN(n59016) );
  CLKNAND2HSV0 U60924 ( .A1(n59161), .A2(n59029), .ZN(n59020) );
  NAND2HSV0 U60925 ( .A1(n59918), .A2(n59328), .ZN(n59160) );
  NAND2HSV0 U60926 ( .A1(n59680), .A2(n59029), .ZN(n59158) );
  NAND2HSV0 U60927 ( .A1(n59177), .A2(n58715), .ZN(n59154) );
  CLKNAND2HSV1 U60928 ( .A1(n59030), .A2(n49098), .ZN(n59152) );
  NAND2HSV0 U60929 ( .A1(n53113), .A2(n59031), .ZN(n59150) );
  CLKNAND2HSV0 U60930 ( .A1(n59179), .A2(\pe6/got [15]), .ZN(n59148) );
  NAND2HSV0 U60931 ( .A1(n59032), .A2(n58811), .ZN(n59143) );
  NAND2HSV0 U60932 ( .A1(n59033), .A2(n33039), .ZN(n59141) );
  CLKNHSV0 U60933 ( .I(n59181), .ZN(n59035) );
  INAND2HSV0 U60934 ( .A1(n59035), .B1(n59034), .ZN(n59139) );
  NAND2HSV0 U60935 ( .A1(n59036), .A2(\pe6/got [10]), .ZN(n59137) );
  CLKNAND2HSV0 U60936 ( .A1(n49829), .A2(n59037), .ZN(n59135) );
  NAND2HSV0 U60937 ( .A1(n26109), .A2(\pe6/got [8]), .ZN(n59133) );
  NAND2HSV0 U60938 ( .A1(n59678), .A2(n58723), .ZN(n59129) );
  NAND2HSV0 U60939 ( .A1(n59597), .A2(n59292), .ZN(n59127) );
  NAND2HSV0 U60940 ( .A1(n59038), .A2(n59235), .ZN(n59120) );
  NAND2HSV0 U60941 ( .A1(n36108), .A2(n59039), .ZN(n59119) );
  NAND2HSV0 U60942 ( .A1(n58336), .A2(n59040), .ZN(n59043) );
  NAND2HSV0 U60943 ( .A1(n59041), .A2(n31555), .ZN(n59042) );
  XOR2HSV0 U60944 ( .A1(n59043), .A2(n59042), .Z(n59049) );
  NAND2HSV0 U60945 ( .A1(n32172), .A2(\pe6/aot [10]), .ZN(n59047) );
  NAND2HSV0 U60946 ( .A1(n59045), .A2(n59044), .ZN(n59046) );
  XOR2HSV0 U60947 ( .A1(n59047), .A2(n59046), .Z(n59048) );
  XOR2HSV0 U60948 ( .A1(n59049), .A2(n59048), .Z(n59060) );
  NAND2HSV0 U60949 ( .A1(n59050), .A2(\pe6/aot [7]), .ZN(n59053) );
  NAND2HSV0 U60950 ( .A1(n59051), .A2(n53115), .ZN(n59052) );
  XOR2HSV0 U60951 ( .A1(n59053), .A2(n59052), .Z(n59058) );
  NAND2HSV0 U60952 ( .A1(\pe6/bq[25] ), .A2(n58665), .ZN(n59056) );
  NAND2HSV0 U60953 ( .A1(n59054), .A2(n58449), .ZN(n59055) );
  XOR2HSV0 U60954 ( .A1(n59056), .A2(n59055), .Z(n59057) );
  XOR2HSV0 U60955 ( .A1(n59058), .A2(n59057), .Z(n59059) );
  XOR2HSV0 U60956 ( .A1(n59060), .A2(n59059), .Z(n59083) );
  NAND2HSV0 U60957 ( .A1(n59062), .A2(n59061), .ZN(n59064) );
  NAND2HSV0 U60958 ( .A1(\pe6/bq[8] ), .A2(\pe6/aot [23]), .ZN(n59063) );
  XOR2HSV0 U60959 ( .A1(n59064), .A2(n59063), .Z(n59070) );
  NAND2HSV0 U60960 ( .A1(n59066), .A2(n59065), .ZN(n59068) );
  NAND2HSV0 U60961 ( .A1(n59251), .A2(n58353), .ZN(n59067) );
  XOR2HSV0 U60962 ( .A1(n59068), .A2(n59067), .Z(n59069) );
  XOR2HSV0 U60963 ( .A1(n59070), .A2(n59069), .Z(n59081) );
  NAND2HSV0 U60964 ( .A1(n58731), .A2(n59272), .ZN(n59073) );
  NAND2HSV0 U60965 ( .A1(n59071), .A2(\pe6/aot [1]), .ZN(n59072) );
  XOR2HSV0 U60966 ( .A1(n59073), .A2(n59072), .Z(n59079) );
  NAND2HSV0 U60967 ( .A1(n59267), .A2(n58459), .ZN(n59077) );
  NAND2HSV0 U60968 ( .A1(n59075), .A2(n59074), .ZN(n59076) );
  XOR2HSV0 U60969 ( .A1(n59077), .A2(n59076), .Z(n59078) );
  XOR2HSV0 U60970 ( .A1(n59079), .A2(n59078), .Z(n59080) );
  XOR2HSV0 U60971 ( .A1(n59081), .A2(n59080), .Z(n59082) );
  XOR2HSV0 U60972 ( .A1(n59083), .A2(n59082), .Z(n59117) );
  NAND2HSV0 U60973 ( .A1(n59084), .A2(\pe6/aot [22]), .ZN(n59086) );
  NAND2HSV0 U60974 ( .A1(\pe6/bq[11] ), .A2(n59264), .ZN(n59085) );
  XOR2HSV0 U60975 ( .A1(n59086), .A2(n59085), .Z(n59093) );
  NAND2HSV0 U60976 ( .A1(n48038), .A2(n59087), .ZN(n59091) );
  NAND2HSV0 U60977 ( .A1(n59089), .A2(n59088), .ZN(n59090) );
  XOR2HSV0 U60978 ( .A1(n59091), .A2(n59090), .Z(n59092) );
  XOR2HSV0 U60979 ( .A1(n59093), .A2(n59092), .Z(n59104) );
  NOR2HSV0 U60980 ( .A1(n59094), .A2(n46637), .ZN(n59096) );
  NAND2HSV0 U60981 ( .A1(n58668), .A2(\pe6/aot [17]), .ZN(n59095) );
  XOR2HSV0 U60982 ( .A1(n59096), .A2(n59095), .Z(n59102) );
  NAND2HSV0 U60983 ( .A1(n59100), .A2(\pe6/aot [11]), .ZN(n59187) );
  XNOR2HSV1 U60984 ( .A1(n59102), .A2(n59101), .ZN(n59103) );
  XNOR2HSV1 U60985 ( .A1(n59104), .A2(n59103), .ZN(n59115) );
  NOR2HSV0 U60986 ( .A1(n59105), .A2(n44396), .ZN(n59198) );
  XOR2HSV0 U60987 ( .A1(n59111), .A2(n59110), .Z(n59112) );
  XNOR2HSV1 U60988 ( .A1(n59113), .A2(n59112), .ZN(n59114) );
  XNOR2HSV1 U60989 ( .A1(n59115), .A2(n59114), .ZN(n59116) );
  XNOR2HSV1 U60990 ( .A1(n59117), .A2(n59116), .ZN(n59118) );
  XOR3HSV2 U60991 ( .A1(n59120), .A2(n59119), .A3(n59118), .Z(n59123) );
  NAND2HSV0 U60992 ( .A1(n59121), .A2(\pe6/got [3]), .ZN(n59122) );
  XNOR2HSV1 U60993 ( .A1(n59123), .A2(n59122), .ZN(n59125) );
  CLKNAND2HSV1 U60994 ( .A1(n59295), .A2(n58479), .ZN(n59124) );
  XNOR2HSV1 U60995 ( .A1(n59125), .A2(n59124), .ZN(n59126) );
  XNOR2HSV1 U60996 ( .A1(n59127), .A2(n59126), .ZN(n59128) );
  XNOR2HSV1 U60997 ( .A1(n59129), .A2(n59128), .ZN(n59131) );
  NAND2HSV0 U60998 ( .A1(n59917), .A2(\pe6/got [7]), .ZN(n59130) );
  XNOR2HSV1 U60999 ( .A1(n59131), .A2(n59130), .ZN(n59132) );
  XNOR2HSV1 U61000 ( .A1(n59133), .A2(n59132), .ZN(n59134) );
  XNOR2HSV1 U61001 ( .A1(n59135), .A2(n59134), .ZN(n59136) );
  XNOR2HSV1 U61002 ( .A1(n59137), .A2(n59136), .ZN(n59138) );
  XNOR2HSV1 U61003 ( .A1(n59139), .A2(n59138), .ZN(n59140) );
  XNOR2HSV1 U61004 ( .A1(n59141), .A2(n59140), .ZN(n59142) );
  XNOR2HSV1 U61005 ( .A1(n59143), .A2(n59142), .ZN(n59146) );
  CLKNAND2HSV0 U61006 ( .A1(n59144), .A2(n49741), .ZN(n59145) );
  XNOR2HSV1 U61007 ( .A1(n59146), .A2(n59145), .ZN(n59147) );
  XNOR2HSV1 U61008 ( .A1(n59148), .A2(n59147), .ZN(n59149) );
  XNOR2HSV1 U61009 ( .A1(n59150), .A2(n59149), .ZN(n59151) );
  XNOR2HSV1 U61010 ( .A1(n59152), .A2(n59151), .ZN(n59153) );
  XNOR2HSV1 U61011 ( .A1(n59154), .A2(n59153), .ZN(n59156) );
  NAND2HSV0 U61012 ( .A1(n59915), .A2(n58807), .ZN(n59155) );
  XNOR2HSV1 U61013 ( .A1(n59156), .A2(n59155), .ZN(n59157) );
  XNOR2HSV1 U61014 ( .A1(n59158), .A2(n59157), .ZN(n59159) );
  XNOR2HSV1 U61015 ( .A1(n59160), .A2(n59159), .ZN(n59163) );
  CLKNAND2HSV0 U61016 ( .A1(n59161), .A2(n59175), .ZN(n59162) );
  XOR2HSV0 U61017 ( .A1(n59163), .A2(n59162), .Z(n59164) );
  NAND2HSV0 U61018 ( .A1(n59918), .A2(n59174), .ZN(n59334) );
  NAND2HSV0 U61019 ( .A1(n59680), .A2(n59175), .ZN(n59332) );
  NAND2HSV0 U61020 ( .A1(n59177), .A2(n59176), .ZN(n59327) );
  NAND2HSV0 U61021 ( .A1(n59916), .A2(n35922), .ZN(n59325) );
  NAND2HSV0 U61022 ( .A1(n58664), .A2(n36104), .ZN(n59323) );
  NAND2HSV0 U61023 ( .A1(n59179), .A2(n59178), .ZN(n59321) );
  CLKNAND2HSV0 U61024 ( .A1(n58722), .A2(\pe6/got [15]), .ZN(n59315) );
  NAND2HSV0 U61025 ( .A1(n59033), .A2(n58810), .ZN(n59313) );
  NAND2HSV0 U61026 ( .A1(n59363), .A2(n59180), .ZN(n59309) );
  NAND2HSV0 U61027 ( .A1(n32165), .A2(n59181), .ZN(n59307) );
  NAND2HSV0 U61028 ( .A1(n26109), .A2(\pe6/got [10]), .ZN(n59305) );
  NAND2HSV0 U61029 ( .A1(n59678), .A2(n59182), .ZN(n59301) );
  NAND2HSV0 U61030 ( .A1(n59183), .A2(n58562), .ZN(n59299) );
  NAND2HSV0 U61031 ( .A1(n59594), .A2(n46173), .ZN(n59185) );
  NAND2HSV0 U61032 ( .A1(n32286), .A2(n58527), .ZN(n59184) );
  XOR2HSV0 U61033 ( .A1(n59185), .A2(n59184), .Z(n59291) );
  XOR2HSV0 U61034 ( .A1(n59187), .A2(n59186), .Z(n59213) );
  CLKNHSV0 U61035 ( .I(n59188), .ZN(n59192) );
  AOI22HSV0 U61036 ( .A1(\pe6/bq[17] ), .A2(n59189), .B1(\pe6/aot [19]), .B2(
        n58668), .ZN(n59190) );
  AOI21HSV0 U61037 ( .A1(n59192), .A2(n59191), .B(n59190), .ZN(n59200) );
  NOR2HSV0 U61038 ( .A1(n59194), .A2(n59193), .ZN(n59197) );
  OAI22HSV0 U61039 ( .A1(n59198), .A2(n59197), .B1(n59196), .B2(n59195), .ZN(
        n59199) );
  XOR2HSV0 U61040 ( .A1(n59200), .A2(n59199), .Z(n59212) );
  NAND2HSV0 U61041 ( .A1(n59201), .A2(\pe6/pq ), .ZN(n59204) );
  NAND2HSV0 U61042 ( .A1(n59202), .A2(n58488), .ZN(n59203) );
  XOR2HSV0 U61043 ( .A1(n59204), .A2(n59203), .Z(n59210) );
  NOR2HSV0 U61044 ( .A1(n59205), .A2(n49188), .ZN(n59208) );
  NAND2HSV0 U61045 ( .A1(n59206), .A2(n35632), .ZN(n59207) );
  XOR2HSV0 U61046 ( .A1(n59208), .A2(n59207), .Z(n59209) );
  XOR2HSV0 U61047 ( .A1(n59210), .A2(n59209), .Z(n59211) );
  XOR3HSV2 U61048 ( .A1(n59213), .A2(n59212), .A3(n59211), .Z(n59289) );
  NAND2HSV0 U61049 ( .A1(n58405), .A2(n32588), .ZN(n59215) );
  NAND2HSV0 U61050 ( .A1(n58833), .A2(\pe6/aot [17]), .ZN(n59214) );
  XOR2HSV0 U61051 ( .A1(n59215), .A2(n59214), .Z(n59221) );
  NAND2HSV0 U61052 ( .A1(n59216), .A2(n59040), .ZN(n59219) );
  NAND2HSV0 U61053 ( .A1(n59217), .A2(\pe6/aot [7]), .ZN(n59218) );
  XOR2HSV0 U61054 ( .A1(n59219), .A2(n59218), .Z(n59220) );
  XOR2HSV0 U61055 ( .A1(n59221), .A2(n59220), .Z(n59230) );
  NAND2HSV0 U61056 ( .A1(n33005), .A2(\pe6/aot [13]), .ZN(n59223) );
  NAND2HSV0 U61057 ( .A1(n58452), .A2(n58991), .ZN(n59222) );
  XOR2HSV0 U61058 ( .A1(n59223), .A2(n59222), .Z(n59228) );
  NAND2HSV0 U61059 ( .A1(n46210), .A2(n49831), .ZN(n59226) );
  NAND2HSV0 U61060 ( .A1(n59224), .A2(n49208), .ZN(n59225) );
  XOR2HSV0 U61061 ( .A1(n59226), .A2(n59225), .Z(n59227) );
  XNOR2HSV1 U61062 ( .A1(n59228), .A2(n59227), .ZN(n59229) );
  XNOR2HSV1 U61063 ( .A1(n59230), .A2(n59229), .ZN(n59233) );
  NAND2HSV0 U61064 ( .A1(n44426), .A2(n59231), .ZN(n59232) );
  XNOR2HSV1 U61065 ( .A1(n59233), .A2(n59232), .ZN(n59288) );
  NAND2HSV0 U61066 ( .A1(n49106), .A2(n59234), .ZN(n59238) );
  NAND2HSV0 U61067 ( .A1(n59236), .A2(n59235), .ZN(n59237) );
  XOR2HSV0 U61068 ( .A1(n59238), .A2(n59237), .Z(n59244) );
  NAND2HSV0 U61069 ( .A1(\pe6/bq[9] ), .A2(n59239), .ZN(n59242) );
  NAND2HSV0 U61070 ( .A1(n59240), .A2(\pe6/aot [21]), .ZN(n59241) );
  XOR2HSV0 U61071 ( .A1(n59242), .A2(n59241), .Z(n59243) );
  XOR2HSV0 U61072 ( .A1(n59244), .A2(n59243), .Z(n59258) );
  NAND2HSV0 U61073 ( .A1(n59246), .A2(n59245), .ZN(n59249) );
  NAND2HSV0 U61074 ( .A1(n59247), .A2(n58459), .ZN(n59248) );
  XOR2HSV0 U61075 ( .A1(n59249), .A2(n59248), .Z(n59256) );
  NAND2HSV0 U61076 ( .A1(n59251), .A2(n59250), .ZN(n59254) );
  NAND2HSV0 U61077 ( .A1(n35740), .A2(n59252), .ZN(n59253) );
  XOR2HSV0 U61078 ( .A1(n59254), .A2(n59253), .Z(n59255) );
  XOR2HSV0 U61079 ( .A1(n59256), .A2(n59255), .Z(n59257) );
  XOR2HSV0 U61080 ( .A1(n59258), .A2(n59257), .Z(n59286) );
  NAND2HSV0 U61081 ( .A1(n59259), .A2(\pe6/aot [1]), .ZN(n59263) );
  NAND2HSV0 U61082 ( .A1(n59261), .A2(n59260), .ZN(n59262) );
  XOR2HSV0 U61083 ( .A1(n59263), .A2(n59262), .Z(n59271) );
  NAND2HSV0 U61084 ( .A1(n59265), .A2(n59264), .ZN(n59269) );
  NAND2HSV0 U61085 ( .A1(n59267), .A2(n59266), .ZN(n59268) );
  XOR2HSV0 U61086 ( .A1(n59269), .A2(n59268), .Z(n59270) );
  XOR2HSV0 U61087 ( .A1(n59271), .A2(n59270), .Z(n59284) );
  NAND2HSV0 U61088 ( .A1(n59273), .A2(n59272), .ZN(n59275) );
  NAND2HSV0 U61089 ( .A1(n58962), .A2(n36153), .ZN(n59274) );
  XOR2HSV0 U61090 ( .A1(n59275), .A2(n59274), .Z(n59282) );
  NAND2HSV0 U61091 ( .A1(n59277), .A2(n59276), .ZN(n59280) );
  NAND2HSV0 U61092 ( .A1(\pe6/bq[2] ), .A2(n59278), .ZN(n59279) );
  XOR2HSV0 U61093 ( .A1(n59280), .A2(n59279), .Z(n59281) );
  XOR2HSV0 U61094 ( .A1(n59282), .A2(n59281), .Z(n59283) );
  XOR2HSV0 U61095 ( .A1(n59284), .A2(n59283), .Z(n59285) );
  XOR2HSV0 U61096 ( .A1(n59286), .A2(n59285), .Z(n59287) );
  XOR3HSV2 U61097 ( .A1(n59289), .A2(n59288), .A3(n59287), .Z(n59290) );
  XOR2HSV0 U61098 ( .A1(n59291), .A2(n59290), .Z(n59294) );
  NAND2HSV0 U61099 ( .A1(n59670), .A2(n59292), .ZN(n59293) );
  XNOR2HSV1 U61100 ( .A1(n59294), .A2(n59293), .ZN(n59297) );
  CLKNAND2HSV1 U61101 ( .A1(n59295), .A2(n58723), .ZN(n59296) );
  XNOR2HSV1 U61102 ( .A1(n59297), .A2(n59296), .ZN(n59298) );
  XNOR2HSV1 U61103 ( .A1(n59299), .A2(n59298), .ZN(n59300) );
  XNOR2HSV1 U61104 ( .A1(n59301), .A2(n59300), .ZN(n59303) );
  NAND2HSV0 U61105 ( .A1(n59917), .A2(n59037), .ZN(n59302) );
  XNOR2HSV1 U61106 ( .A1(n59303), .A2(n59302), .ZN(n59304) );
  XNOR2HSV1 U61107 ( .A1(n59305), .A2(n59304), .ZN(n59306) );
  XNOR2HSV1 U61108 ( .A1(n59307), .A2(n59306), .ZN(n59308) );
  XNOR2HSV1 U61109 ( .A1(n59309), .A2(n59308), .ZN(n59310) );
  XOR2HSV0 U61110 ( .A1(n59311), .A2(n59310), .Z(n59312) );
  XNOR2HSV1 U61111 ( .A1(n59313), .A2(n59312), .ZN(n59314) );
  XNOR2HSV1 U61112 ( .A1(n59315), .A2(n59314), .ZN(n59319) );
  NAND2HSV0 U61113 ( .A1(n59317), .A2(n59316), .ZN(n59318) );
  XNOR2HSV1 U61114 ( .A1(n59319), .A2(n59318), .ZN(n59320) );
  XNOR2HSV1 U61115 ( .A1(n59321), .A2(n59320), .ZN(n59322) );
  XNOR2HSV1 U61116 ( .A1(n59323), .A2(n59322), .ZN(n59324) );
  XNOR2HSV1 U61117 ( .A1(n59325), .A2(n59324), .ZN(n59326) );
  XNOR2HSV1 U61118 ( .A1(n59327), .A2(n59326), .ZN(n59330) );
  NAND2HSV0 U61119 ( .A1(n59915), .A2(n59328), .ZN(n59329) );
  XNOR2HSV1 U61120 ( .A1(n59330), .A2(n59329), .ZN(n59331) );
  XNOR2HSV1 U61121 ( .A1(n59332), .A2(n59331), .ZN(n59333) );
  XNOR2HSV1 U61122 ( .A1(n59334), .A2(n59333), .ZN(n59337) );
  NAND2HSV0 U61123 ( .A1(n59335), .A2(n32970), .ZN(n59336) );
endmodule

