
module topcell ( clk, ctr, rst, ai, gi, bi, po );
  input [8:1] ai;
  input [8:1] gi;
  input [8:1] bi;
  output [1:8] po;
  input clk, ctr, rst;
  wire   po1, ctro1, po2, ctro2, po3, ctro3, po4, ctro4, po5, ctro5, po6,
         ctro6, \pov7[5] , po7, ctro7, po8, ctro8, po9, ctro9, po10, ctro10,
         po11, ctro11, po12, ctro12, po13, ctro13, \pov14[7] , po14, ctro14,
         \pov15[4] , po15, ctro15, po16, ctro16, po17, ctro17, po18, ctro18,
         \pov19[7] , po19, ctro19, po20, ctro20, po21, ctro21, \pe1/ti_7[7] ,
         \pe1/ti_7[6] , \pe1/ti_7[5] , \pe1/ti_7[3] , \pe1/ti_7[2] ,
         \pe1/bq[1] , \pe1/bq[2] , \pe1/bq[3] , \pe1/bq[4] , \pe1/bq[5] ,
         \pe1/bq[6] , \pe1/bq[7] , \pe1/bq[8] , \pe1/ctrq , \pe2/ti_7[5] ,
         \pe2/ti_7[3] , \pe2/ti_7[1] , \pe2/ti_1 , \pe2/ti_1t , \pe2/bq[1] ,
         \pe2/bq[2] , \pe2/bq[3] , \pe2/bq[4] , \pe2/bq[5] , \pe2/bq[6] ,
         \pe2/bq[7] , \pe2/bq[8] , \pe2/ctrq , \pe2/pq , \pe3/ti_7[5] ,
         \pe3/ti_7[1] , \pe3/ti_1 , \pe3/ti_1t , \pe3/bq[1] , \pe3/bq[2] ,
         \pe3/bq[3] , \pe3/bq[4] , \pe3/bq[5] , \pe3/bq[6] , \pe3/bq[7] ,
         \pe3/bq[8] , \pe3/ctrq , \pe3/pq , \pe4/ti_7[1] , \pe4/ti_1 ,
         \pe4/ti_1t , \pe4/bq[1] , \pe4/bq[2] , \pe4/bq[3] , \pe4/bq[4] ,
         \pe4/bq[5] , \pe4/bq[6] , \pe4/bq[7] , \pe4/bq[8] , \pe4/bqt[7] ,
         \pe4/ctrq , \pe4/pq , \pe5/ti_7[7] , \pe5/ti_1 , \pe5/ti_1t ,
         \pe5/bq[1] , \pe5/bq[2] , \pe5/bq[3] , \pe5/bq[4] , \pe5/bq[5] ,
         \pe5/bq[6] , \pe5/bq[7] , \pe5/bq[8] , \pe5/ctrq , \pe5/pq ,
         \pe6/ti_7[5] , \pe6/ti_1 , \pe6/ti_1t , \pe6/bq[1] , \pe6/bq[2] ,
         \pe6/bq[3] , \pe6/bq[4] , \pe6/bq[5] , \pe6/bq[6] , \pe6/bq[7] ,
         \pe6/bq[8] , \pe6/ctrq , \pe6/pq , \pe7/ti_7[5] , \pe7/ti_7[1] ,
         \pe7/ti_1 , \pe7/ti_1t , \pe7/bq[1] , \pe7/bq[2] , \pe7/bq[3] ,
         \pe7/bq[4] , \pe7/bq[5] , \pe7/bq[6] , \pe7/bq[7] , \pe7/bq[8] ,
         \pe7/ctrq , \pe7/pq , \pe8/ti_7[1] , \pe8/ti_1 , \pe8/ti_1t ,
         \pe8/bq[1] , \pe8/bq[2] , \pe8/bq[3] , \pe8/bq[4] , \pe8/bq[5] ,
         \pe8/bq[6] , \pe8/bq[7] , \pe8/bq[8] , \pe8/ctrq , \pe8/pq ,
         \pe9/ti_7[1] , \pe9/ti_1 , \pe9/ti_1t , \pe9/bq[1] , \pe9/bq[2] ,
         \pe9/bq[3] , \pe9/bq[4] , \pe9/bq[5] , \pe9/bq[6] , \pe9/bq[7] ,
         \pe9/bq[8] , \pe9/ctrq , \pe9/pq , \pe10/ti_7[6] , \pe10/ti_7[5] ,
         \pe10/ti_1 , \pe10/ti_1t , \pe10/bq[1] , \pe10/bq[2] , \pe10/bq[3] ,
         \pe10/bq[4] , \pe10/bq[5] , \pe10/bq[6] , \pe10/bq[7] , \pe10/bq[8] ,
         \pe10/ctrq , \pe10/pq , \pe11/ti_7[5] , \pe11/ti_7[1] , \pe11/ti_1 ,
         \pe11/ti_1t , \pe11/bq[1] , \pe11/bq[2] , \pe11/bq[3] , \pe11/bq[4] ,
         \pe11/bq[5] , \pe11/bq[6] , \pe11/bq[7] , \pe11/bq[8] , \pe11/ctrq ,
         \pe11/pq , \pe12/ti_7[3] , \pe12/ti_7[1] , \pe12/ti_1 , \pe12/ti_1t ,
         \pe12/bq[1] , \pe12/bq[2] , \pe12/bq[3] , \pe12/bq[4] , \pe12/bq[5] ,
         \pe12/bq[6] , \pe12/bq[7] , \pe12/bq[8] , \pe12/ctrq , \pe12/pq ,
         \pe13/ti_7[4] , \pe13/ti_7[1] , \pe13/ti_1 , \pe13/ti_1t ,
         \pe13/bq[1] , \pe13/bq[2] , \pe13/bq[3] , \pe13/bq[4] , \pe13/bq[5] ,
         \pe13/bq[6] , \pe13/bq[7] , \pe13/bq[8] , \pe13/ctrq , \pe13/pq ,
         \pe14/ti_7[5] , \pe14/ti_7[3] , \pe14/ti_1 , \pe14/ti_1t ,
         \pe14/bq[1] , \pe14/bq[2] , \pe14/bq[3] , \pe14/bq[4] , \pe14/bq[5] ,
         \pe14/bq[6] , \pe14/bq[7] , \pe14/bq[8] , \pe14/ctrq , \pe14/pq ,
         \pe15/ti_7[5] , \pe15/ti_7[3] , \pe15/ti_1 , \pe15/ti_1t ,
         \pe15/bq[1] , \pe15/bq[2] , \pe15/bq[3] , \pe15/bq[4] , \pe15/bq[5] ,
         \pe15/bq[6] , \pe15/bq[7] , \pe15/bq[8] , \pe15/ctrq , \pe15/pq ,
         \pe16/ti_7[7] , \pe16/ti_7[3] , \pe16/ti_7[1] , \pe16/ti_1 ,
         \pe16/ti_1t , \pe16/bq[1] , \pe16/bq[2] , \pe16/bq[3] , \pe16/bq[4] ,
         \pe16/bq[5] , \pe16/bq[6] , \pe16/bq[7] , \pe16/bq[8] , \pe16/ctrq ,
         \pe16/pq , \pe17/ti_7[7] , \pe17/ti_7[3] , \pe17/ti_7[1] ,
         \pe17/ti_1 , \pe17/ti_1t , \pe17/bq[1] , \pe17/bq[2] , \pe17/bq[3] ,
         \pe17/bq[4] , \pe17/bq[5] , \pe17/bq[6] , \pe17/bq[7] , \pe17/bq[8] ,
         \pe17/ctrq , \pe17/pq , \pe18/ti_7[5] , \pe18/ti_7[1] , \pe18/ti_1 ,
         \pe18/ti_1t , \pe18/bq[1] , \pe18/bq[2] , \pe18/bq[3] , \pe18/bq[4] ,
         \pe18/bq[5] , \pe18/bq[6] , \pe18/bq[7] , \pe18/bq[8] , \pe18/ctrq ,
         \pe18/pq , \pe19/ti_7[1] , \pe19/ti_1 , \pe19/ti_1t , \pe19/bq[1] ,
         \pe19/bq[2] , \pe19/bq[3] , \pe19/bq[4] , \pe19/bq[5] , \pe19/bq[6] ,
         \pe19/bq[7] , \pe19/bq[8] , \pe19/ctrq , \pe19/pq , \pe20/ti_7[5] ,
         \pe20/ti_1 , \pe20/ti_1t , \pe20/bq[1] , \pe20/bq[2] , \pe20/bq[3] ,
         \pe20/bq[4] , \pe20/bq[5] , \pe20/bq[6] , \pe20/bq[7] , \pe20/bq[8] ,
         \pe20/ctrq , \pe20/pq , \pe21/ti_7[5] , \pe21/ti_7[3] ,
         \pe21/ti_7[1] , \pe21/ti_1 , \pe21/ti_1t , \pe21/bq[1] , \pe21/bq[2] ,
         \pe21/bq[3] , \pe21/bq[4] , \pe21/bq[5] , \pe21/bq[6] , \pe21/bq[7] ,
         \pe21/bq[8] , \pe21/ctrq , \pe21/pq , n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295;
  wire   [8:1] ao1;
  wire   [8:1] go1;
  wire   [8:1] bo1;
  wire   [1:7] poh1;
  wire   [1:7] pov1;
  wire   [8:1] ao2;
  wire   [8:1] go2;
  wire   [8:1] bo2;
  wire   [1:7] poh2;
  wire   [8:1] ao3;
  wire   [8:1] go3;
  wire   [8:1] bo3;
  wire   [1:7] poh3;
  wire   [8:1] ao4;
  wire   [8:1] go4;
  wire   [8:1] bo4;
  wire   [1:7] poh4;
  wire   [8:1] ao5;
  wire   [8:1] go5;
  wire   [8:1] bo5;
  wire   [1:7] poh5;
  wire   [8:1] ao6;
  wire   [8:1] go6;
  wire   [8:1] bo6;
  wire   [1:7] poh6;
  wire   [8:1] ao7;
  wire   [8:1] go7;
  wire   [8:1] bo7;
  wire   [1:7] poh7;
  wire   [8:1] ao8;
  wire   [8:1] go8;
  wire   [8:1] bo8;
  wire   [1:7] poh8;
  wire   [8:1] ao9;
  wire   [8:1] go9;
  wire   [8:1] bo9;
  wire   [1:7] poh9;
  wire   [1:7] pov9;
  wire   [8:1] ao10;
  wire   [8:1] go10;
  wire   [8:1] bo10;
  wire   [1:7] poh10;
  wire   [8:1] ao11;
  wire   [8:1] go11;
  wire   [8:1] bo11;
  wire   [1:7] poh11;
  wire   [8:1] ao12;
  wire   [8:1] go12;
  wire   [8:1] bo12;
  wire   [1:7] poh12;
  wire   [8:1] ao13;
  wire   [8:1] go13;
  wire   [8:1] bo13;
  wire   [1:7] poh13;
  wire   [8:1] ao14;
  wire   [8:1] go14;
  wire   [8:1] bo14;
  wire   [1:7] poh14;
  wire   [8:1] ao15;
  wire   [8:1] go15;
  wire   [8:1] bo15;
  wire   [1:7] poh15;
  wire   [8:1] ao16;
  wire   [8:1] go16;
  wire   [8:1] bo16;
  wire   [1:7] poh16;
  wire   [8:1] ao17;
  wire   [8:1] go17;
  wire   [8:1] bo17;
  wire   [1:7] poh17;
  wire   [8:1] ao18;
  wire   [8:1] go18;
  wire   [8:1] bo18;
  wire   [1:7] poh18;
  wire   [8:1] ao19;
  wire   [8:1] go19;
  wire   [8:1] bo19;
  wire   [1:7] poh19;
  wire   [8:1] ao20;
  wire   [8:1] go20;
  wire   [8:1] bo20;
  wire   [1:7] poh20;
  wire   [8:1] bo21;
  wire   [1:7] poh21;
  wire   [1:7] \pe1/poht ;
  wire   [8:1] \pe1/got ;
  wire   [8:1] \pe1/aot ;
  wire   [1:7] \pe1/ti_7t ;
  wire   [1:7] \pe2/poht ;
  wire   [8:1] \pe2/got ;
  wire   [8:1] \pe2/aot ;
  wire   [1:7] \pe2/ti_7t ;
  wire   [1:7] \pe2/phq ;
  wire   [1:7] \pe2/pvq ;
  wire   [1:7] \pe3/poht ;
  wire   [8:1] \pe3/got ;
  wire   [8:1] \pe3/aot ;
  wire   [1:7] \pe3/ti_7t ;
  wire   [1:7] \pe3/phq ;
  wire   [1:7] \pe3/pvq ;
  wire   [1:7] \pe4/poht ;
  wire   [8:1] \pe4/got ;
  wire   [8:1] \pe4/aot ;
  wire   [1:7] \pe4/ti_7t ;
  wire   [1:7] \pe4/phq ;
  wire   [1:7] \pe4/pvq ;
  wire   [1:7] \pe5/poht ;
  wire   [8:1] \pe5/got ;
  wire   [8:1] \pe5/aot ;
  wire   [1:7] \pe5/ti_7t ;
  wire   [1:7] \pe5/phq ;
  wire   [1:7] \pe5/pvq ;
  wire   [1:7] \pe6/poht ;
  wire   [8:1] \pe6/got ;
  wire   [8:1] \pe6/aot ;
  wire   [1:7] \pe6/ti_7t ;
  wire   [1:7] \pe6/phq ;
  wire   [1:7] \pe6/pvq ;
  wire   [1:7] \pe7/poht ;
  wire   [8:1] \pe7/got ;
  wire   [8:1] \pe7/aot ;
  wire   [1:7] \pe7/ti_7t ;
  wire   [1:7] \pe7/phq ;
  wire   [1:7] \pe7/pvq ;
  wire   [1:7] \pe8/poht ;
  wire   [8:1] \pe8/got ;
  wire   [8:1] \pe8/aot ;
  wire   [1:7] \pe8/ti_7t ;
  wire   [1:7] \pe8/phq ;
  wire   [1:7] \pe8/pvq ;
  wire   [1:7] \pe9/poht ;
  wire   [8:1] \pe9/got ;
  wire   [8:1] \pe9/aot ;
  wire   [1:7] \pe9/ti_7t ;
  wire   [1:7] \pe9/phq ;
  wire   [1:7] \pe9/pvq ;
  wire   [1:7] \pe10/poht ;
  wire   [8:1] \pe10/got ;
  wire   [8:1] \pe10/aot ;
  wire   [1:7] \pe10/ti_7t ;
  wire   [1:7] \pe10/phq ;
  wire   [1:7] \pe10/pvq ;
  wire   [1:7] \pe11/poht ;
  wire   [8:1] \pe11/got ;
  wire   [8:1] \pe11/aot ;
  wire   [1:7] \pe11/ti_7t ;
  wire   [1:7] \pe11/phq ;
  wire   [1:7] \pe11/pvq ;
  wire   [1:7] \pe12/poht ;
  wire   [8:1] \pe12/got ;
  wire   [8:1] \pe12/aot ;
  wire   [1:7] \pe12/ti_7t ;
  wire   [1:7] \pe12/phq ;
  wire   [1:7] \pe12/pvq ;
  wire   [1:7] \pe13/poht ;
  wire   [8:1] \pe13/got ;
  wire   [8:1] \pe13/aot ;
  wire   [1:7] \pe13/ti_7t ;
  wire   [1:7] \pe13/phq ;
  wire   [1:7] \pe13/pvq ;
  wire   [1:7] \pe14/poht ;
  wire   [8:1] \pe14/got ;
  wire   [8:1] \pe14/aot ;
  wire   [1:7] \pe14/ti_7t ;
  wire   [1:7] \pe14/phq ;
  wire   [1:7] \pe14/pvq ;
  wire   [1:7] \pe15/poht ;
  wire   [8:1] \pe15/got ;
  wire   [8:1] \pe15/aot ;
  wire   [1:7] \pe15/ti_7t ;
  wire   [1:7] \pe15/phq ;
  wire   [1:7] \pe15/pvq ;
  wire   [1:7] \pe16/poht ;
  wire   [8:1] \pe16/got ;
  wire   [8:1] \pe16/aot ;
  wire   [1:7] \pe16/ti_7t ;
  wire   [1:7] \pe16/phq ;
  wire   [1:7] \pe16/pvq ;
  wire   [1:7] \pe17/poht ;
  wire   [8:1] \pe17/got ;
  wire   [8:1] \pe17/aot ;
  wire   [1:7] \pe17/ti_7t ;
  wire   [1:7] \pe17/phq ;
  wire   [1:7] \pe17/pvq ;
  wire   [1:7] \pe18/poht ;
  wire   [8:1] \pe18/got ;
  wire   [8:1] \pe18/aot ;
  wire   [1:7] \pe18/ti_7t ;
  wire   [1:7] \pe18/phq ;
  wire   [1:7] \pe18/pvq ;
  wire   [1:7] \pe19/poht ;
  wire   [8:1] \pe19/got ;
  wire   [8:1] \pe19/aot ;
  wire   [1:7] \pe19/ti_7t ;
  wire   [1:7] \pe19/phq ;
  wire   [1:7] \pe19/pvq ;
  wire   [1:7] \pe20/poht ;
  wire   [8:1] \pe20/got ;
  wire   [8:1] \pe20/aot ;
  wire   [1:7] \pe20/ti_7t ;
  wire   [1:7] \pe20/phq ;
  wire   [1:7] \pe20/pvq ;
  wire   [1:7] \pe21/poht ;
  wire   [8:1] \pe21/got ;
  wire   [8:1] \pe21/aot ;
  wire   [1:7] \pe21/ti_7t ;
  wire   [1:7] \pe21/phq ;
  wire   [1:7] \pe21/pvq ;

  DRNQHSV4 \pe1/delaycell1/q_reg[8]  ( .D(ai[1]), .CK(clk), .RDN(n14832), .Q(
        \pe1/aot [1]) );
  DRNQHSV4 \pe1/delaycell1/q_reg[7]  ( .D(ai[2]), .CK(clk), .RDN(n14801), .Q(
        \pe1/aot [2]) );
  DRNQHSV4 \pe1/delaycell1/q_reg[6]  ( .D(ai[3]), .CK(clk), .RDN(rst), .Q(
        \pe1/aot [3]) );
  DRNQHSV4 \pe1/delaycell1/q_reg[5]  ( .D(ai[4]), .CK(clk), .RDN(n14789), .Q(
        \pe1/aot [4]) );
  DRNQHSV4 \pe1/delaycell1/q_reg[4]  ( .D(ai[5]), .CK(clk), .RDN(n14726), .Q(
        \pe1/aot [5]) );
  DRNQHSV4 \pe1/delaycell1/q_reg[2]  ( .D(ai[7]), .CK(clk), .RDN(n15173), .Q(
        \pe1/aot [7]) );
  DRNQHSV4 \pe1/delaycell2/q_reg[6]  ( .D(gi[3]), .CK(clk), .RDN(n14801), .Q(
        \pe1/got [3]) );
  DRNQHSV4 \pe1/delaycell2/q_reg[5]  ( .D(gi[4]), .CK(clk), .RDN(rst), .Q(
        \pe1/got [4]) );
  DRNQHSV4 \pe1/delaycell2/q_reg[4]  ( .D(gi[5]), .CK(clk), .RDN(rst), .Q(
        \pe1/got [5]) );
  DRNQHSV4 \pe1/delaycell2/q_reg[3]  ( .D(gi[6]), .CK(clk), .RDN(rst), .Q(
        \pe1/got [6]) );
  DRNQHSV4 \pe1/delaycell2/q_reg[2]  ( .D(gi[7]), .CK(clk), .RDN(rst), .Q(
        \pe1/got [7]) );
  DRNQHSV4 \pe1/delaycell2/q_reg[1]  ( .D(gi[8]), .CK(clk), .RDN(n14807), .Q(
        \pe1/got [8]) );
  DRNQHSV4 \pe1/delaycell8/q_reg  ( .D(\pe1/ctrq ), .CK(clk), .RDN(n14719), 
        .Q(ctro1) );
  DRNQHSV4 \pe1/delaycell19/q_reg[7]  ( .D(n14967), .CK(clk), .RDN(n14755), 
        .Q(\pe1/bq[2] ) );
  DRNQHSV4 \pe1/delaycell19/q_reg[6]  ( .D(n15008), .CK(clk), .RDN(n14729), 
        .Q(\pe1/bq[3] ) );
  DRNQHSV4 \pe1/delaycell19/q_reg[5]  ( .D(n14971), .CK(clk), .RDN(n14766), 
        .Q(\pe1/bq[4] ) );
  DRNQHSV4 \pe1/delaycell19/q_reg[4]  ( .D(n14997), .CK(clk), .RDN(n14766), 
        .Q(\pe1/bq[5] ) );
  DRNQHSV4 \pe1/delaycell19/q_reg[3]  ( .D(n15064), .CK(clk), .RDN(n14764), 
        .Q(\pe1/bq[6] ) );
  DRNQHSV4 \pe1/delaycell19/q_reg[2]  ( .D(n14975), .CK(clk), .RDN(n14797), 
        .Q(\pe1/bq[7] ) );
  DRNQHSV4 \pe1/delaycell19/q_reg[1]  ( .D(n14974), .CK(clk), .RDN(n14718), 
        .Q(\pe1/bq[8] ) );
  DRNQHSV4 \pe1/delaycell21/q_reg[3]  ( .D(\pe1/ti_7[3] ), .CK(clk), .RDN(
        n14871), .Q(\pe1/ti_7t [3]) );
  DRNQHSV4 \pe2/delaycell1/q_reg[8]  ( .D(ao1[1]), .CK(clk), .RDN(n14723), .Q(
        \pe2/aot [1]) );
  DRNQHSV4 \pe2/delaycell1/q_reg[7]  ( .D(ao1[2]), .CK(clk), .RDN(n14718), .Q(
        \pe2/aot [2]) );
  DRNQHSV4 \pe2/delaycell1/q_reg[6]  ( .D(ao1[3]), .CK(clk), .RDN(n14745), .Q(
        \pe2/aot [3]) );
  DRNQHSV4 \pe2/delaycell1/q_reg[5]  ( .D(ao1[4]), .CK(clk), .RDN(n14786), .Q(
        \pe2/aot [4]) );
  DRNQHSV4 \pe2/delaycell1/q_reg[4]  ( .D(ao1[5]), .CK(clk), .RDN(n14778), .Q(
        \pe2/aot [5]) );
  DRNQHSV4 \pe2/delaycell1/q_reg[3]  ( .D(ao1[6]), .CK(clk), .RDN(n14720), .Q(
        \pe2/aot [6]) );
  DRNQHSV4 \pe2/delaycell1/q_reg[2]  ( .D(ao1[7]), .CK(clk), .RDN(n14720), .Q(
        \pe2/aot [7]) );
  DRNQHSV4 \pe2/delaycell1/q_reg[1]  ( .D(ao1[8]), .CK(clk), .RDN(n14814), .Q(
        \pe2/aot [8]) );
  DRNQHSV4 \pe2/delaycell2/q_reg[8]  ( .D(go1[1]), .CK(clk), .RDN(n14800), .Q(
        \pe2/got [1]) );
  DRNQHSV4 \pe2/delaycell2/q_reg[7]  ( .D(go1[2]), .CK(clk), .RDN(n14757), .Q(
        \pe2/got [2]) );
  DRNQHSV4 \pe2/delaycell2/q_reg[6]  ( .D(go1[3]), .CK(clk), .RDN(n14747), .Q(
        \pe2/got [3]) );
  DRNQHSV4 \pe2/delaycell2/q_reg[5]  ( .D(go1[4]), .CK(clk), .RDN(n14756), .Q(
        \pe2/got [4]) );
  DRNQHSV4 \pe2/delaycell2/q_reg[4]  ( .D(go1[5]), .CK(clk), .RDN(n15173), .Q(
        \pe2/got [5]) );
  DRNQHSV4 \pe2/delaycell2/q_reg[2]  ( .D(go1[7]), .CK(clk), .RDN(n14714), .Q(
        \pe2/got [7]) );
  DRNQHSV4 \pe2/delaycell2/q_reg[1]  ( .D(go1[8]), .CK(clk), .RDN(n14726), .Q(
        \pe2/got [8]) );
  DRNQHSV4 \pe2/delaycell5/q_reg[6]  ( .D(pov1[6]), .CK(clk), .RDN(n14721), 
        .Q(\pe2/pvq [6]) );
  DRNQHSV4 \pe2/delaycell5/q_reg[4]  ( .D(n15295), .CK(clk), .RDN(n14720), .Q(
        \pe2/pvq [4]) );
  DRNQHSV4 \pe2/delaycell5/q_reg[2]  ( .D(pov1[2]), .CK(clk), .RDN(n14716), 
        .Q(\pe2/pvq [2]) );
  DRNQHSV4 \pe2/delaycell5/q_reg[1]  ( .D(n14956), .CK(clk), .RDN(n14732), .Q(
        \pe2/pvq [1]) );
  DRNQHSV4 \pe2/delaycell6/q_reg[7]  ( .D(poh1[7]), .CK(clk), .RDN(n14796), 
        .Q(\pe2/phq [7]) );
  DRNQHSV4 \pe2/delaycell6/q_reg[6]  ( .D(poh1[6]), .CK(clk), .RDN(n14796), 
        .Q(\pe2/phq [6]) );
  DRNQHSV4 \pe2/delaycell6/q_reg[5]  ( .D(poh1[5]), .CK(clk), .RDN(n14765), 
        .Q(\pe2/phq [5]) );
  DRNQHSV4 \pe2/delaycell6/q_reg[4]  ( .D(poh1[4]), .CK(clk), .RDN(n14717), 
        .Q(\pe2/phq [4]) );
  DRNQHSV4 \pe2/delaycell6/q_reg[3]  ( .D(poh1[3]), .CK(clk), .RDN(n14773), 
        .Q(\pe2/phq [3]) );
  DRNQHSV4 \pe2/delaycell6/q_reg[2]  ( .D(poh1[2]), .CK(clk), .RDN(n14774), 
        .Q(\pe2/phq [2]) );
  DRNQHSV4 \pe2/delaycell6/q_reg[1]  ( .D(poh1[1]), .CK(clk), .RDN(n14871), 
        .Q(\pe2/phq [1]) );
  DRNQHSV4 \pe2/delaycell7/q_reg  ( .D(n14868), .CK(clk), .RDN(n14749), .Q(
        \pe2/ctrq ) );
  DRNQHSV4 \pe2/delaycell19/q_reg[8]  ( .D(n14983), .CK(clk), .RDN(n14787), 
        .Q(\pe2/bq[1] ) );
  DRNQHSV4 \pe2/delaycell19/q_reg[7]  ( .D(n14999), .CK(clk), .RDN(n14744), 
        .Q(\pe2/bq[2] ) );
  DRNQHSV4 \pe2/delaycell19/q_reg[6]  ( .D(n14966), .CK(clk), .RDN(n14757), 
        .Q(\pe2/bq[3] ) );
  DRNQHSV4 \pe2/delaycell19/q_reg[5]  ( .D(n14970), .CK(clk), .RDN(n14794), 
        .Q(\pe2/bq[4] ) );
  DRNQHSV4 \pe2/delaycell19/q_reg[4]  ( .D(n15004), .CK(clk), .RDN(n14787), 
        .Q(\pe2/bq[5] ) );
  DRNQHSV4 \pe2/delaycell19/q_reg[3]  ( .D(n14984), .CK(clk), .RDN(n14720), 
        .Q(\pe2/bq[6] ) );
  DRNQHSV4 \pe2/delaycell19/q_reg[2]  ( .D(n14976), .CK(clk), .RDN(n14745), 
        .Q(\pe2/bq[7] ) );
  DRNQHSV4 \pe2/delaycell19/q_reg[1]  ( .D(n15047), .CK(clk), .RDN(n14763), 
        .Q(\pe2/bq[8] ) );
  DRNQHSV4 \pe2/delaycell20/q_reg  ( .D(\pe2/ti_1t ), .CK(clk), .RDN(n14744), 
        .Q(\pe2/ti_1 ) );
  DRNQHSV4 \pe2/delaycell21/q_reg[3]  ( .D(\pe2/ti_7[3] ), .CK(clk), .RDN(
        n14770), .Q(\pe2/ti_7t [3]) );
  DRNQHSV4 \pe3/delaycell1/q_reg[8]  ( .D(ao2[1]), .CK(clk), .RDN(n14748), .Q(
        \pe3/aot [1]) );
  DRNQHSV4 \pe3/delaycell1/q_reg[7]  ( .D(ao2[2]), .CK(clk), .RDN(n14780), .Q(
        \pe3/aot [2]) );
  DRNQHSV4 \pe3/delaycell1/q_reg[6]  ( .D(ao2[3]), .CK(clk), .RDN(n14781), .Q(
        \pe3/aot [3]) );
  DRNQHSV4 \pe3/delaycell1/q_reg[5]  ( .D(ao2[4]), .CK(clk), .RDN(n14792), .Q(
        \pe3/aot [4]) );
  DRNQHSV4 \pe3/delaycell1/q_reg[4]  ( .D(ao2[5]), .CK(clk), .RDN(n14797), .Q(
        \pe3/aot [5]) );
  DRNQHSV4 \pe3/delaycell1/q_reg[3]  ( .D(ao2[6]), .CK(clk), .RDN(n14722), .Q(
        \pe3/aot [6]) );
  DRNQHSV4 \pe3/delaycell1/q_reg[2]  ( .D(ao2[7]), .CK(clk), .RDN(n14767), .Q(
        \pe3/aot [7]) );
  DRNQHSV4 \pe3/delaycell2/q_reg[8]  ( .D(go2[1]), .CK(clk), .RDN(n14714), .Q(
        \pe3/got [1]) );
  DRNQHSV4 \pe3/delaycell2/q_reg[7]  ( .D(go2[2]), .CK(clk), .RDN(n14751), .Q(
        \pe3/got [2]) );
  DRNQHSV4 \pe3/delaycell2/q_reg[6]  ( .D(go2[3]), .CK(clk), .RDN(n14711), .Q(
        \pe3/got [3]) );
  DRNQHSV4 \pe3/delaycell2/q_reg[5]  ( .D(go2[4]), .CK(clk), .RDN(n14776), .Q(
        \pe3/got [4]) );
  DRNQHSV4 \pe3/delaycell2/q_reg[4]  ( .D(go2[5]), .CK(clk), .RDN(n14803), .Q(
        \pe3/got [5]) );
  DRNQHSV4 \pe3/delaycell2/q_reg[3]  ( .D(go2[6]), .CK(clk), .RDN(n14730), .Q(
        \pe3/got [6]) );
  DRNQHSV4 \pe3/delaycell2/q_reg[2]  ( .D(go2[7]), .CK(clk), .RDN(n14748), .Q(
        \pe3/got [7]) );
  DRNQHSV4 \pe3/delaycell2/q_reg[1]  ( .D(go2[8]), .CK(clk), .RDN(n14766), .Q(
        \pe3/got [8]) );
  DRNQHSV4 \pe3/delaycell5/q_reg[6]  ( .D(n15291), .CK(clk), .RDN(n14785), .Q(
        \pe3/pvq [6]) );
  DRNQHSV4 \pe3/delaycell5/q_reg[2]  ( .D(n15294), .CK(clk), .RDN(n14833), .Q(
        \pe3/pvq [2]) );
  DRNQHSV4 \pe3/delaycell6/q_reg[5]  ( .D(poh2[5]), .CK(clk), .RDN(n14871), 
        .Q(\pe3/phq [5]) );
  DRNQHSV4 \pe3/delaycell6/q_reg[4]  ( .D(poh2[4]), .CK(clk), .RDN(n14726), 
        .Q(\pe3/phq [4]) );
  DRNQHSV4 \pe3/delaycell6/q_reg[3]  ( .D(poh2[3]), .CK(clk), .RDN(n14788), 
        .Q(\pe3/phq [3]) );
  DRNQHSV4 \pe3/delaycell6/q_reg[2]  ( .D(poh2[2]), .CK(clk), .RDN(rst), .Q(
        \pe3/phq [2]) );
  DRNQHSV4 \pe3/delaycell6/q_reg[1]  ( .D(poh2[1]), .CK(clk), .RDN(n14808), 
        .Q(\pe3/phq [1]) );
  DRNQHSV4 \pe3/delaycell7/q_reg  ( .D(n9358), .CK(clk), .RDN(n14808), .Q(
        \pe3/ctrq ) );
  DRNQHSV4 \pe3/delaycell19/q_reg[8]  ( .D(n15101), .CK(clk), .RDN(n14762), 
        .Q(\pe3/bq[1] ) );
  DRNQHSV4 \pe3/delaycell19/q_reg[7]  ( .D(n15102), .CK(clk), .RDN(n14764), 
        .Q(\pe3/bq[2] ) );
  DRNQHSV4 \pe3/delaycell19/q_reg[6]  ( .D(n15045), .CK(clk), .RDN(n14766), 
        .Q(\pe3/bq[3] ) );
  DRNQHSV4 \pe3/delaycell19/q_reg[5]  ( .D(n15044), .CK(clk), .RDN(n14753), 
        .Q(\pe3/bq[4] ) );
  DRNQHSV4 \pe3/delaycell19/q_reg[4]  ( .D(n15043), .CK(clk), .RDN(n14783), 
        .Q(\pe3/bq[5] ) );
  DRNQHSV4 \pe3/delaycell19/q_reg[3]  ( .D(n15100), .CK(clk), .RDN(n15173), 
        .Q(\pe3/bq[6] ) );
  DRNQHSV4 \pe3/delaycell19/q_reg[2]  ( .D(n15042), .CK(clk), .RDN(n14719), 
        .Q(\pe3/bq[7] ) );
  DRNQHSV4 \pe4/delaycell1/q_reg[8]  ( .D(ao3[1]), .CK(clk), .RDN(n14871), .Q(
        \pe4/aot [1]) );
  DRNQHSV4 \pe4/delaycell1/q_reg[7]  ( .D(ao3[2]), .CK(clk), .RDN(n14766), .Q(
        \pe4/aot [2]) );
  DRNQHSV4 \pe4/delaycell1/q_reg[6]  ( .D(ao3[3]), .CK(clk), .RDN(n14769), .Q(
        \pe4/aot [3]) );
  DRNQHSV4 \pe4/delaycell1/q_reg[5]  ( .D(ao3[4]), .CK(clk), .RDN(n14773), .Q(
        \pe4/aot [4]) );
  DRNQHSV4 \pe4/delaycell1/q_reg[3]  ( .D(ao3[6]), .CK(clk), .RDN(n14813), .Q(
        \pe4/aot [6]) );
  DRNQHSV4 \pe4/delaycell2/q_reg[8]  ( .D(go3[1]), .CK(clk), .RDN(n14806), .Q(
        \pe4/got [1]) );
  DRNQHSV4 \pe4/delaycell2/q_reg[7]  ( .D(go3[2]), .CK(clk), .RDN(n14810), .Q(
        \pe4/got [2]) );
  DRNQHSV4 \pe4/delaycell2/q_reg[6]  ( .D(go3[3]), .CK(clk), .RDN(n14753), .Q(
        \pe4/got [3]) );
  DRNQHSV4 \pe4/delaycell2/q_reg[5]  ( .D(go3[4]), .CK(clk), .RDN(n14754), .Q(
        \pe4/got [4]) );
  DRNQHSV4 \pe4/delaycell2/q_reg[4]  ( .D(go3[5]), .CK(clk), .RDN(n14871), .Q(
        \pe4/got [5]) );
  DRNQHSV4 \pe4/delaycell2/q_reg[3]  ( .D(go3[6]), .CK(clk), .RDN(n14716), .Q(
        \pe4/got [6]) );
  DRNQHSV4 \pe4/delaycell2/q_reg[2]  ( .D(go3[7]), .CK(clk), .RDN(n14812), .Q(
        \pe4/got [7]) );
  DRNQHSV4 \pe4/delaycell5/q_reg[6]  ( .D(n15286), .CK(clk), .RDN(n14754), .Q(
        \pe4/pvq [6]) );
  DRNQHSV4 \pe4/delaycell5/q_reg[4]  ( .D(n14825), .CK(clk), .RDN(n14749), .Q(
        \pe4/pvq [4]) );
  DRNQHSV4 \pe4/delaycell5/q_reg[2]  ( .D(n15289), .CK(clk), .RDN(n14815), .Q(
        \pe4/pvq [2]) );
  DRNQHSV4 \pe4/delaycell6/q_reg[7]  ( .D(poh3[7]), .CK(clk), .RDN(n14762), 
        .Q(\pe4/phq [7]) );
  DRNQHSV4 \pe4/delaycell6/q_reg[6]  ( .D(poh3[6]), .CK(clk), .RDN(n14766), 
        .Q(\pe4/phq [6]) );
  DRNQHSV4 \pe4/delaycell6/q_reg[5]  ( .D(poh3[5]), .CK(clk), .RDN(n14727), 
        .Q(\pe4/phq [5]) );
  DRNQHSV4 \pe4/delaycell6/q_reg[4]  ( .D(poh3[4]), .CK(clk), .RDN(n8938), .Q(
        \pe4/phq [4]) );
  DRNQHSV4 \pe4/delaycell6/q_reg[3]  ( .D(poh3[3]), .CK(clk), .RDN(n14710), 
        .Q(\pe4/phq [3]) );
  DRNQHSV4 \pe4/delaycell6/q_reg[2]  ( .D(poh3[2]), .CK(clk), .RDN(n14798), 
        .Q(\pe4/phq [2]) );
  DRNQHSV4 \pe4/delaycell6/q_reg[1]  ( .D(poh3[1]), .CK(clk), .RDN(n14833), 
        .Q(\pe4/phq [1]) );
  DRNQHSV4 \pe4/delaycell19/q_reg[8]  ( .D(n15041), .CK(clk), .RDN(n14817), 
        .Q(\pe4/bq[1] ) );
  DRNQHSV4 \pe4/delaycell19/q_reg[7]  ( .D(n15040), .CK(clk), .RDN(n14817), 
        .Q(\pe4/bq[2] ) );
  DRNQHSV4 \pe4/delaycell19/q_reg[6]  ( .D(n15106), .CK(clk), .RDN(n14788), 
        .Q(\pe4/bq[3] ) );
  DRNQHSV4 \pe4/delaycell19/q_reg[5]  ( .D(n15107), .CK(clk), .RDN(n14718), 
        .Q(\pe4/bq[4] ) );
  DRNQHSV4 \pe4/delaycell19/q_reg[4]  ( .D(n15105), .CK(clk), .RDN(n14804), 
        .Q(\pe4/bq[5] ) );
  DRNQHSV4 \pe4/delaycell19/q_reg[3]  ( .D(n15104), .CK(clk), .RDN(rst), .Q(
        \pe4/bq[6] ) );
  DRNQHSV4 \pe4/delaycell19/q_reg[2]  ( .D(\pe4/bqt[7] ), .CK(clk), .RDN(
        n14800), .Q(\pe4/bq[7] ) );
  DRNQHSV4 \pe4/delaycell20/q_reg  ( .D(\pe4/ti_1t ), .CK(clk), .RDN(n14783), 
        .Q(\pe4/ti_1 ) );
  DRNQHSV4 \pe5/delaycell1/q_reg[8]  ( .D(ao4[1]), .CK(clk), .RDN(n14726), .Q(
        \pe5/aot [1]) );
  DRNQHSV4 \pe5/delaycell1/q_reg[7]  ( .D(ao4[2]), .CK(clk), .RDN(n14815), .Q(
        \pe5/aot [2]) );
  DRNQHSV4 \pe5/delaycell1/q_reg[6]  ( .D(ao4[3]), .CK(clk), .RDN(n14756), .Q(
        \pe5/aot [3]) );
  DRNQHSV4 \pe5/delaycell1/q_reg[5]  ( .D(ao4[4]), .CK(clk), .RDN(n14717), .Q(
        \pe5/aot [4]) );
  DRNQHSV4 \pe5/delaycell1/q_reg[4]  ( .D(ao4[5]), .CK(clk), .RDN(n14721), .Q(
        \pe5/aot [5]) );
  DRNQHSV4 \pe5/delaycell1/q_reg[3]  ( .D(ao4[6]), .CK(clk), .RDN(n14768), .Q(
        \pe5/aot [6]) );
  DRNQHSV4 \pe5/delaycell1/q_reg[2]  ( .D(ao4[7]), .CK(clk), .RDN(n14799), .Q(
        \pe5/aot [7]) );
  DRNQHSV4 \pe5/delaycell2/q_reg[8]  ( .D(go4[1]), .CK(clk), .RDN(n15173), .Q(
        \pe5/got [1]) );
  DRNQHSV4 \pe5/delaycell2/q_reg[7]  ( .D(go4[2]), .CK(clk), .RDN(n14721), .Q(
        \pe5/got [2]) );
  DRNQHSV4 \pe5/delaycell2/q_reg[6]  ( .D(go4[3]), .CK(clk), .RDN(n14775), .Q(
        \pe5/got [3]) );
  DRNQHSV4 \pe5/delaycell2/q_reg[5]  ( .D(go4[4]), .CK(clk), .RDN(n14801), .Q(
        \pe5/got [4]) );
  DRNQHSV4 \pe5/delaycell2/q_reg[4]  ( .D(go4[5]), .CK(clk), .RDN(n14808), .Q(
        \pe5/got [5]) );
  DRNQHSV4 \pe5/delaycell2/q_reg[3]  ( .D(go4[6]), .CK(clk), .RDN(n14793), .Q(
        \pe5/got [6]) );
  DRNQHSV4 \pe5/delaycell2/q_reg[2]  ( .D(go4[7]), .CK(clk), .RDN(n14801), .Q(
        \pe5/got [7]) );
  DRNQHSV4 \pe5/delaycell2/q_reg[1]  ( .D(go4[8]), .CK(clk), .RDN(n14752), .Q(
        \pe5/got [8]) );
  DRNQHSV4 \pe5/delaycell5/q_reg[6]  ( .D(n15281), .CK(clk), .RDN(n14778), .Q(
        \pe5/pvq [6]) );
  DRNQHSV4 \pe5/delaycell5/q_reg[2]  ( .D(n15284), .CK(clk), .RDN(n14714), .Q(
        \pe5/pvq [2]) );
  DRNQHSV4 \pe5/delaycell6/q_reg[7]  ( .D(poh4[7]), .CK(clk), .RDN(n14761), 
        .Q(\pe5/phq [7]) );
  DRNQHSV4 \pe5/delaycell6/q_reg[6]  ( .D(poh4[6]), .CK(clk), .RDN(n14793), 
        .Q(\pe5/phq [6]) );
  DRNQHSV4 \pe5/delaycell6/q_reg[5]  ( .D(poh4[5]), .CK(clk), .RDN(n14778), 
        .Q(\pe5/phq [5]) );
  DRNQHSV4 \pe5/delaycell6/q_reg[4]  ( .D(poh4[4]), .CK(clk), .RDN(n14788), 
        .Q(\pe5/phq [4]) );
  DRNQHSV4 \pe5/delaycell6/q_reg[3]  ( .D(poh4[3]), .CK(clk), .RDN(n14778), 
        .Q(\pe5/phq [3]) );
  DRNQHSV4 \pe5/delaycell6/q_reg[2]  ( .D(poh4[2]), .CK(clk), .RDN(n14812), 
        .Q(\pe5/phq [2]) );
  DRNQHSV4 \pe5/delaycell6/q_reg[1]  ( .D(poh4[1]), .CK(clk), .RDN(n14770), 
        .Q(\pe5/phq [1]) );
  DRNQHSV4 \pe5/delaycell7/q_reg  ( .D(n14861), .CK(clk), .RDN(n14753), .Q(
        \pe5/ctrq ) );
  DRNQHSV4 \pe5/delaycell19/q_reg[8]  ( .D(n15039), .CK(clk), .RDN(n14714), 
        .Q(\pe5/bq[1] ) );
  DRNQHSV4 \pe5/delaycell19/q_reg[7]  ( .D(n15038), .CK(clk), .RDN(n14766), 
        .Q(\pe5/bq[2] ) );
  DRNQHSV4 \pe5/delaycell19/q_reg[6]  ( .D(n15112), .CK(clk), .RDN(n14725), 
        .Q(\pe5/bq[3] ) );
  DRNQHSV4 \pe5/delaycell19/q_reg[5]  ( .D(n15113), .CK(clk), .RDN(n14773), 
        .Q(\pe5/bq[4] ) );
  DRNQHSV4 \pe5/delaycell19/q_reg[4]  ( .D(n15109), .CK(clk), .RDN(n14710), 
        .Q(\pe5/bq[5] ) );
  DRNQHSV4 \pe5/delaycell19/q_reg[3]  ( .D(n15111), .CK(clk), .RDN(n14723), 
        .Q(\pe5/bq[6] ) );
  DRNQHSV4 \pe5/delaycell19/q_reg[2]  ( .D(n15110), .CK(clk), .RDN(n14717), 
        .Q(\pe5/bq[7] ) );
  DRNQHSV4 \pe5/delaycell19/q_reg[1]  ( .D(n15108), .CK(clk), .RDN(n14832), 
        .Q(\pe5/bq[8] ) );
  DRNQHSV4 \pe5/delaycell20/q_reg  ( .D(\pe5/ti_1t ), .CK(clk), .RDN(n14754), 
        .Q(\pe5/ti_1 ) );
  DRNQHSV4 \pe6/delaycell1/q_reg[8]  ( .D(ao5[1]), .CK(clk), .RDN(n14806), .Q(
        \pe6/aot [1]) );
  DRNQHSV4 \pe6/delaycell1/q_reg[7]  ( .D(ao5[2]), .CK(clk), .RDN(n14713), .Q(
        \pe6/aot [2]) );
  DRNQHSV4 \pe6/delaycell1/q_reg[6]  ( .D(ao5[3]), .CK(clk), .RDN(n14808), .Q(
        \pe6/aot [3]) );
  DRNQHSV4 \pe6/delaycell1/q_reg[5]  ( .D(ao5[4]), .CK(clk), .RDN(n14754), .Q(
        \pe6/aot [4]) );
  DRNQHSV4 \pe6/delaycell1/q_reg[4]  ( .D(ao5[5]), .CK(clk), .RDN(n14802), .Q(
        \pe6/aot [5]) );
  DRNQHSV4 \pe6/delaycell1/q_reg[2]  ( .D(ao5[7]), .CK(clk), .RDN(n14763), .Q(
        \pe6/aot [7]) );
  DRNQHSV4 \pe6/delaycell2/q_reg[8]  ( .D(go5[1]), .CK(clk), .RDN(n15174), .Q(
        \pe6/got [1]) );
  DRNQHSV4 \pe6/delaycell2/q_reg[7]  ( .D(go5[2]), .CK(clk), .RDN(n8938), .Q(
        \pe6/got [2]) );
  DRNQHSV4 \pe6/delaycell2/q_reg[6]  ( .D(go5[3]), .CK(clk), .RDN(n14797), .Q(
        \pe6/got [3]) );
  DRNQHSV4 \pe6/delaycell2/q_reg[5]  ( .D(go5[4]), .CK(clk), .RDN(n14811), .Q(
        \pe6/got [4]) );
  DRNQHSV4 \pe6/delaycell2/q_reg[4]  ( .D(go5[5]), .CK(clk), .RDN(rst), .Q(
        \pe6/got [5]) );
  DRNQHSV4 \pe6/delaycell2/q_reg[3]  ( .D(go5[6]), .CK(clk), .RDN(n14747), .Q(
        \pe6/got [6]) );
  DRNQHSV4 \pe6/delaycell2/q_reg[2]  ( .D(go5[7]), .CK(clk), .RDN(n14746), .Q(
        \pe6/got [7]) );
  DRNQHSV4 \pe6/delaycell3/q_reg[7]  ( .D(bo5[2]), .CK(clk), .RDN(n15174), .Q(
        bo6[2]) );
  DRNQHSV4 \pe6/delaycell5/q_reg[4]  ( .D(n15277), .CK(clk), .RDN(n14722), .Q(
        \pe6/pvq [4]) );
  DRNQHSV4 \pe6/delaycell5/q_reg[2]  ( .D(n15279), .CK(clk), .RDN(n14815), .Q(
        \pe6/pvq [2]) );
  DRNQHSV4 \pe6/delaycell6/q_reg[7]  ( .D(poh5[7]), .CK(clk), .RDN(n14761), 
        .Q(\pe6/phq [7]) );
  DRNQHSV4 \pe6/delaycell6/q_reg[6]  ( .D(poh5[6]), .CK(clk), .RDN(n14789), 
        .Q(\pe6/phq [6]) );
  DRNQHSV4 \pe6/delaycell6/q_reg[5]  ( .D(poh5[5]), .CK(clk), .RDN(n14723), 
        .Q(\pe6/phq [5]) );
  DRNQHSV4 \pe6/delaycell6/q_reg[4]  ( .D(poh5[4]), .CK(clk), .RDN(n14804), 
        .Q(\pe6/phq [4]) );
  DRNQHSV4 \pe6/delaycell6/q_reg[3]  ( .D(poh5[3]), .CK(clk), .RDN(n14754), 
        .Q(\pe6/phq [3]) );
  DRNQHSV4 \pe6/delaycell6/q_reg[2]  ( .D(poh5[2]), .CK(clk), .RDN(n14719), 
        .Q(\pe6/phq [2]) );
  DRNQHSV4 \pe6/delaycell6/q_reg[1]  ( .D(poh5[1]), .CK(clk), .RDN(n14725), 
        .Q(\pe6/phq [1]) );
  DRNQHSV4 \pe6/delaycell19/q_reg[8]  ( .D(n15118), .CK(clk), .RDN(n14780), 
        .Q(\pe6/bq[1] ) );
  DRNQHSV4 \pe6/delaycell19/q_reg[7]  ( .D(n15120), .CK(clk), .RDN(n14749), 
        .Q(\pe6/bq[2] ) );
  DRNQHSV4 \pe6/delaycell19/q_reg[6]  ( .D(n15119), .CK(clk), .RDN(n14789), 
        .Q(\pe6/bq[3] ) );
  DRNQHSV4 \pe6/delaycell19/q_reg[5]  ( .D(n15117), .CK(clk), .RDN(n14721), 
        .Q(\pe6/bq[4] ) );
  DRNQHSV4 \pe6/delaycell19/q_reg[4]  ( .D(n15116), .CK(clk), .RDN(n14833), 
        .Q(\pe6/bq[5] ) );
  DRNQHSV4 \pe6/delaycell19/q_reg[2]  ( .D(n8919), .CK(clk), .RDN(n14713), .Q(
        \pe6/bq[7] ) );
  DRNQHSV4 \pe6/delaycell20/q_reg  ( .D(\pe6/ti_1t ), .CK(clk), .RDN(n14731), 
        .Q(\pe6/ti_1 ) );
  DRNQHSV4 \pe7/delaycell1/q_reg[8]  ( .D(ao6[1]), .CK(clk), .RDN(n14784), .Q(
        \pe7/aot [1]) );
  DRNQHSV4 \pe7/delaycell1/q_reg[7]  ( .D(ao6[2]), .CK(clk), .RDN(n14777), .Q(
        \pe7/aot [2]) );
  DRNQHSV4 \pe7/delaycell1/q_reg[6]  ( .D(ao6[3]), .CK(clk), .RDN(n14871), .Q(
        \pe7/aot [3]) );
  DRNQHSV4 \pe7/delaycell1/q_reg[5]  ( .D(ao6[4]), .CK(clk), .RDN(n14762), .Q(
        \pe7/aot [4]) );
  DRNQHSV4 \pe7/delaycell1/q_reg[4]  ( .D(ao6[5]), .CK(clk), .RDN(n14728), .Q(
        \pe7/aot [5]) );
  DRNQHSV4 \pe7/delaycell1/q_reg[3]  ( .D(ao6[6]), .CK(clk), .RDN(n14796), .Q(
        \pe7/aot [6]) );
  DRNQHSV4 \pe7/delaycell1/q_reg[2]  ( .D(ao6[7]), .CK(clk), .RDN(n14787), .Q(
        \pe7/aot [7]) );
  DRNQHSV4 \pe7/delaycell1/q_reg[1]  ( .D(ao6[8]), .CK(clk), .RDN(n14814), .Q(
        \pe7/aot [8]) );
  DRNQHSV4 \pe7/delaycell2/q_reg[8]  ( .D(go6[1]), .CK(clk), .RDN(n14716), .Q(
        \pe7/got [1]) );
  DRNQHSV4 \pe7/delaycell2/q_reg[7]  ( .D(go6[2]), .CK(clk), .RDN(n14719), .Q(
        \pe7/got [2]) );
  DRNQHSV4 \pe7/delaycell2/q_reg[6]  ( .D(go6[3]), .CK(clk), .RDN(n14803), .Q(
        \pe7/got [3]) );
  DRNQHSV4 \pe7/delaycell2/q_reg[5]  ( .D(go6[4]), .CK(clk), .RDN(n14711), .Q(
        \pe7/got [4]) );
  DRNQHSV4 \pe7/delaycell2/q_reg[4]  ( .D(go6[5]), .CK(clk), .RDN(n14730), .Q(
        \pe7/got [5]) );
  DRNQHSV4 \pe7/delaycell2/q_reg[3]  ( .D(go6[6]), .CK(clk), .RDN(n14812), .Q(
        \pe7/got [6]) );
  DRNQHSV4 \pe7/delaycell2/q_reg[2]  ( .D(go6[7]), .CK(clk), .RDN(n14775), .Q(
        \pe7/got [7]) );
  DRNQHSV4 \pe7/delaycell2/q_reg[1]  ( .D(go6[8]), .CK(clk), .RDN(n14784), .Q(
        \pe7/got [8]) );
  DRNQHSV4 \pe7/delaycell3/q_reg[8]  ( .D(bo6[1]), .CK(clk), .RDN(n14731), .Q(
        bo7[1]) );
  DRNQHSV4 \pe7/delaycell3/q_reg[7]  ( .D(bo6[2]), .CK(clk), .RDN(n14730), .Q(
        bo7[2]) );
  DRNQHSV4 \pe7/delaycell5/q_reg[4]  ( .D(n15197), .CK(clk), .RDN(n14833), .Q(
        \pe7/pvq [4]) );
  DRNQHSV4 \pe7/delaycell6/q_reg[7]  ( .D(poh6[7]), .CK(clk), .RDN(n14716), 
        .Q(\pe7/phq [7]) );
  DRNQHSV4 \pe7/delaycell6/q_reg[6]  ( .D(poh6[6]), .CK(clk), .RDN(n14713), 
        .Q(\pe7/phq [6]) );
  DRNQHSV4 \pe7/delaycell6/q_reg[5]  ( .D(poh6[5]), .CK(clk), .RDN(n14715), 
        .Q(\pe7/phq [5]) );
  DRNQHSV4 \pe7/delaycell6/q_reg[4]  ( .D(poh6[4]), .CK(clk), .RDN(n14711), 
        .Q(\pe7/phq [4]) );
  DRNQHSV4 \pe7/delaycell6/q_reg[3]  ( .D(poh6[3]), .CK(clk), .RDN(n14806), 
        .Q(\pe7/phq [3]) );
  DRNQHSV4 \pe7/delaycell6/q_reg[2]  ( .D(poh6[2]), .CK(clk), .RDN(n14773), 
        .Q(\pe7/phq [2]) );
  DRNQHSV4 \pe7/delaycell6/q_reg[1]  ( .D(poh6[1]), .CK(clk), .RDN(n14756), 
        .Q(\pe7/phq [1]) );
  DRNQHSV4 \pe7/delaycell7/q_reg  ( .D(n15088), .CK(clk), .RDN(n14784), .Q(
        \pe7/ctrq ) );
  DRNQHSV4 \pe7/delaycell8/q_reg  ( .D(n12067), .CK(clk), .RDN(n14800), .Q(
        ctro7) );
  DRNQHSV4 \pe7/delaycell19/q_reg[8]  ( .D(n15037), .CK(clk), .RDN(n14774), 
        .Q(\pe7/bq[1] ) );
  DRNQHSV4 \pe7/delaycell19/q_reg[7]  ( .D(n15036), .CK(clk), .RDN(n8938), .Q(
        \pe7/bq[2] ) );
  DRNQHSV4 \pe7/delaycell19/q_reg[6]  ( .D(n15125), .CK(clk), .RDN(n14772), 
        .Q(\pe7/bq[3] ) );
  DRNQHSV4 \pe7/delaycell19/q_reg[5]  ( .D(n15126), .CK(clk), .RDN(n14763), 
        .Q(\pe7/bq[4] ) );
  DRNQHSV4 \pe7/delaycell19/q_reg[4]  ( .D(n15122), .CK(clk), .RDN(n14780), 
        .Q(\pe7/bq[5] ) );
  DRNQHSV4 \pe7/delaycell19/q_reg[3]  ( .D(n15124), .CK(clk), .RDN(n8938), .Q(
        \pe7/bq[6] ) );
  DRNQHSV4 \pe7/delaycell19/q_reg[2]  ( .D(n15123), .CK(clk), .RDN(n14833), 
        .Q(\pe7/bq[7] ) );
  DRNQHSV4 \pe7/delaycell19/q_reg[1]  ( .D(n15121), .CK(clk), .RDN(n14871), 
        .Q(\pe7/bq[8] ) );
  DRNQHSV4 \pe7/delaycell20/q_reg  ( .D(\pe7/ti_1t ), .CK(clk), .RDN(n14726), 
        .Q(\pe7/ti_1 ) );
  DRNQHSV4 \pe8/delaycell1/q_reg[8]  ( .D(ao7[1]), .CK(clk), .RDN(n14773), .Q(
        \pe8/aot [1]) );
  DRNQHSV4 \pe8/delaycell1/q_reg[7]  ( .D(ao7[2]), .CK(clk), .RDN(n14780), .Q(
        \pe8/aot [2]) );
  DRNQHSV4 \pe8/delaycell1/q_reg[6]  ( .D(ao7[3]), .CK(clk), .RDN(n14712), .Q(
        \pe8/aot [3]) );
  DRNQHSV4 \pe8/delaycell1/q_reg[5]  ( .D(ao7[4]), .CK(clk), .RDN(n14802), .Q(
        \pe8/aot [4]) );
  DRNQHSV4 \pe8/delaycell1/q_reg[4]  ( .D(ao7[5]), .CK(clk), .RDN(n14712), .Q(
        \pe8/aot [5]) );
  DRNQHSV4 \pe8/delaycell1/q_reg[3]  ( .D(ao7[6]), .CK(clk), .RDN(n14793), .Q(
        \pe8/aot [6]) );
  DRNQHSV4 \pe8/delaycell1/q_reg[2]  ( .D(ao7[7]), .CK(clk), .RDN(n14776), .Q(
        \pe8/aot [7]) );
  DRNQHSV4 \pe8/delaycell2/q_reg[8]  ( .D(go7[1]), .CK(clk), .RDN(n14712), .Q(
        \pe8/got [1]) );
  DRNQHSV4 \pe8/delaycell2/q_reg[7]  ( .D(go7[2]), .CK(clk), .RDN(n14815), .Q(
        \pe8/got [2]) );
  DRNQHSV4 \pe8/delaycell2/q_reg[6]  ( .D(go7[3]), .CK(clk), .RDN(n14721), .Q(
        \pe8/got [3]) );
  DRNQHSV4 \pe8/delaycell2/q_reg[5]  ( .D(go7[4]), .CK(clk), .RDN(n14721), .Q(
        \pe8/got [4]) );
  DRNQHSV4 \pe8/delaycell2/q_reg[4]  ( .D(go7[5]), .CK(clk), .RDN(n14727), .Q(
        \pe8/got [5]) );
  DRNQHSV4 \pe8/delaycell2/q_reg[2]  ( .D(go7[7]), .CK(clk), .RDN(n14718), .Q(
        \pe8/got [7]) );
  DRNQHSV4 \pe8/delaycell2/q_reg[1]  ( .D(go7[8]), .CK(clk), .RDN(n14812), .Q(
        \pe8/got [8]) );
  DRNQHSV4 \pe8/delaycell3/q_reg[6]  ( .D(bo7[3]), .CK(clk), .RDN(n14783), .Q(
        bo8[3]) );
  DRNQHSV4 \pe8/delaycell5/q_reg[6]  ( .D(n15270), .CK(clk), .RDN(n14785), .Q(
        \pe8/pvq [6]) );
  DRNQHSV4 \pe8/delaycell5/q_reg[2]  ( .D(n15272), .CK(clk), .RDN(n14717), .Q(
        \pe8/pvq [2]) );
  DRNQHSV4 \pe8/delaycell6/q_reg[7]  ( .D(poh7[7]), .CK(clk), .RDN(n14804), 
        .Q(\pe8/phq [7]) );
  DRNQHSV4 \pe8/delaycell6/q_reg[6]  ( .D(poh7[6]), .CK(clk), .RDN(n14786), 
        .Q(\pe8/phq [6]) );
  DRNQHSV4 \pe8/delaycell6/q_reg[5]  ( .D(poh7[5]), .CK(clk), .RDN(n14804), 
        .Q(\pe8/phq [5]) );
  DRNQHSV4 \pe8/delaycell6/q_reg[4]  ( .D(poh7[4]), .CK(clk), .RDN(n14814), 
        .Q(\pe8/phq [4]) );
  DRNQHSV4 \pe8/delaycell6/q_reg[3]  ( .D(poh7[3]), .CK(clk), .RDN(n14730), 
        .Q(\pe8/phq [3]) );
  DRNQHSV4 \pe8/delaycell6/q_reg[2]  ( .D(poh7[2]), .CK(clk), .RDN(n14757), 
        .Q(\pe8/phq [2]) );
  DRNQHSV4 \pe8/delaycell6/q_reg[1]  ( .D(poh7[1]), .CK(clk), .RDN(n14753), 
        .Q(\pe8/phq [1]) );
  DRNQHSV4 \pe8/delaycell7/q_reg  ( .D(n12309), .CK(clk), .RDN(n14833), .Q(
        \pe8/ctrq ) );
  DRNQHSV4 \pe8/delaycell19/q_reg[8]  ( .D(n15131), .CK(clk), .RDN(n14771), 
        .Q(\pe8/bq[1] ) );
  DRNQHSV4 \pe8/delaycell19/q_reg[7]  ( .D(n15035), .CK(clk), .RDN(n14759), 
        .Q(\pe8/bq[2] ) );
  DRNQHSV4 \pe8/delaycell19/q_reg[6]  ( .D(n15058), .CK(clk), .RDN(n15173), 
        .Q(\pe8/bq[3] ) );
  DRNQHSV4 \pe8/delaycell19/q_reg[5]  ( .D(n14996), .CK(clk), .RDN(n14752), 
        .Q(\pe8/bq[4] ) );
  DRNQHSV4 \pe8/delaycell19/q_reg[4]  ( .D(n14986), .CK(clk), .RDN(n14730), 
        .Q(\pe8/bq[5] ) );
  DRNQHSV4 \pe8/delaycell19/q_reg[3]  ( .D(n15130), .CK(clk), .RDN(n14806), 
        .Q(\pe8/bq[6] ) );
  DRNQHSV4 \pe8/delaycell19/q_reg[1]  ( .D(n15128), .CK(clk), .RDN(n14751), 
        .Q(\pe8/bq[8] ) );
  DRNQHSV4 \pe9/delaycell1/q_reg[8]  ( .D(ao8[1]), .CK(clk), .RDN(n14785), .Q(
        \pe9/aot [1]) );
  DRNQHSV4 \pe9/delaycell1/q_reg[7]  ( .D(ao8[2]), .CK(clk), .RDN(n14767), .Q(
        \pe9/aot [2]) );
  DRNQHSV4 \pe9/delaycell1/q_reg[6]  ( .D(ao8[3]), .CK(clk), .RDN(n14794), .Q(
        \pe9/aot [3]) );
  DRNQHSV4 \pe9/delaycell1/q_reg[5]  ( .D(ao8[4]), .CK(clk), .RDN(n14814), .Q(
        \pe9/aot [4]) );
  DRNQHSV4 \pe9/delaycell1/q_reg[4]  ( .D(ao8[5]), .CK(clk), .RDN(n14796), .Q(
        \pe9/aot [5]) );
  DRNQHSV4 \pe9/delaycell1/q_reg[3]  ( .D(ao8[6]), .CK(clk), .RDN(n14724), .Q(
        \pe9/aot [6]) );
  DRNQHSV4 \pe9/delaycell1/q_reg[2]  ( .D(ao8[7]), .CK(clk), .RDN(n14754), .Q(
        \pe9/aot [7]) );
  DRNQHSV4 \pe9/delaycell1/q_reg[1]  ( .D(ao8[8]), .CK(clk), .RDN(n14747), .Q(
        \pe9/aot [8]) );
  DRNQHSV4 \pe9/delaycell2/q_reg[8]  ( .D(go8[1]), .CK(clk), .RDN(n14777), .Q(
        \pe9/got [1]) );
  DRNQHSV4 \pe9/delaycell2/q_reg[7]  ( .D(go8[2]), .CK(clk), .RDN(n14799), .Q(
        \pe9/got [2]) );
  DRNQHSV4 \pe9/delaycell2/q_reg[6]  ( .D(go8[3]), .CK(clk), .RDN(n14811), .Q(
        \pe9/got [3]) );
  DRNQHSV4 \pe9/delaycell2/q_reg[5]  ( .D(go8[4]), .CK(clk), .RDN(n14719), .Q(
        \pe9/got [4]) );
  DRNQHSV4 \pe9/delaycell2/q_reg[4]  ( .D(go8[5]), .CK(clk), .RDN(n14832), .Q(
        \pe9/got [5]) );
  DRNQHSV4 \pe9/delaycell2/q_reg[3]  ( .D(go8[6]), .CK(clk), .RDN(n14812), .Q(
        \pe9/got [6]) );
  DRNQHSV4 \pe9/delaycell2/q_reg[2]  ( .D(go8[7]), .CK(clk), .RDN(n14753), .Q(
        \pe9/got [7]) );
  DRNQHSV4 \pe9/delaycell2/q_reg[1]  ( .D(go8[8]), .CK(clk), .RDN(n15174), .Q(
        \pe9/got [8]) );
  DRNQHSV4 \pe9/delaycell3/q_reg[7]  ( .D(bo8[2]), .CK(clk), .RDN(n14776), .Q(
        bo9[2]) );
  DRNQHSV4 \pe9/delaycell3/q_reg[6]  ( .D(bo8[3]), .CK(clk), .RDN(n14817), .Q(
        bo9[3]) );
  DRNQHSV4 \pe9/delaycell5/q_reg[6]  ( .D(n15203), .CK(clk), .RDN(n14713), .Q(
        \pe9/pvq [6]) );
  DRNQHSV4 \pe9/delaycell5/q_reg[5]  ( .D(n15204), .CK(clk), .RDN(n14729), .Q(
        \pe9/pvq [5]) );
  DRNQHSV4 \pe9/delaycell5/q_reg[4]  ( .D(n15266), .CK(clk), .RDN(n14767), .Q(
        \pe9/pvq [4]) );
  DRNQHSV4 \pe9/delaycell5/q_reg[2]  ( .D(n15268), .CK(clk), .RDN(n14761), .Q(
        \pe9/pvq [2]) );
  DRNQHSV4 \pe9/delaycell6/q_reg[7]  ( .D(poh8[7]), .CK(clk), .RDN(n14730), 
        .Q(\pe9/phq [7]) );
  DRNQHSV4 \pe9/delaycell6/q_reg[6]  ( .D(poh8[6]), .CK(clk), .RDN(n14729), 
        .Q(\pe9/phq [6]) );
  DRNQHSV4 \pe9/delaycell6/q_reg[5]  ( .D(poh8[5]), .CK(clk), .RDN(n14778), 
        .Q(\pe9/phq [5]) );
  DRNQHSV4 \pe9/delaycell6/q_reg[4]  ( .D(poh8[4]), .CK(clk), .RDN(n14786), 
        .Q(\pe9/phq [4]) );
  DRNQHSV4 \pe9/delaycell6/q_reg[3]  ( .D(poh8[3]), .CK(clk), .RDN(n14730), 
        .Q(\pe9/phq [3]) );
  DRNQHSV4 \pe9/delaycell6/q_reg[2]  ( .D(poh8[2]), .CK(clk), .RDN(n14786), 
        .Q(\pe9/phq [2]) );
  DRNQHSV4 \pe9/delaycell6/q_reg[1]  ( .D(poh8[1]), .CK(clk), .RDN(n14774), 
        .Q(\pe9/phq [1]) );
  DRNQHSV4 \pe9/delaycell19/q_reg[8]  ( .D(n15138), .CK(clk), .RDN(n15094), 
        .Q(\pe9/bq[1] ) );
  DRNQHSV4 \pe9/delaycell19/q_reg[7]  ( .D(n15034), .CK(clk), .RDN(n14754), 
        .Q(\pe9/bq[2] ) );
  DRNQHSV4 \pe9/delaycell19/q_reg[6]  ( .D(n15137), .CK(clk), .RDN(n14770), 
        .Q(\pe9/bq[3] ) );
  DRNQHSV4 \pe9/delaycell19/q_reg[5]  ( .D(n15059), .CK(clk), .RDN(n14755), 
        .Q(\pe9/bq[4] ) );
  DRNQHSV4 \pe9/delaycell19/q_reg[4]  ( .D(n15136), .CK(clk), .RDN(n14724), 
        .Q(\pe9/bq[5] ) );
  DRNQHSV4 \pe9/delaycell19/q_reg[3]  ( .D(n15135), .CK(clk), .RDN(n14730), 
        .Q(\pe9/bq[6] ) );
  DRNQHSV4 \pe9/delaycell19/q_reg[2]  ( .D(n8918), .CK(clk), .RDN(n15174), .Q(
        \pe9/bq[7] ) );
  DRNQHSV4 \pe9/delaycell20/q_reg  ( .D(\pe9/ti_1t ), .CK(clk), .RDN(n14796), 
        .Q(\pe9/ti_1 ) );
  DRNQHSV4 \pe10/delaycell1/q_reg[8]  ( .D(ao9[1]), .CK(clk), .RDN(n14817), 
        .Q(\pe10/aot [1]) );
  DRNQHSV4 \pe10/delaycell1/q_reg[7]  ( .D(ao9[2]), .CK(clk), .RDN(n14789), 
        .Q(\pe10/aot [2]) );
  DRNQHSV4 \pe10/delaycell1/q_reg[6]  ( .D(ao9[3]), .CK(clk), .RDN(n15094), 
        .Q(\pe10/aot [3]) );
  DRNQHSV4 \pe10/delaycell1/q_reg[5]  ( .D(ao9[4]), .CK(clk), .RDN(n14724), 
        .Q(\pe10/aot [4]) );
  DRNQHSV4 \pe10/delaycell1/q_reg[4]  ( .D(ao9[5]), .CK(clk), .RDN(n15094), 
        .Q(\pe10/aot [5]) );
  DRNQHSV4 \pe10/delaycell1/q_reg[2]  ( .D(ao9[7]), .CK(clk), .RDN(n14787), 
        .Q(\pe10/aot [7]) );
  DRNQHSV4 \pe10/delaycell1/q_reg[1]  ( .D(ao9[8]), .CK(clk), .RDN(n14754), 
        .Q(\pe10/aot [8]) );
  DRNQHSV4 \pe10/delaycell2/q_reg[8]  ( .D(go9[1]), .CK(clk), .RDN(n14753), 
        .Q(\pe10/got [1]) );
  DRNQHSV4 \pe10/delaycell2/q_reg[7]  ( .D(go9[2]), .CK(clk), .RDN(n14745), 
        .Q(\pe10/got [2]) );
  DRNQHSV4 \pe10/delaycell2/q_reg[6]  ( .D(go9[3]), .CK(clk), .RDN(n14760), 
        .Q(\pe10/got [3]) );
  DRNQHSV4 \pe10/delaycell2/q_reg[5]  ( .D(go9[4]), .CK(clk), .RDN(n14756), 
        .Q(\pe10/got [4]) );
  DRNQHSV4 \pe10/delaycell2/q_reg[4]  ( .D(go9[5]), .CK(clk), .RDN(n14810), 
        .Q(\pe10/got [5]) );
  DRNQHSV4 \pe10/delaycell3/q_reg[7]  ( .D(bo9[2]), .CK(clk), .RDN(n14731), 
        .Q(bo10[2]) );
  DRNQHSV4 \pe10/delaycell3/q_reg[6]  ( .D(bo9[3]), .CK(clk), .RDN(n14720), 
        .Q(bo10[3]) );
  DRNQHSV4 \pe10/delaycell5/q_reg[5]  ( .D(pov9[5]), .CK(clk), .RDN(n14731), 
        .Q(\pe10/pvq [5]) );
  DRNQHSV4 \pe10/delaycell5/q_reg[2]  ( .D(n15265), .CK(clk), .RDN(n14724), 
        .Q(\pe10/pvq [2]) );
  DRNQHSV4 \pe10/delaycell6/q_reg[7]  ( .D(poh9[7]), .CK(clk), .RDN(n14716), 
        .Q(\pe10/phq [7]) );
  DRNQHSV4 \pe10/delaycell6/q_reg[5]  ( .D(poh9[5]), .CK(clk), .RDN(n14816), 
        .Q(\pe10/phq [5]) );
  DRNQHSV4 \pe10/delaycell6/q_reg[4]  ( .D(poh9[4]), .CK(clk), .RDN(n14808), 
        .Q(\pe10/phq [4]) );
  DRNQHSV4 \pe10/delaycell6/q_reg[3]  ( .D(poh9[3]), .CK(clk), .RDN(n14816), 
        .Q(\pe10/phq [3]) );
  DRNQHSV4 \pe10/delaycell6/q_reg[2]  ( .D(poh9[2]), .CK(clk), .RDN(n14718), 
        .Q(\pe10/phq [2]) );
  DRNQHSV4 \pe10/delaycell6/q_reg[1]  ( .D(poh9[1]), .CK(clk), .RDN(n14723), 
        .Q(\pe10/phq [1]) );
  DRNQHSV4 \pe10/delaycell7/q_reg  ( .D(n9790), .CK(clk), .RDN(n14728), .Q(
        \pe10/ctrq ) );
  DRNQHSV4 \pe10/delaycell19/q_reg[8]  ( .D(n15033), .CK(clk), .RDN(n14722), 
        .Q(\pe10/bq[1] ) );
  DRNQHSV4 \pe10/delaycell19/q_reg[7]  ( .D(n15032), .CK(clk), .RDN(n14813), 
        .Q(\pe10/bq[2] ) );
  DRNQHSV4 \pe10/delaycell19/q_reg[6]  ( .D(n15031), .CK(clk), .RDN(n14812), 
        .Q(\pe10/bq[3] ) );
  DRNQHSV4 \pe10/delaycell19/q_reg[5]  ( .D(n15030), .CK(clk), .RDN(n14810), 
        .Q(\pe10/bq[4] ) );
  DRNQHSV4 \pe10/delaycell19/q_reg[4]  ( .D(n14989), .CK(clk), .RDN(n14724), 
        .Q(\pe10/bq[5] ) );
  DRNQHSV4 \pe10/delaycell19/q_reg[3]  ( .D(n15029), .CK(clk), .RDN(n14744), 
        .Q(\pe10/bq[6] ) );
  DRNQHSV4 \pe10/delaycell19/q_reg[2]  ( .D(n15053), .CK(clk), .RDN(n14817), 
        .Q(\pe10/bq[7] ) );
  DRNQHSV4 \pe10/delaycell19/q_reg[1]  ( .D(n15028), .CK(clk), .RDN(n14757), 
        .Q(\pe10/bq[8] ) );
  DRNQHSV4 \pe11/delaycell1/q_reg[8]  ( .D(ao10[1]), .CK(clk), .RDN(n14813), 
        .Q(\pe11/aot [1]) );
  DRNQHSV4 \pe11/delaycell1/q_reg[7]  ( .D(ao10[2]), .CK(clk), .RDN(n14781), 
        .Q(\pe11/aot [2]) );
  DRNQHSV4 \pe11/delaycell1/q_reg[6]  ( .D(ao10[3]), .CK(clk), .RDN(n14712), 
        .Q(\pe11/aot [3]) );
  DRNQHSV4 \pe11/delaycell1/q_reg[5]  ( .D(ao10[4]), .CK(clk), .RDN(n14722), 
        .Q(\pe11/aot [4]) );
  DRNQHSV4 \pe11/delaycell1/q_reg[4]  ( .D(ao10[5]), .CK(clk), .RDN(n14808), 
        .Q(\pe11/aot [5]) );
  DRNQHSV4 \pe11/delaycell1/q_reg[3]  ( .D(ao10[6]), .CK(clk), .RDN(n14776), 
        .Q(\pe11/aot [6]) );
  DRNQHSV4 \pe11/delaycell2/q_reg[8]  ( .D(go10[1]), .CK(clk), .RDN(n15174), 
        .Q(\pe11/got [1]) );
  DRNQHSV4 \pe11/delaycell2/q_reg[7]  ( .D(go10[2]), .CK(clk), .RDN(n14816), 
        .Q(\pe11/got [2]) );
  DRNQHSV4 \pe11/delaycell2/q_reg[6]  ( .D(go10[3]), .CK(clk), .RDN(n14778), 
        .Q(\pe11/got [3]) );
  DRNQHSV4 \pe11/delaycell2/q_reg[5]  ( .D(go10[4]), .CK(clk), .RDN(n14764), 
        .Q(\pe11/got [4]) );
  DRNQHSV4 \pe11/delaycell2/q_reg[4]  ( .D(go10[5]), .CK(clk), .RDN(n14802), 
        .Q(\pe11/got [5]) );
  DRNQHSV4 \pe11/delaycell2/q_reg[2]  ( .D(go10[7]), .CK(clk), .RDN(n14725), 
        .Q(\pe11/got [7]) );
  DRNQHSV4 \pe11/delaycell2/q_reg[1]  ( .D(go10[8]), .CK(clk), .RDN(n15174), 
        .Q(\pe11/got [8]) );
  DRNQHSV4 \pe11/delaycell3/q_reg[7]  ( .D(bo10[2]), .CK(clk), .RDN(n14804), 
        .Q(bo11[2]) );
  DRNQHSV4 \pe11/delaycell3/q_reg[6]  ( .D(bo10[3]), .CK(clk), .RDN(n14746), 
        .Q(bo11[3]) );
  DRNQHSV4 \pe11/delaycell3/q_reg[4]  ( .D(bo10[5]), .CK(clk), .RDN(n14765), 
        .Q(bo11[5]) );
  DRNQHSV4 \pe11/delaycell5/q_reg[2]  ( .D(n15263), .CK(clk), .RDN(n14786), 
        .Q(\pe11/pvq [2]) );
  DRNQHSV4 \pe11/delaycell6/q_reg[7]  ( .D(poh10[7]), .CK(clk), .RDN(n14725), 
        .Q(\pe11/phq [7]) );
  DRNQHSV4 \pe11/delaycell6/q_reg[6]  ( .D(poh10[6]), .CK(clk), .RDN(n14768), 
        .Q(\pe11/phq [6]) );
  DRNQHSV4 \pe11/delaycell6/q_reg[5]  ( .D(poh10[5]), .CK(clk), .RDN(n14773), 
        .Q(\pe11/phq [5]) );
  DRNQHSV4 \pe11/delaycell6/q_reg[4]  ( .D(poh10[4]), .CK(clk), .RDN(n14756), 
        .Q(\pe11/phq [4]) );
  DRNQHSV4 \pe11/delaycell6/q_reg[3]  ( .D(poh10[3]), .CK(clk), .RDN(n14721), 
        .Q(\pe11/phq [3]) );
  DRNQHSV4 \pe11/delaycell6/q_reg[2]  ( .D(poh10[2]), .CK(clk), .RDN(n14760), 
        .Q(\pe11/phq [2]) );
  DRNQHSV4 \pe11/delaycell6/q_reg[1]  ( .D(poh10[1]), .CK(clk), .RDN(n14774), 
        .Q(\pe11/phq [1]) );
  DRNQHSV4 \pe11/delaycell7/q_reg  ( .D(n14828), .CK(clk), .RDN(n14787), .Q(
        \pe11/ctrq ) );
  DRNQHSV4 \pe11/delaycell19/q_reg[8]  ( .D(n15145), .CK(clk), .RDN(n14797), 
        .Q(\pe11/bq[1] ) );
  DRNQHSV4 \pe11/delaycell19/q_reg[7]  ( .D(n15143), .CK(clk), .RDN(n14726), 
        .Q(\pe11/bq[2] ) );
  DRNQHSV4 \pe11/delaycell19/q_reg[6]  ( .D(n15144), .CK(clk), .RDN(n14753), 
        .Q(\pe11/bq[3] ) );
  DRNQHSV4 \pe11/delaycell19/q_reg[5]  ( .D(n15027), .CK(clk), .RDN(n14732), 
        .Q(\pe11/bq[4] ) );
  DRNQHSV4 \pe11/delaycell19/q_reg[4]  ( .D(n15141), .CK(clk), .RDN(n14728), 
        .Q(\pe11/bq[5] ) );
  DRNQHSV4 \pe11/delaycell19/q_reg[3]  ( .D(n15142), .CK(clk), .RDN(n14764), 
        .Q(\pe11/bq[6] ) );
  DRNQHSV4 \pe11/delaycell19/q_reg[2]  ( .D(n14995), .CK(clk), .RDN(n14744), 
        .Q(\pe11/bq[7] ) );
  DRNQHSV4 \pe11/delaycell20/q_reg  ( .D(\pe11/ti_1t ), .CK(clk), .RDN(n14724), 
        .Q(\pe11/ti_1 ) );
  DRNQHSV4 \pe12/delaycell1/q_reg[8]  ( .D(ao11[1]), .CK(clk), .RDN(n14772), 
        .Q(\pe12/aot [1]) );
  DRNQHSV4 \pe12/delaycell1/q_reg[7]  ( .D(ao11[2]), .CK(clk), .RDN(n14744), 
        .Q(\pe12/aot [2]) );
  DRNQHSV4 \pe12/delaycell1/q_reg[6]  ( .D(ao11[3]), .CK(clk), .RDN(n14724), 
        .Q(\pe12/aot [3]) );
  DRNQHSV4 \pe12/delaycell1/q_reg[5]  ( .D(ao11[4]), .CK(clk), .RDN(n14728), 
        .Q(\pe12/aot [4]) );
  DRNQHSV4 \pe12/delaycell1/q_reg[4]  ( .D(ao11[5]), .CK(clk), .RDN(n14804), 
        .Q(\pe12/aot [5]) );
  DRNQHSV4 \pe12/delaycell1/q_reg[3]  ( .D(ao11[6]), .CK(clk), .RDN(n14752), 
        .Q(\pe12/aot [6]) );
  DRNQHSV4 \pe12/delaycell1/q_reg[2]  ( .D(ao11[7]), .CK(clk), .RDN(n14744), 
        .Q(\pe12/aot [7]) );
  DRNQHSV4 \pe12/delaycell1/q_reg[1]  ( .D(ao11[8]), .CK(clk), .RDN(n14761), 
        .Q(\pe12/aot [8]) );
  DRNQHSV4 \pe12/delaycell2/q_reg[8]  ( .D(go11[1]), .CK(clk), .RDN(n14780), 
        .Q(\pe12/got [1]) );
  DRNQHSV4 \pe12/delaycell2/q_reg[7]  ( .D(go11[2]), .CK(clk), .RDN(n14745), 
        .Q(\pe12/got [2]) );
  DRNQHSV4 \pe12/delaycell2/q_reg[6]  ( .D(go11[3]), .CK(clk), .RDN(n14809), 
        .Q(\pe12/got [3]) );
  DRNQHSV4 \pe12/delaycell2/q_reg[5]  ( .D(go11[4]), .CK(clk), .RDN(n14725), 
        .Q(\pe12/got [4]) );
  DRNQHSV4 \pe12/delaycell2/q_reg[4]  ( .D(go11[5]), .CK(clk), .RDN(n14746), 
        .Q(\pe12/got [5]) );
  DRNQHSV4 \pe12/delaycell2/q_reg[3]  ( .D(go11[6]), .CK(clk), .RDN(n14792), 
        .Q(\pe12/got [6]) );
  DRNQHSV4 \pe12/delaycell2/q_reg[2]  ( .D(go11[7]), .CK(clk), .RDN(n14769), 
        .Q(\pe12/got [7]) );
  DRNQHSV4 \pe12/delaycell2/q_reg[1]  ( .D(go11[8]), .CK(clk), .RDN(n14778), 
        .Q(\pe12/got [8]) );
  DRNQHSV4 \pe12/delaycell3/q_reg[7]  ( .D(bo11[2]), .CK(clk), .RDN(n14755), 
        .Q(bo12[2]) );
  DRNQHSV4 \pe12/delaycell3/q_reg[6]  ( .D(bo11[3]), .CK(clk), .RDN(n14811), 
        .Q(bo12[3]) );
  DRNQHSV4 \pe12/delaycell3/q_reg[4]  ( .D(bo11[5]), .CK(clk), .RDN(n14720), 
        .Q(bo12[5]) );
  DRNQHSV4 \pe12/delaycell3/q_reg[3]  ( .D(bo11[6]), .CK(clk), .RDN(n14792), 
        .Q(bo12[6]) );
  DRNQHSV4 \pe12/delaycell5/q_reg[2]  ( .D(n15259), .CK(clk), .RDN(n14807), 
        .Q(\pe12/pvq [2]) );
  DRNQHSV4 \pe12/delaycell6/q_reg[7]  ( .D(poh11[7]), .CK(clk), .RDN(n14871), 
        .Q(\pe12/phq [7]) );
  DRNQHSV4 \pe12/delaycell6/q_reg[6]  ( .D(poh11[6]), .CK(clk), .RDN(n15173), 
        .Q(\pe12/phq [6]) );
  DRNQHSV4 \pe12/delaycell6/q_reg[5]  ( .D(poh11[5]), .CK(clk), .RDN(n14781), 
        .Q(\pe12/phq [5]) );
  DRNQHSV4 \pe12/delaycell6/q_reg[4]  ( .D(poh11[4]), .CK(clk), .RDN(n14744), 
        .Q(\pe12/phq [4]) );
  DRNQHSV4 \pe12/delaycell6/q_reg[3]  ( .D(poh11[3]), .CK(clk), .RDN(n14770), 
        .Q(\pe12/phq [3]) );
  DRNQHSV4 \pe12/delaycell6/q_reg[2]  ( .D(poh11[2]), .CK(clk), .RDN(n14770), 
        .Q(\pe12/phq [2]) );
  DRNQHSV4 \pe12/delaycell6/q_reg[1]  ( .D(poh11[1]), .CK(clk), .RDN(n14747), 
        .Q(\pe12/phq [1]) );
  DRNQHSV4 \pe12/delaycell7/q_reg  ( .D(n15090), .CK(clk), .RDN(n14760), .Q(
        \pe12/ctrq ) );
  DRNQHSV4 \pe12/delaycell19/q_reg[8]  ( .D(n14982), .CK(clk), .RDN(n14747), 
        .Q(\pe12/bq[1] ) );
  DRNQHSV4 \pe12/delaycell19/q_reg[7]  ( .D(n14994), .CK(clk), .RDN(n14779), 
        .Q(\pe12/bq[2] ) );
  DRNQHSV4 \pe12/delaycell19/q_reg[6]  ( .D(n14998), .CK(clk), .RDN(n14798), 
        .Q(\pe12/bq[3] ) );
  DRNQHSV4 \pe12/delaycell19/q_reg[5]  ( .D(n14985), .CK(clk), .RDN(n14772), 
        .Q(\pe12/bq[4] ) );
  DRNQHSV4 \pe12/delaycell19/q_reg[4]  ( .D(n15003), .CK(clk), .RDN(n14728), 
        .Q(\pe12/bq[5] ) );
  DRNQHSV4 \pe12/delaycell19/q_reg[3]  ( .D(n15002), .CK(clk), .RDN(n14727), 
        .Q(\pe12/bq[6] ) );
  DRNQHSV4 \pe12/delaycell19/q_reg[2]  ( .D(n15062), .CK(clk), .RDN(n14712), 
        .Q(\pe12/bq[7] ) );
  DRNQHSV4 \pe12/delaycell19/q_reg[1]  ( .D(n14979), .CK(clk), .RDN(n14749), 
        .Q(\pe12/bq[8] ) );
  DRNQHSV4 \pe12/delaycell20/q_reg  ( .D(\pe12/ti_1t ), .CK(clk), .RDN(n14746), 
        .Q(\pe12/ti_1 ) );
  DRNQHSV4 \pe13/delaycell1/q_reg[8]  ( .D(ao12[1]), .CK(clk), .RDN(n14767), 
        .Q(\pe13/aot [1]) );
  DRNQHSV4 \pe13/delaycell1/q_reg[7]  ( .D(ao12[2]), .CK(clk), .RDN(n14723), 
        .Q(\pe13/aot [2]) );
  DRNQHSV4 \pe13/delaycell1/q_reg[6]  ( .D(ao12[3]), .CK(clk), .RDN(n14731), 
        .Q(\pe13/aot [3]) );
  DRNQHSV4 \pe13/delaycell1/q_reg[5]  ( .D(ao12[4]), .CK(clk), .RDN(n14800), 
        .Q(\pe13/aot [4]) );
  DRNQHSV4 \pe13/delaycell1/q_reg[4]  ( .D(ao12[5]), .CK(clk), .RDN(n14778), 
        .Q(\pe13/aot [5]) );
  DRNQHSV4 \pe13/delaycell1/q_reg[3]  ( .D(ao12[6]), .CK(clk), .RDN(n14713), 
        .Q(\pe13/aot [6]) );
  DRNQHSV4 \pe13/delaycell1/q_reg[2]  ( .D(ao12[7]), .CK(clk), .RDN(n14772), 
        .Q(\pe13/aot [7]) );
  DRNQHSV4 \pe13/delaycell1/q_reg[1]  ( .D(ao12[8]), .CK(clk), .RDN(n14783), 
        .Q(\pe13/aot [8]) );
  DRNQHSV4 \pe13/delaycell2/q_reg[8]  ( .D(go12[1]), .CK(clk), .RDN(n14732), 
        .Q(\pe13/got [1]) );
  DRNQHSV4 \pe13/delaycell2/q_reg[7]  ( .D(go12[2]), .CK(clk), .RDN(n14800), 
        .Q(\pe13/got [2]) );
  DRNQHSV4 \pe13/delaycell2/q_reg[6]  ( .D(go12[3]), .CK(clk), .RDN(n14780), 
        .Q(\pe13/got [3]) );
  DRNQHSV4 \pe13/delaycell2/q_reg[5]  ( .D(go12[4]), .CK(clk), .RDN(n14807), 
        .Q(\pe13/got [4]) );
  DRNQHSV4 \pe13/delaycell2/q_reg[4]  ( .D(go12[5]), .CK(clk), .RDN(n14800), 
        .Q(\pe13/got [5]) );
  DRNQHSV4 \pe13/delaycell2/q_reg[3]  ( .D(go12[6]), .CK(clk), .RDN(n14764), 
        .Q(\pe13/got [6]) );
  DRNQHSV4 \pe13/delaycell2/q_reg[2]  ( .D(go12[7]), .CK(clk), .RDN(n14722), 
        .Q(\pe13/got [7]) );
  DRNQHSV4 \pe13/delaycell2/q_reg[1]  ( .D(go12[8]), .CK(clk), .RDN(n14762), 
        .Q(\pe13/got [8]) );
  DRNQHSV4 \pe13/delaycell3/q_reg[8]  ( .D(bo12[1]), .CK(clk), .RDN(n14715), 
        .Q(bo13[1]) );
  DRNQHSV4 \pe13/delaycell3/q_reg[7]  ( .D(bo12[2]), .CK(clk), .RDN(n14756), 
        .Q(bo13[2]) );
  DRNQHSV4 \pe13/delaycell3/q_reg[6]  ( .D(bo12[3]), .CK(clk), .RDN(n14794), 
        .Q(bo13[3]) );
  DRNQHSV4 \pe13/delaycell3/q_reg[3]  ( .D(bo12[6]), .CK(clk), .RDN(n14715), 
        .Q(bo13[6]) );
  DRNQHSV4 \pe13/delaycell5/q_reg[2]  ( .D(n15252), .CK(clk), .RDN(n14812), 
        .Q(\pe13/pvq [2]) );
  DRNQHSV4 \pe13/delaycell6/q_reg[7]  ( .D(poh12[7]), .CK(clk), .RDN(rst), .Q(
        \pe13/phq [7]) );
  DRNQHSV4 \pe13/delaycell6/q_reg[6]  ( .D(poh12[6]), .CK(clk), .RDN(n14786), 
        .Q(\pe13/phq [6]) );
  DRNQHSV4 \pe13/delaycell6/q_reg[5]  ( .D(poh12[5]), .CK(clk), .RDN(n14768), 
        .Q(\pe13/phq [5]) );
  DRNQHSV4 \pe13/delaycell6/q_reg[4]  ( .D(poh12[4]), .CK(clk), .RDN(n14765), 
        .Q(\pe13/phq [4]) );
  DRNQHSV4 \pe13/delaycell6/q_reg[3]  ( .D(poh12[3]), .CK(clk), .RDN(n14772), 
        .Q(\pe13/phq [3]) );
  DRNQHSV4 \pe13/delaycell6/q_reg[2]  ( .D(poh12[2]), .CK(clk), .RDN(n14769), 
        .Q(\pe13/phq [2]) );
  DRNQHSV4 \pe13/delaycell6/q_reg[1]  ( .D(poh12[1]), .CK(clk), .RDN(n14781), 
        .Q(\pe13/phq [1]) );
  DRNQHSV4 \pe13/delaycell7/q_reg  ( .D(n14831), .CK(clk), .RDN(n14798), .Q(
        \pe13/ctrq ) );
  DRNQHSV4 \pe13/delaycell8/q_reg  ( .D(n14795), .CK(clk), .RDN(n14755), .Q(
        ctro13) );
  DRNQHSV4 \pe13/delaycell19/q_reg[8]  ( .D(n15026), .CK(clk), .RDN(n14710), 
        .Q(\pe13/bq[1] ) );
  DRNQHSV4 \pe13/delaycell19/q_reg[7]  ( .D(n14981), .CK(clk), .RDN(n14773), 
        .Q(\pe13/bq[2] ) );
  DRNQHSV4 \pe13/delaycell19/q_reg[6]  ( .D(n15152), .CK(clk), .RDN(n14713), 
        .Q(\pe13/bq[3] ) );
  DRNQHSV4 \pe13/delaycell19/q_reg[5]  ( .D(n15149), .CK(clk), .RDN(n14751), 
        .Q(\pe13/bq[4] ) );
  DRNQHSV4 \pe13/delaycell19/q_reg[4]  ( .D(n15151), .CK(clk), .RDN(n14782), 
        .Q(\pe13/bq[5] ) );
  DRNQHSV4 \pe13/delaycell19/q_reg[3]  ( .D(n15150), .CK(clk), .RDN(n14755), 
        .Q(\pe13/bq[6] ) );
  DRNQHSV4 \pe13/delaycell19/q_reg[2]  ( .D(n15148), .CK(clk), .RDN(n14712), 
        .Q(\pe13/bq[7] ) );
  DRNQHSV4 \pe13/delaycell19/q_reg[1]  ( .D(n15147), .CK(clk), .RDN(n14781), 
        .Q(\pe13/bq[8] ) );
  DRNQHSV4 \pe13/delaycell20/q_reg  ( .D(\pe13/ti_1t ), .CK(clk), .RDN(n14715), 
        .Q(\pe13/ti_1 ) );
  DRNQHSV4 \pe14/delaycell1/q_reg[8]  ( .D(ao13[1]), .CK(clk), .RDN(n14784), 
        .Q(\pe14/aot [1]) );
  DRNQHSV4 \pe14/delaycell1/q_reg[7]  ( .D(ao13[2]), .CK(clk), .RDN(n14787), 
        .Q(\pe14/aot [2]) );
  DRNQHSV4 \pe14/delaycell1/q_reg[6]  ( .D(ao13[3]), .CK(clk), .RDN(n14757), 
        .Q(\pe14/aot [3]) );
  DRNQHSV4 \pe14/delaycell1/q_reg[5]  ( .D(ao13[4]), .CK(clk), .RDN(n14780), 
        .Q(\pe14/aot [4]) );
  DRNQHSV4 \pe14/delaycell1/q_reg[4]  ( .D(ao13[5]), .CK(clk), .RDN(n14756), 
        .Q(\pe14/aot [5]) );
  DRNQHSV4 \pe14/delaycell1/q_reg[3]  ( .D(ao13[6]), .CK(clk), .RDN(n14716), 
        .Q(\pe14/aot [6]) );
  DRNQHSV4 \pe14/delaycell1/q_reg[2]  ( .D(ao13[7]), .CK(clk), .RDN(n14799), 
        .Q(\pe14/aot [7]) );
  DRNQHSV4 \pe14/delaycell1/q_reg[1]  ( .D(ao13[8]), .CK(clk), .RDN(n14776), 
        .Q(\pe14/aot [8]) );
  DRNQHSV4 \pe14/delaycell2/q_reg[8]  ( .D(go13[1]), .CK(clk), .RDN(n14714), 
        .Q(\pe14/got [1]) );
  DRNQHSV4 \pe14/delaycell2/q_reg[7]  ( .D(go13[2]), .CK(clk), .RDN(n14776), 
        .Q(\pe14/got [2]) );
  DRNQHSV4 \pe14/delaycell2/q_reg[6]  ( .D(go13[3]), .CK(clk), .RDN(n14782), 
        .Q(\pe14/got [3]) );
  DRNQHSV4 \pe14/delaycell2/q_reg[5]  ( .D(go13[4]), .CK(clk), .RDN(n14745), 
        .Q(\pe14/got [4]) );
  DRNQHSV4 \pe14/delaycell2/q_reg[4]  ( .D(go13[5]), .CK(clk), .RDN(n8938), 
        .Q(\pe14/got [5]) );
  DRNQHSV4 \pe14/delaycell2/q_reg[3]  ( .D(go13[6]), .CK(clk), .RDN(n14731), 
        .Q(\pe14/got [6]) );
  DRNQHSV4 \pe14/delaycell2/q_reg[2]  ( .D(go13[7]), .CK(clk), .RDN(n14800), 
        .Q(\pe14/got [7]) );
  DRNQHSV4 \pe14/delaycell2/q_reg[1]  ( .D(go13[8]), .CK(clk), .RDN(n14779), 
        .Q(\pe14/got [8]) );
  DRNQHSV4 \pe14/delaycell3/q_reg[8]  ( .D(bo13[1]), .CK(clk), .RDN(n14775), 
        .Q(bo14[1]) );
  DRNQHSV4 \pe14/delaycell3/q_reg[7]  ( .D(bo13[2]), .CK(clk), .RDN(n14780), 
        .Q(bo14[2]) );
  DRNQHSV4 \pe14/delaycell3/q_reg[6]  ( .D(bo13[3]), .CK(clk), .RDN(n14723), 
        .Q(bo14[3]) );
  DRNQHSV4 \pe14/delaycell3/q_reg[5]  ( .D(bo13[4]), .CK(clk), .RDN(n14798), 
        .Q(bo14[4]) );
  DRNQHSV4 \pe14/delaycell3/q_reg[3]  ( .D(bo13[6]), .CK(clk), .RDN(n14788), 
        .Q(bo14[6]) );
  DRNQHSV4 \pe14/delaycell3/q_reg[2]  ( .D(bo13[7]), .CK(clk), .RDN(n14792), 
        .Q(bo14[7]) );
  DRNQHSV4 \pe14/delaycell5/q_reg[2]  ( .D(n15245), .CK(clk), .RDN(n14728), 
        .Q(\pe14/pvq [2]) );
  DRNQHSV4 \pe14/delaycell6/q_reg[7]  ( .D(poh13[7]), .CK(clk), .RDN(n14728), 
        .Q(\pe14/phq [7]) );
  DRNQHSV4 \pe14/delaycell6/q_reg[6]  ( .D(poh13[6]), .CK(clk), .RDN(n14810), 
        .Q(\pe14/phq [6]) );
  DRNQHSV4 \pe14/delaycell6/q_reg[5]  ( .D(poh13[5]), .CK(clk), .RDN(n14809), 
        .Q(\pe14/phq [5]) );
  DRNQHSV4 \pe14/delaycell6/q_reg[4]  ( .D(poh13[4]), .CK(clk), .RDN(n14809), 
        .Q(\pe14/phq [4]) );
  DRNQHSV4 \pe14/delaycell6/q_reg[3]  ( .D(poh13[3]), .CK(clk), .RDN(n14779), 
        .Q(\pe14/phq [3]) );
  DRNQHSV4 \pe14/delaycell6/q_reg[2]  ( .D(poh13[2]), .CK(clk), .RDN(n14779), 
        .Q(\pe14/phq [2]) );
  DRNQHSV4 \pe14/delaycell6/q_reg[1]  ( .D(poh13[1]), .CK(clk), .RDN(n14716), 
        .Q(\pe14/phq [1]) );
  DRNQHSV4 \pe14/delaycell7/q_reg  ( .D(n15087), .CK(clk), .RDN(n14766), .Q(
        \pe14/ctrq ) );
  DRNQHSV4 \pe14/delaycell19/q_reg[8]  ( .D(n15154), .CK(clk), .RDN(n14777), 
        .Q(\pe14/bq[1] ) );
  DRNQHSV4 \pe14/delaycell19/q_reg[7]  ( .D(n15025), .CK(clk), .RDN(n14712), 
        .Q(\pe14/bq[2] ) );
  DRNQHSV4 \pe14/delaycell19/q_reg[6]  ( .D(n15052), .CK(clk), .RDN(n14798), 
        .Q(\pe14/bq[3] ) );
  DRNQHSV4 \pe14/delaycell19/q_reg[5]  ( .D(n15153), .CK(clk), .RDN(n14731), 
        .Q(\pe14/bq[4] ) );
  DRNQHSV4 \pe14/delaycell19/q_reg[4]  ( .D(n15024), .CK(clk), .RDN(n14720), 
        .Q(\pe14/bq[5] ) );
  DRNQHSV4 \pe14/delaycell19/q_reg[3]  ( .D(n14993), .CK(clk), .RDN(n15173), 
        .Q(\pe14/bq[6] ) );
  DRNQHSV4 \pe14/delaycell19/q_reg[2]  ( .D(n15006), .CK(clk), .RDN(n14776), 
        .Q(\pe14/bq[7] ) );
  DRNQHSV4 \pe14/delaycell19/q_reg[1]  ( .D(n14977), .CK(clk), .RDN(rst), .Q(
        \pe14/bq[8] ) );
  DRNQHSV4 \pe14/delaycell20/q_reg  ( .D(\pe14/ti_1t ), .CK(clk), .RDN(n14718), 
        .Q(\pe14/ti_1 ) );
  DRNQHSV4 \pe15/delaycell1/q_reg[8]  ( .D(ao14[1]), .CK(clk), .RDN(n14773), 
        .Q(\pe15/aot [1]) );
  DRNQHSV4 \pe15/delaycell1/q_reg[7]  ( .D(ao14[2]), .CK(clk), .RDN(n14755), 
        .Q(\pe15/aot [2]) );
  DRNQHSV4 \pe15/delaycell1/q_reg[6]  ( .D(ao14[3]), .CK(clk), .RDN(n14799), 
        .Q(\pe15/aot [3]) );
  DRNQHSV4 \pe15/delaycell1/q_reg[5]  ( .D(ao14[4]), .CK(clk), .RDN(n14801), 
        .Q(\pe15/aot [4]) );
  DRNQHSV4 \pe15/delaycell1/q_reg[4]  ( .D(ao14[5]), .CK(clk), .RDN(n14766), 
        .Q(\pe15/aot [5]) );
  DRNQHSV4 \pe15/delaycell1/q_reg[3]  ( .D(ao14[6]), .CK(clk), .RDN(n14777), 
        .Q(\pe15/aot [6]) );
  DRNQHSV4 \pe15/delaycell1/q_reg[2]  ( .D(ao14[7]), .CK(clk), .RDN(n14803), 
        .Q(\pe15/aot [7]) );
  DRNQHSV4 \pe15/delaycell2/q_reg[8]  ( .D(go14[1]), .CK(clk), .RDN(n14779), 
        .Q(\pe15/got [1]) );
  DRNQHSV4 \pe15/delaycell2/q_reg[7]  ( .D(go14[2]), .CK(clk), .RDN(n14744), 
        .Q(\pe15/got [2]) );
  DRNQHSV4 \pe15/delaycell2/q_reg[6]  ( .D(go14[3]), .CK(clk), .RDN(n14729), 
        .Q(\pe15/got [3]) );
  DRNQHSV4 \pe15/delaycell2/q_reg[5]  ( .D(go14[4]), .CK(clk), .RDN(n14785), 
        .Q(\pe15/got [4]) );
  DRNQHSV4 \pe15/delaycell2/q_reg[4]  ( .D(go14[5]), .CK(clk), .RDN(n14777), 
        .Q(\pe15/got [5]) );
  DRNQHSV4 \pe15/delaycell2/q_reg[3]  ( .D(go14[6]), .CK(clk), .RDN(n14765), 
        .Q(\pe15/got [6]) );
  DRNQHSV4 \pe15/delaycell2/q_reg[2]  ( .D(go14[7]), .CK(clk), .RDN(n14787), 
        .Q(\pe15/got [7]) );
  DRNQHSV4 \pe15/delaycell2/q_reg[1]  ( .D(go14[8]), .CK(clk), .RDN(n14817), 
        .Q(\pe15/got [8]) );
  DRNQHSV4 \pe15/delaycell3/q_reg[8]  ( .D(bo14[1]), .CK(clk), .RDN(n14777), 
        .Q(bo15[1]) );
  DRNQHSV4 \pe15/delaycell3/q_reg[7]  ( .D(bo14[2]), .CK(clk), .RDN(n14724), 
        .Q(bo15[2]) );
  DRNQHSV4 \pe15/delaycell3/q_reg[6]  ( .D(bo14[3]), .CK(clk), .RDN(n14774), 
        .Q(bo15[3]) );
  DRNQHSV4 \pe15/delaycell3/q_reg[5]  ( .D(bo14[4]), .CK(clk), .RDN(n14748), 
        .Q(bo15[4]) );
  DRNQHSV4 \pe15/delaycell3/q_reg[3]  ( .D(bo14[6]), .CK(clk), .RDN(n14793), 
        .Q(bo15[6]) );
  DRNQHSV4 \pe15/delaycell3/q_reg[2]  ( .D(bo14[7]), .CK(clk), .RDN(n14745), 
        .Q(bo15[7]) );
  DRNQHSV4 \pe15/delaycell3/q_reg[1]  ( .D(bo14[8]), .CK(clk), .RDN(n14789), 
        .Q(bo15[8]) );
  DRNQHSV4 \pe15/delaycell6/q_reg[7]  ( .D(poh14[7]), .CK(clk), .RDN(n14746), 
        .Q(\pe15/phq [7]) );
  DRNQHSV4 \pe15/delaycell6/q_reg[6]  ( .D(poh14[6]), .CK(clk), .RDN(n14817), 
        .Q(\pe15/phq [6]) );
  DRNQHSV4 \pe15/delaycell6/q_reg[5]  ( .D(poh14[5]), .CK(clk), .RDN(n14765), 
        .Q(\pe15/phq [5]) );
  DRNQHSV4 \pe15/delaycell6/q_reg[4]  ( .D(poh14[4]), .CK(clk), .RDN(n14727), 
        .Q(\pe15/phq [4]) );
  DRNQHSV4 \pe15/delaycell6/q_reg[3]  ( .D(poh14[3]), .CK(clk), .RDN(n14793), 
        .Q(\pe15/phq [3]) );
  DRNQHSV4 \pe15/delaycell6/q_reg[2]  ( .D(poh14[2]), .CK(clk), .RDN(n14783), 
        .Q(\pe15/phq [2]) );
  DRNQHSV4 \pe15/delaycell6/q_reg[1]  ( .D(poh14[1]), .CK(clk), .RDN(n14770), 
        .Q(\pe15/phq [1]) );
  DRNQHSV4 \pe15/delaycell7/q_reg  ( .D(n14702), .CK(clk), .RDN(n14725), .Q(
        \pe15/ctrq ) );
  DRNQHSV4 \pe15/delaycell19/q_reg[8]  ( .D(n15159), .CK(clk), .RDN(n14726), 
        .Q(\pe15/bq[1] ) );
  DRNQHSV4 \pe15/delaycell19/q_reg[7]  ( .D(n15023), .CK(clk), .RDN(n14723), 
        .Q(\pe15/bq[2] ) );
  DRNQHSV4 \pe15/delaycell19/q_reg[6]  ( .D(n15161), .CK(clk), .RDN(n14719), 
        .Q(\pe15/bq[3] ) );
  DRNQHSV4 \pe15/delaycell19/q_reg[5]  ( .D(n15022), .CK(clk), .RDN(n14715), 
        .Q(\pe15/bq[4] ) );
  DRNQHSV4 \pe15/delaycell19/q_reg[4]  ( .D(n15158), .CK(clk), .RDN(n14777), 
        .Q(\pe15/bq[5] ) );
  DRNQHSV4 \pe15/delaycell19/q_reg[3]  ( .D(n15156), .CK(clk), .RDN(n14730), 
        .Q(\pe15/bq[6] ) );
  DRNQHSV4 \pe15/delaycell19/q_reg[2]  ( .D(n15157), .CK(clk), .RDN(n14721), 
        .Q(\pe15/bq[7] ) );
  DRNQHSV4 \pe15/delaycell19/q_reg[1]  ( .D(n15155), .CK(clk), .RDN(n14772), 
        .Q(\pe15/bq[8] ) );
  DRNQHSV4 \pe15/delaycell20/q_reg  ( .D(\pe15/ti_1t ), .CK(clk), .RDN(n14783), 
        .Q(\pe15/ti_1 ) );
  DRNQHSV4 \pe16/delaycell1/q_reg[8]  ( .D(ao15[1]), .CK(clk), .RDN(n14718), 
        .Q(\pe16/aot [1]) );
  DRNQHSV4 \pe16/delaycell1/q_reg[7]  ( .D(ao15[2]), .CK(clk), .RDN(n14718), 
        .Q(\pe16/aot [2]) );
  DRNQHSV4 \pe16/delaycell1/q_reg[6]  ( .D(ao15[3]), .CK(clk), .RDN(n14815), 
        .Q(\pe16/aot [3]) );
  DRNQHSV4 \pe16/delaycell1/q_reg[5]  ( .D(ao15[4]), .CK(clk), .RDN(n14800), 
        .Q(\pe16/aot [4]) );
  DRNQHSV4 \pe16/delaycell1/q_reg[4]  ( .D(ao15[5]), .CK(clk), .RDN(n14797), 
        .Q(\pe16/aot [5]) );
  DRNQHSV4 \pe16/delaycell1/q_reg[3]  ( .D(ao15[6]), .CK(clk), .RDN(n14810), 
        .Q(\pe16/aot [6]) );
  DRNQHSV4 \pe16/delaycell1/q_reg[2]  ( .D(ao15[7]), .CK(clk), .RDN(n14817), 
        .Q(\pe16/aot [7]) );
  DRNQHSV4 \pe16/delaycell1/q_reg[1]  ( .D(ao15[8]), .CK(clk), .RDN(n14760), 
        .Q(\pe16/aot [8]) );
  DRNQHSV4 \pe16/delaycell2/q_reg[8]  ( .D(go15[1]), .CK(clk), .RDN(n14724), 
        .Q(\pe16/got [1]) );
  DRNQHSV4 \pe16/delaycell2/q_reg[7]  ( .D(go15[2]), .CK(clk), .RDN(n14800), 
        .Q(\pe16/got [2]) );
  DRNQHSV4 \pe16/delaycell2/q_reg[6]  ( .D(go15[3]), .CK(clk), .RDN(n14777), 
        .Q(\pe16/got [3]) );
  DRNQHSV4 \pe16/delaycell2/q_reg[5]  ( .D(go15[4]), .CK(clk), .RDN(n14781), 
        .Q(\pe16/got [4]) );
  DRNQHSV4 \pe16/delaycell2/q_reg[4]  ( .D(go15[5]), .CK(clk), .RDN(n8938), 
        .Q(\pe16/got [5]) );
  DRNQHSV4 \pe16/delaycell2/q_reg[3]  ( .D(go15[6]), .CK(clk), .RDN(n14806), 
        .Q(\pe16/got [6]) );
  DRNQHSV4 \pe16/delaycell2/q_reg[2]  ( .D(go15[7]), .CK(clk), .RDN(n14792), 
        .Q(\pe16/got [7]) );
  DRNQHSV4 \pe16/delaycell2/q_reg[1]  ( .D(go15[8]), .CK(clk), .RDN(n14782), 
        .Q(\pe16/got [8]) );
  DRNQHSV4 \pe16/delaycell3/q_reg[8]  ( .D(bo15[1]), .CK(clk), .RDN(n14726), 
        .Q(bo16[1]) );
  DRNQHSV4 \pe16/delaycell3/q_reg[7]  ( .D(bo15[2]), .CK(clk), .RDN(n14814), 
        .Q(bo16[2]) );
  DRNQHSV4 \pe16/delaycell3/q_reg[6]  ( .D(bo15[3]), .CK(clk), .RDN(n14794), 
        .Q(bo16[3]) );
  DRNQHSV4 \pe16/delaycell3/q_reg[5]  ( .D(bo15[4]), .CK(clk), .RDN(n14782), 
        .Q(bo16[4]) );
  DRNQHSV4 \pe16/delaycell3/q_reg[4]  ( .D(bo15[5]), .CK(clk), .RDN(n14779), 
        .Q(bo16[5]) );
  DRNQHSV4 \pe16/delaycell3/q_reg[3]  ( .D(bo15[6]), .CK(clk), .RDN(n14729), 
        .Q(bo16[6]) );
  DRNQHSV4 \pe16/delaycell3/q_reg[2]  ( .D(bo15[7]), .CK(clk), .RDN(n14727), 
        .Q(bo16[7]) );
  DRNQHSV4 \pe16/delaycell3/q_reg[1]  ( .D(bo15[8]), .CK(clk), .RDN(n14770), 
        .Q(bo16[8]) );
  DRNQHSV4 \pe16/delaycell5/q_reg[6]  ( .D(n15202), .CK(clk), .RDN(n14714), 
        .Q(\pe16/pvq [6]) );
  DRNQHSV4 \pe16/delaycell5/q_reg[4]  ( .D(\pov15[4] ), .CK(clk), .RDN(n14770), 
        .Q(\pe16/pvq [4]) );
  DRNQHSV4 \pe16/delaycell5/q_reg[2]  ( .D(n15234), .CK(clk), .RDN(n14765), 
        .Q(\pe16/pvq [2]) );
  DRNQHSV4 \pe16/delaycell6/q_reg[7]  ( .D(poh15[7]), .CK(clk), .RDN(n14724), 
        .Q(\pe16/phq [7]) );
  DRNQHSV4 \pe16/delaycell6/q_reg[6]  ( .D(poh15[6]), .CK(clk), .RDN(n14718), 
        .Q(\pe16/phq [6]) );
  DRNQHSV4 \pe16/delaycell6/q_reg[5]  ( .D(poh15[5]), .CK(clk), .RDN(n14755), 
        .Q(\pe16/phq [5]) );
  DRNQHSV4 \pe16/delaycell6/q_reg[4]  ( .D(poh15[4]), .CK(clk), .RDN(n14752), 
        .Q(\pe16/phq [4]) );
  DRNQHSV4 \pe16/delaycell6/q_reg[3]  ( .D(poh15[3]), .CK(clk), .RDN(n14794), 
        .Q(\pe16/phq [3]) );
  DRNQHSV4 \pe16/delaycell6/q_reg[2]  ( .D(poh15[2]), .CK(clk), .RDN(n14727), 
        .Q(\pe16/phq [2]) );
  DRNQHSV4 \pe16/delaycell6/q_reg[1]  ( .D(poh15[1]), .CK(clk), .RDN(n14807), 
        .Q(\pe16/phq [1]) );
  DRNQHSV4 \pe16/delaycell7/q_reg  ( .D(n14704), .CK(clk), .RDN(n14772), .Q(
        \pe16/ctrq ) );
  DRNQHSV4 \pe16/delaycell8/q_reg  ( .D(n14743), .CK(clk), .RDN(n14728), .Q(
        ctro16) );
  DRNQHSV4 \pe16/delaycell19/q_reg[8]  ( .D(n15021), .CK(clk), .RDN(n14730), 
        .Q(\pe16/bq[1] ) );
  DRNQHSV4 \pe16/delaycell19/q_reg[7]  ( .D(n14992), .CK(clk), .RDN(n14752), 
        .Q(\pe16/bq[2] ) );
  DRNQHSV4 \pe16/delaycell19/q_reg[6]  ( .D(n15163), .CK(clk), .RDN(n14719), 
        .Q(\pe16/bq[3] ) );
  DRNQHSV4 \pe16/delaycell19/q_reg[5]  ( .D(n15162), .CK(clk), .RDN(n14832), 
        .Q(\pe16/bq[4] ) );
  DRNQHSV4 \pe16/delaycell19/q_reg[4]  ( .D(n14991), .CK(clk), .RDN(n14722), 
        .Q(\pe16/bq[5] ) );
  DRNQHSV4 \pe16/delaycell19/q_reg[3]  ( .D(n15001), .CK(clk), .RDN(n14713), 
        .Q(\pe16/bq[6] ) );
  DRNQHSV4 \pe16/delaycell19/q_reg[2]  ( .D(n15051), .CK(clk), .RDN(n14715), 
        .Q(\pe16/bq[7] ) );
  DRNQHSV4 \pe16/delaycell19/q_reg[1]  ( .D(n15056), .CK(clk), .RDN(n14785), 
        .Q(\pe16/bq[8] ) );
  DRNQHSV4 \pe16/delaycell20/q_reg  ( .D(\pe16/ti_1t ), .CK(clk), .RDN(n14720), 
        .Q(\pe16/ti_1 ) );
  DRNQHSV4 \pe17/delaycell1/q_reg[8]  ( .D(ao16[1]), .CK(clk), .RDN(n14784), 
        .Q(\pe17/aot [1]) );
  DRNQHSV4 \pe17/delaycell1/q_reg[7]  ( .D(ao16[2]), .CK(clk), .RDN(n14718), 
        .Q(\pe17/aot [2]) );
  DRNQHSV4 \pe17/delaycell1/q_reg[6]  ( .D(ao16[3]), .CK(clk), .RDN(n14715), 
        .Q(\pe17/aot [3]) );
  DRNQHSV4 \pe17/delaycell1/q_reg[5]  ( .D(ao16[4]), .CK(clk), .RDN(n14780), 
        .Q(\pe17/aot [4]) );
  DRNQHSV4 \pe17/delaycell1/q_reg[4]  ( .D(ao16[5]), .CK(clk), .RDN(n14832), 
        .Q(\pe17/aot [5]) );
  DRNQHSV4 \pe17/delaycell1/q_reg[3]  ( .D(ao16[6]), .CK(clk), .RDN(n14715), 
        .Q(\pe17/aot [6]) );
  DRNQHSV4 \pe17/delaycell1/q_reg[2]  ( .D(ao16[7]), .CK(clk), .RDN(n14766), 
        .Q(\pe17/aot [7]) );
  DRNQHSV4 \pe17/delaycell1/q_reg[1]  ( .D(ao16[8]), .CK(clk), .RDN(n14711), 
        .Q(\pe17/aot [8]) );
  DRNQHSV4 \pe17/delaycell2/q_reg[8]  ( .D(go16[1]), .CK(clk), .RDN(n8938), 
        .Q(\pe17/got [1]) );
  DRNQHSV4 \pe17/delaycell2/q_reg[7]  ( .D(go16[2]), .CK(clk), .RDN(n14710), 
        .Q(\pe17/got [2]) );
  DRNQHSV4 \pe17/delaycell2/q_reg[6]  ( .D(go16[3]), .CK(clk), .RDN(n14748), 
        .Q(\pe17/got [3]) );
  DRNQHSV4 \pe17/delaycell2/q_reg[5]  ( .D(go16[4]), .CK(clk), .RDN(n14771), 
        .Q(\pe17/got [4]) );
  DRNQHSV4 \pe17/delaycell2/q_reg[4]  ( .D(go16[5]), .CK(clk), .RDN(n14803), 
        .Q(\pe17/got [5]) );
  DRNQHSV4 \pe17/delaycell2/q_reg[3]  ( .D(go16[6]), .CK(clk), .RDN(n14792), 
        .Q(\pe17/got [6]) );
  DRNQHSV4 \pe17/delaycell2/q_reg[2]  ( .D(go16[7]), .CK(clk), .RDN(n14729), 
        .Q(\pe17/got [7]) );
  DRNQHSV4 \pe17/delaycell2/q_reg[1]  ( .D(go16[8]), .CK(clk), .RDN(n14801), 
        .Q(\pe17/got [8]) );
  DRNQHSV4 \pe17/delaycell3/q_reg[8]  ( .D(bo16[1]), .CK(clk), .RDN(n14711), 
        .Q(bo17[1]) );
  DRNQHSV4 \pe17/delaycell3/q_reg[7]  ( .D(bo16[2]), .CK(clk), .RDN(n14759), 
        .Q(bo17[2]) );
  DRNQHSV4 \pe17/delaycell3/q_reg[6]  ( .D(bo16[3]), .CK(clk), .RDN(n14810), 
        .Q(bo17[3]) );
  DRNQHSV4 \pe17/delaycell3/q_reg[5]  ( .D(bo16[4]), .CK(clk), .RDN(n14722), 
        .Q(bo17[4]) );
  DRNQHSV4 \pe17/delaycell3/q_reg[4]  ( .D(bo16[5]), .CK(clk), .RDN(n14751), 
        .Q(bo17[5]) );
  DRNQHSV4 \pe17/delaycell3/q_reg[3]  ( .D(bo16[6]), .CK(clk), .RDN(n14748), 
        .Q(bo17[6]) );
  DRNQHSV4 \pe17/delaycell3/q_reg[2]  ( .D(bo16[7]), .CK(clk), .RDN(n14803), 
        .Q(bo17[7]) );
  DRNQHSV4 \pe17/delaycell3/q_reg[1]  ( .D(bo16[8]), .CK(clk), .RDN(n14767), 
        .Q(bo17[8]) );
  DRNQHSV4 \pe17/delaycell5/q_reg[6]  ( .D(n15227), .CK(clk), .RDN(n14771), 
        .Q(\pe17/pvq [6]) );
  DRNQHSV4 \pe17/delaycell5/q_reg[2]  ( .D(n15230), .CK(clk), .RDN(n14732), 
        .Q(\pe17/pvq [2]) );
  DRNQHSV4 \pe17/delaycell6/q_reg[7]  ( .D(poh16[7]), .CK(clk), .RDN(n14732), 
        .Q(\pe17/phq [7]) );
  DRNQHSV4 \pe17/delaycell6/q_reg[6]  ( .D(poh16[6]), .CK(clk), .RDN(n14798), 
        .Q(\pe17/phq [6]) );
  DRNQHSV4 \pe17/delaycell6/q_reg[5]  ( .D(poh16[5]), .CK(clk), .RDN(n14729), 
        .Q(\pe17/phq [5]) );
  DRNQHSV4 \pe17/delaycell6/q_reg[4]  ( .D(poh16[4]), .CK(clk), .RDN(n14773), 
        .Q(\pe17/phq [4]) );
  DRNQHSV4 \pe17/delaycell6/q_reg[3]  ( .D(poh16[3]), .CK(clk), .RDN(n14725), 
        .Q(\pe17/phq [3]) );
  DRNQHSV4 \pe17/delaycell6/q_reg[2]  ( .D(poh16[2]), .CK(clk), .RDN(n14784), 
        .Q(\pe17/phq [2]) );
  DRNQHSV4 \pe17/delaycell6/q_reg[1]  ( .D(poh16[1]), .CK(clk), .RDN(n14710), 
        .Q(\pe17/phq [1]) );
  DRNQHSV4 \pe17/delaycell7/q_reg  ( .D(n10689), .CK(clk), .RDN(n14784), .Q(
        \pe17/ctrq ) );
  DRNQHSV4 \pe17/delaycell8/q_reg  ( .D(n14892), .CK(clk), .RDN(n14811), .Q(
        ctro17) );
  DRNQHSV4 \pe17/delaycell19/q_reg[8]  ( .D(n15005), .CK(clk), .RDN(n14771), 
        .Q(\pe17/bq[1] ) );
  DRNQHSV4 \pe17/delaycell19/q_reg[7]  ( .D(n15166), .CK(clk), .RDN(n14732), 
        .Q(\pe17/bq[2] ) );
  DRNQHSV4 \pe17/delaycell19/q_reg[6]  ( .D(n14987), .CK(clk), .RDN(n14749), 
        .Q(\pe17/bq[3] ) );
  DRNQHSV4 \pe17/delaycell19/q_reg[5]  ( .D(n15020), .CK(clk), .RDN(n14751), 
        .Q(\pe17/bq[4] ) );
  DRNQHSV4 \pe17/delaycell19/q_reg[4]  ( .D(n15165), .CK(clk), .RDN(n14710), 
        .Q(\pe17/bq[5] ) );
  DRNQHSV4 \pe17/delaycell19/q_reg[3]  ( .D(n15000), .CK(clk), .RDN(n14752), 
        .Q(\pe17/bq[6] ) );
  DRNQHSV4 \pe17/delaycell19/q_reg[2]  ( .D(n15164), .CK(clk), .RDN(n14808), 
        .Q(\pe17/bq[7] ) );
  DRNQHSV4 \pe17/delaycell19/q_reg[1]  ( .D(n15057), .CK(clk), .RDN(n14778), 
        .Q(\pe17/bq[8] ) );
  DRNQHSV4 \pe17/delaycell20/q_reg  ( .D(\pe17/ti_1t ), .CK(clk), .RDN(n14833), 
        .Q(\pe17/ti_1 ) );
  DRNQHSV4 \pe18/delaycell1/q_reg[8]  ( .D(ao17[1]), .CK(clk), .RDN(n14797), 
        .Q(\pe18/aot [1]) );
  DRNQHSV4 \pe18/delaycell1/q_reg[7]  ( .D(ao17[2]), .CK(clk), .RDN(n14770), 
        .Q(\pe18/aot [2]) );
  DRNQHSV4 \pe18/delaycell1/q_reg[6]  ( .D(ao17[3]), .CK(clk), .RDN(n14815), 
        .Q(\pe18/aot [3]) );
  DRNQHSV4 \pe18/delaycell1/q_reg[5]  ( .D(ao17[4]), .CK(clk), .RDN(n14810), 
        .Q(\pe18/aot [4]) );
  DRNQHSV4 \pe18/delaycell1/q_reg[4]  ( .D(ao17[5]), .CK(clk), .RDN(n14712), 
        .Q(\pe18/aot [5]) );
  DRNQHSV4 \pe18/delaycell1/q_reg[3]  ( .D(ao17[6]), .CK(clk), .RDN(n14755), 
        .Q(\pe18/aot [6]) );
  DRNQHSV4 \pe18/delaycell1/q_reg[2]  ( .D(ao17[7]), .CK(clk), .RDN(n14768), 
        .Q(\pe18/aot [7]) );
  DRNQHSV4 \pe18/delaycell1/q_reg[1]  ( .D(ao17[8]), .CK(clk), .RDN(n14762), 
        .Q(\pe18/aot [8]) );
  DRNQHSV4 \pe18/delaycell2/q_reg[8]  ( .D(go17[1]), .CK(clk), .RDN(n14814), 
        .Q(\pe18/got [1]) );
  DRNQHSV4 \pe18/delaycell2/q_reg[7]  ( .D(go17[2]), .CK(clk), .RDN(n14811), 
        .Q(\pe18/got [2]) );
  DRNQHSV4 \pe18/delaycell2/q_reg[6]  ( .D(go17[3]), .CK(clk), .RDN(n14814), 
        .Q(\pe18/got [3]) );
  DRNQHSV4 \pe18/delaycell2/q_reg[5]  ( .D(go17[4]), .CK(clk), .RDN(n14748), 
        .Q(\pe18/got [4]) );
  DRNQHSV4 \pe18/delaycell2/q_reg[4]  ( .D(go17[5]), .CK(clk), .RDN(n14782), 
        .Q(\pe18/got [5]) );
  DRNQHSV4 \pe18/delaycell2/q_reg[3]  ( .D(go17[6]), .CK(clk), .RDN(n14806), 
        .Q(\pe18/got [6]) );
  DRNQHSV4 \pe18/delaycell2/q_reg[2]  ( .D(go17[7]), .CK(clk), .RDN(n14724), 
        .Q(\pe18/got [7]) );
  DRNQHSV4 \pe18/delaycell2/q_reg[1]  ( .D(go17[8]), .CK(clk), .RDN(n14786), 
        .Q(\pe18/got [8]) );
  DRNQHSV4 \pe18/delaycell3/q_reg[8]  ( .D(bo17[1]), .CK(clk), .RDN(n14731), 
        .Q(bo18[1]) );
  DRNQHSV4 \pe18/delaycell3/q_reg[7]  ( .D(bo17[2]), .CK(clk), .RDN(n14810), 
        .Q(bo18[2]) );
  DRNQHSV4 \pe18/delaycell3/q_reg[6]  ( .D(bo17[3]), .CK(clk), .RDN(n14723), 
        .Q(bo18[3]) );
  DRNQHSV4 \pe18/delaycell3/q_reg[5]  ( .D(bo17[4]), .CK(clk), .RDN(n14809), 
        .Q(bo18[4]) );
  DRNQHSV4 \pe18/delaycell3/q_reg[4]  ( .D(bo17[5]), .CK(clk), .RDN(n14746), 
        .Q(bo18[5]) );
  DRNQHSV4 \pe18/delaycell3/q_reg[3]  ( .D(bo17[6]), .CK(clk), .RDN(n14746), 
        .Q(bo18[6]) );
  DRNQHSV4 \pe18/delaycell3/q_reg[2]  ( .D(bo17[7]), .CK(clk), .RDN(n14764), 
        .Q(bo18[7]) );
  DRNQHSV4 \pe18/delaycell3/q_reg[1]  ( .D(bo17[8]), .CK(clk), .RDN(n14783), 
        .Q(bo18[8]) );
  DRNQHSV4 \pe18/delaycell5/q_reg[6]  ( .D(n15221), .CK(clk), .RDN(n14793), 
        .Q(\pe18/pvq [6]) );
  DRNQHSV4 \pe18/delaycell5/q_reg[2]  ( .D(n15224), .CK(clk), .RDN(n14728), 
        .Q(\pe18/pvq [2]) );
  DRNQHSV4 \pe18/delaycell6/q_reg[7]  ( .D(poh17[7]), .CK(clk), .RDN(n14784), 
        .Q(\pe18/phq [7]) );
  DRNQHSV4 \pe18/delaycell6/q_reg[6]  ( .D(poh17[6]), .CK(clk), .RDN(n14732), 
        .Q(\pe18/phq [6]) );
  DRNQHSV4 \pe18/delaycell6/q_reg[5]  ( .D(poh17[5]), .CK(clk), .RDN(n14711), 
        .Q(\pe18/phq [5]) );
  DRNQHSV4 \pe18/delaycell6/q_reg[4]  ( .D(poh17[4]), .CK(clk), .RDN(n14744), 
        .Q(\pe18/phq [4]) );
  DRNQHSV4 \pe18/delaycell6/q_reg[3]  ( .D(poh17[3]), .CK(clk), .RDN(n14728), 
        .Q(\pe18/phq [3]) );
  DRNQHSV4 \pe18/delaycell6/q_reg[2]  ( .D(poh17[2]), .CK(clk), .RDN(n14799), 
        .Q(\pe18/phq [2]) );
  DRNQHSV4 \pe18/delaycell6/q_reg[1]  ( .D(poh17[1]), .CK(clk), .RDN(n14756), 
        .Q(\pe18/phq [1]) );
  DRNQHSV4 \pe18/delaycell7/q_reg  ( .D(n14013), .CK(clk), .RDN(n14809), .Q(
        \pe18/ctrq ) );
  DRNQHSV4 \pe18/delaycell19/q_reg[8]  ( .D(n14973), .CK(clk), .RDN(n14793), 
        .Q(\pe18/bq[1] ) );
  DRNQHSV4 \pe18/delaycell19/q_reg[7]  ( .D(n15019), .CK(clk), .RDN(n14724), 
        .Q(\pe18/bq[2] ) );
  DRNQHSV4 \pe18/delaycell19/q_reg[6]  ( .D(n14969), .CK(clk), .RDN(n14760), 
        .Q(\pe18/bq[3] ) );
  DRNQHSV4 \pe18/delaycell19/q_reg[5]  ( .D(n15018), .CK(clk), .RDN(n14812), 
        .Q(\pe18/bq[4] ) );
  DRNQHSV4 \pe18/delaycell19/q_reg[4]  ( .D(n15050), .CK(clk), .RDN(n14749), 
        .Q(\pe18/bq[5] ) );
  DRNQHSV4 \pe18/delaycell19/q_reg[3]  ( .D(n15017), .CK(clk), .RDN(n14771), 
        .Q(\pe18/bq[6] ) );
  DRNQHSV4 \pe18/delaycell19/q_reg[2]  ( .D(n14990), .CK(clk), .RDN(n14748), 
        .Q(\pe18/bq[7] ) );
  DRNQHSV4 \pe18/delaycell19/q_reg[1]  ( .D(n14988), .CK(clk), .RDN(n14771), 
        .Q(\pe18/bq[8] ) );
  DRNQHSV4 \pe18/delaycell20/q_reg  ( .D(\pe18/ti_1t ), .CK(clk), .RDN(rst), 
        .Q(\pe18/ti_1 ) );
  DRNQHSV4 \pe19/delaycell1/q_reg[8]  ( .D(ao18[1]), .CK(clk), .RDN(n14714), 
        .Q(\pe19/aot [1]) );
  DRNQHSV4 \pe19/delaycell1/q_reg[7]  ( .D(ao18[2]), .CK(clk), .RDN(n14748), 
        .Q(\pe19/aot [2]) );
  DRNQHSV4 \pe19/delaycell1/q_reg[6]  ( .D(ao18[3]), .CK(clk), .RDN(n14775), 
        .Q(\pe19/aot [3]) );
  DRNQHSV4 \pe19/delaycell1/q_reg[5]  ( .D(ao18[4]), .CK(clk), .RDN(n14711), 
        .Q(\pe19/aot [4]) );
  DRNQHSV4 \pe19/delaycell1/q_reg[4]  ( .D(ao18[5]), .CK(clk), .RDN(n14793), 
        .Q(\pe19/aot [5]) );
  DRNQHSV4 \pe19/delaycell1/q_reg[3]  ( .D(ao18[6]), .CK(clk), .RDN(n14784), 
        .Q(\pe19/aot [6]) );
  DRNQHSV4 \pe19/delaycell1/q_reg[2]  ( .D(ao18[7]), .CK(clk), .RDN(n14811), 
        .Q(\pe19/aot [7]) );
  DRNQHSV4 \pe19/delaycell1/q_reg[1]  ( .D(ao18[8]), .CK(clk), .RDN(n14711), 
        .Q(\pe19/aot [8]) );
  DRNQHSV4 \pe19/delaycell2/q_reg[8]  ( .D(go18[1]), .CK(clk), .RDN(n14809), 
        .Q(\pe19/got [1]) );
  DRNQHSV4 \pe19/delaycell2/q_reg[7]  ( .D(go18[2]), .CK(clk), .RDN(n14719), 
        .Q(\pe19/got [2]) );
  DRNQHSV4 \pe19/delaycell2/q_reg[6]  ( .D(go18[3]), .CK(clk), .RDN(n14770), 
        .Q(\pe19/got [3]) );
  DRNQHSV4 \pe19/delaycell2/q_reg[5]  ( .D(go18[4]), .CK(clk), .RDN(n14786), 
        .Q(\pe19/got [4]) );
  DRNQHSV4 \pe19/delaycell2/q_reg[4]  ( .D(go18[5]), .CK(clk), .RDN(n14761), 
        .Q(\pe19/got [5]) );
  DRNQHSV4 \pe19/delaycell2/q_reg[3]  ( .D(go18[6]), .CK(clk), .RDN(n14800), 
        .Q(\pe19/got [6]) );
  DRNQHSV4 \pe19/delaycell2/q_reg[2]  ( .D(go18[7]), .CK(clk), .RDN(n14871), 
        .Q(\pe19/got [7]) );
  DRNQHSV4 \pe19/delaycell2/q_reg[1]  ( .D(go18[8]), .CK(clk), .RDN(n14713), 
        .Q(\pe19/got [8]) );
  DRNQHSV4 \pe19/delaycell3/q_reg[8]  ( .D(bo18[1]), .CK(clk), .RDN(n14782), 
        .Q(bo19[1]) );
  DRNQHSV4 \pe19/delaycell3/q_reg[7]  ( .D(bo18[2]), .CK(clk), .RDN(n14754), 
        .Q(bo19[2]) );
  DRNQHSV4 \pe19/delaycell3/q_reg[6]  ( .D(bo18[3]), .CK(clk), .RDN(n14775), 
        .Q(bo19[3]) );
  DRNQHSV4 \pe19/delaycell3/q_reg[5]  ( .D(bo18[4]), .CK(clk), .RDN(n14789), 
        .Q(bo19[4]) );
  DRNQHSV4 \pe19/delaycell3/q_reg[4]  ( .D(bo18[5]), .CK(clk), .RDN(n14710), 
        .Q(bo19[5]) );
  DRNQHSV4 \pe19/delaycell3/q_reg[3]  ( .D(bo18[6]), .CK(clk), .RDN(n14768), 
        .Q(bo19[6]) );
  DRNQHSV4 \pe19/delaycell3/q_reg[2]  ( .D(bo18[7]), .CK(clk), .RDN(n14780), 
        .Q(bo19[7]) );
  DRNQHSV4 \pe19/delaycell3/q_reg[1]  ( .D(bo18[8]), .CK(clk), .RDN(n14774), 
        .Q(bo19[8]) );
  DRNQHSV4 \pe19/delaycell5/q_reg[2]  ( .D(n15219), .CK(clk), .RDN(rst), .Q(
        \pe19/pvq [2]) );
  DRNQHSV4 \pe19/delaycell6/q_reg[7]  ( .D(poh18[7]), .CK(clk), .RDN(n14816), 
        .Q(\pe19/phq [7]) );
  DRNQHSV4 \pe19/delaycell6/q_reg[6]  ( .D(poh18[6]), .CK(clk), .RDN(n14816), 
        .Q(\pe19/phq [6]) );
  DRNQHSV4 \pe19/delaycell6/q_reg[5]  ( .D(poh18[5]), .CK(clk), .RDN(n14815), 
        .Q(\pe19/phq [5]) );
  DRNQHSV4 \pe19/delaycell6/q_reg[4]  ( .D(poh18[4]), .CK(clk), .RDN(n14815), 
        .Q(\pe19/phq [4]) );
  DRNQHSV4 \pe19/delaycell6/q_reg[3]  ( .D(poh18[3]), .CK(clk), .RDN(n14782), 
        .Q(\pe19/phq [3]) );
  DRNQHSV4 \pe19/delaycell6/q_reg[2]  ( .D(poh18[2]), .CK(clk), .RDN(n14792), 
        .Q(\pe19/phq [2]) );
  DRNQHSV4 \pe19/delaycell6/q_reg[1]  ( .D(poh18[1]), .CK(clk), .RDN(n14772), 
        .Q(\pe19/phq [1]) );
  DRNQHSV4 \pe19/delaycell7/q_reg  ( .D(n13143), .CK(clk), .RDN(n14815), .Q(
        \pe19/ctrq ) );
  DRNQHSV4 \pe19/delaycell8/q_reg  ( .D(n14501), .CK(clk), .RDN(n14731), .Q(
        ctro19) );
  DRNQHSV4 \pe19/delaycell19/q_reg[8]  ( .D(n14968), .CK(clk), .RDN(n14773), 
        .Q(\pe19/bq[1] ) );
  DRNQHSV4 \pe19/delaycell19/q_reg[7]  ( .D(n14972), .CK(clk), .RDN(n14815), 
        .Q(\pe19/bq[2] ) );
  DRNQHSV4 \pe19/delaycell19/q_reg[6]  ( .D(n15016), .CK(clk), .RDN(n14871), 
        .Q(\pe19/bq[3] ) );
  DRNQHSV4 \pe19/delaycell19/q_reg[5]  ( .D(n15015), .CK(clk), .RDN(n14792), 
        .Q(\pe19/bq[4] ) );
  DRNQHSV4 \pe19/delaycell19/q_reg[4]  ( .D(n15055), .CK(clk), .RDN(n14773), 
        .Q(\pe19/bq[5] ) );
  DRNQHSV4 \pe19/delaycell19/q_reg[3]  ( .D(n15014), .CK(clk), .RDN(n14719), 
        .Q(\pe19/bq[6] ) );
  DRNQHSV4 \pe19/delaycell19/q_reg[2]  ( .D(n15061), .CK(clk), .RDN(n14722), 
        .Q(\pe19/bq[7] ) );
  DRNQHSV4 \pe19/delaycell19/q_reg[1]  ( .D(n14978), .CK(clk), .RDN(n14714), 
        .Q(\pe19/bq[8] ) );
  DRNQHSV4 \pe19/delaycell20/q_reg  ( .D(\pe19/ti_1t ), .CK(clk), .RDN(n14802), 
        .Q(\pe19/ti_1 ) );
  DRNQHSV4 \pe20/delaycell1/q_reg[8]  ( .D(ao19[1]), .CK(clk), .RDN(n14768), 
        .Q(\pe20/aot [1]) );
  DRNQHSV4 \pe20/delaycell1/q_reg[7]  ( .D(ao19[2]), .CK(clk), .RDN(n14713), 
        .Q(\pe20/aot [2]) );
  DRNQHSV4 \pe20/delaycell1/q_reg[6]  ( .D(ao19[3]), .CK(clk), .RDN(n14796), 
        .Q(\pe20/aot [3]) );
  DRNQHSV4 \pe20/delaycell1/q_reg[5]  ( .D(ao19[4]), .CK(clk), .RDN(n14803), 
        .Q(\pe20/aot [4]) );
  DRNQHSV4 \pe20/delaycell1/q_reg[4]  ( .D(ao19[5]), .CK(clk), .RDN(n14789), 
        .Q(\pe20/aot [5]) );
  DRNQHSV4 \pe20/delaycell1/q_reg[3]  ( .D(ao19[6]), .CK(clk), .RDN(n14714), 
        .Q(\pe20/aot [6]) );
  DRNQHSV4 \pe20/delaycell1/q_reg[2]  ( .D(ao19[7]), .CK(clk), .RDN(n14803), 
        .Q(\pe20/aot [7]) );
  DRNQHSV4 \pe20/delaycell2/q_reg[8]  ( .D(go19[1]), .CK(clk), .RDN(n14808), 
        .Q(\pe20/got [1]) );
  DRNQHSV4 \pe20/delaycell2/q_reg[7]  ( .D(go19[2]), .CK(clk), .RDN(n14808), 
        .Q(\pe20/got [2]) );
  DRNQHSV4 \pe20/delaycell2/q_reg[6]  ( .D(go19[3]), .CK(clk), .RDN(n14762), 
        .Q(\pe20/got [3]) );
  DRNQHSV4 \pe20/delaycell2/q_reg[5]  ( .D(go19[4]), .CK(clk), .RDN(n14762), 
        .Q(\pe20/got [4]) );
  DRNQHSV4 \pe20/delaycell2/q_reg[4]  ( .D(go19[5]), .CK(clk), .RDN(n14794), 
        .Q(\pe20/got [5]) );
  DRNQHSV4 \pe20/delaycell2/q_reg[3]  ( .D(go19[6]), .CK(clk), .RDN(n14802), 
        .Q(\pe20/got [6]) );
  DRNQHSV4 \pe20/delaycell2/q_reg[2]  ( .D(go19[7]), .CK(clk), .RDN(n14713), 
        .Q(\pe20/got [7]) );
  DRNQHSV4 \pe20/delaycell2/q_reg[1]  ( .D(go19[8]), .CK(clk), .RDN(n14732), 
        .Q(\pe20/got [8]) );
  DRNQHSV4 \pe20/delaycell3/q_reg[8]  ( .D(bo19[1]), .CK(clk), .RDN(n14787), 
        .Q(bo20[1]) );
  DRNQHSV4 \pe20/delaycell3/q_reg[7]  ( .D(bo19[2]), .CK(clk), .RDN(n14802), 
        .Q(bo20[2]) );
  DRNQHSV4 \pe20/delaycell3/q_reg[6]  ( .D(bo19[3]), .CK(clk), .RDN(n14833), 
        .Q(bo20[3]) );
  DRNQHSV4 \pe20/delaycell3/q_reg[5]  ( .D(bo19[4]), .CK(clk), .RDN(n14723), 
        .Q(bo20[4]) );
  DRNQHSV4 \pe20/delaycell3/q_reg[4]  ( .D(bo19[5]), .CK(clk), .RDN(n14723), 
        .Q(bo20[5]) );
  DRNQHSV4 \pe20/delaycell3/q_reg[3]  ( .D(bo19[6]), .CK(clk), .RDN(n14722), 
        .Q(bo20[6]) );
  DRNQHSV4 \pe20/delaycell3/q_reg[2]  ( .D(bo19[7]), .CK(clk), .RDN(n14775), 
        .Q(bo20[7]) );
  DRNQHSV4 \pe20/delaycell3/q_reg[1]  ( .D(bo19[8]), .CK(clk), .RDN(n14788), 
        .Q(bo20[8]) );
  DRNQHSV4 \pe20/delaycell5/q_reg[5]  ( .D(n15210), .CK(clk), .RDN(n14788), 
        .Q(\pe20/pvq [5]) );
  DRNQHSV4 \pe20/delaycell5/q_reg[2]  ( .D(n15213), .CK(clk), .RDN(n14727), 
        .Q(\pe20/pvq [2]) );
  DRNQHSV4 \pe20/delaycell5/q_reg[1]  ( .D(n9500), .CK(clk), .RDN(n14744), .Q(
        \pe20/pvq [1]) );
  DRNQHSV4 \pe20/delaycell6/q_reg[7]  ( .D(poh19[7]), .CK(clk), .RDN(n14722), 
        .Q(\pe20/phq [7]) );
  DRNQHSV4 \pe20/delaycell6/q_reg[6]  ( .D(poh19[6]), .CK(clk), .RDN(n14801), 
        .Q(\pe20/phq [6]) );
  DRNQHSV4 \pe20/delaycell6/q_reg[5]  ( .D(poh19[5]), .CK(clk), .RDN(n14761), 
        .Q(\pe20/phq [5]) );
  DRNQHSV4 \pe20/delaycell6/q_reg[4]  ( .D(poh19[4]), .CK(clk), .RDN(n14775), 
        .Q(\pe20/phq [4]) );
  DRNQHSV4 \pe20/delaycell6/q_reg[3]  ( .D(poh19[3]), .CK(clk), .RDN(n14760), 
        .Q(\pe20/phq [3]) );
  DRNQHSV4 \pe20/delaycell6/q_reg[2]  ( .D(poh19[2]), .CK(clk), .RDN(n14814), 
        .Q(\pe20/phq [2]) );
  DRNQHSV4 \pe20/delaycell6/q_reg[1]  ( .D(poh19[1]), .CK(clk), .RDN(n14808), 
        .Q(\pe20/phq [1]) );
  DRNQHSV4 \pe20/delaycell7/q_reg  ( .D(n14700), .CK(clk), .RDN(n14804), .Q(
        \pe20/ctrq ) );
  DRNQHSV4 \pe20/delaycell19/q_reg[8]  ( .D(n15013), .CK(clk), .RDN(n14771), 
        .Q(\pe20/bq[1] ) );
  DRNQHSV4 \pe20/delaycell19/q_reg[7]  ( .D(n15012), .CK(clk), .RDN(n14801), 
        .Q(\pe20/bq[2] ) );
  DRNQHSV4 \pe20/delaycell19/q_reg[6]  ( .D(n15171), .CK(clk), .RDN(n14755), 
        .Q(\pe20/bq[3] ) );
  DRNQHSV4 \pe20/delaycell19/q_reg[5]  ( .D(n15170), .CK(clk), .RDN(n14753), 
        .Q(\pe20/bq[4] ) );
  DRNQHSV4 \pe20/delaycell19/q_reg[4]  ( .D(n15011), .CK(clk), .RDN(n14809), 
        .Q(\pe20/bq[5] ) );
  DRNQHSV4 \pe20/delaycell19/q_reg[3]  ( .D(n15010), .CK(clk), .RDN(n14751), 
        .Q(\pe20/bq[6] ) );
  DRNQHSV4 \pe20/delaycell19/q_reg[2]  ( .D(n15169), .CK(clk), .RDN(n14807), 
        .Q(\pe20/bq[7] ) );
  DRNQHSV4 \pe21/delaycell1/q_reg[8]  ( .D(ao20[1]), .CK(clk), .RDN(n14772), 
        .Q(\pe21/aot [1]) );
  DRNQHSV4 \pe21/delaycell1/q_reg[7]  ( .D(ao20[2]), .CK(clk), .RDN(n14760), 
        .Q(\pe21/aot [2]) );
  DRNQHSV4 \pe21/delaycell1/q_reg[6]  ( .D(ao20[3]), .CK(clk), .RDN(n14729), 
        .Q(\pe21/aot [3]) );
  DRNQHSV4 \pe21/delaycell1/q_reg[5]  ( .D(ao20[4]), .CK(clk), .RDN(n14724), 
        .Q(\pe21/aot [4]) );
  DRNQHSV4 \pe21/delaycell1/q_reg[4]  ( .D(ao20[5]), .CK(clk), .RDN(n14712), 
        .Q(\pe21/aot [5]) );
  DRNQHSV4 \pe21/delaycell1/q_reg[3]  ( .D(ao20[6]), .CK(clk), .RDN(n14745), 
        .Q(\pe21/aot [6]) );
  DRNQHSV4 \pe21/delaycell1/q_reg[2]  ( .D(ao20[7]), .CK(clk), .RDN(n14759), 
        .Q(\pe21/aot [7]) );
  DRNQHSV4 \pe21/delaycell1/q_reg[1]  ( .D(ao20[8]), .CK(clk), .RDN(n14731), 
        .Q(\pe21/aot [8]) );
  DRNQHSV4 \pe21/delaycell2/q_reg[8]  ( .D(go20[1]), .CK(clk), .RDN(n14765), 
        .Q(\pe21/got [1]) );
  DRNQHSV4 \pe21/delaycell2/q_reg[7]  ( .D(go20[2]), .CK(clk), .RDN(n15094), 
        .Q(\pe21/got [2]) );
  DRNQHSV4 \pe21/delaycell2/q_reg[6]  ( .D(go20[3]), .CK(clk), .RDN(n14796), 
        .Q(\pe21/got [3]) );
  DRNQHSV4 \pe21/delaycell2/q_reg[5]  ( .D(go20[4]), .CK(clk), .RDN(n14731), 
        .Q(\pe21/got [4]) );
  DRNQHSV4 \pe21/delaycell2/q_reg[4]  ( .D(go20[5]), .CK(clk), .RDN(n14754), 
        .Q(\pe21/got [5]) );
  DRNQHSV4 \pe21/delaycell2/q_reg[3]  ( .D(go20[6]), .CK(clk), .RDN(n14725), 
        .Q(\pe21/got [6]) );
  DRNQHSV4 \pe21/delaycell2/q_reg[2]  ( .D(go20[7]), .CK(clk), .RDN(n15174), 
        .Q(\pe21/got [7]) );
  DRNQHSV4 \pe21/delaycell2/q_reg[1]  ( .D(go20[8]), .CK(clk), .RDN(n14765), 
        .Q(\pe21/got [8]) );
  DRNQHSV4 \pe21/delaycell3/q_reg[6]  ( .D(bo20[3]), .CK(clk), .RDN(n14763), 
        .Q(bo21[3]) );
  DRNQHSV4 \pe21/delaycell3/q_reg[5]  ( .D(bo20[4]), .CK(clk), .RDN(n14799), 
        .Q(bo21[4]) );
  DRNQHSV4 \pe21/delaycell3/q_reg[2]  ( .D(bo20[7]), .CK(clk), .RDN(n14799), 
        .Q(bo21[7]) );
  DRNQHSV4 \pe21/delaycell5/q_reg[6]  ( .D(n15207), .CK(clk), .RDN(n14732), 
        .Q(\pe21/pvq [6]) );
  DRNQHSV4 \pe21/delaycell5/q_reg[2]  ( .D(n15209), .CK(clk), .RDN(n14763), 
        .Q(\pe21/pvq [2]) );
  DRNQHSV4 \pe21/delaycell6/q_reg[7]  ( .D(poh20[7]), .CK(clk), .RDN(n14799), 
        .Q(\pe21/phq [7]) );
  DRNQHSV4 \pe21/delaycell6/q_reg[6]  ( .D(poh20[6]), .CK(clk), .RDN(n14763), 
        .Q(\pe21/phq [6]) );
  DRNQHSV4 \pe21/delaycell6/q_reg[5]  ( .D(poh20[5]), .CK(clk), .RDN(n14710), 
        .Q(\pe21/phq [5]) );
  DRNQHSV4 \pe21/delaycell6/q_reg[4]  ( .D(poh20[4]), .CK(clk), .RDN(n14763), 
        .Q(\pe21/phq [4]) );
  DRNQHSV4 \pe21/delaycell6/q_reg[3]  ( .D(poh20[3]), .CK(clk), .RDN(n14770), 
        .Q(\pe21/phq [3]) );
  DRNQHSV4 \pe21/delaycell6/q_reg[2]  ( .D(poh20[2]), .CK(clk), .RDN(n14732), 
        .Q(\pe21/phq [2]) );
  DRNQHSV4 \pe21/delaycell6/q_reg[1]  ( .D(poh20[1]), .CK(clk), .RDN(n14801), 
        .Q(\pe21/phq [1]) );
  DRNQHSV4 \pe21/delaycell7/q_reg  ( .D(n15177), .CK(clk), .RDN(n14719), .Q(
        \pe21/ctrq ) );
  DRNQHSV4 \pe21/delaycell19/q_reg[8]  ( .D(n15009), .CK(clk), .RDN(n14781), 
        .Q(\pe21/bq[1] ) );
  DRNQHSV4 \pe21/delaycell19/q_reg[7]  ( .D(n15060), .CK(clk), .RDN(n14782), 
        .Q(\pe21/bq[2] ) );
  DRNQHSV4 \pe21/delaycell19/q_reg[6]  ( .D(n15048), .CK(clk), .RDN(n14796), 
        .Q(\pe21/bq[3] ) );
  DRNQHSV4 \pe21/delaycell19/q_reg[5]  ( .D(n15063), .CK(clk), .RDN(n14711), 
        .Q(\pe21/bq[4] ) );
  DRNQHSV4 \pe21/delaycell19/q_reg[4]  ( .D(n15172), .CK(clk), .RDN(n14726), 
        .Q(\pe21/bq[5] ) );
  DRNQHSV4 \pe21/delaycell19/q_reg[3]  ( .D(n15007), .CK(clk), .RDN(n14769), 
        .Q(\pe21/bq[6] ) );
  DRNQHSV4 \pe21/delaycell19/q_reg[2]  ( .D(n15049), .CK(clk), .RDN(n14721), 
        .Q(\pe21/bq[7] ) );
  DRNQHSV4 \pe21/delaycell19/q_reg[1]  ( .D(n8917), .CK(clk), .RDN(n14715), 
        .Q(\pe21/bq[8] ) );
  DRNQHSV4 \pe21/delaycell20/q_reg  ( .D(\pe21/ti_1t ), .CK(clk), .RDN(n14811), 
        .Q(\pe21/ti_1 ) );
  DRNQHSV4 \pe21/delaycell21/q_reg[2]  ( .D(n10876), .CK(clk), .RDN(n14759), 
        .Q(\pe21/ti_7t [2]) );
  DRNQHSV1 \pe5/delaycell21/q_reg[4]  ( .D(n12780), .CK(clk), .RDN(n14786), 
        .Q(\pe5/ti_7t [4]) );
  DRNQHSV1 \pe3/delaycell21/q_reg[6]  ( .D(n14941), .CK(clk), .RDN(n14730), 
        .Q(\pe3/ti_7t [6]) );
  DRNQHSV1 \pe3/delaycell21/q_reg[2]  ( .D(n14872), .CK(clk), .RDN(n14732), 
        .Q(\pe3/ti_7t [2]) );
  DRNQHSV1 \pe15/delaycell21/q_reg[2]  ( .D(n5946), .CK(clk), .RDN(n14727), 
        .Q(\pe15/ti_7t [2]) );
  DRNQHSV1 \pe4/delaycell21/q_reg[4]  ( .D(n14933), .CK(clk), .RDN(n14813), 
        .Q(\pe4/ti_7t [4]) );
  DRNQHSV1 \pe4/delaycell21/q_reg[2]  ( .D(n14733), .CK(clk), .RDN(n14799), 
        .Q(\pe4/ti_7t [2]) );
  DRNQHSV1 \pe15/delaycell21/q_reg[1]  ( .D(n15072), .CK(clk), .RDN(n14812), 
        .Q(\pe15/ti_7t [1]) );
  DRNQHSV1 \pe20/delaycell21/q_reg[7]  ( .D(n14709), .CK(clk), .RDN(n14798), 
        .Q(\pe20/ti_7t [7]) );
  DRNQHSV1 \pe9/delaycell21/q_reg[2]  ( .D(n14896), .CK(clk), .RDN(n14757), 
        .Q(\pe9/ti_7t [2]) );
  DRNQHSV1 \pe13/delaycell21/q_reg[4]  ( .D(\pe13/ti_7[4] ), .CK(clk), .RDN(
        n14723), .Q(\pe13/ti_7t [4]) );
  DRNQHSV1 \pe21/delaycell21/q_reg[4]  ( .D(n15175), .CK(clk), .RDN(n14759), 
        .Q(\pe21/ti_7t [4]) );
  DRNQHSV1 \pe21/delaycell21/q_reg[7]  ( .D(n15085), .CK(clk), .RDN(n14787), 
        .Q(\pe21/ti_7t [7]) );
  DRNQHSV1 \pe14/delaycell21/q_reg[7]  ( .D(n14930), .CK(clk), .RDN(n14746), 
        .Q(\pe14/ti_7t [7]) );
  DRNQHSV2 \pe5/delaycell24/q_reg[2]  ( .D(\pe5/poht [2]), .CK(clk), .RDN(
        n14753), .Q(poh5[2]) );
  DRNQHSV2 \pe21/delaycell21/q_reg[5]  ( .D(\pe21/ti_7[5] ), .CK(clk), .RDN(
        n14760), .Q(\pe21/ti_7t [5]) );
  DRNQHSV2 \pe21/delaycell21/q_reg[6]  ( .D(n7519), .CK(clk), .RDN(n15173), 
        .Q(\pe21/ti_7t [6]) );
  DRNQHSV1 \pe1/delaycell21/q_reg[7]  ( .D(n8947), .CK(clk), .RDN(n14797), .Q(
        \pe1/ti_7t [7]) );
  DRNQHSV2 \pe21/delaycell3/q_reg[4]  ( .D(bo20[5]), .CK(clk), .RDN(n14767), 
        .Q(bo21[5]) );
  DRNQHSV2 \pe21/delaycell3/q_reg[1]  ( .D(bo20[8]), .CK(clk), .RDN(n14799), 
        .Q(bo21[8]) );
  DRNQHSV2 \pe21/delaycell3/q_reg[8]  ( .D(bo20[1]), .CK(clk), .RDN(n14810), 
        .Q(bo21[1]) );
  DRNQHSV2 \pe21/delaycell3/q_reg[7]  ( .D(bo20[2]), .CK(clk), .RDN(n14769), 
        .Q(bo21[2]) );
  DRNQHSV2 \pe21/delaycell3/q_reg[3]  ( .D(bo20[6]), .CK(clk), .RDN(n14776), 
        .Q(bo21[6]) );
  DRNQHSV1 \pe2/delaycell21/q_reg[7]  ( .D(n14957), .CK(clk), .RDN(n14766), 
        .Q(\pe2/ti_7t [7]) );
  DRNQHSV1 \pe13/delaycell21/q_reg[7]  ( .D(n14961), .CK(clk), .RDN(n14765), 
        .Q(\pe13/ti_7t [7]) );
  DRNQHSV1 \pe1/delaycell21/q_reg[6]  ( .D(\pe1/ti_7[6] ), .CK(clk), .RDN(
        n15174), .Q(\pe1/ti_7t [6]) );
  DRNQHSV1 \pe5/delaycell21/q_reg[6]  ( .D(n15193), .CK(clk), .RDN(n14808), 
        .Q(\pe5/ti_7t [6]) );
  DRNQHSV1 \pe7/delaycell21/q_reg[7]  ( .D(n14852), .CK(clk), .RDN(n14720), 
        .Q(\pe7/ti_7t [7]) );
  DRNQHSV1 \pe18/delaycell21/q_reg[7]  ( .D(n14683), .CK(clk), .RDN(n14777), 
        .Q(\pe18/ti_7t [7]) );
  DRNQHSV1 \pe19/delaycell21/q_reg[7]  ( .D(n14862), .CK(clk), .RDN(n14751), 
        .Q(\pe19/ti_7t [7]) );
  DRNQHSV1 \pe1/delaycell22/q_reg[8]  ( .D(\pe1/aot [1]), .CK(clk), .RDN(
        n14762), .Q(ao1[1]) );
  DRNQHSV1 \pe1/delaycell22/q_reg[7]  ( .D(\pe1/aot [2]), .CK(clk), .RDN(
        n14762), .Q(ao1[2]) );
  DRNQHSV1 \pe1/delaycell22/q_reg[6]  ( .D(\pe1/aot [3]), .CK(clk), .RDN(
        n14776), .Q(ao1[3]) );
  DRNQHSV1 \pe1/delaycell22/q_reg[5]  ( .D(\pe1/aot [4]), .CK(clk), .RDN(
        n14816), .Q(ao1[4]) );
  DRNQHSV1 \pe1/delaycell22/q_reg[4]  ( .D(\pe1/aot [5]), .CK(clk), .RDN(
        n14764), .Q(ao1[5]) );
  DRNQHSV1 \pe1/delaycell22/q_reg[3]  ( .D(\pe1/aot [6]), .CK(clk), .RDN(
        n14832), .Q(ao1[6]) );
  DRNQHSV1 \pe1/delaycell22/q_reg[2]  ( .D(\pe1/aot [7]), .CK(clk), .RDN(
        n14764), .Q(ao1[7]) );
  DRNQHSV1 \pe1/delaycell22/q_reg[1]  ( .D(\pe1/aot [8]), .CK(clk), .RDN(
        n14751), .Q(ao1[8]) );
  DRNQHSV1 \pe1/delaycell23/q_reg[8]  ( .D(\pe1/got [1]), .CK(clk), .RDN(
        n14759), .Q(go1[1]) );
  DRNQHSV1 \pe1/delaycell23/q_reg[7]  ( .D(\pe1/got [2]), .CK(clk), .RDN(
        n14753), .Q(go1[2]) );
  DRNQHSV1 \pe1/delaycell23/q_reg[6]  ( .D(\pe1/got [3]), .CK(clk), .RDN(
        n14747), .Q(go1[3]) );
  DRNQHSV1 \pe1/delaycell23/q_reg[5]  ( .D(\pe1/got [4]), .CK(clk), .RDN(
        n14763), .Q(go1[4]) );
  DRNQHSV1 \pe1/delaycell23/q_reg[4]  ( .D(\pe1/got [5]), .CK(clk), .RDN(
        n14753), .Q(go1[5]) );
  DRNQHSV1 \pe1/delaycell23/q_reg[3]  ( .D(\pe1/got [6]), .CK(clk), .RDN(
        n14768), .Q(go1[6]) );
  DRNQHSV1 \pe1/delaycell23/q_reg[2]  ( .D(n14703), .CK(clk), .RDN(n15173), 
        .Q(go1[7]) );
  DRNQHSV1 \pe1/delaycell23/q_reg[1]  ( .D(\pe1/got [8]), .CK(clk), .RDN(
        n14723), .Q(go1[8]) );
  DRNQHSV2 \pe1/delaycell24/q_reg[6]  ( .D(\pe1/poht [6]), .CK(clk), .RDN(
        n14775), .Q(poh1[6]) );
  DRNQHSV2 \pe1/delaycell24/q_reg[3]  ( .D(\pe1/poht [3]), .CK(clk), .RDN(
        n14730), .Q(poh1[3]) );
  DRNQHSV2 \pe1/delaycell24/q_reg[2]  ( .D(\pe1/poht [2]), .CK(clk), .RDN(
        n14747), .Q(poh1[2]) );
  DRNQHSV2 \pe1/delaycell24/q_reg[1]  ( .D(\pe1/poht [1]), .CK(clk), .RDN(
        n14785), .Q(poh1[1]) );
  DRNQHSV1 \pe2/delaycell22/q_reg[8]  ( .D(\pe2/aot [1]), .CK(clk), .RDN(
        n14793), .Q(ao2[1]) );
  DRNQHSV1 \pe2/delaycell22/q_reg[7]  ( .D(\pe2/aot [2]), .CK(clk), .RDN(
        n14712), .Q(ao2[2]) );
  DRNQHSV1 \pe2/delaycell22/q_reg[6]  ( .D(\pe2/aot [3]), .CK(clk), .RDN(
        n14745), .Q(ao2[3]) );
  DRNQHSV1 \pe2/delaycell22/q_reg[5]  ( .D(\pe2/aot [4]), .CK(clk), .RDN(
        n14807), .Q(ao2[4]) );
  DRNQHSV1 \pe2/delaycell22/q_reg[4]  ( .D(\pe2/aot [5]), .CK(clk), .RDN(
        n14766), .Q(ao2[5]) );
  DRNQHSV1 \pe2/delaycell22/q_reg[3]  ( .D(n14741), .CK(clk), .RDN(n14751), 
        .Q(ao2[6]) );
  DRNQHSV1 \pe2/delaycell22/q_reg[2]  ( .D(\pe2/aot [7]), .CK(clk), .RDN(
        n14724), .Q(ao2[7]) );
  DRNQHSV1 \pe2/delaycell22/q_reg[1]  ( .D(n14858), .CK(clk), .RDN(n14778), 
        .Q(ao2[8]) );
  DRNQHSV1 \pe2/delaycell23/q_reg[8]  ( .D(\pe2/got [1]), .CK(clk), .RDN(
        n15094), .Q(go2[1]) );
  DRNQHSV1 \pe2/delaycell23/q_reg[7]  ( .D(\pe2/got [2]), .CK(clk), .RDN(
        n14816), .Q(go2[2]) );
  DRNQHSV1 \pe2/delaycell23/q_reg[6]  ( .D(\pe2/got [3]), .CK(clk), .RDN(
        n14784), .Q(go2[3]) );
  DRNQHSV1 \pe2/delaycell23/q_reg[5]  ( .D(\pe2/got [4]), .CK(clk), .RDN(
        n14797), .Q(go2[4]) );
  DRNQHSV1 \pe2/delaycell23/q_reg[4]  ( .D(n6721), .CK(clk), .RDN(n14814), .Q(
        go2[5]) );
  DRNQHSV1 \pe2/delaycell23/q_reg[3]  ( .D(n14822), .CK(clk), .RDN(n14725), 
        .Q(go2[6]) );
  DRNQHSV1 \pe2/delaycell23/q_reg[2]  ( .D(\pe2/got [7]), .CK(clk), .RDN(
        n14745), .Q(go2[7]) );
  DRNQHSV1 \pe2/delaycell23/q_reg[1]  ( .D(n14818), .CK(clk), .RDN(n15174), 
        .Q(go2[8]) );
  DRNQHSV2 \pe2/delaycell24/q_reg[7]  ( .D(\pe2/poht [7]), .CK(clk), .RDN(
        n14798), .Q(poh2[7]) );
  DRNQHSV2 \pe2/delaycell24/q_reg[6]  ( .D(\pe2/poht [6]), .CK(clk), .RDN(
        n14749), .Q(poh2[6]) );
  DRNQHSV2 \pe2/delaycell24/q_reg[4]  ( .D(\pe2/poht [4]), .CK(clk), .RDN(
        n14769), .Q(poh2[4]) );
  DRNQHSV2 \pe2/delaycell24/q_reg[3]  ( .D(\pe2/poht [3]), .CK(clk), .RDN(
        n14802), .Q(poh2[3]) );
  DRNQHSV1 \pe3/delaycell22/q_reg[8]  ( .D(\pe3/aot [1]), .CK(clk), .RDN(
        n14769), .Q(ao3[1]) );
  DRNQHSV1 \pe3/delaycell22/q_reg[7]  ( .D(\pe3/aot [2]), .CK(clk), .RDN(
        n14721), .Q(ao3[2]) );
  DRNQHSV1 \pe3/delaycell22/q_reg[6]  ( .D(\pe3/aot [3]), .CK(clk), .RDN(
        n14784), .Q(ao3[3]) );
  DRNQHSV1 \pe3/delaycell22/q_reg[5]  ( .D(\pe3/aot [4]), .CK(clk), .RDN(
        n14763), .Q(ao3[4]) );
  DRNQHSV1 \pe3/delaycell22/q_reg[4]  ( .D(\pe3/aot [5]), .CK(clk), .RDN(
        n14766), .Q(ao3[5]) );
  DRNQHSV1 \pe3/delaycell22/q_reg[3]  ( .D(\pe3/aot [6]), .CK(clk), .RDN(
        n14757), .Q(ao3[6]) );
  DRNQHSV1 \pe3/delaycell22/q_reg[2]  ( .D(n14738), .CK(clk), .RDN(n14731), 
        .Q(ao3[7]) );
  DRNQHSV1 \pe3/delaycell22/q_reg[1]  ( .D(n14953), .CK(clk), .RDN(n14717), 
        .Q(ao3[8]) );
  DRNQHSV1 \pe3/delaycell23/q_reg[8]  ( .D(\pe3/got [1]), .CK(clk), .RDN(
        n14797), .Q(go3[1]) );
  DRNQHSV1 \pe3/delaycell23/q_reg[7]  ( .D(\pe3/got [2]), .CK(clk), .RDN(
        n14771), .Q(go3[2]) );
  DRNQHSV1 \pe3/delaycell23/q_reg[6]  ( .D(\pe3/got [3]), .CK(clk), .RDN(
        n14814), .Q(go3[3]) );
  DRNQHSV1 \pe3/delaycell23/q_reg[5]  ( .D(\pe3/got [4]), .CK(clk), .RDN(
        n14814), .Q(go3[4]) );
  DRNQHSV1 \pe3/delaycell23/q_reg[4]  ( .D(\pe3/got [5]), .CK(clk), .RDN(
        n14771), .Q(go3[5]) );
  DRNQHSV1 \pe3/delaycell23/q_reg[3]  ( .D(\pe3/got [6]), .CK(clk), .RDN(
        n15174), .Q(go3[6]) );
  DRNQHSV1 \pe3/delaycell23/q_reg[2]  ( .D(n14931), .CK(clk), .RDN(n14749), 
        .Q(go3[7]) );
  DRNQHSV1 \pe3/delaycell23/q_reg[1]  ( .D(n15180), .CK(clk), .RDN(n14763), 
        .Q(go3[8]) );
  DRNQHSV2 \pe3/delaycell24/q_reg[7]  ( .D(\pe3/poht [7]), .CK(clk), .RDN(
        n15094), .Q(poh3[7]) );
  DRNQHSV2 \pe3/delaycell24/q_reg[6]  ( .D(\pe3/poht [6]), .CK(clk), .RDN(
        n14720), .Q(poh3[6]) );
  DRNQHSV1 \pe4/delaycell22/q_reg[8]  ( .D(\pe4/aot [1]), .CK(clk), .RDN(
        n14752), .Q(ao4[1]) );
  DRNQHSV1 \pe4/delaycell22/q_reg[7]  ( .D(\pe4/aot [2]), .CK(clk), .RDN(
        n14833), .Q(ao4[2]) );
  DRNQHSV1 \pe4/delaycell22/q_reg[6]  ( .D(\pe4/aot [3]), .CK(clk), .RDN(
        n14833), .Q(ao4[3]) );
  DRNQHSV1 \pe4/delaycell22/q_reg[5]  ( .D(\pe4/aot [4]), .CK(clk), .RDN(
        n14780), .Q(ao4[4]) );
  DRNQHSV1 \pe4/delaycell22/q_reg[3]  ( .D(\pe4/aot [6]), .CK(clk), .RDN(
        n14794), .Q(ao4[6]) );
  DRNQHSV1 \pe4/delaycell22/q_reg[1]  ( .D(n14843), .CK(clk), .RDN(n8938), .Q(
        ao4[8]) );
  DRNQHSV1 \pe4/delaycell23/q_reg[8]  ( .D(\pe4/got [1]), .CK(clk), .RDN(rst), 
        .Q(go4[1]) );
  DRNQHSV1 \pe4/delaycell23/q_reg[7]  ( .D(\pe4/got [2]), .CK(clk), .RDN(
        n14785), .Q(go4[2]) );
  DRNQHSV1 \pe4/delaycell23/q_reg[6]  ( .D(\pe4/got [3]), .CK(clk), .RDN(
        n14762), .Q(go4[3]) );
  DRNQHSV1 \pe4/delaycell23/q_reg[5]  ( .D(\pe4/got [4]), .CK(clk), .RDN(
        n14768), .Q(go4[4]) );
  DRNQHSV1 \pe4/delaycell23/q_reg[4]  ( .D(\pe4/got [5]), .CK(clk), .RDN(
        n14786), .Q(go4[5]) );
  DRNQHSV1 \pe4/delaycell23/q_reg[3]  ( .D(\pe4/got [6]), .CK(clk), .RDN(
        n14799), .Q(go4[6]) );
  DRNQHSV1 \pe4/delaycell23/q_reg[2]  ( .D(\pe4/got [7]), .CK(clk), .RDN(
        n14748), .Q(go4[7]) );
  DRNQHSV1 \pe4/delaycell24/q_reg[7]  ( .D(\pe4/poht [7]), .CK(clk), .RDN(
        n14794), .Q(poh4[7]) );
  DRNQHSV1 \pe4/delaycell24/q_reg[3]  ( .D(\pe4/poht [3]), .CK(clk), .RDN(
        n14794), .Q(poh4[3]) );
  DRNQHSV1 \pe5/delaycell22/q_reg[8]  ( .D(\pe5/aot [1]), .CK(clk), .RDN(
        n14812), .Q(ao5[1]) );
  DRNQHSV1 \pe5/delaycell22/q_reg[7]  ( .D(\pe5/aot [2]), .CK(clk), .RDN(
        n14753), .Q(ao5[2]) );
  DRNQHSV1 \pe5/delaycell22/q_reg[6]  ( .D(\pe5/aot [3]), .CK(clk), .RDN(
        n14871), .Q(ao5[3]) );
  DRNQHSV1 \pe5/delaycell22/q_reg[5]  ( .D(\pe5/aot [4]), .CK(clk), .RDN(
        n14814), .Q(ao5[4]) );
  DRNQHSV1 \pe5/delaycell22/q_reg[4]  ( .D(\pe5/aot [5]), .CK(clk), .RDN(
        n15094), .Q(ao5[5]) );
  DRNQHSV1 \pe5/delaycell22/q_reg[3]  ( .D(\pe5/aot [6]), .CK(clk), .RDN(
        n14770), .Q(ao5[6]) );
  DRNQHSV1 \pe5/delaycell22/q_reg[2]  ( .D(\pe5/aot [7]), .CK(clk), .RDN(
        n14763), .Q(ao5[7]) );
  DRNQHSV1 \pe5/delaycell23/q_reg[8]  ( .D(\pe5/got [1]), .CK(clk), .RDN(
        n14778), .Q(go5[1]) );
  DRNQHSV1 \pe5/delaycell23/q_reg[7]  ( .D(\pe5/got [2]), .CK(clk), .RDN(
        n14787), .Q(go5[2]) );
  DRNQHSV1 \pe5/delaycell23/q_reg[6]  ( .D(\pe5/got [3]), .CK(clk), .RDN(
        n14714), .Q(go5[3]) );
  DRNQHSV1 \pe5/delaycell23/q_reg[5]  ( .D(\pe5/got [4]), .CK(clk), .RDN(
        n14711), .Q(go5[4]) );
  DRNQHSV1 \pe5/delaycell23/q_reg[4]  ( .D(\pe5/got [5]), .CK(clk), .RDN(
        n14747), .Q(go5[5]) );
  DRNQHSV1 \pe5/delaycell23/q_reg[3]  ( .D(\pe5/got [6]), .CK(clk), .RDN(
        n15174), .Q(go5[6]) );
  DRNQHSV1 \pe5/delaycell23/q_reg[2]  ( .D(\pe5/got [7]), .CK(clk), .RDN(
        n14764), .Q(go5[7]) );
  DRNQHSV1 \pe5/delaycell23/q_reg[1]  ( .D(n15067), .CK(clk), .RDN(n14721), 
        .Q(go5[8]) );
  DRNQHSV2 \pe5/delaycell24/q_reg[7]  ( .D(\pe5/poht [7]), .CK(clk), .RDN(
        n14767), .Q(poh5[7]) );
  DRNQHSV2 \pe5/delaycell24/q_reg[6]  ( .D(\pe5/poht [6]), .CK(clk), .RDN(
        n14797), .Q(poh5[6]) );
  DRNQHSV2 \pe5/delaycell24/q_reg[5]  ( .D(\pe5/poht [5]), .CK(clk), .RDN(
        n14767), .Q(poh5[5]) );
  DRNQHSV2 \pe5/delaycell24/q_reg[4]  ( .D(\pe5/poht [4]), .CK(clk), .RDN(
        n14759), .Q(poh5[4]) );
  DRNQHSV2 \pe5/delaycell24/q_reg[3]  ( .D(\pe5/poht [3]), .CK(clk), .RDN(
        n14801), .Q(poh5[3]) );
  DRNQHSV2 \pe5/delaycell24/q_reg[1]  ( .D(\pe5/poht [1]), .CK(clk), .RDN(rst), 
        .Q(poh5[1]) );
  DRNQHSV1 \pe6/delaycell22/q_reg[8]  ( .D(\pe6/aot [1]), .CK(clk), .RDN(
        n14763), .Q(ao6[1]) );
  DRNQHSV1 \pe6/delaycell22/q_reg[7]  ( .D(\pe6/aot [2]), .CK(clk), .RDN(
        n14715), .Q(ao6[2]) );
  DRNQHSV1 \pe6/delaycell22/q_reg[6]  ( .D(\pe6/aot [3]), .CK(clk), .RDN(
        n14760), .Q(ao6[3]) );
  DRNQHSV1 \pe6/delaycell22/q_reg[5]  ( .D(\pe6/aot [4]), .CK(clk), .RDN(
        n14720), .Q(ao6[4]) );
  DRNQHSV1 \pe6/delaycell22/q_reg[4]  ( .D(\pe6/aot [5]), .CK(clk), .RDN(
        n14813), .Q(ao6[5]) );
  DRNQHSV1 \pe6/delaycell22/q_reg[3]  ( .D(n14849), .CK(clk), .RDN(n14816), 
        .Q(ao6[6]) );
  DRNQHSV1 \pe6/delaycell22/q_reg[2]  ( .D(\pe6/aot [7]), .CK(clk), .RDN(
        n14786), .Q(ao6[7]) );
  DRNQHSV1 \pe6/delaycell23/q_reg[8]  ( .D(\pe6/got [1]), .CK(clk), .RDN(
        n14717), .Q(go6[1]) );
  DRNQHSV1 \pe6/delaycell23/q_reg[7]  ( .D(\pe6/got [2]), .CK(clk), .RDN(
        n14817), .Q(go6[2]) );
  DRNQHSV1 \pe6/delaycell23/q_reg[6]  ( .D(\pe6/got [3]), .CK(clk), .RDN(
        n14787), .Q(go6[3]) );
  DRNQHSV1 \pe6/delaycell23/q_reg[5]  ( .D(\pe6/got [4]), .CK(clk), .RDN(
        n14759), .Q(go6[4]) );
  DRNQHSV1 \pe6/delaycell23/q_reg[4]  ( .D(\pe6/got [5]), .CK(clk), .RDN(
        n14787), .Q(go6[5]) );
  DRNQHSV1 \pe6/delaycell23/q_reg[3]  ( .D(\pe6/got [6]), .CK(clk), .RDN(
        n14785), .Q(go6[6]) );
  DRNQHSV1 \pe6/delaycell23/q_reg[2]  ( .D(n5977), .CK(clk), .RDN(n14731), .Q(
        go6[7]) );
  DRNQHSV1 \pe6/delaycell23/q_reg[1]  ( .D(\pe6/got [8]), .CK(clk), .RDN(
        n14747), .Q(go6[8]) );
  DRNQHSV2 \pe6/delaycell24/q_reg[2]  ( .D(\pe6/poht [2]), .CK(clk), .RDN(
        n14806), .Q(poh6[2]) );
  DRNQHSV2 \pe6/delaycell24/q_reg[1]  ( .D(\pe6/poht [1]), .CK(clk), .RDN(
        n15174), .Q(poh6[1]) );
  DRNQHSV1 \pe7/delaycell22/q_reg[8]  ( .D(\pe7/aot [1]), .CK(clk), .RDN(
        n14787), .Q(ao7[1]) );
  DRNQHSV1 \pe7/delaycell22/q_reg[7]  ( .D(\pe7/aot [2]), .CK(clk), .RDN(
        n14782), .Q(ao7[2]) );
  DRNQHSV1 \pe7/delaycell22/q_reg[6]  ( .D(\pe7/aot [3]), .CK(clk), .RDN(
        n14759), .Q(ao7[3]) );
  DRNQHSV1 \pe7/delaycell22/q_reg[5]  ( .D(\pe7/aot [4]), .CK(clk), .RDN(
        n14807), .Q(ao7[4]) );
  DRNQHSV1 \pe7/delaycell22/q_reg[4]  ( .D(\pe7/aot [5]), .CK(clk), .RDN(
        n14723), .Q(ao7[5]) );
  DRNQHSV1 \pe7/delaycell22/q_reg[3]  ( .D(n14705), .CK(clk), .RDN(n14764), 
        .Q(ao7[6]) );
  DRNQHSV1 \pe7/delaycell22/q_reg[2]  ( .D(n8940), .CK(clk), .RDN(n14725), .Q(
        ao7[7]) );
  DRNQHSV1 \pe7/delaycell22/q_reg[1]  ( .D(\pe7/aot [8]), .CK(clk), .RDN(
        n14764), .Q(ao7[8]) );
  DRNQHSV1 \pe7/delaycell23/q_reg[8]  ( .D(\pe7/got [1]), .CK(clk), .RDN(
        n14797), .Q(go7[1]) );
  DRNQHSV1 \pe7/delaycell23/q_reg[7]  ( .D(\pe7/got [2]), .CK(clk), .RDN(
        n14756), .Q(go7[2]) );
  DRNQHSV1 \pe7/delaycell23/q_reg[6]  ( .D(\pe7/got [3]), .CK(clk), .RDN(
        n14749), .Q(go7[3]) );
  DRNQHSV1 \pe7/delaycell23/q_reg[5]  ( .D(n6038), .CK(clk), .RDN(n14761), .Q(
        go7[4]) );
  DRNQHSV1 \pe7/delaycell23/q_reg[4]  ( .D(\pe7/got [5]), .CK(clk), .RDN(
        n14807), .Q(go7[5]) );
  DRNQHSV1 \pe7/delaycell23/q_reg[3]  ( .D(\pe7/got [6]), .CK(clk), .RDN(
        n14726), .Q(go7[6]) );
  DRNQHSV1 \pe7/delaycell23/q_reg[2]  ( .D(n14829), .CK(clk), .RDN(n14748), 
        .Q(go7[7]) );
  DRNQHSV1 \pe7/delaycell23/q_reg[1]  ( .D(n5967), .CK(clk), .RDN(n14760), .Q(
        go7[8]) );
  DRNQHSV1 \pe7/delaycell24/q_reg[7]  ( .D(\pe7/poht [7]), .CK(clk), .RDN(
        n14788), .Q(poh7[7]) );
  DRNQHSV1 \pe7/delaycell24/q_reg[6]  ( .D(\pe7/poht [6]), .CK(clk), .RDN(
        n14832), .Q(poh7[6]) );
  DRNQHSV2 \pe7/delaycell24/q_reg[5]  ( .D(\pe7/poht [5]), .CK(clk), .RDN(
        n14780), .Q(poh7[5]) );
  DRNQHSV2 \pe7/delaycell24/q_reg[3]  ( .D(\pe7/poht [3]), .CK(clk), .RDN(
        n14721), .Q(poh7[3]) );
  DRNQHSV2 \pe7/delaycell24/q_reg[1]  ( .D(\pe7/poht [1]), .CK(clk), .RDN(
        n14777), .Q(poh7[1]) );
  DRNQHSV1 \pe8/delaycell22/q_reg[8]  ( .D(\pe8/aot [1]), .CK(clk), .RDN(
        n14759), .Q(ao8[1]) );
  DRNQHSV1 \pe8/delaycell22/q_reg[7]  ( .D(\pe8/aot [2]), .CK(clk), .RDN(
        n14716), .Q(ao8[2]) );
  DRNQHSV1 \pe8/delaycell22/q_reg[6]  ( .D(\pe8/aot [3]), .CK(clk), .RDN(
        n14747), .Q(ao8[3]) );
  DRNQHSV1 \pe8/delaycell22/q_reg[5]  ( .D(\pe8/aot [4]), .CK(clk), .RDN(
        n14744), .Q(ao8[4]) );
  DRNQHSV1 \pe8/delaycell22/q_reg[4]  ( .D(n5948), .CK(clk), .RDN(n14769), .Q(
        ao8[5]) );
  DRNQHSV1 \pe8/delaycell22/q_reg[3]  ( .D(n14947), .CK(clk), .RDN(n14761), 
        .Q(ao8[6]) );
  DRNQHSV1 \pe8/delaycell22/q_reg[2]  ( .D(\pe8/aot [7]), .CK(clk), .RDN(
        n14806), .Q(ao8[7]) );
  DRNQHSV1 \pe8/delaycell22/q_reg[1]  ( .D(n14950), .CK(clk), .RDN(n14757), 
        .Q(ao8[8]) );
  DRNQHSV1 \pe8/delaycell23/q_reg[8]  ( .D(\pe8/got [1]), .CK(clk), .RDN(
        n14728), .Q(go8[1]) );
  DRNQHSV1 \pe8/delaycell23/q_reg[7]  ( .D(\pe8/got [2]), .CK(clk), .RDN(
        n14727), .Q(go8[2]) );
  DRNQHSV1 \pe8/delaycell23/q_reg[6]  ( .D(\pe8/got [3]), .CK(clk), .RDN(
        n14714), .Q(go8[3]) );
  DRNQHSV1 \pe8/delaycell23/q_reg[5]  ( .D(\pe8/got [4]), .CK(clk), .RDN(
        n14777), .Q(go8[4]) );
  DRNQHSV1 \pe8/delaycell23/q_reg[4]  ( .D(\pe8/got [5]), .CK(clk), .RDN(
        n14772), .Q(go8[5]) );
  DRNQHSV1 \pe8/delaycell23/q_reg[2]  ( .D(\pe8/got [7]), .CK(clk), .RDN(
        n14769), .Q(go8[7]) );
  DRNQHSV1 \pe8/delaycell23/q_reg[1]  ( .D(\pe8/got [8]), .CK(clk), .RDN(
        n14762), .Q(go8[8]) );
  DRNQHSV2 \pe8/delaycell24/q_reg[7]  ( .D(\pe8/poht [7]), .CK(clk), .RDN(
        n14871), .Q(poh8[7]) );
  DRNQHSV2 \pe8/delaycell24/q_reg[5]  ( .D(\pe8/poht [5]), .CK(clk), .RDN(
        n14801), .Q(poh8[5]) );
  DRNQHSV2 \pe8/delaycell24/q_reg[4]  ( .D(\pe8/poht [4]), .CK(clk), .RDN(
        n14765), .Q(poh8[4]) );
  DRNQHSV2 \pe8/delaycell24/q_reg[3]  ( .D(\pe8/poht [3]), .CK(clk), .RDN(
        n14774), .Q(poh8[3]) );
  DRNQHSV1 \pe9/delaycell22/q_reg[8]  ( .D(\pe9/aot [1]), .CK(clk), .RDN(
        n14729), .Q(ao9[1]) );
  DRNQHSV1 \pe9/delaycell22/q_reg[7]  ( .D(\pe9/aot [2]), .CK(clk), .RDN(
        n14767), .Q(ao9[2]) );
  DRNQHSV1 \pe9/delaycell22/q_reg[6]  ( .D(\pe9/aot [3]), .CK(clk), .RDN(
        n14765), .Q(ao9[3]) );
  DRNQHSV1 \pe9/delaycell22/q_reg[5]  ( .D(\pe9/aot [4]), .CK(clk), .RDN(
        n14751), .Q(ao9[4]) );
  DRNQHSV1 \pe9/delaycell22/q_reg[4]  ( .D(n8950), .CK(clk), .RDN(n14800), .Q(
        ao9[5]) );
  DRNQHSV1 \pe9/delaycell22/q_reg[3]  ( .D(\pe9/aot [6]), .CK(clk), .RDN(
        n14752), .Q(ao9[6]) );
  DRNQHSV1 \pe9/delaycell22/q_reg[2]  ( .D(\pe9/aot [7]), .CK(clk), .RDN(
        n14713), .Q(ao9[7]) );
  DRNQHSV1 \pe9/delaycell22/q_reg[1]  ( .D(n14942), .CK(clk), .RDN(n15174), 
        .Q(ao9[8]) );
  DRNQHSV1 \pe9/delaycell23/q_reg[8]  ( .D(\pe9/got [1]), .CK(clk), .RDN(
        n14776), .Q(go9[1]) );
  DRNQHSV1 \pe9/delaycell23/q_reg[7]  ( .D(\pe9/got [2]), .CK(clk), .RDN(
        n14715), .Q(go9[2]) );
  DRNQHSV1 \pe9/delaycell23/q_reg[6]  ( .D(\pe9/got [3]), .CK(clk), .RDN(
        n14813), .Q(go9[3]) );
  DRNQHSV1 \pe9/delaycell23/q_reg[5]  ( .D(\pe9/got [4]), .CK(clk), .RDN(
        n14726), .Q(go9[4]) );
  DRNQHSV1 \pe9/delaycell23/q_reg[4]  ( .D(\pe9/got [5]), .CK(clk), .RDN(
        n14730), .Q(go9[5]) );
  DRNQHSV1 \pe9/delaycell23/q_reg[3]  ( .D(\pe9/got [6]), .CK(clk), .RDN(
        n14727), .Q(go9[6]) );
  DRNQHSV1 \pe9/delaycell23/q_reg[2]  ( .D(\pe9/got [7]), .CK(clk), .RDN(
        n14712), .Q(go9[7]) );
  DRNQHSV1 \pe9/delaycell23/q_reg[1]  ( .D(n9420), .CK(clk), .RDN(rst), .Q(
        go9[8]) );
  DRNQHSV1 \pe10/delaycell22/q_reg[8]  ( .D(\pe10/aot [1]), .CK(clk), .RDN(
        n14814), .Q(ao10[1]) );
  DRNQHSV1 \pe10/delaycell22/q_reg[7]  ( .D(\pe10/aot [2]), .CK(clk), .RDN(
        n14726), .Q(ao10[2]) );
  DRNQHSV1 \pe10/delaycell22/q_reg[6]  ( .D(\pe10/aot [3]), .CK(clk), .RDN(
        n14769), .Q(ao10[3]) );
  DRNQHSV1 \pe10/delaycell22/q_reg[5]  ( .D(\pe10/aot [4]), .CK(clk), .RDN(
        n14871), .Q(ao10[4]) );
  DRNQHSV1 \pe10/delaycell22/q_reg[4]  ( .D(\pe10/aot [5]), .CK(clk), .RDN(
        n14748), .Q(ao10[5]) );
  DRNQHSV1 \pe10/delaycell22/q_reg[2]  ( .D(n14844), .CK(clk), .RDN(n14787), 
        .Q(ao10[7]) );
  DRNQHSV1 \pe10/delaycell22/q_reg[1]  ( .D(n14951), .CK(clk), .RDN(n14768), 
        .Q(ao10[8]) );
  DRNQHSV1 \pe10/delaycell23/q_reg[8]  ( .D(\pe10/got [1]), .CK(clk), .RDN(
        n14788), .Q(go10[1]) );
  DRNQHSV1 \pe10/delaycell23/q_reg[7]  ( .D(\pe10/got [2]), .CK(clk), .RDN(
        n14716), .Q(go10[2]) );
  DRNQHSV1 \pe10/delaycell23/q_reg[6]  ( .D(\pe10/got [3]), .CK(clk), .RDN(
        n14807), .Q(go10[3]) );
  DRNQHSV1 \pe10/delaycell23/q_reg[5]  ( .D(\pe10/got [4]), .CK(clk), .RDN(
        n14811), .Q(go10[4]) );
  DRNQHSV1 \pe10/delaycell23/q_reg[4]  ( .D(\pe10/got [5]), .CK(clk), .RDN(
        n14746), .Q(go10[5]) );
  DRNQHSV1 \pe10/delaycell23/q_reg[2]  ( .D(\pe10/got [7]), .CK(clk), .RDN(
        n14816), .Q(go10[7]) );
  DRNQHSV1 \pe10/delaycell23/q_reg[1]  ( .D(\pe10/got [8]), .CK(clk), .RDN(
        n14783), .Q(go10[8]) );
  DRNQHSV2 \pe10/delaycell24/q_reg[4]  ( .D(\pe10/poht [4]), .CK(clk), .RDN(
        n14784), .Q(poh10[4]) );
  DRNQHSV2 \pe10/delaycell24/q_reg[3]  ( .D(\pe10/poht [3]), .CK(clk), .RDN(
        n14788), .Q(poh10[3]) );
  DRNQHSV2 \pe10/delaycell24/q_reg[2]  ( .D(\pe10/poht [2]), .CK(clk), .RDN(
        n14767), .Q(poh10[2]) );
  DRNQHSV1 \pe11/delaycell22/q_reg[8]  ( .D(\pe11/aot [1]), .CK(clk), .RDN(
        n14778), .Q(ao11[1]) );
  DRNQHSV1 \pe11/delaycell22/q_reg[7]  ( .D(\pe11/aot [2]), .CK(clk), .RDN(
        n14746), .Q(ao11[2]) );
  DRNQHSV1 \pe11/delaycell22/q_reg[6]  ( .D(\pe11/aot [3]), .CK(clk), .RDN(
        n14729), .Q(ao11[3]) );
  DRNQHSV1 \pe11/delaycell22/q_reg[5]  ( .D(\pe11/aot [4]), .CK(clk), .RDN(
        n14765), .Q(ao11[4]) );
  DRNQHSV1 \pe11/delaycell22/q_reg[4]  ( .D(\pe11/aot [5]), .CK(clk), .RDN(rst), .Q(ao11[5]) );
  DRNQHSV1 \pe11/delaycell22/q_reg[3]  ( .D(\pe11/aot [6]), .CK(clk), .RDN(
        n14775), .Q(ao11[6]) );
  DRNQHSV1 \pe11/delaycell22/q_reg[2]  ( .D(n14837), .CK(clk), .RDN(n14833), 
        .Q(ao11[7]) );
  DRNQHSV1 \pe11/delaycell23/q_reg[8]  ( .D(\pe11/got [1]), .CK(clk), .RDN(
        n14799), .Q(go11[1]) );
  DRNQHSV1 \pe11/delaycell23/q_reg[7]  ( .D(\pe11/got [2]), .CK(clk), .RDN(
        n14785), .Q(go11[2]) );
  DRNQHSV1 \pe11/delaycell23/q_reg[6]  ( .D(\pe11/got [3]), .CK(clk), .RDN(
        n14764), .Q(go11[3]) );
  DRNQHSV1 \pe11/delaycell23/q_reg[5]  ( .D(\pe11/got [4]), .CK(clk), .RDN(
        n14751), .Q(go11[4]) );
  DRNQHSV1 \pe11/delaycell23/q_reg[4]  ( .D(\pe11/got [5]), .CK(clk), .RDN(
        n14713), .Q(go11[5]) );
  DRNQHSV1 \pe11/delaycell23/q_reg[2]  ( .D(\pe11/got [7]), .CK(clk), .RDN(
        n14788), .Q(go11[7]) );
  DRNQHSV1 \pe11/delaycell23/q_reg[1]  ( .D(n15179), .CK(clk), .RDN(n14788), 
        .Q(go11[8]) );
  DRNQHSV1 \pe11/delaycell24/q_reg[7]  ( .D(\pe11/poht [7]), .CK(clk), .RDN(
        n14722), .Q(poh11[7]) );
  DRNQHSV1 \pe12/delaycell22/q_reg[8]  ( .D(\pe12/aot [1]), .CK(clk), .RDN(
        n14785), .Q(ao12[1]) );
  DRNQHSV1 \pe12/delaycell22/q_reg[7]  ( .D(\pe12/aot [2]), .CK(clk), .RDN(
        n14779), .Q(ao12[2]) );
  DRNQHSV1 \pe12/delaycell22/q_reg[6]  ( .D(\pe12/aot [3]), .CK(clk), .RDN(
        n14802), .Q(ao12[3]) );
  DRNQHSV1 \pe12/delaycell22/q_reg[5]  ( .D(\pe12/aot [4]), .CK(clk), .RDN(
        n14746), .Q(ao12[4]) );
  DRNQHSV1 \pe12/delaycell22/q_reg[4]  ( .D(\pe12/aot [5]), .CK(clk), .RDN(
        n14800), .Q(ao12[5]) );
  DRNQHSV1 \pe12/delaycell22/q_reg[3]  ( .D(\pe12/aot [6]), .CK(clk), .RDN(
        n14716), .Q(ao12[6]) );
  DRNQHSV1 \pe12/delaycell22/q_reg[2]  ( .D(n14948), .CK(clk), .RDN(n14783), 
        .Q(ao12[7]) );
  DRNQHSV1 \pe12/delaycell22/q_reg[1]  ( .D(n14876), .CK(clk), .RDN(n14757), 
        .Q(ao12[8]) );
  DRNQHSV1 \pe12/delaycell23/q_reg[8]  ( .D(\pe12/got [1]), .CK(clk), .RDN(
        n14716), .Q(go12[1]) );
  DRNQHSV1 \pe12/delaycell23/q_reg[7]  ( .D(\pe12/got [2]), .CK(clk), .RDN(
        n14804), .Q(go12[2]) );
  DRNQHSV1 \pe12/delaycell23/q_reg[6]  ( .D(\pe12/got [3]), .CK(clk), .RDN(
        n14807), .Q(go12[3]) );
  DRNQHSV1 \pe12/delaycell23/q_reg[5]  ( .D(\pe12/got [4]), .CK(clk), .RDN(
        n14781), .Q(go12[4]) );
  DRNQHSV1 \pe12/delaycell23/q_reg[4]  ( .D(\pe12/got [5]), .CK(clk), .RDN(
        n14780), .Q(go12[5]) );
  DRNQHSV1 \pe12/delaycell23/q_reg[3]  ( .D(\pe12/got [6]), .CK(clk), .RDN(
        n8938), .Q(go12[6]) );
  DRNQHSV1 \pe12/delaycell23/q_reg[2]  ( .D(\pe12/got [7]), .CK(clk), .RDN(
        n14812), .Q(go12[7]) );
  DRNQHSV1 \pe12/delaycell23/q_reg[1]  ( .D(n5958), .CK(clk), .RDN(n14744), 
        .Q(go12[8]) );
  DRNQHSV1 \pe12/delaycell24/q_reg[7]  ( .D(\pe12/poht [7]), .CK(clk), .RDN(
        n14793), .Q(poh12[7]) );
  DRNQHSV1 \pe12/delaycell24/q_reg[6]  ( .D(\pe12/poht [6]), .CK(clk), .RDN(
        n14802), .Q(poh12[6]) );
  DRNQHSV2 \pe12/delaycell24/q_reg[4]  ( .D(\pe12/poht [4]), .CK(clk), .RDN(
        n14803), .Q(poh12[4]) );
  DRNQHSV2 \pe12/delaycell24/q_reg[3]  ( .D(\pe12/poht [3]), .CK(clk), .RDN(
        n14767), .Q(poh12[3]) );
  DRNQHSV2 \pe12/delaycell24/q_reg[2]  ( .D(\pe12/poht [2]), .CK(clk), .RDN(
        n14749), .Q(poh12[2]) );
  DRNQHSV1 \pe13/delaycell22/q_reg[8]  ( .D(\pe13/aot [1]), .CK(clk), .RDN(
        n14788), .Q(ao13[1]) );
  DRNQHSV1 \pe13/delaycell22/q_reg[7]  ( .D(\pe13/aot [2]), .CK(clk), .RDN(
        n14769), .Q(ao13[2]) );
  DRNQHSV1 \pe13/delaycell22/q_reg[6]  ( .D(\pe13/aot [3]), .CK(clk), .RDN(
        n14804), .Q(ao13[3]) );
  DRNQHSV1 \pe13/delaycell22/q_reg[5]  ( .D(\pe13/aot [4]), .CK(clk), .RDN(
        n14715), .Q(ao13[4]) );
  DRNQHSV1 \pe13/delaycell22/q_reg[4]  ( .D(\pe13/aot [5]), .CK(clk), .RDN(
        n14797), .Q(ao13[5]) );
  DRNQHSV1 \pe13/delaycell22/q_reg[3]  ( .D(\pe13/aot [6]), .CK(clk), .RDN(
        n14778), .Q(ao13[6]) );
  DRNQHSV1 \pe13/delaycell22/q_reg[2]  ( .D(\pe13/aot [7]), .CK(clk), .RDN(
        n14782), .Q(ao13[7]) );
  DRNQHSV1 \pe13/delaycell22/q_reg[1]  ( .D(n14939), .CK(clk), .RDN(n14729), 
        .Q(ao13[8]) );
  DRNQHSV1 \pe13/delaycell23/q_reg[8]  ( .D(\pe13/got [1]), .CK(clk), .RDN(
        n14759), .Q(go13[1]) );
  DRNQHSV1 \pe13/delaycell23/q_reg[7]  ( .D(\pe13/got [2]), .CK(clk), .RDN(
        n14725), .Q(go13[2]) );
  DRNQHSV1 \pe13/delaycell23/q_reg[6]  ( .D(\pe13/got [3]), .CK(clk), .RDN(
        n14767), .Q(go13[3]) );
  DRNQHSV1 \pe13/delaycell23/q_reg[5]  ( .D(\pe13/got [4]), .CK(clk), .RDN(
        n14716), .Q(go13[4]) );
  DRNQHSV1 \pe13/delaycell23/q_reg[4]  ( .D(\pe13/got [5]), .CK(clk), .RDN(
        n14783), .Q(go13[5]) );
  DRNQHSV1 \pe13/delaycell23/q_reg[3]  ( .D(\pe13/got [6]), .CK(clk), .RDN(
        n14725), .Q(go13[6]) );
  DRNQHSV1 \pe13/delaycell23/q_reg[2]  ( .D(\pe13/got [7]), .CK(clk), .RDN(
        n14766), .Q(go13[7]) );
  DRNQHSV1 \pe13/delaycell23/q_reg[1]  ( .D(n14750), .CK(clk), .RDN(n14721), 
        .Q(go13[8]) );
  DRNQHSV2 \pe13/delaycell24/q_reg[7]  ( .D(\pe13/poht [7]), .CK(clk), .RDN(
        n15174), .Q(poh13[7]) );
  DRNQHSV1 \pe13/delaycell24/q_reg[6]  ( .D(\pe13/poht [6]), .CK(clk), .RDN(
        n14809), .Q(poh13[6]) );
  DRNQHSV1 \pe13/delaycell24/q_reg[3]  ( .D(\pe13/poht [3]), .CK(clk), .RDN(
        n14833), .Q(poh13[3]) );
  DRNQHSV1 \pe13/delaycell24/q_reg[1]  ( .D(\pe13/poht [1]), .CK(clk), .RDN(
        n14806), .Q(poh13[1]) );
  DRNQHSV1 \pe14/delaycell22/q_reg[8]  ( .D(\pe14/aot [1]), .CK(clk), .RDN(
        n14811), .Q(ao14[1]) );
  DRNQHSV1 \pe14/delaycell22/q_reg[7]  ( .D(\pe14/aot [2]), .CK(clk), .RDN(
        n14747), .Q(ao14[2]) );
  DRNQHSV1 \pe14/delaycell22/q_reg[6]  ( .D(\pe14/aot [3]), .CK(clk), .RDN(
        n14727), .Q(ao14[3]) );
  DRNQHSV1 \pe14/delaycell22/q_reg[5]  ( .D(\pe14/aot [4]), .CK(clk), .RDN(
        n14753), .Q(ao14[4]) );
  DRNQHSV1 \pe14/delaycell22/q_reg[4]  ( .D(\pe14/aot [5]), .CK(clk), .RDN(
        n14785), .Q(ao14[5]) );
  DRNQHSV1 \pe14/delaycell22/q_reg[3]  ( .D(n14889), .CK(clk), .RDN(n14832), 
        .Q(ao14[6]) );
  DRNQHSV1 \pe14/delaycell22/q_reg[2]  ( .D(n14706), .CK(clk), .RDN(n14804), 
        .Q(ao14[7]) );
  DRNQHSV1 \pe14/delaycell22/q_reg[1]  ( .D(n14891), .CK(clk), .RDN(n14789), 
        .Q(ao14[8]) );
  DRNQHSV1 \pe14/delaycell23/q_reg[8]  ( .D(\pe14/got [1]), .CK(clk), .RDN(
        n14772), .Q(go14[1]) );
  DRNQHSV1 \pe14/delaycell23/q_reg[7]  ( .D(\pe14/got [2]), .CK(clk), .RDN(
        n14815), .Q(go14[2]) );
  DRNQHSV1 \pe14/delaycell23/q_reg[6]  ( .D(\pe14/got [3]), .CK(clk), .RDN(
        n14793), .Q(go14[3]) );
  DRNQHSV1 \pe14/delaycell23/q_reg[5]  ( .D(\pe14/got [4]), .CK(clk), .RDN(
        n14732), .Q(go14[4]) );
  DRNQHSV1 \pe14/delaycell23/q_reg[4]  ( .D(\pe14/got [5]), .CK(clk), .RDN(
        n14779), .Q(go14[5]) );
  DRNQHSV1 \pe14/delaycell23/q_reg[3]  ( .D(\pe14/got [6]), .CK(clk), .RDN(
        n14722), .Q(go14[6]) );
  DRNQHSV1 \pe14/delaycell23/q_reg[2]  ( .D(\pe14/got [7]), .CK(clk), .RDN(
        n14761), .Q(go14[7]) );
  DRNQHSV1 \pe14/delaycell23/q_reg[1]  ( .D(n8955), .CK(clk), .RDN(n14789), 
        .Q(go14[8]) );
  DRNQHSV2 \pe14/delaycell24/q_reg[7]  ( .D(\pe14/poht [7]), .CK(clk), .RDN(
        n14727), .Q(poh14[7]) );
  DRNQHSV2 \pe14/delaycell24/q_reg[6]  ( .D(\pe14/poht [6]), .CK(clk), .RDN(
        n14751), .Q(poh14[6]) );
  DRNQHSV2 \pe14/delaycell24/q_reg[3]  ( .D(\pe14/poht [3]), .CK(clk), .RDN(
        n14765), .Q(poh14[3]) );
  DRNQHSV2 \pe14/delaycell24/q_reg[1]  ( .D(n15199), .CK(clk), .RDN(n14786), 
        .Q(poh14[1]) );
  DRNQHSV1 \pe15/delaycell22/q_reg[8]  ( .D(\pe15/aot [1]), .CK(clk), .RDN(
        n14804), .Q(ao15[1]) );
  DRNQHSV1 \pe15/delaycell22/q_reg[7]  ( .D(\pe15/aot [2]), .CK(clk), .RDN(
        n14780), .Q(ao15[2]) );
  DRNQHSV1 \pe15/delaycell22/q_reg[6]  ( .D(\pe15/aot [3]), .CK(clk), .RDN(
        n14812), .Q(ao15[3]) );
  DRNQHSV1 \pe15/delaycell22/q_reg[5]  ( .D(\pe15/aot [4]), .CK(clk), .RDN(
        n14759), .Q(ao15[4]) );
  DRNQHSV1 \pe15/delaycell22/q_reg[4]  ( .D(\pe15/aot [5]), .CK(clk), .RDN(
        n14832), .Q(ao15[5]) );
  DRNQHSV1 \pe15/delaycell22/q_reg[3]  ( .D(n14739), .CK(clk), .RDN(n14722), 
        .Q(ao15[6]) );
  DRNQHSV1 \pe15/delaycell22/q_reg[2]  ( .D(n14936), .CK(clk), .RDN(n14763), 
        .Q(ao15[7]) );
  DRNQHSV1 \pe15/delaycell22/q_reg[1]  ( .D(n14937), .CK(clk), .RDN(n14812), 
        .Q(ao15[8]) );
  DRNQHSV1 \pe15/delaycell23/q_reg[8]  ( .D(\pe15/got [1]), .CK(clk), .RDN(
        n14779), .Q(go15[1]) );
  DRNQHSV1 \pe15/delaycell23/q_reg[7]  ( .D(\pe15/got [2]), .CK(clk), .RDN(rst), .Q(go15[2]) );
  DRNQHSV1 \pe15/delaycell23/q_reg[6]  ( .D(\pe15/got [3]), .CK(clk), .RDN(
        n14871), .Q(go15[3]) );
  DRNQHSV1 \pe15/delaycell23/q_reg[5]  ( .D(\pe15/got [4]), .CK(clk), .RDN(
        n14716), .Q(go15[4]) );
  DRNQHSV1 \pe15/delaycell23/q_reg[4]  ( .D(\pe15/got [5]), .CK(clk), .RDN(
        n14755), .Q(go15[5]) );
  DRNQHSV1 \pe15/delaycell23/q_reg[2]  ( .D(n14864), .CK(clk), .RDN(n14806), 
        .Q(go15[7]) );
  DRNQHSV1 \pe15/delaycell23/q_reg[1]  ( .D(n15178), .CK(clk), .RDN(n14773), 
        .Q(go15[8]) );
  DRNQHSV2 \pe15/delaycell24/q_reg[7]  ( .D(\pe15/poht [7]), .CK(clk), .RDN(
        n14718), .Q(poh15[7]) );
  DRNQHSV2 \pe15/delaycell24/q_reg[6]  ( .D(\pe15/poht [6]), .CK(clk), .RDN(
        n14783), .Q(poh15[6]) );
  DRNQHSV2 \pe15/delaycell24/q_reg[3]  ( .D(\pe15/poht [3]), .CK(clk), .RDN(
        n15094), .Q(poh15[3]) );
  DRNQHSV2 \pe15/delaycell24/q_reg[1]  ( .D(\pe15/poht [1]), .CK(clk), .RDN(
        n14719), .Q(poh15[1]) );
  DRNQHSV1 \pe16/delaycell22/q_reg[8]  ( .D(\pe16/aot [1]), .CK(clk), .RDN(
        n14796), .Q(ao16[1]) );
  DRNQHSV1 \pe16/delaycell22/q_reg[7]  ( .D(\pe16/aot [2]), .CK(clk), .RDN(
        n14781), .Q(ao16[2]) );
  DRNQHSV1 \pe16/delaycell22/q_reg[6]  ( .D(\pe16/aot [3]), .CK(clk), .RDN(
        n14798), .Q(ao16[3]) );
  DRNQHSV1 \pe16/delaycell22/q_reg[5]  ( .D(\pe16/aot [4]), .CK(clk), .RDN(
        n14784), .Q(ao16[4]) );
  DRNQHSV1 \pe16/delaycell22/q_reg[4]  ( .D(\pe16/aot [5]), .CK(clk), .RDN(
        n14783), .Q(ao16[5]) );
  DRNQHSV1 \pe16/delaycell22/q_reg[3]  ( .D(n14932), .CK(clk), .RDN(n14777), 
        .Q(ao16[6]) );
  DRNQHSV1 \pe16/delaycell22/q_reg[2]  ( .D(\pe16/aot [7]), .CK(clk), .RDN(
        n14745), .Q(ao16[7]) );
  DRNQHSV1 \pe16/delaycell22/q_reg[1]  ( .D(\pe16/aot [8]), .CK(clk), .RDN(rst), .Q(ao16[8]) );
  DRNQHSV1 \pe16/delaycell23/q_reg[8]  ( .D(\pe16/got [1]), .CK(clk), .RDN(
        n14729), .Q(go16[1]) );
  DRNQHSV1 \pe16/delaycell23/q_reg[7]  ( .D(\pe16/got [2]), .CK(clk), .RDN(
        n14718), .Q(go16[2]) );
  DRNQHSV1 \pe16/delaycell23/q_reg[5]  ( .D(\pe16/got [4]), .CK(clk), .RDN(
        n14711), .Q(go16[4]) );
  DRNQHSV1 \pe16/delaycell23/q_reg[4]  ( .D(\pe16/got [5]), .CK(clk), .RDN(
        n14779), .Q(go16[5]) );
  DRNQHSV1 \pe16/delaycell23/q_reg[3]  ( .D(\pe16/got [6]), .CK(clk), .RDN(
        n14787), .Q(go16[6]) );
  DRNQHSV1 \pe16/delaycell23/q_reg[2]  ( .D(n14873), .CK(clk), .RDN(n14796), 
        .Q(go16[7]) );
  DRNQHSV1 \pe16/delaycell23/q_reg[1]  ( .D(n11179), .CK(clk), .RDN(n14798), 
        .Q(go16[8]) );
  DRNQHSV1 \pe16/delaycell24/q_reg[2]  ( .D(\pe16/poht [2]), .CK(clk), .RDN(
        n14798), .Q(poh16[2]) );
  DRNQHSV2 \pe16/delaycell24/q_reg[1]  ( .D(\pe16/poht [1]), .CK(clk), .RDN(
        n14798), .Q(poh16[1]) );
  DRNQHSV1 \pe17/delaycell22/q_reg[8]  ( .D(\pe17/aot [1]), .CK(clk), .RDN(
        n14723), .Q(ao17[1]) );
  DRNQHSV1 \pe17/delaycell22/q_reg[7]  ( .D(\pe17/aot [2]), .CK(clk), .RDN(
        n14785), .Q(ao17[2]) );
  DRNQHSV1 \pe17/delaycell22/q_reg[6]  ( .D(\pe17/aot [3]), .CK(clk), .RDN(
        n14802), .Q(ao17[3]) );
  DRNQHSV1 \pe17/delaycell22/q_reg[5]  ( .D(\pe17/aot [4]), .CK(clk), .RDN(
        n14802), .Q(ao17[4]) );
  DRNQHSV1 \pe17/delaycell22/q_reg[4]  ( .D(\pe17/aot [5]), .CK(clk), .RDN(
        n14798), .Q(ao17[5]) );
  DRNQHSV1 \pe17/delaycell22/q_reg[2]  ( .D(\pe17/aot [7]), .CK(clk), .RDN(
        n14783), .Q(ao17[7]) );
  DRNQHSV1 \pe17/delaycell23/q_reg[8]  ( .D(\pe17/got [1]), .CK(clk), .RDN(
        n14753), .Q(go17[1]) );
  DRNQHSV1 \pe17/delaycell23/q_reg[7]  ( .D(\pe17/got [2]), .CK(clk), .RDN(
        n14810), .Q(go17[2]) );
  DRNQHSV1 \pe17/delaycell23/q_reg[6]  ( .D(\pe17/got [3]), .CK(clk), .RDN(
        n14775), .Q(go17[3]) );
  DRNQHSV1 \pe17/delaycell23/q_reg[5]  ( .D(\pe17/got [4]), .CK(clk), .RDN(
        n14727), .Q(go17[4]) );
  DRNQHSV1 \pe17/delaycell23/q_reg[4]  ( .D(\pe17/got [5]), .CK(clk), .RDN(
        n14789), .Q(go17[5]) );
  DRNQHSV1 \pe17/delaycell23/q_reg[3]  ( .D(\pe17/got [6]), .CK(clk), .RDN(
        n14770), .Q(go17[6]) );
  DRNQHSV1 \pe17/delaycell23/q_reg[2]  ( .D(\pe17/got [7]), .CK(clk), .RDN(
        n14769), .Q(go17[7]) );
  DRNQHSV1 \pe17/delaycell23/q_reg[1]  ( .D(\pe17/got [8]), .CK(clk), .RDN(
        n15094), .Q(go17[8]) );
  DRNQHSV2 \pe17/delaycell24/q_reg[4]  ( .D(\pe17/poht [4]), .CK(clk), .RDN(
        n14711), .Q(poh17[4]) );
  DRNQHSV1 \pe18/delaycell22/q_reg[8]  ( .D(\pe18/aot [1]), .CK(clk), .RDN(
        n14786), .Q(ao18[1]) );
  DRNQHSV1 \pe18/delaycell22/q_reg[7]  ( .D(\pe18/aot [2]), .CK(clk), .RDN(
        n14774), .Q(ao18[2]) );
  DRNQHSV1 \pe18/delaycell22/q_reg[6]  ( .D(\pe18/aot [3]), .CK(clk), .RDN(
        n14793), .Q(ao18[3]) );
  DRNQHSV1 \pe18/delaycell22/q_reg[5]  ( .D(\pe18/aot [4]), .CK(clk), .RDN(
        n14759), .Q(ao18[4]) );
  DRNQHSV1 \pe18/delaycell22/q_reg[4]  ( .D(\pe18/aot [5]), .CK(clk), .RDN(
        n14796), .Q(ao18[5]) );
  DRNQHSV1 \pe18/delaycell22/q_reg[3]  ( .D(n14894), .CK(clk), .RDN(n14753), 
        .Q(ao18[6]) );
  DRNQHSV1 \pe18/delaycell22/q_reg[2]  ( .D(\pe18/aot [7]), .CK(clk), .RDN(
        n14766), .Q(ao18[7]) );
  DRNQHSV1 \pe18/delaycell22/q_reg[1]  ( .D(n11988), .CK(clk), .RDN(n14789), 
        .Q(ao18[8]) );
  DRNQHSV1 \pe18/delaycell23/q_reg[8]  ( .D(\pe18/got [1]), .CK(clk), .RDN(
        n14788), .Q(go18[1]) );
  DRNQHSV1 \pe18/delaycell23/q_reg[7]  ( .D(\pe18/got [2]), .CK(clk), .RDN(
        n14832), .Q(go18[2]) );
  DRNQHSV1 \pe18/delaycell23/q_reg[6]  ( .D(\pe18/got [3]), .CK(clk), .RDN(
        n14712), .Q(go18[3]) );
  DRNQHSV1 \pe18/delaycell23/q_reg[5]  ( .D(\pe18/got [4]), .CK(clk), .RDN(rst), .Q(go18[4]) );
  DRNQHSV1 \pe18/delaycell23/q_reg[4]  ( .D(\pe18/got [5]), .CK(clk), .RDN(
        n14798), .Q(go18[5]) );
  DRNQHSV1 \pe18/delaycell23/q_reg[3]  ( .D(n6039), .CK(clk), .RDN(n14798), 
        .Q(go18[6]) );
  DRNQHSV1 \pe18/delaycell23/q_reg[2]  ( .D(\pe18/got [7]), .CK(clk), .RDN(
        n8938), .Q(go18[7]) );
  DRNQHSV1 \pe18/delaycell23/q_reg[1]  ( .D(n5997), .CK(clk), .RDN(n14727), 
        .Q(go18[8]) );
  DRNQHSV1 \pe19/delaycell22/q_reg[8]  ( .D(\pe19/aot [1]), .CK(clk), .RDN(
        n14803), .Q(ao19[1]) );
  DRNQHSV1 \pe19/delaycell22/q_reg[7]  ( .D(\pe19/aot [2]), .CK(clk), .RDN(
        n14747), .Q(ao19[2]) );
  DRNQHSV1 \pe19/delaycell22/q_reg[6]  ( .D(\pe19/aot [3]), .CK(clk), .RDN(
        n14771), .Q(ao19[3]) );
  DRNQHSV1 \pe19/delaycell22/q_reg[5]  ( .D(\pe19/aot [4]), .CK(clk), .RDN(
        n14810), .Q(ao19[4]) );
  DRNQHSV1 \pe19/delaycell22/q_reg[3]  ( .D(\pe19/aot [6]), .CK(clk), .RDN(
        n14714), .Q(ao19[6]) );
  DRNQHSV1 \pe19/delaycell22/q_reg[1]  ( .D(n14915), .CK(clk), .RDN(n14792), 
        .Q(ao19[8]) );
  DRNQHSV1 \pe19/delaycell23/q_reg[8]  ( .D(\pe19/got [1]), .CK(clk), .RDN(
        n14773), .Q(go19[1]) );
  DRNQHSV1 \pe19/delaycell23/q_reg[7]  ( .D(\pe19/got [2]), .CK(clk), .RDN(
        n14752), .Q(go19[2]) );
  DRNQHSV1 \pe19/delaycell23/q_reg[6]  ( .D(\pe19/got [3]), .CK(clk), .RDN(
        n14710), .Q(go19[3]) );
  DRNQHSV1 \pe19/delaycell23/q_reg[5]  ( .D(\pe19/got [4]), .CK(clk), .RDN(
        n14716), .Q(go19[4]) );
  DRNQHSV1 \pe19/delaycell23/q_reg[4]  ( .D(\pe19/got [5]), .CK(clk), .RDN(
        n14833), .Q(go19[5]) );
  DRNQHSV1 \pe19/delaycell23/q_reg[2]  ( .D(n14841), .CK(clk), .RDN(n14751), 
        .Q(go19[7]) );
  DRNQHSV1 \pe19/delaycell23/q_reg[1]  ( .D(n14859), .CK(clk), .RDN(n14767), 
        .Q(go19[8]) );
  DRNQHSV1 \pe19/delaycell24/q_reg[7]  ( .D(\pe19/poht [7]), .CK(clk), .RDN(
        n14808), .Q(poh19[7]) );
  DRNQHSV1 \pe19/delaycell24/q_reg[6]  ( .D(\pe19/poht [6]), .CK(clk), .RDN(
        n14804), .Q(poh19[6]) );
  DRNQHSV1 \pe19/delaycell24/q_reg[5]  ( .D(\pe19/poht [5]), .CK(clk), .RDN(
        n14779), .Q(poh19[5]) );
  DRNQHSV1 \pe19/delaycell24/q_reg[4]  ( .D(\pe19/poht [4]), .CK(clk), .RDN(
        n14754), .Q(poh19[4]) );
  DRNQHSV1 \pe19/delaycell24/q_reg[3]  ( .D(\pe19/poht [3]), .CK(clk), .RDN(
        n14803), .Q(poh19[3]) );
  DRNQHSV1 \pe19/delaycell24/q_reg[2]  ( .D(\pe19/poht [2]), .CK(clk), .RDN(
        n14775), .Q(poh19[2]) );
  DRNQHSV1 \pe19/delaycell24/q_reg[1]  ( .D(\pe19/poht [1]), .CK(clk), .RDN(
        n14729), .Q(poh19[1]) );
  DRNQHSV1 \pe20/delaycell22/q_reg[8]  ( .D(\pe20/aot [1]), .CK(clk), .RDN(
        n14817), .Q(ao20[1]) );
  DRNQHSV1 \pe20/delaycell22/q_reg[7]  ( .D(\pe20/aot [2]), .CK(clk), .RDN(
        n14772), .Q(ao20[2]) );
  DRNQHSV1 \pe20/delaycell22/q_reg[6]  ( .D(\pe20/aot [3]), .CK(clk), .RDN(
        n14748), .Q(ao20[3]) );
  DRNQHSV1 \pe20/delaycell22/q_reg[5]  ( .D(\pe20/aot [4]), .CK(clk), .RDN(
        n14760), .Q(ao20[4]) );
  DRNQHSV1 \pe20/delaycell22/q_reg[4]  ( .D(\pe20/aot [5]), .CK(clk), .RDN(
        n14801), .Q(ao20[5]) );
  DRNQHSV1 \pe20/delaycell22/q_reg[3]  ( .D(n14946), .CK(clk), .RDN(n14730), 
        .Q(ao20[6]) );
  DRNQHSV1 \pe20/delaycell22/q_reg[2]  ( .D(n8937), .CK(clk), .RDN(n14759), 
        .Q(ao20[7]) );
  DRNQHSV1 \pe20/delaycell23/q_reg[8]  ( .D(\pe20/got [1]), .CK(clk), .RDN(
        n14785), .Q(go20[1]) );
  DRNQHSV1 \pe20/delaycell23/q_reg[7]  ( .D(\pe20/got [2]), .CK(clk), .RDN(
        n15173), .Q(go20[2]) );
  DRNQHSV1 \pe20/delaycell23/q_reg[6]  ( .D(\pe20/got [3]), .CK(clk), .RDN(
        n14746), .Q(go20[3]) );
  DRNQHSV1 \pe20/delaycell23/q_reg[5]  ( .D(\pe20/got [4]), .CK(clk), .RDN(
        n14719), .Q(go20[4]) );
  DRNQHSV1 \pe20/delaycell23/q_reg[4]  ( .D(\pe20/got [5]), .CK(clk), .RDN(
        n14794), .Q(go20[5]) );
  DRNQHSV1 \pe20/delaycell23/q_reg[3]  ( .D(\pe20/got [6]), .CK(clk), .RDN(
        n14757), .Q(go20[6]) );
  DRNQHSV1 \pe20/delaycell23/q_reg[1]  ( .D(n14865), .CK(clk), .RDN(n14756), 
        .Q(go20[8]) );
  DRNQHSV1 \pe20/delaycell24/q_reg[3]  ( .D(\pe20/poht [3]), .CK(clk), .RDN(
        n14771), .Q(poh20[3]) );
  DRNQHSV1 \pe13/delaycell21/q_reg[6]  ( .D(n15188), .CK(clk), .RDN(n14776), 
        .Q(\pe13/ti_7t [6]) );
  DRNQHSV1 \pe2/delaycell21/q_reg[6]  ( .D(n6170), .CK(clk), .RDN(n14762), .Q(
        \pe2/ti_7t [6]) );
  DRNQHSV1 \pe21/delaycell24/q_reg[7]  ( .D(\pe21/poht [7]), .CK(clk), .RDN(
        n14806), .Q(poh21[7]) );
  DRNQHSV1 \pe1/delaycell21/q_reg[5]  ( .D(\pe1/ti_7[5] ), .CK(clk), .RDN(
        n14816), .Q(\pe1/ti_7t [5]) );
  DRNQHSV1 \pe4/delaycell21/q_reg[7]  ( .D(n6706), .CK(clk), .RDN(n14810), .Q(
        \pe4/ti_7t [7]) );
  DRNQHSV1 \pe10/delaycell21/q_reg[7]  ( .D(n15187), .CK(clk), .RDN(n14756), 
        .Q(\pe10/ti_7t [7]) );
  DRNQHSV1 \pe11/delaycell21/q_reg[6]  ( .D(n14830), .CK(clk), .RDN(n14832), 
        .Q(\pe11/ti_7t [6]) );
  DRNQHSV1 \pe12/delaycell21/q_reg[4]  ( .D(n14943), .CK(clk), .RDN(n14764), 
        .Q(\pe12/ti_7t [4]) );
  DRNQHSV1 \pe12/delaycell21/q_reg[6]  ( .D(n15190), .CK(clk), .RDN(n8938), 
        .Q(\pe12/ti_7t [6]) );
  DRNQHSV1 \pe14/delaycell21/q_reg[6]  ( .D(n14855), .CK(clk), .RDN(n14748), 
        .Q(\pe14/ti_7t [6]) );
  DRNQHSV1 \pe15/delaycell21/q_reg[6]  ( .D(n14914), .CK(clk), .RDN(n14710), 
        .Q(\pe15/ti_7t [6]) );
  DRNQHSV1 \pe18/delaycell21/q_reg[6]  ( .D(n15168), .CK(clk), .RDN(n14817), 
        .Q(\pe18/ti_7t [6]) );
  DRNQHSV1 \pe19/delaycell21/q_reg[5]  ( .D(n15084), .CK(clk), .RDN(n14780), 
        .Q(\pe19/ti_7t [5]) );
  DRNQHSV2 \pe1/delaycell3/q_reg[2]  ( .D(bi[7]), .CK(clk), .RDN(rst), .Q(
        bo1[7]) );
  DRNQHSV2 \pe2/delaycell3/q_reg[8]  ( .D(bo1[1]), .CK(clk), .RDN(n14799), .Q(
        bo2[1]) );
  DRNQHSV2 \pe2/delaycell3/q_reg[7]  ( .D(bo1[2]), .CK(clk), .RDN(n14719), .Q(
        bo2[2]) );
  DRNQHSV2 \pe2/delaycell3/q_reg[6]  ( .D(bo1[3]), .CK(clk), .RDN(n14801), .Q(
        bo2[3]) );
  DRNQHSV2 \pe2/delaycell3/q_reg[5]  ( .D(bo1[4]), .CK(clk), .RDN(n14794), .Q(
        bo2[4]) );
  DRNQHSV2 \pe2/delaycell3/q_reg[4]  ( .D(bo1[5]), .CK(clk), .RDN(n14802), .Q(
        bo2[5]) );
  DRNQHSV2 \pe2/delaycell3/q_reg[3]  ( .D(bo1[6]), .CK(clk), .RDN(n14782), .Q(
        bo2[6]) );
  DRNQHSV2 \pe2/delaycell3/q_reg[2]  ( .D(bo1[7]), .CK(clk), .RDN(n14768), .Q(
        bo2[7]) );
  DRNQHSV2 \pe2/delaycell3/q_reg[1]  ( .D(bo1[8]), .CK(clk), .RDN(n14800), .Q(
        bo2[8]) );
  DRNQHSV2 \pe3/delaycell3/q_reg[6]  ( .D(bo2[3]), .CK(clk), .RDN(n14720), .Q(
        bo3[3]) );
  DRNQHSV2 \pe3/delaycell3/q_reg[5]  ( .D(bo2[4]), .CK(clk), .RDN(n14809), .Q(
        bo3[4]) );
  DRNQHSV2 \pe3/delaycell3/q_reg[4]  ( .D(bo2[5]), .CK(clk), .RDN(n14769), .Q(
        bo3[5]) );
  DRNQHSV2 \pe3/delaycell3/q_reg[2]  ( .D(bo2[7]), .CK(clk), .RDN(n14781), .Q(
        bo3[7]) );
  DRNQHSV2 \pe3/delaycell3/q_reg[1]  ( .D(bo2[8]), .CK(clk), .RDN(n14725), .Q(
        bo3[8]) );
  DRNQHSV1 \pe5/delaycell21/q_reg[7]  ( .D(\pe5/ti_7[7] ), .CK(clk), .RDN(
        n14761), .Q(\pe5/ti_7t [7]) );
  DRNQHSV2 \pe3/delaycell3/q_reg[8]  ( .D(bo2[1]), .CK(clk), .RDN(n14811), .Q(
        bo3[1]) );
  DRNQHSV2 \pe3/delaycell3/q_reg[7]  ( .D(bo2[2]), .CK(clk), .RDN(n14814), .Q(
        bo3[2]) );
  DRNQHSV2 \pe3/delaycell3/q_reg[3]  ( .D(bo2[6]), .CK(clk), .RDN(n14817), .Q(
        bo3[6]) );
  DRNQHSV2 \pe4/delaycell3/q_reg[6]  ( .D(bo3[3]), .CK(clk), .RDN(n14779), .Q(
        bo4[3]) );
  DRNQHSV2 \pe4/delaycell3/q_reg[5]  ( .D(bo3[4]), .CK(clk), .RDN(n14765), .Q(
        bo4[4]) );
  DRNQHSV2 \pe4/delaycell3/q_reg[4]  ( .D(bo3[5]), .CK(clk), .RDN(n14775), .Q(
        bo4[5]) );
  DRNQHSV2 \pe4/delaycell3/q_reg[3]  ( .D(bo3[6]), .CK(clk), .RDN(n14794), .Q(
        bo4[6]) );
  DRNQHSV2 \pe4/delaycell3/q_reg[2]  ( .D(bo3[7]), .CK(clk), .RDN(n14782), .Q(
        bo4[7]) );
  DRNQHSV2 \pe4/delaycell3/q_reg[1]  ( .D(bo3[8]), .CK(clk), .RDN(n14808), .Q(
        bo4[8]) );
  DRNQHSV2 \pe5/delaycell3/q_reg[6]  ( .D(bo4[3]), .CK(clk), .RDN(n15094), .Q(
        bo5[3]) );
  DRNQHSV2 \pe5/delaycell3/q_reg[5]  ( .D(bo4[4]), .CK(clk), .RDN(n15173), .Q(
        bo5[4]) );
  DRNQHSV2 \pe5/delaycell3/q_reg[4]  ( .D(bo4[5]), .CK(clk), .RDN(n14812), .Q(
        bo5[5]) );
  DRNQHSV2 \pe5/delaycell3/q_reg[3]  ( .D(bo4[6]), .CK(clk), .RDN(n14803), .Q(
        bo5[6]) );
  DRNQHSV2 \pe5/delaycell3/q_reg[2]  ( .D(bo4[7]), .CK(clk), .RDN(n14748), .Q(
        bo5[7]) );
  DRNQHSV2 \pe5/delaycell3/q_reg[1]  ( .D(bo4[8]), .CK(clk), .RDN(n14813), .Q(
        bo5[8]) );
  DRNQHSV2 \pe6/delaycell3/q_reg[5]  ( .D(bo5[4]), .CK(clk), .RDN(n14751), .Q(
        bo6[4]) );
  DRNQHSV2 \pe6/delaycell3/q_reg[4]  ( .D(bo5[5]), .CK(clk), .RDN(n15094), .Q(
        bo6[5]) );
  DRNQHSV2 \pe6/delaycell3/q_reg[3]  ( .D(bo5[6]), .CK(clk), .RDN(n14810), .Q(
        bo6[6]) );
  DRNQHSV2 \pe6/delaycell3/q_reg[2]  ( .D(bo5[7]), .CK(clk), .RDN(n14768), .Q(
        bo6[7]) );
  DRNQHSV2 \pe6/delaycell3/q_reg[1]  ( .D(bo5[8]), .CK(clk), .RDN(n14757), .Q(
        bo6[8]) );
  DRNQHSV2 \pe7/delaycell3/q_reg[4]  ( .D(bo6[5]), .CK(clk), .RDN(n14787), .Q(
        bo7[5]) );
  DRNQHSV2 \pe7/delaycell3/q_reg[3]  ( .D(bo6[6]), .CK(clk), .RDN(n14788), .Q(
        bo7[6]) );
  DRNQHSV2 \pe7/delaycell3/q_reg[2]  ( .D(bo6[7]), .CK(clk), .RDN(n14710), .Q(
        bo7[7]) );
  DRNQHSV2 \pe7/delaycell3/q_reg[1]  ( .D(bo6[8]), .CK(clk), .RDN(n14745), .Q(
        bo7[8]) );
  DRNQHSV2 \pe8/delaycell3/q_reg[8]  ( .D(bo7[1]), .CK(clk), .RDN(n14814), .Q(
        bo8[1]) );
  DRNQHSV2 \pe8/delaycell3/q_reg[3]  ( .D(bo7[6]), .CK(clk), .RDN(n14792), .Q(
        bo8[6]) );
  DRNQHSV2 \pe8/delaycell3/q_reg[2]  ( .D(bo7[7]), .CK(clk), .RDN(n14746), .Q(
        bo8[7]) );
  DRNQHSV2 \pe8/delaycell3/q_reg[1]  ( .D(bo7[8]), .CK(clk), .RDN(n15173), .Q(
        bo8[8]) );
  DRNQHSV2 \pe9/delaycell3/q_reg[8]  ( .D(bo8[1]), .CK(clk), .RDN(n14765), .Q(
        bo9[1]) );
  DRNQHSV2 \pe9/delaycell3/q_reg[3]  ( .D(bo8[6]), .CK(clk), .RDN(n14726), .Q(
        bo9[6]) );
  DRNQHSV2 \pe9/delaycell3/q_reg[2]  ( .D(bo8[7]), .CK(clk), .RDN(n14752), .Q(
        bo9[7]) );
  DRNQHSV2 \pe9/delaycell3/q_reg[1]  ( .D(bo8[8]), .CK(clk), .RDN(n14807), .Q(
        bo9[8]) );
  DRNQHSV2 \pe13/delaycell3/q_reg[4]  ( .D(bo12[5]), .CK(clk), .RDN(n14800), 
        .Q(bo13[5]) );
  DRNQHSV1 \pe3/delaycell21/q_reg[7]  ( .D(n14819), .CK(clk), .RDN(n14803), 
        .Q(\pe3/ti_7t [7]) );
  DRNQHSV1 \pe11/delaycell21/q_reg[7]  ( .D(n14257), .CK(clk), .RDN(n14754), 
        .Q(\pe11/ti_7t [7]) );
  DRNQHSV1 \pe3/delaycell21/q_reg[5]  ( .D(\pe3/ti_7[5] ), .CK(clk), .RDN(
        n14725), .Q(\pe3/ti_7t [5]) );
  DRNQHSV1 \pe8/delaycell21/q_reg[7]  ( .D(n15091), .CK(clk), .RDN(n14775), 
        .Q(\pe8/ti_7t [7]) );
  DRNQHSV1 \pe14/delaycell21/q_reg[4]  ( .D(n15195), .CK(clk), .RDN(n14720), 
        .Q(\pe14/ti_7t [4]) );
  DRNQHSV1 \pe16/delaycell21/q_reg[5]  ( .D(n14835), .CK(clk), .RDN(n14775), 
        .Q(\pe16/ti_7t [5]) );
  DRNQHSV1 \pe17/delaycell21/q_reg[5]  ( .D(n14824), .CK(clk), .RDN(n14762), 
        .Q(\pe17/ti_7t [5]) );
  DRNQHSV1 \pe16/delaycell21/q_reg[7]  ( .D(\pe16/ti_7[7] ), .CK(clk), .RDN(
        rst), .Q(\pe16/ti_7t [7]) );
  DRNQHSV1 \pe20/delaycell21/q_reg[5]  ( .D(\pe20/ti_7[5] ), .CK(clk), .RDN(
        n14781), .Q(\pe20/ti_7t [5]) );
  DRNQHSV1 \pe10/delaycell21/q_reg[4]  ( .D(n15191), .CK(clk), .RDN(n14797), 
        .Q(\pe10/ti_7t [4]) );
  DRNQHSV1 \pe18/delaycell21/q_reg[5]  ( .D(\pe18/ti_7[5] ), .CK(clk), .RDN(
        n14751), .Q(\pe18/ti_7t [5]) );
  DRNQHSV1 \pe15/delaycell21/q_reg[5]  ( .D(\pe15/ti_7[5] ), .CK(clk), .RDN(
        n14772), .Q(\pe15/ti_7t [5]) );
  DRNQHSV1 \pe6/delaycell21/q_reg[5]  ( .D(\pe6/ti_7[5] ), .CK(clk), .RDN(
        n14807), .Q(\pe6/ti_7t [5]) );
  DRNQHSV2 \delaycell/q_reg  ( .D(po21), .CK(clk), .RDN(n14718), .Q(po[1]) );
  DRNQHSV1 \pe2/delaycell21/q_reg[5]  ( .D(\pe2/ti_7[5] ), .CK(clk), .RDN(
        n14744), .Q(\pe2/ti_7t [5]) );
  DRNQHSV1 \pe11/delaycell21/q_reg[5]  ( .D(\pe11/ti_7[5] ), .CK(clk), .RDN(
        n14727), .Q(\pe11/ti_7t [5]) );
  DRNQHSV1 \pe12/delaycell21/q_reg[5]  ( .D(n14701), .CK(clk), .RDN(n14781), 
        .Q(\pe12/ti_7t [5]) );
  DRNQHSV1 \pe14/delaycell21/q_reg[5]  ( .D(\pe14/ti_7[5] ), .CK(clk), .RDN(
        n14752), .Q(\pe14/ti_7t [5]) );
  DRNQHSV1 \pe17/delaycell21/q_reg[7]  ( .D(\pe17/ti_7[7] ), .CK(clk), .RDN(
        n14786), .Q(\pe17/ti_7t [7]) );
  DRNQHSV1 \pe1/delaycell21/q_reg[1]  ( .D(n10242), .CK(clk), .RDN(n14767), 
        .Q(\pe1/ti_7t [1]) );
  DRNQHSV1 \pe2/delaycell21/q_reg[1]  ( .D(\pe2/ti_7[1] ), .CK(clk), .RDN(
        n14808), .Q(\pe2/ti_7t [1]) );
  DRNQHSV1 \pe3/delaycell21/q_reg[1]  ( .D(n5949), .CK(clk), .RDN(n14783), .Q(
        \pe3/ti_7t [1]) );
  DRNQHSV1 \pe5/delaycell21/q_reg[1]  ( .D(n10346), .CK(clk), .RDN(n14729), 
        .Q(\pe5/ti_7t [1]) );
  DRNQHSV1 \pe7/delaycell21/q_reg[1]  ( .D(\pe7/ti_7[1] ), .CK(clk), .RDN(
        n14756), .Q(\pe7/ti_7t [1]) );
  DRNQHSV1 \pe11/delaycell21/q_reg[1]  ( .D(\pe11/ti_7[1] ), .CK(clk), .RDN(
        n14779), .Q(\pe11/ti_7t [1]) );
  DRNQHSV1 \pe11/delaycell21/q_reg[3]  ( .D(n14366), .CK(clk), .RDN(n14789), 
        .Q(\pe11/ti_7t [3]) );
  DRNQHSV1 \pe12/delaycell21/q_reg[1]  ( .D(\pe12/ti_7[1] ), .CK(clk), .RDN(
        n14804), .Q(\pe12/ti_7t [1]) );
  DRNQHSV1 \pe13/delaycell21/q_reg[1]  ( .D(\pe13/ti_7[1] ), .CK(clk), .RDN(
        n14806), .Q(\pe13/ti_7t [1]) );
  DRNQHSV1 \pe16/delaycell21/q_reg[1]  ( .D(\pe16/ti_7[1] ), .CK(clk), .RDN(
        n14760), .Q(\pe16/ti_7t [1]) );
  DRNQHSV1 \pe17/delaycell21/q_reg[1]  ( .D(\pe17/ti_7[1] ), .CK(clk), .RDN(
        n14801), .Q(\pe17/ti_7t [1]) );
  DRNQHSV1 \pe19/delaycell21/q_reg[1]  ( .D(\pe19/ti_7[1] ), .CK(clk), .RDN(
        n14809), .Q(\pe19/ti_7t [1]) );
  DRNQHSV1 \pe20/delaycell21/q_reg[1]  ( .D(n7465), .CK(clk), .RDN(n14768), 
        .Q(\pe20/ti_7t [1]) );
  DRNQHSV1 \pe20/delaycell21/q_reg[3]  ( .D(n11854), .CK(clk), .RDN(n14794), 
        .Q(\pe20/ti_7t [3]) );
  DRNQHSV1 \pe21/delaycell5/q_reg[4]  ( .D(n14821), .CK(clk), .RDN(n14763), 
        .Q(\pe21/pvq [4]) );
  DRNQHSV1 \pe6/delaycell5/q_reg[7]  ( .D(n15275), .CK(clk), .RDN(n14803), .Q(
        \pe6/pvq [7]) );
  DRNQHSV1 \pe6/delaycell5/q_reg[5]  ( .D(n15276), .CK(clk), .RDN(n14801), .Q(
        \pe6/pvq [5]) );
  DRNQHSV1 \pe6/delaycell5/q_reg[3]  ( .D(n15278), .CK(clk), .RDN(n14813), .Q(
        \pe6/pvq [3]) );
  DRNQHSV1 \pe8/delaycell21/q_reg[3]  ( .D(n14857), .CK(clk), .RDN(n14786), 
        .Q(\pe8/ti_7t [3]) );
  DRNQHSV2 \pe14/delaycell5/q_reg[7]  ( .D(n15240), .CK(clk), .RDN(n14717), 
        .Q(\pe14/pvq [7]) );
  DRNQHSV1 \pe14/delaycell5/q_reg[6]  ( .D(n15241), .CK(clk), .RDN(n14712), 
        .Q(\pe14/pvq [6]) );
  DRNQHSV1 \pe14/delaycell5/q_reg[5]  ( .D(n15242), .CK(clk), .RDN(n14721), 
        .Q(\pe14/pvq [5]) );
  DRNQHSV1 \pe14/delaycell5/q_reg[4]  ( .D(n15243), .CK(clk), .RDN(n14746), 
        .Q(\pe14/pvq [4]) );
  DRNQHSV1 \pe14/delaycell5/q_reg[3]  ( .D(n15244), .CK(clk), .RDN(n14718), 
        .Q(\pe14/pvq [3]) );
  DRNQHSV1 \pe2/delaycell21/q_reg[2]  ( .D(n14934), .CK(clk), .RDN(n14768), 
        .Q(\pe2/ti_7t [2]) );
  DRNQHSV1 \pe5/delaycell21/q_reg[3]  ( .D(n14916), .CK(clk), .RDN(n14785), 
        .Q(\pe5/ti_7t [3]) );
  DRNQHSV1 \pe18/delaycell21/q_reg[2]  ( .D(n11996), .CK(clk), .RDN(n14788), 
        .Q(\pe18/ti_7t [2]) );
  DRNQHSV1 \pe1/delaycell21/q_reg[2]  ( .D(n6027), .CK(clk), .RDN(n14797), .Q(
        \pe1/ti_7t [2]) );
  DRNQHSV1 \pe1/delaycell21/q_reg[4]  ( .D(n14847), .CK(clk), .RDN(n14748), 
        .Q(\pe1/ti_7t [4]) );
  DRNQHSV2 \pe2/delaycell5/q_reg[7]  ( .D(pov1[7]), .CK(clk), .RDN(n14721), 
        .Q(\pe2/pvq [7]) );
  DRNQHSV1 \pe2/delaycell5/q_reg[5]  ( .D(pov1[5]), .CK(clk), .RDN(n14760), 
        .Q(\pe2/pvq [5]) );
  DRNQHSV1 \pe2/delaycell21/q_reg[4]  ( .D(n14935), .CK(clk), .RDN(n14775), 
        .Q(\pe2/ti_7t [4]) );
  DRNQHSV2 \pe3/delaycell5/q_reg[7]  ( .D(n15290), .CK(clk), .RDN(n15094), .Q(
        \pe3/pvq [7]) );
  DRNQHSV1 \pe3/delaycell5/q_reg[5]  ( .D(n15292), .CK(clk), .RDN(n15174), .Q(
        \pe3/pvq [5]) );
  DRNQHSV1 \pe3/delaycell5/q_reg[4]  ( .D(n15070), .CK(clk), .RDN(n14754), .Q(
        \pe3/pvq [4]) );
  DRNQHSV1 \pe3/delaycell5/q_reg[3]  ( .D(n15293), .CK(clk), .RDN(n14761), .Q(
        \pe3/pvq [3]) );
  DRNQHSV1 \pe3/delaycell21/q_reg[4]  ( .D(n6326), .CK(clk), .RDN(n14727), .Q(
        \pe3/ti_7t [4]) );
  DRNQHSV2 \pe4/delaycell5/q_reg[7]  ( .D(n15285), .CK(clk), .RDN(n14717), .Q(
        \pe4/pvq [7]) );
  DRNQHSV1 \pe4/delaycell5/q_reg[5]  ( .D(n15287), .CK(clk), .RDN(n14731), .Q(
        \pe4/pvq [5]) );
  DRNQHSV1 \pe4/delaycell5/q_reg[3]  ( .D(n15288), .CK(clk), .RDN(n14766), .Q(
        \pe4/pvq [3]) );
  DRNQHSV2 \pe5/delaycell5/q_reg[7]  ( .D(n15280), .CK(clk), .RDN(n14815), .Q(
        \pe5/pvq [7]) );
  DRNQHSV1 \pe5/delaycell5/q_reg[3]  ( .D(n15283), .CK(clk), .RDN(n14789), .Q(
        \pe5/pvq [3]) );
  DRNQHSV2 \pe7/delaycell5/q_reg[7]  ( .D(n15274), .CK(clk), .RDN(n14786), .Q(
        \pe7/pvq [7]) );
  DRNQHSV1 \pe7/delaycell5/q_reg[5]  ( .D(n15198), .CK(clk), .RDN(n14801), .Q(
        \pe7/pvq [5]) );
  DRNQHSV1 \pe8/delaycell5/q_reg[7]  ( .D(n15269), .CK(clk), .RDN(n14726), .Q(
        \pe8/pvq [7]) );
  DRNQHSV1 \pe8/delaycell5/q_reg[3]  ( .D(n15271), .CK(clk), .RDN(n14794), .Q(
        \pe8/pvq [3]) );
  DRNQHSV1 \pe8/delaycell21/q_reg[4]  ( .D(n15066), .CK(clk), .RDN(n14773), 
        .Q(\pe8/ti_7t [4]) );
  DRNQHSV1 \pe9/delaycell5/q_reg[7]  ( .D(n15076), .CK(clk), .RDN(n14748), .Q(
        \pe9/pvq [7]) );
  DRNQHSV1 \pe9/delaycell21/q_reg[1]  ( .D(\pe9/ti_7[1] ), .CK(clk), .RDN(
        n14761), .Q(\pe9/ti_7t [1]) );
  DRNQHSV2 \pe10/delaycell5/q_reg[7]  ( .D(pov9[7]), .CK(clk), .RDN(n14725), 
        .Q(\pe10/pvq [7]) );
  DRNQHSV1 \pe10/delaycell5/q_reg[6]  ( .D(n6737), .CK(clk), .RDN(n14710), .Q(
        \pe10/pvq [6]) );
  DRNQHSV1 \pe10/delaycell5/q_reg[4]  ( .D(n15069), .CK(clk), .RDN(n14781), 
        .Q(\pe10/pvq [4]) );
  DRNQHSV1 \pe10/delaycell5/q_reg[3]  ( .D(n7881), .CK(clk), .RDN(n14781), .Q(
        \pe10/pvq [3]) );
  DRNQHSV1 \pe10/delaycell21/q_reg[2]  ( .D(n14940), .CK(clk), .RDN(n14765), 
        .Q(\pe10/ti_7t [2]) );
  DRNQHSV1 \pe11/delaycell5/q_reg[7]  ( .D(n15201), .CK(clk), .RDN(n14749), 
        .Q(\pe11/pvq [7]) );
  DRNQHSV1 \pe11/delaycell5/q_reg[5]  ( .D(n15262), .CK(clk), .RDN(n14757), 
        .Q(\pe11/pvq [5]) );
  DRNQHSV1 \pe11/delaycell5/q_reg[4]  ( .D(n15200), .CK(clk), .RDN(n14832), 
        .Q(\pe11/pvq [4]) );
  DRNQHSV1 \pe11/delaycell21/q_reg[4]  ( .D(n14737), .CK(clk), .RDN(n14803), 
        .Q(\pe11/ti_7t [4]) );
  DRNQHSV2 \pe12/delaycell5/q_reg[7]  ( .D(n15254), .CK(clk), .RDN(n8938), .Q(
        \pe12/pvq [7]) );
  DRNQHSV1 \pe12/delaycell5/q_reg[6]  ( .D(n15255), .CK(clk), .RDN(n14777), 
        .Q(\pe12/pvq [6]) );
  DRNQHSV1 \pe12/delaycell5/q_reg[5]  ( .D(n15256), .CK(clk), .RDN(n14792), 
        .Q(\pe12/pvq [5]) );
  DRNQHSV1 \pe12/delaycell5/q_reg[3]  ( .D(n15258), .CK(clk), .RDN(n14804), 
        .Q(\pe12/pvq [3]) );
  DRNQHSV2 \pe13/delaycell5/q_reg[7]  ( .D(n15247), .CK(clk), .RDN(n14793), 
        .Q(\pe13/pvq [7]) );
  DRNQHSV1 \pe13/delaycell5/q_reg[6]  ( .D(n15248), .CK(clk), .RDN(n14715), 
        .Q(\pe13/pvq [6]) );
  DRNQHSV1 \pe13/delaycell5/q_reg[5]  ( .D(n15249), .CK(clk), .RDN(n14729), 
        .Q(\pe13/pvq [5]) );
  DRNQHSV1 \pe13/delaycell5/q_reg[3]  ( .D(n15251), .CK(clk), .RDN(n14811), 
        .Q(\pe13/pvq [3]) );
  DRNQHSV1 \pe13/delaycell21/q_reg[2]  ( .D(n9882), .CK(clk), .RDN(n14717), 
        .Q(\pe13/ti_7t [2]) );
  DRNQHSV2 \pe15/delaycell5/q_reg[7]  ( .D(\pov14[7] ), .CK(clk), .RDN(n14761), 
        .Q(\pe15/pvq [7]) );
  DRNQHSV1 \pe15/delaycell5/q_reg[6]  ( .D(n6771), .CK(clk), .RDN(n14809), .Q(
        \pe15/pvq [6]) );
  DRNQHSV1 \pe15/delaycell5/q_reg[5]  ( .D(n15236), .CK(clk), .RDN(n14811), 
        .Q(\pe15/pvq [5]) );
  DRNQHSV1 \pe15/delaycell5/q_reg[4]  ( .D(n15237), .CK(clk), .RDN(n15173), 
        .Q(\pe15/pvq [4]) );
  DRNQHSV1 \pe15/delaycell5/q_reg[1]  ( .D(n9103), .CK(clk), .RDN(n14747), .Q(
        \pe15/pvq [1]) );
  DRNQHSV1 \pe15/delaycell21/q_reg[4]  ( .D(n7127), .CK(clk), .RDN(n14815), 
        .Q(\pe15/ti_7t [4]) );
  DRNQHSV1 \pe16/delaycell5/q_reg[7]  ( .D(n15231), .CK(clk), .RDN(n14755), 
        .Q(\pe16/pvq [7]) );
  DRNQHSV2 \pe17/delaycell5/q_reg[5]  ( .D(n15228), .CK(clk), .RDN(n14716), 
        .Q(\pe17/pvq [5]) );
  DRNQHSV1 \pe17/delaycell5/q_reg[4]  ( .D(n15185), .CK(clk), .RDN(n14784), 
        .Q(\pe17/pvq [4]) );
  DRNQHSV1 \pe17/delaycell5/q_reg[3]  ( .D(n15229), .CK(clk), .RDN(n14773), 
        .Q(\pe17/pvq [3]) );
  DRNQHSV1 \pe17/delaycell21/q_reg[2]  ( .D(n14962), .CK(clk), .RDN(n14751), 
        .Q(\pe17/ti_7t [2]) );
  DRNQHSV1 \pe18/delaycell5/q_reg[7]  ( .D(n15220), .CK(clk), .RDN(n14756), 
        .Q(\pe18/pvq [7]) );
  DRNQHSV1 \pe18/delaycell5/q_reg[5]  ( .D(n15222), .CK(clk), .RDN(n14789), 
        .Q(\pe18/pvq [5]) );
  DRNQHSV1 \pe18/delaycell5/q_reg[4]  ( .D(n12107), .CK(clk), .RDN(n14771), 
        .Q(\pe18/pvq [4]) );
  DRNQHSV1 \pe18/delaycell5/q_reg[3]  ( .D(n15223), .CK(clk), .RDN(n14759), 
        .Q(\pe18/pvq [3]) );
  DRNQHSV1 \pe18/delaycell21/q_reg[4]  ( .D(n14851), .CK(clk), .RDN(n14779), 
        .Q(\pe18/ti_7t [4]) );
  DRNQHSV2 \pe19/delaycell5/q_reg[7]  ( .D(n15214), .CK(clk), .RDN(n15173), 
        .Q(\pe19/pvq [7]) );
  DRNQHSV1 \pe19/delaycell5/q_reg[6]  ( .D(n15215), .CK(clk), .RDN(n14778), 
        .Q(\pe19/pvq [6]) );
  DRNQHSV1 \pe19/delaycell5/q_reg[3]  ( .D(n15218), .CK(clk), .RDN(n14751), 
        .Q(\pe19/pvq [3]) );
  DRNQHSV1 \pe19/delaycell5/q_reg[1]  ( .D(n14826), .CK(clk), .RDN(n14815), 
        .Q(\pe19/pvq [1]) );
  DRNQHSV2 \pe20/delaycell5/q_reg[7]  ( .D(\pov19[7] ), .CK(clk), .RDN(n14761), 
        .Q(\pe20/pvq [7]) );
  DRNQHSV1 \pe20/delaycell5/q_reg[6]  ( .D(n15073), .CK(clk), .RDN(n14775), 
        .Q(\pe20/pvq [6]) );
  DRNQHSV1 \pe20/delaycell5/q_reg[4]  ( .D(n15211), .CK(clk), .RDN(n14803), 
        .Q(\pe20/pvq [4]) );
  DRNQHSV1 \pe20/delaycell21/q_reg[4]  ( .D(n15184), .CK(clk), .RDN(n14786), 
        .Q(\pe20/ti_7t [4]) );
  DRNQHSV2 \pe21/delaycell5/q_reg[7]  ( .D(n15206), .CK(clk), .RDN(n14710), 
        .Q(\pe21/pvq [7]) );
  DRNQHSV1 \pe21/delaycell5/q_reg[5]  ( .D(n15208), .CK(clk), .RDN(n14764), 
        .Q(\pe21/pvq [5]) );
  DRNQHSV1 \pe21/delaycell5/q_reg[3]  ( .D(n10409), .CK(clk), .RDN(n14764), 
        .Q(\pe21/pvq [3]) );
  DRNQHSV1 \pe21/delaycell21/q_reg[1]  ( .D(\pe21/ti_7[1] ), .CK(clk), .RDN(
        n14783), .Q(\pe21/ti_7t [1]) );
  DRNQHSV1 \pe14/delaycell21/q_reg[2]  ( .D(n14944), .CK(clk), .RDN(n14760), 
        .Q(\pe14/ti_7t [2]) );
  DRNQHSV1 \pe19/delaycell21/q_reg[2]  ( .D(n9581), .CK(clk), .RDN(n14725), 
        .Q(\pe19/ti_7t [2]) );
  DRNQHSV1 \pe20/delaycell21/q_reg[2]  ( .D(n6026), .CK(clk), .RDN(n14794), 
        .Q(\pe20/ti_7t [2]) );
  DRNQHSV1 \pe21/delaycell21/q_reg[3]  ( .D(\pe21/ti_7[3] ), .CK(clk), .RDN(
        n14777), .Q(\pe21/ti_7t [3]) );
  DRNQHSV2 \pe2/delaycell4/q_reg  ( .D(po1), .CK(clk), .RDN(n14714), .Q(
        \pe2/pq ) );
  DRNQHSV2 \pe3/delaycell4/q_reg  ( .D(po2), .CK(clk), .RDN(n14809), .Q(
        \pe3/pq ) );
  DRNQHSV1 \pe4/delaycell21/q_reg[3]  ( .D(n15086), .CK(clk), .RDN(n14754), 
        .Q(\pe4/ti_7t [3]) );
  DRNQHSV1 \pe5/delaycell4/q_reg  ( .D(po4), .CK(clk), .RDN(n14799), .Q(
        \pe5/pq ) );
  DRNQHSV2 \pe8/delaycell4/q_reg  ( .D(po7), .CK(clk), .RDN(n14757), .Q(
        \pe8/pq ) );
  DRNQHSV2 \pe9/delaycell4/q_reg  ( .D(po8), .CK(clk), .RDN(n14789), .Q(
        \pe9/pq ) );
  DRNQHSV1 \pe9/delaycell21/q_reg[3]  ( .D(n10443), .CK(clk), .RDN(n14814), 
        .Q(\pe9/ti_7t [3]) );
  DRNQHSV2 \pe11/delaycell4/q_reg  ( .D(po10), .CK(clk), .RDN(n14776), .Q(
        \pe11/pq ) );
  DRNQHSV2 \pe13/delaycell4/q_reg  ( .D(po12), .CK(clk), .RDN(n14720), .Q(
        \pe13/pq ) );
  DRNQHSV1 \pe18/delaycell21/q_reg[3]  ( .D(n15194), .CK(clk), .RDN(n14762), 
        .Q(\pe18/ti_7t [3]) );
  DRNQHSV1 \pe20/delaycell4/q_reg  ( .D(po19), .CK(clk), .RDN(n14722), .Q(
        \pe20/pq ) );
  DRNQHSV1 \pe16/delaycell21/q_reg[3]  ( .D(\pe16/ti_7[3] ), .CK(clk), .RDN(
        n14720), .Q(\pe16/ti_7t [3]) );
  DRNQHSV1 \pe17/delaycell21/q_reg[3]  ( .D(\pe17/ti_7[3] ), .CK(clk), .RDN(
        n14768), .Q(\pe17/ti_7t [3]) );
  DRNQHSV2 \pe8/delaycell5/q_reg[1]  ( .D(n15273), .CK(clk), .RDN(n14832), .Q(
        \pe8/pvq [1]) );
  DRNQHSV1 \pe7/delaycell21/q_reg[3]  ( .D(n15183), .CK(clk), .RDN(n14817), 
        .Q(\pe7/ti_7t [3]) );
  DRNQHSV1 \pe12/delaycell21/q_reg[3]  ( .D(\pe12/ti_7[3] ), .CK(clk), .RDN(
        n14776), .Q(\pe12/ti_7t [3]) );
  DRNQHSV1 \pe8/delaycell21/q_reg[1]  ( .D(\pe8/ti_7[1] ), .CK(clk), .RDN(
        n14774), .Q(\pe8/ti_7t [1]) );
  DRNQHSV1 \pe16/delaycell21/q_reg[4]  ( .D(n14827), .CK(clk), .RDN(n14807), 
        .Q(\pe16/ti_7t [4]) );
  DRNQHSV1 \pe13/delaycell21/q_reg[3]  ( .D(n15065), .CK(clk), .RDN(n14726), 
        .Q(\pe13/ti_7t [3]) );
  DRNQHSV1 \pe19/delaycell21/q_reg[3]  ( .D(n12148), .CK(clk), .RDN(n14816), 
        .Q(\pe19/ti_7t [3]) );
  DRNQHSV1 \pe5/delaycell8/q_reg  ( .D(\pe5/ctrq ), .CK(clk), .RDN(n14804), 
        .Q(ctro5) );
  DRNQHSV2 \pe1/delaycell2/q_reg[8]  ( .D(gi[1]), .CK(clk), .RDN(rst), .Q(
        \pe1/got [1]) );
  DRNQHSV2 \pe1/delaycell2/q_reg[7]  ( .D(gi[2]), .CK(clk), .RDN(rst), .Q(
        \pe1/got [2]) );
  DRNQHSV2 \pe6/delaycell3/q_reg[6]  ( .D(bo5[3]), .CK(clk), .RDN(n14777), .Q(
        bo6[3]) );
  DRNQHSV2 \pe4/delaycell3/q_reg[8]  ( .D(bo3[1]), .CK(clk), .RDN(n14796), .Q(
        bo4[1]) );
  DRNQHSV2 \pe4/delaycell3/q_reg[7]  ( .D(bo3[2]), .CK(clk), .RDN(n14832), .Q(
        bo4[2]) );
  DRNQHSV2 \pe5/delaycell3/q_reg[8]  ( .D(bo4[1]), .CK(clk), .RDN(n14832), .Q(
        bo5[1]) );
  DRNQHSV2 \pe5/delaycell3/q_reg[7]  ( .D(bo4[2]), .CK(clk), .RDN(n14811), .Q(
        bo5[2]) );
  DRNQHSV2 \pe8/delaycell3/q_reg[5]  ( .D(bo7[4]), .CK(clk), .RDN(n15094), .Q(
        bo8[4]) );
  DRNQHSV2 \pe8/delaycell3/q_reg[4]  ( .D(bo7[5]), .CK(clk), .RDN(n14810), .Q(
        bo8[5]) );
  DRNQHSV2 \pe9/delaycell3/q_reg[5]  ( .D(bo8[4]), .CK(clk), .RDN(n14745), .Q(
        bo9[4]) );
  DRNQHSV2 \pe10/delaycell3/q_reg[8]  ( .D(bo9[1]), .CK(clk), .RDN(n14799), 
        .Q(bo10[1]) );
  DRNQHSV2 \pe10/delaycell3/q_reg[5]  ( .D(bo9[4]), .CK(clk), .RDN(n14719), 
        .Q(bo10[4]) );
  DRNQHSV2 \pe10/delaycell3/q_reg[3]  ( .D(bo9[6]), .CK(clk), .RDN(n14780), 
        .Q(bo10[6]) );
  DRNQHSV2 \pe10/delaycell3/q_reg[2]  ( .D(bo9[7]), .CK(clk), .RDN(n14809), 
        .Q(bo10[7]) );
  DRNQHSV2 \pe10/delaycell3/q_reg[1]  ( .D(bo9[8]), .CK(clk), .RDN(n14806), 
        .Q(bo10[8]) );
  DRNQHSV2 \pe11/delaycell3/q_reg[5]  ( .D(bo10[4]), .CK(clk), .RDN(n14732), 
        .Q(bo11[4]) );
  DRNQHSV2 \pe11/delaycell3/q_reg[2]  ( .D(bo10[7]), .CK(clk), .RDN(n14769), 
        .Q(bo11[7]) );
  DRNQHSV2 \pe11/delaycell3/q_reg[1]  ( .D(bo10[8]), .CK(clk), .RDN(n14782), 
        .Q(bo11[8]) );
  DRNQHSV2 \pe12/delaycell3/q_reg[5]  ( .D(bo11[4]), .CK(clk), .RDN(n14811), 
        .Q(bo12[4]) );
  DRNQHSV2 \pe12/delaycell3/q_reg[2]  ( .D(bo11[7]), .CK(clk), .RDN(n14711), 
        .Q(bo12[7]) );
  DRNQHSV2 \pe12/delaycell3/q_reg[1]  ( .D(bo11[8]), .CK(clk), .RDN(n14792), 
        .Q(bo12[8]) );
  DRNQHSV2 \pe14/delaycell3/q_reg[4]  ( .D(bo13[5]), .CK(clk), .RDN(n14746), 
        .Q(bo14[5]) );
  DRNQHSV2 \pe6/delaycell3/q_reg[8]  ( .D(bo5[1]), .CK(clk), .RDN(n14802), .Q(
        bo6[1]) );
  DRNQHSV2 \pe7/delaycell3/q_reg[6]  ( .D(bo6[3]), .CK(clk), .RDN(n14715), .Q(
        bo7[3]) );
  DRNQHSV2 \pe9/delaycell3/q_reg[4]  ( .D(bo8[5]), .CK(clk), .RDN(n14717), .Q(
        bo9[5]) );
  DRNQHSV2 \pe11/delaycell3/q_reg[8]  ( .D(bo10[1]), .CK(clk), .RDN(n14767), 
        .Q(bo11[1]) );
  DRNQHSV2 \pe11/delaycell3/q_reg[3]  ( .D(bo10[6]), .CK(clk), .RDN(n14759), 
        .Q(bo11[6]) );
  DRNQHSV2 \pe13/delaycell3/q_reg[5]  ( .D(bo12[4]), .CK(clk), .RDN(n14813), 
        .Q(bo13[4]) );
  DRNQHSV2 \pe13/delaycell3/q_reg[2]  ( .D(bo12[7]), .CK(clk), .RDN(n14710), 
        .Q(bo13[7]) );
  DRNQHSV2 \pe13/delaycell3/q_reg[1]  ( .D(bo12[8]), .CK(clk), .RDN(n15094), 
        .Q(bo13[8]) );
  DRNQHSV2 \pe15/delaycell3/q_reg[4]  ( .D(bo14[5]), .CK(clk), .RDN(n14756), 
        .Q(bo15[5]) );
  DRNQHSV2 \pe14/delaycell21/q_reg[3]  ( .D(n5969), .CK(clk), .RDN(n14744), 
        .Q(\pe14/ti_7t [3]) );
  DRNQHSV4 \pe8/delaycell5/q_reg[4]  ( .D(n14823), .CK(clk), .RDN(n14833), .Q(
        \pe8/pvq [4]) );
  DRNQHSV2 \pe5/delaycell5/q_reg[5]  ( .D(n15282), .CK(clk), .RDN(n14817), .Q(
        \pe5/pvq [5]) );
  DRNQHSV1 \pe7/delaycell21/q_reg[6]  ( .D(n15189), .CK(clk), .RDN(n14723), 
        .Q(\pe7/ti_7t [6]) );
  DRNQHSV2 \pe6/delaycell21/q_reg[1]  ( .D(n14895), .CK(clk), .RDN(n15094), 
        .Q(\pe6/ti_7t [1]) );
  DRNQHSV4 \pe7/delaycell21/q_reg[5]  ( .D(\pe7/ti_7[5] ), .CK(clk), .RDN(
        n14794), .Q(\pe7/ti_7t [5]) );
  DRNQHSV4 \pe15/delaycell4/q_reg  ( .D(po14), .CK(clk), .RDN(n14785), .Q(
        \pe15/pq ) );
  DRNQHSV1 \pe12/delaycell21/q_reg[7]  ( .D(n14959), .CK(clk), .RDN(n14717), 
        .Q(\pe12/ti_7t [7]) );
  DRNQHSV2 \pe12/delaycell24/q_reg[1]  ( .D(\pe12/poht [1]), .CK(clk), .RDN(
        n14816), .Q(poh12[1]) );
  DRNQHSV4 \pe3/delaycell8/q_reg  ( .D(n12357), .CK(clk), .RDN(n14745), .Q(
        ctro3) );
  DRNQHSV2 \pe10/delaycell21/q_reg[3]  ( .D(n14856), .CK(clk), .RDN(n14782), 
        .Q(\pe10/ti_7t [3]) );
  DRNQHSV4 \pe9/delaycell21/q_reg[4]  ( .D(n6209), .CK(clk), .RDN(n14732), .Q(
        \pe9/ti_7t [4]) );
  DRNQHSV1 \pe16/delaycell24/q_reg[6]  ( .D(\pe16/poht [6]), .CK(clk), .RDN(
        n14806), .Q(poh16[6]) );
  DRNQHSV1 \pe3/delaycell24/q_reg[2]  ( .D(\pe3/poht [2]), .CK(clk), .RDN(
        n14807), .Q(poh3[2]) );
  DRNQHSV1 \pe3/delaycell24/q_reg[4]  ( .D(\pe3/poht [4]), .CK(clk), .RDN(
        n14757), .Q(poh3[4]) );
  DRNQHSV1 \pe16/delaycell24/q_reg[7]  ( .D(\pe16/poht [7]), .CK(clk), .RDN(
        n14796), .Q(poh16[7]) );
  DRNQHSV1 \pe12/delaycell24/q_reg[5]  ( .D(\pe12/poht [5]), .CK(clk), .RDN(
        n14804), .Q(poh12[5]) );
  DRNQHSV1 \pe2/delaycell24/q_reg[1]  ( .D(\pe2/poht [1]), .CK(clk), .RDN(
        n14745), .Q(poh2[1]) );
  DRNQHSV1 \pe10/delaycell24/q_reg[7]  ( .D(\pe10/poht [7]), .CK(clk), .RDN(
        n14812), .Q(poh10[7]) );
  DRNQHSV1 \pe13/delaycell24/q_reg[2]  ( .D(\pe13/poht [2]), .CK(clk), .RDN(
        n14710), .Q(poh13[2]) );
  DRNQHSV1 \pe8/delaycell24/q_reg[6]  ( .D(\pe8/poht [6]), .CK(clk), .RDN(
        n14717), .Q(poh8[6]) );
  DRNQHSV1 \pe1/delaycell24/q_reg[7]  ( .D(\pe1/poht [7]), .CK(clk), .RDN(
        n14871), .Q(poh1[7]) );
  DRNQHSV1 \pe10/delaycell24/q_reg[1]  ( .D(\pe10/poht [1]), .CK(clk), .RDN(
        n14749), .Q(poh10[1]) );
  DRNQHSV1 \pe11/delaycell24/q_reg[5]  ( .D(\pe11/poht [5]), .CK(clk), .RDN(
        n8938), .Q(poh11[5]) );
  DRNQHSV1 \pe11/delaycell24/q_reg[1]  ( .D(\pe11/poht [1]), .CK(clk), .RDN(
        n14778), .Q(poh11[1]) );
  DRNQHSV2 \pe21/delaycell24/q_reg[2]  ( .D(\pe21/poht [2]), .CK(clk), .RDN(
        n14755), .Q(poh21[2]) );
  DRNQHSV4 \pe3/delaycell5/q_reg[1]  ( .D(n14707), .CK(clk), .RDN(n15173), .Q(
        \pe3/pvq [1]) );
  DRNQHSV1 \pe19/delaycell4/q_reg  ( .D(po18), .CK(clk), .RDN(n14717), .Q(
        \pe19/pq ) );
  DRNQHSV2 \pe9/delaycell5/q_reg[3]  ( .D(n15267), .CK(clk), .RDN(n14777), .Q(
        \pe9/pvq [3]) );
  DRNQHSV4 \pe15/delaycell8/q_reg  ( .D(n15160), .CK(clk), .RDN(n14833), .Q(
        ctro15) );
  DRNQHSV1 \pe18/delaycell24/q_reg[5]  ( .D(\pe18/poht [5]), .CK(clk), .RDN(
        n14784), .Q(poh18[5]) );
  DRNQHSV2 \pe16/delaycell24/q_reg[4]  ( .D(\pe16/poht [4]), .CK(clk), .RDN(
        n14744), .Q(poh16[4]) );
  DRNQHSV1 \pe10/delaycell24/q_reg[5]  ( .D(\pe10/poht [5]), .CK(clk), .RDN(
        n14806), .Q(poh10[5]) );
  DRNQHSV1 \pe10/delaycell24/q_reg[6]  ( .D(\pe10/poht [6]), .CK(clk), .RDN(
        n14732), .Q(poh10[6]) );
  DRNQHSV1 \pe4/delaycell24/q_reg[4]  ( .D(\pe4/poht [4]), .CK(clk), .RDN(
        n14749), .Q(poh4[4]) );
  DRNQHSV1 \pe18/delaycell24/q_reg[3]  ( .D(\pe18/poht [3]), .CK(clk), .RDN(
        n14813), .Q(poh18[3]) );
  DRNQHSV1 \pe3/delaycell24/q_reg[5]  ( .D(\pe3/poht [5]), .CK(clk), .RDN(
        n14749), .Q(poh3[5]) );
  DRNQHSV1 \pe9/delaycell21/q_reg[7]  ( .D(n7875), .CK(clk), .RDN(rst), .Q(
        \pe9/ti_7t [7]) );
  DSNHSV4 \pe10/delaycell5/q_reg[1]  ( .D(n14927), .CK(clk), .SDN(n14779), .Q(
        n14929), .QN(\pe10/pvq [1]) );
  DSNHSV4 \pe9/delaycell7/q_reg  ( .D(n15082), .CK(clk), .SDN(n14717), .Q(
        n14926), .QN(\pe9/ctrq ) );
  DSNHSV4 \pe9/delaycell5/q_reg[1]  ( .D(n14925), .CK(clk), .SDN(n14871), .QN(
        \pe9/pvq [1]) );
  DRNQHSV1 \pe8/delaycell24/q_reg[2]  ( .D(\pe8/poht [2]), .CK(clk), .RDN(rst), 
        .Q(poh8[2]) );
  DSNHSV4 \pe8/delaycell20/q_reg  ( .D(\pe8/ti_1t ), .CK(clk), .SDN(n14776), 
        .Q(n15127), .QN(\pe8/ti_1 ) );
  DRNQHSV1 \pe18/delaycell24/q_reg[4]  ( .D(\pe18/poht [4]), .CK(clk), .RDN(
        rst), .Q(poh18[4]) );
  DRNQHSV1 \pe18/delaycell24/q_reg[1]  ( .D(\pe18/poht [1]), .CK(clk), .RDN(
        n14798), .Q(poh18[1]) );
  DSNHSV4 \pe11/delaycell19/q_reg[1]  ( .D(n14980), .CK(clk), .SDN(n14762), 
        .Q(n14854), .QN(\pe11/bq[8] ) );
  DSNHSV4 \pe11/delaycell21/q_reg[2]  ( .D(n14924), .CK(clk), .SDN(n14792), 
        .QN(\pe11/ti_7t [2]) );
  DSNHSV4 \pe11/delaycell1/q_reg[2]  ( .D(n14923), .CK(clk), .SDN(n14746), .Q(
        n14836), .QN(\pe11/aot [7]) );
  DSNHSV4 \pe11/delaycell1/q_reg[1]  ( .D(n14921), .CK(clk), .SDN(n14792), .Q(
        n14922), .QN(\pe11/aot [8]) );
  DSNHSV4 \pe4/delaycell1/q_reg[2]  ( .D(n14919), .CK(clk), .SDN(n14812), .Q(
        n14920), .QN(\pe4/aot [7]) );
  DSNHSV4 \pe8/delaycell2/q_reg[3]  ( .D(n14918), .CK(clk), .SDN(rst), .Q(
        n15134), .QN(\pe8/got [6]) );
  DRNQHSV1 \pe21/delaycell4/q_reg  ( .D(po20), .CK(clk), .RDN(n14807), .Q(
        \pe21/pq ) );
  DSNHSV4 \pe20/delaycell19/q_reg[1]  ( .D(n8916), .CK(clk), .SDN(n14747), .Q(
        n14954), .QN(\pe20/bq[8] ) );
  DRNQHSV2 \pe8/delaycell24/q_reg[1]  ( .D(\pe8/poht [1]), .CK(clk), .RDN(
        n14771), .Q(poh8[1]) );
  DSNHSV4 \pe8/delaycell21/q_reg[2]  ( .D(n15079), .CK(clk), .SDN(n14768), 
        .QN(\pe8/ti_7t [2]) );
  DSNHSV4 \pe8/delaycell1/q_reg[1]  ( .D(n14917), .CK(clk), .SDN(rst), .Q(
        n14838), .QN(\pe8/aot [8]) );
  DSNHSV4 \pe8/delaycell19/q_reg[2]  ( .D(n15129), .CK(clk), .SDN(n14802), .Q(
        n15132), .QN(\pe8/bq[7] ) );
  DSNHSV4 \pe10/delaycell20/q_reg  ( .D(\pe10/ti_1t ), .CK(clk), .SDN(n14802), 
        .Q(n15139), .QN(\pe10/ti_1 ) );
  DSNHSV1 \pe10/delaycell23/q_reg[3]  ( .D(n15097), .CK(clk), .SDN(n14775), 
        .Q(n14913) );
  DSNHSV4 \pe10/delaycell2/q_reg[3]  ( .D(n14912), .CK(clk), .SDN(n14714), .Q(
        n15097), .QN(\pe10/got [6]) );
  DSNHSV4 \pe10/delaycell2/q_reg[1]  ( .D(n14911), .CK(clk), .SDN(n14752), .Q(
        n15098), .QN(\pe10/got [8]) );
  DSNHSV4 \pe10/delaycell2/q_reg[2]  ( .D(n14910), .CK(clk), .SDN(n14717), .Q(
        n15140), .QN(\pe10/got [7]) );
  DRNQHSV1 \pe20/delaycell24/q_reg[1]  ( .D(\pe20/poht [1]), .CK(clk), .RDN(
        n14723), .Q(poh20[1]) );
  DSNHSV4 \pe21/delaycell5/q_reg[1]  ( .D(n14909), .CK(clk), .SDN(n14769), 
        .QN(\pe21/pvq [1]) );
  DSNHSV4 \pe20/delaycell20/q_reg  ( .D(\pe20/ti_1t ), .CK(clk), .SDN(n8938), 
        .Q(n14839), .QN(\pe20/ti_1 ) );
  DSNHSV4 \pe20/delaycell1/q_reg[1]  ( .D(n14907), .CK(clk), .SDN(n14752), .Q(
        n14908), .QN(\pe20/aot [8]) );
  DSNHSV4 \pe10/delaycell1/q_reg[3]  ( .D(n14905), .CK(clk), .SDN(n14785), .Q(
        n14906), .QN(\pe10/aot [6]) );
  DSNHSV4 \pe4/delaycell8/q_reg  ( .D(n14904), .CK(clk), .SDN(n14816), .Q(
        n14955), .QN(ctro4) );
  DSNHSV4 \pe4/delaycell7/q_reg  ( .D(n10789), .CK(clk), .SDN(n14782), .Q(
        n14904), .QN(\pe4/ctrq ) );
  DSNHSV4 \pe9/delaycell19/q_reg[1]  ( .D(n15133), .CK(clk), .SDN(n14764), .Q(
        n15093), .QN(\pe9/bq[8] ) );
  DSNHSV4 \pe11/delaycell2/q_reg[3]  ( .D(n14913), .CK(clk), .SDN(n14760), .Q(
        n15146), .QN(\pe11/got [6]) );
  DSNHSV4 \pe9/delaycell8/q_reg  ( .D(n14926), .CK(clk), .SDN(n14797), .Q(
        n15074), .QN(ctro9) );
  DSNHSV4 \pe15/delaycell1/q_reg[1]  ( .D(n14903), .CK(clk), .SDN(n14774), 
        .QN(\pe15/aot [8]) );
  DRNQHSV1 \pe21/delaycell24/q_reg[6]  ( .D(\pe21/poht [6]), .CK(clk), .RDN(
        n14763), .Q(poh21[6]) );
  DSNHSV4 \pe5/delaycell5/q_reg[4]  ( .D(n14902), .CK(clk), .SDN(n14767), .QN(
        \pe5/pvq [4]) );
  DSNHSV4 \pe4/delaycell19/q_reg[1]  ( .D(n15103), .CK(clk), .SDN(n14716), .Q(
        n14875), .QN(\pe4/bq[8] ) );
  DSNHSV4 \pe5/delaycell5/q_reg[1]  ( .D(n14901), .CK(clk), .SDN(n14807), .QN(
        \pe5/pvq [1]) );
  DSNHSV4 \pe4/delaycell5/q_reg[1]  ( .D(n14900), .CK(clk), .SDN(n14719), .QN(
        \pe4/pvq [1]) );
  DSNHSV4 \pe4/delaycell2/q_reg[1]  ( .D(n14928), .CK(clk), .SDN(n14747), .Q(
        n15083), .QN(\pe4/got [8]) );
  DSNHSV4 \pe4/delaycell1/q_reg[1]  ( .D(n14899), .CK(clk), .SDN(n14797), .Q(
        n14842), .QN(\pe4/aot [8]) );
  DSNHSV4 \pe4/delaycell1/q_reg[4]  ( .D(n14897), .CK(clk), .SDN(n14754), .Q(
        n14898), .QN(\pe4/aot [5]) );
  DRNQHSV1 \pe21/delaycell24/q_reg[1]  ( .D(\pe21/poht [1]), .CK(clk), .RDN(
        n14802), .Q(poh21[1]) );
  DRNQHSV1 \pe21/delaycell24/q_reg[4]  ( .D(\pe21/poht [4]), .CK(clk), .RDN(
        n14774), .Q(poh21[4]) );
  DRNQHSV1 \pe3/delaycell24/q_reg[1]  ( .D(\pe3/poht [1]), .CK(clk), .RDN(
        n14776), .Q(poh3[1]) );
  DRNQHSV2 \pe18/delaycell24/q_reg[2]  ( .D(\pe18/poht [2]), .CK(clk), .RDN(
        n14796), .Q(poh18[2]) );
  DRNQHSV2 \pe17/delaycell5/q_reg[1]  ( .D(n14736), .CK(clk), .RDN(rst), .Q(
        \pe17/pvq [1]) );
  DRNQHSV1 \pe16/delaycell24/q_reg[3]  ( .D(\pe16/poht [3]), .CK(clk), .RDN(
        n14711), .Q(poh16[3]) );
  DSNHSV4 \pe3/delaycell1/q_reg[1]  ( .D(n14888), .CK(clk), .SDN(n14717), .QN(
        \pe3/aot [8]) );
  DSNHSV4 \pe3/delaycell19/q_reg[1]  ( .D(n15054), .CK(clk), .SDN(n14762), .Q(
        n14834), .QN(\pe3/bq[8] ) );
  DSNHSV4 \pe3/delaycell20/q_reg  ( .D(\pe3/ti_1t ), .CK(clk), .SDN(n15173), 
        .Q(n8924), .QN(\pe3/ti_1 ) );
  DSNHSV4 \pe7/delaycell5/q_reg[3]  ( .D(n14887), .CK(clk), .SDN(n14761), .QN(
        \pe7/pvq [3]) );
  DRNQHSV1 \pe7/delaycell4/q_reg  ( .D(po6), .CK(clk), .RDN(n14763), .Q(
        \pe7/pq ) );
  DSNHSV4 \pe6/delaycell1/q_reg[1]  ( .D(n14884), .CK(clk), .SDN(n14788), .Q(
        n14885), .QN(\pe6/aot [8]) );
  DRNQHSV2 \pe6/delaycell24/q_reg[3]  ( .D(\pe6/poht [3]), .CK(clk), .RDN(
        n14771), .Q(poh6[3]) );
  DSNHSV4 \pe6/delaycell19/q_reg[1]  ( .D(n15114), .CK(clk), .SDN(n14715), .Q(
        n14863), .QN(\pe6/bq[8] ) );
  DSNHSV4 \pe6/delaycell1/q_reg[3]  ( .D(n14883), .CK(clk), .SDN(n15173), .Q(
        n14848), .QN(\pe6/aot [6]) );
  DSNHSV4 \pe6/delaycell2/q_reg[1]  ( .D(n14882), .CK(clk), .SDN(n14783), .Q(
        n15095), .QN(\pe6/got [8]) );
  DSNHSV4 \pe6/delaycell19/q_reg[3]  ( .D(n15115), .CK(clk), .SDN(rst), .Q(
        n14845), .QN(\pe6/bq[6] ) );
  DSNHSV4 \pe7/delaycell5/q_reg[1]  ( .D(n14734), .CK(clk), .SDN(n14749), .QN(
        \pe7/pvq [1]) );
  DSNHSV4 \pe6/delaycell5/q_reg[1]  ( .D(n14881), .CK(clk), .SDN(n14789), .QN(
        \pe6/pvq [1]) );
  DSNHSV4 \pe6/delaycell7/q_reg  ( .D(n10307), .CK(clk), .SDN(rst), .Q(n14869), 
        .QN(\pe6/ctrq ) );
  DSNHSV4 \pe6/delaycell21/q_reg[2]  ( .D(n14880), .CK(clk), .SDN(n14749), 
        .QN(\pe6/ti_7t [2]) );
  DRNQHSV2 \pe6/delaycell4/q_reg  ( .D(po5), .CK(clk), .RDN(n14776), .Q(
        \pe6/pq ) );
  DSNHSV4 \pe5/delaycell1/q_reg[1]  ( .D(n14878), .CK(clk), .SDN(n14716), .Q(
        n14879), .QN(\pe5/aot [8]) );
  DSNHSV4 \pe6/delaycell21/q_reg[3]  ( .D(n14877), .CK(clk), .SDN(n14811), 
        .QN(\pe6/ti_7t [3]) );
  DRNQHSV4 \pe8/delaycell8/q_reg  ( .D(n14758), .CK(clk), .RDN(n14752), .Q(
        ctro8) );
  DRNQHSV4 \pe20/delaycell8/q_reg  ( .D(n12362), .CK(clk), .RDN(n14793), .Q(
        ctro20) );
  DRNQHSV2 \pe19/delaycell22/q_reg[2]  ( .D(n14945), .CK(clk), .RDN(n14796), 
        .Q(ao19[7]) );
  DRNQHSV2 \pe17/delaycell21/q_reg[6]  ( .D(n7039), .CK(clk), .RDN(n14781), 
        .Q(\pe17/ti_7t [6]) );
  DRNQHSV1 \pe17/delaycell22/q_reg[1]  ( .D(n14949), .CK(clk), .RDN(n14810), 
        .Q(ao17[8]) );
  DRNQHSV1 \pe16/delaycell21/q_reg[6]  ( .D(n15186), .CK(clk), .RDN(n14833), 
        .Q(\pe16/ti_7t [6]) );
  DRNQHSV2 \pe8/delaycell3/q_reg[7]  ( .D(bo7[2]), .CK(clk), .RDN(n14813), .Q(
        bo8[2]) );
  DRNQHSV2 \pe6/delaycell24/q_reg[5]  ( .D(\pe6/poht [5]), .CK(clk), .RDN(
        n14807), .Q(poh6[5]) );
  DRNQHSV4 \pe1/delaycell3/q_reg[7]  ( .D(bi[2]), .CK(clk), .RDN(n14809), .Q(
        bo1[2]) );
  DRNQHSV4 \pe1/delaycell3/q_reg[3]  ( .D(bi[6]), .CK(clk), .RDN(n14772), .Q(
        bo1[6]) );
  DRNQHSV2 \pe14/delaycell21/q_reg[1]  ( .D(n14964), .CK(clk), .RDN(n14769), 
        .Q(\pe14/ti_7t [1]) );
  DRNQHSV4 \pe1/delaycell3/q_reg[1]  ( .D(bi[8]), .CK(clk), .RDN(n14813), .Q(
        bo1[8]) );
  DRNQHSV1 \pe11/delaycell24/q_reg[2]  ( .D(\pe11/poht [2]), .CK(clk), .RDN(
        n14712), .Q(poh11[2]) );
  DRNQHSV1 \pe18/delaycell24/q_reg[7]  ( .D(\pe18/poht [7]), .CK(clk), .RDN(
        n14771), .Q(poh18[7]) );
  DRNQHSV4 \pe5/delaycell21/q_reg[2]  ( .D(n14952), .CK(clk), .RDN(n14752), 
        .Q(\pe5/ti_7t [2]) );
  DRNQHSV1 \pe17/delaycell24/q_reg[2]  ( .D(\pe17/poht [2]), .CK(clk), .RDN(
        n14756), .Q(poh17[2]) );
  DRNQHSV1 \pe3/delaycell6/q_reg[7]  ( .D(poh2[7]), .CK(clk), .RDN(n14730), 
        .Q(\pe3/phq [7]) );
  DRNQHSV1 \pe3/delaycell6/q_reg[6]  ( .D(poh2[6]), .CK(clk), .RDN(n14800), 
        .Q(\pe3/phq [6]) );
  DRNQHSV4 \pe1/delaycell3/q_reg[6]  ( .D(bi[3]), .CK(clk), .RDN(n14832), .Q(
        bo1[3]) );
  DRNQHSV4 \pe1/delaycell3/q_reg[8]  ( .D(bi[1]), .CK(clk), .RDN(rst), .Q(
        bo1[1]) );
  DRNQHSV4 \pe1/delaycell3/q_reg[5]  ( .D(bi[4]), .CK(clk), .RDN(rst), .Q(
        bo1[4]) );
  DRNQHSV4 \pe1/delaycell3/q_reg[4]  ( .D(bi[5]), .CK(clk), .RDN(rst), .Q(
        bo1[5]) );
  DRNQHSV4 \pe1/delaycell7/q_reg  ( .D(ctr), .CK(clk), .RDN(n14719), .Q(
        \pe1/ctrq ) );
  DRNQHSV1 \pe4/delaycell21/q_reg[1]  ( .D(\pe4/ti_7[1] ), .CK(clk), .RDN(
        n14761), .Q(\pe4/ti_7t [1]) );
  DRNQHSV2 \pe19/delaycell5/q_reg[5]  ( .D(n15216), .CK(clk), .RDN(n14774), 
        .Q(\pe19/pvq [5]) );
  DRNQHSV4 \pe6/delaycell8/q_reg  ( .D(n14870), .CK(clk), .RDN(n14779), .Q(
        ctro6) );
  DRNQHSV4 \pe12/delaycell8/q_reg  ( .D(n14938), .CK(clk), .RDN(n14771), .Q(
        ctro12) );
  DRNQHSV1 \pe1/delaycell24/q_reg[4]  ( .D(\pe1/poht [4]), .CK(clk), .RDN(
        n14779), .Q(poh1[4]) );
  DRNQHSV1 \pe1/delaycell24/q_reg[5]  ( .D(\pe1/poht [5]), .CK(clk), .RDN(
        n14769), .Q(poh1[5]) );
  DRNQHSV4 \pe1/delaycell19/q_reg[8]  ( .D(n15046), .CK(clk), .RDN(n14764), 
        .Q(\pe1/bq[1] ) );
  DRNQHSV2 \pe16/delaycell21/q_reg[2]  ( .D(n7528), .CK(clk), .RDN(n14755), 
        .Q(\pe16/ti_7t [2]) );
  DSNHSV1 \pe5/delaycell22/q_reg[1]  ( .D(n14879), .CK(clk), .SDN(n14730), .Q(
        n14884) );
  DRNQHSV2 \pe10/delaycell21/q_reg[6]  ( .D(\pe10/ti_7[6] ), .CK(clk), .RDN(
        n14785), .Q(\pe10/ti_7t [6]) );
  DRNQHSV4 \pe6/delaycell21/q_reg[7]  ( .D(n14179), .CK(clk), .RDN(rst), .Q(
        \pe6/ti_7t [7]) );
  DRNQHSV2 \pe15/delaycell21/q_reg[3]  ( .D(\pe15/ti_7[3] ), .CK(clk), .RDN(
        n14712), .Q(\pe15/ti_7t [3]) );
  DRNQHSV2 \pe16/delaycell5/q_reg[1]  ( .D(n15235), .CK(clk), .RDN(n14714), 
        .Q(\pe16/pvq [1]) );
  DRNQHSV4 \pe10/delaycell8/q_reg  ( .D(n14554), .CK(clk), .RDN(n14712), .Q(
        ctro10) );
  DRNQHSV4 \pe11/delaycell5/q_reg[1]  ( .D(n15264), .CK(clk), .RDN(n14757), 
        .Q(\pe11/pvq [1]) );
  DRNQHSV4 \pe6/delaycell21/q_reg[4]  ( .D(n15077), .CK(clk), .RDN(n14813), 
        .Q(\pe6/ti_7t [4]) );
  DRNQHSV2 \pe18/delaycell5/q_reg[1]  ( .D(n15225), .CK(clk), .RDN(n8938), .Q(
        \pe18/pvq [1]) );
  DRNQHSV1 \pe17/delaycell5/q_reg[7]  ( .D(n15226), .CK(clk), .RDN(n14813), 
        .Q(\pe17/pvq [7]) );
  DRNQHSV1 \pe10/delaycell21/q_reg[5]  ( .D(\pe10/ti_7[5] ), .CK(clk), .RDN(
        n14809), .Q(\pe10/ti_7t [5]) );
  DRNQHSV1 \pe9/delaycell21/q_reg[6]  ( .D(n15068), .CK(clk), .RDN(n15174), 
        .Q(\pe9/ti_7t [6]) );
  DRNQHSV1 \pe7/delaycell21/q_reg[4]  ( .D(n15081), .CK(clk), .RDN(n14711), 
        .Q(\pe7/ti_7t [4]) );
  DRNQHSV1 \pe11/delaycell24/q_reg[3]  ( .D(\pe11/poht [3]), .CK(clk), .RDN(
        n14804), .Q(poh11[3]) );
  DRNQHSV1 \pe12/delaycell5/q_reg[4]  ( .D(n15257), .CK(clk), .RDN(n14710), 
        .Q(\pe12/pvq [4]) );
  DRNQHSV1 \pe12/delaycell4/q_reg  ( .D(po11), .CK(clk), .RDN(n14803), .Q(
        \pe12/pq ) );
  DRNQHSV1 \pe9/delaycell24/q_reg[7]  ( .D(\pe9/poht [7]), .CK(clk), .RDN(
        n14757), .Q(poh9[7]) );
  DSNHSV2 \pe7/delaycell5/q_reg[2]  ( .D(n15071), .CK(clk), .SDN(n14754), .QN(
        \pe7/pvq [2]) );
  DRNQHSV1 \pe9/delaycell24/q_reg[1]  ( .D(\pe9/poht [1]), .CK(clk), .RDN(
        n15094), .Q(poh9[1]) );
  DRNQHSV1 \pe10/delaycell4/q_reg  ( .D(po9), .CK(clk), .RDN(n14746), .Q(
        \pe10/pq ) );
  DRNQHSV1 \pe5/delaycell21/q_reg[5]  ( .D(n14846), .CK(clk), .RDN(n14726), 
        .Q(\pe5/ti_7t [5]) );
  DRNQHSV1 \pe7/delaycell21/q_reg[2]  ( .D(n14860), .CK(clk), .RDN(n14761), 
        .Q(\pe7/ti_7t [2]) );
  DRNQHSV1 \pe7/delaycell24/q_reg[2]  ( .D(\pe7/poht [2]), .CK(clk), .RDN(
        n14794), .Q(poh7[2]) );
  DRNQHSV1 \pe11/delaycell24/q_reg[6]  ( .D(\pe11/poht [6]), .CK(clk), .RDN(
        n14745), .Q(poh11[6]) );
  DRNQHSV1 \pe18/delaycell21/q_reg[1]  ( .D(\pe18/ti_7[1] ), .CK(clk), .RDN(
        n14777), .Q(\pe18/ti_7t [1]) );
  DRNQHSV1 \pe21/delaycell24/q_reg[3]  ( .D(\pe21/poht [3]), .CK(clk), .RDN(
        n14774), .Q(poh21[3]) );
  DRNQHSV4 \pe7/delaycell3/q_reg[5]  ( .D(bo6[4]), .CK(clk), .RDN(n14806), .Q(
        bo7[4]) );
  DRNQHSV1 \pe8/delaycell21/q_reg[6]  ( .D(n15182), .CK(clk), .RDN(n14806), 
        .Q(\pe8/ti_7t [6]) );
  DRNQHSV4 \pe18/delaycell8/q_reg  ( .D(n14564), .CK(clk), .RDN(n14816), .Q(
        ctro18) );
  DRNQHSV1 \pe13/delaycell5/q_reg[4]  ( .D(n15250), .CK(clk), .RDN(n14752), 
        .Q(\pe13/pvq [4]) );
  DRNQHSV1 \pe12/delaycell3/q_reg[8]  ( .D(bo11[1]), .CK(clk), .RDN(n14722), 
        .Q(bo12[1]) );
  DRNQHSV4 \pe15/delaycell5/q_reg[3]  ( .D(n15238), .CK(clk), .RDN(n14781), 
        .Q(\pe15/pvq [3]) );
  DRNQHSV1 \pe11/delaycell24/q_reg[4]  ( .D(\pe11/poht [4]), .CK(clk), .RDN(
        n14760), .Q(poh11[4]) );
  DSNHSV2 \pe7/delaycell5/q_reg[6]  ( .D(n14886), .CK(clk), .SDN(rst), .QN(
        \pe7/pvq [6]) );
  DRNQHSV1 \pe15/delaycell5/q_reg[2]  ( .D(n15239), .CK(clk), .RDN(n14747), 
        .Q(\pe15/pvq [2]) );
  DRNQHSV1 \pe4/delaycell21/q_reg[5]  ( .D(n14850), .CK(clk), .RDN(n14774), 
        .Q(\pe4/ti_7t [5]) );
  DRNQHSV1 \pe4/delaycell4/q_reg  ( .D(po3), .CK(clk), .RDN(n14717), .Q(
        \pe4/pq ) );
  DRNQHSV1 \pe21/delaycell24/q_reg[5]  ( .D(\pe21/poht [5]), .CK(clk), .RDN(
        n14731), .Q(poh21[5]) );
  DRNQHSV2 \pe4/delaycell24/q_reg[5]  ( .D(\pe4/poht [5]), .CK(clk), .RDN(
        n14774), .Q(poh4[5]) );
  DRNQHSV2 \pe4/delaycell24/q_reg[6]  ( .D(\pe4/poht [6]), .CK(clk), .RDN(
        n14802), .Q(poh4[6]) );
  DRNQHSV1 \pe4/delaycell24/q_reg[2]  ( .D(\pe4/poht [2]), .CK(clk), .RDN(
        n14757), .Q(poh4[2]) );
  DRNQHSV2 \pe15/delaycell23/q_reg[3]  ( .D(\pe15/got [6]), .CK(clk), .RDN(
        n14728), .Q(go15[6]) );
  DRNQHSV1 \pe15/delaycell21/q_reg[7]  ( .D(n14853), .CK(clk), .RDN(n14728), 
        .Q(\pe15/ti_7t [7]) );
  DRNQHSV1 \pe6/delaycell21/q_reg[6]  ( .D(n15089), .CK(clk), .RDN(n14774), 
        .Q(\pe6/ti_7t [6]) );
  DSNHSV1 \pe10/delaycell22/q_reg[3]  ( .D(n14906), .CK(clk), .SDN(n14812), 
        .QN(ao10[6]) );
  DSNHSV1 \pe20/delaycell22/q_reg[1]  ( .D(n14908), .CK(clk), .SDN(n14801), 
        .QN(ao20[8]) );
  DSNHSV1 \pe11/delaycell22/q_reg[1]  ( .D(n14922), .CK(clk), .SDN(rst), .QN(
        ao11[8]) );
  DSNHSV1 \pe4/delaycell22/q_reg[4]  ( .D(n14898), .CK(clk), .SDN(n14776), 
        .QN(ao4[5]) );
  DSNHSV1 \pe4/delaycell22/q_reg[2]  ( .D(n14920), .CK(clk), .SDN(n14785), 
        .QN(ao4[7]) );
  DSNHSV1 \pe6/delaycell22/q_reg[1]  ( .D(n14885), .CK(clk), .SDN(n14748), 
        .QN(ao6[8]) );
  DSNHSV1 \pe8/delaycell23/q_reg[3]  ( .D(n15134), .CK(clk), .SDN(n14711), 
        .QN(go8[6]) );
  DSNHSV1 \pe11/delaycell23/q_reg[3]  ( .D(n15146), .CK(clk), .SDN(n14732), 
        .QN(go11[6]) );
  DSNHSV1 \pe4/delaycell23/q_reg[1]  ( .D(n15083), .CK(clk), .SDN(n14756), 
        .QN(go4[8]) );
  DRNQHSV1 \pe19/delaycell23/q_reg[3]  ( .D(\pe19/got [6]), .CK(clk), .RDN(
        n14756), .Q(go19[6]) );
  DSNHSV1 \pe19/delaycell22/q_reg[4]  ( .D(n15099), .CK(clk), .SDN(n15174), 
        .QN(ao19[5]) );
  DSNHSV1 \pe17/delaycell21/q_reg[4]  ( .D(n15167), .CK(clk), .SDN(rst), .Q(
        n15080), .QN(\pe17/ti_7t [4]) );
  DRNQHSV1 \pe8/delaycell21/q_reg[5]  ( .D(n14893), .CK(clk), .RDN(rst), .Q(
        \pe8/ti_7t [5]) );
  DRNQHSV4 \pe2/delaycell2/q_reg[3]  ( .D(go1[6]), .CK(clk), .RDN(n14811), .Q(
        n14822) );
  DRNQHSV1 \pe10/delaycell3/q_reg[4]  ( .D(bo9[5]), .CK(clk), .RDN(n14784), 
        .Q(bo10[5]) );
  DRSNHSV1 \pe10/delaycell21/q_reg[1]  ( .D(n6033), .CK(clk), .SDN(1'b1), 
        .RDN(n14807), .Q(\pe10/ti_7t [1]), .QN(n15096) );
  DRNQHSV1 \pe16/delaycell5/q_reg[3]  ( .D(n15233), .CK(clk), .RDN(n14796), 
        .Q(\pe16/pvq [3]) );
  DRNQHSV1 \pe18/delaycell24/q_reg[6]  ( .D(\pe18/poht [6]), .CK(clk), .RDN(
        n14798), .Q(poh18[6]) );
  DRNQHSV2 \pe16/delaycell23/q_reg[6]  ( .D(\pe16/got [3]), .CK(clk), .RDN(
        n14710), .Q(go16[3]) );
  DRNQHSV1 \pe4/delaycell24/q_reg[1]  ( .D(\pe4/poht [1]), .CK(clk), .RDN(
        n14754), .Q(poh4[1]) );
  DRNQHSV1 \pe19/delaycell21/q_reg[4]  ( .D(n11713), .CK(clk), .RDN(n14810), 
        .Q(\pe19/ti_7t [4]) );
  DRNQHSV1 \pe12/delaycell5/q_reg[1]  ( .D(n15260), .CK(clk), .RDN(n14745), 
        .Q(\pe12/pvq [1]) );
  DRNQHSV1 \pe15/delaycell24/q_reg[2]  ( .D(\pe15/poht [2]), .CK(clk), .RDN(
        n14762), .Q(poh15[2]) );
  DRNQHSV1 \pe12/delaycell21/q_reg[2]  ( .D(n14255), .CK(clk), .RDN(n14793), 
        .Q(\pe12/ti_7t [2]) );
  DRNQHSV1 \pe20/delaycell23/q_reg[2]  ( .D(n14890), .CK(clk), .RDN(n14759), 
        .Q(go20[7]) );
  DRNQHSV2 \pe14/delaycell3/q_reg[1]  ( .D(bo13[8]), .CK(clk), .RDN(n14817), 
        .Q(bo14[8]) );
  DRNQHSV1 \pe17/delaycell24/q_reg[6]  ( .D(\pe17/poht [6]), .CK(clk), .RDN(
        n14755), .Q(poh17[6]) );
  DRNQHSV1 \pe14/delaycell8/q_reg  ( .D(n14742), .CK(clk), .RDN(n14802), .Q(
        ctro14) );
  DRNQHSV2 \pe3/delaycell21/q_reg[3]  ( .D(n14820), .CK(clk), .RDN(n14747), 
        .Q(\pe3/ti_7t [3]) );
  DRNQHSV4 \pe11/delaycell8/q_reg  ( .D(n14791), .CK(clk), .RDN(n14792), .Q(
        ctro11) );
  DRNQHSV4 \pe2/delaycell8/q_reg  ( .D(n8946), .CK(clk), .RDN(n14772), .Q(
        ctro2) );
  DRNQHSV4 \pe21/delaycell8/q_reg  ( .D(n6014), .CK(clk), .RDN(n14717), .Q(
        ctro21) );
  DRNQHSV2 \pe15/delaycell24/q_reg[4]  ( .D(\pe15/poht [4]), .CK(clk), .RDN(
        n14749), .Q(poh15[4]) );
  DRNQHSV2 \pe15/delaycell24/q_reg[5]  ( .D(\pe15/poht [5]), .CK(clk), .RDN(
        n14813), .Q(poh15[5]) );
  DRNQHSV2 \pe10/delaycell6/q_reg[6]  ( .D(poh9[6]), .CK(clk), .RDN(n14715), 
        .Q(\pe10/phq [6]) );
  DRNQHSV1 \pe11/delaycell5/q_reg[3]  ( .D(n15075), .CK(clk), .RDN(n14713), 
        .Q(\pe11/pvq [3]) );
  DRNQHSV2 \pe4/delaycell21/q_reg[6]  ( .D(n12602), .CK(clk), .RDN(n14769), 
        .Q(\pe4/ti_7t [6]) );
  DRNQHSV1 \pe13/delaycell21/q_reg[5]  ( .D(n13603), .CK(clk), .RDN(n14792), 
        .Q(\pe13/ti_7t [5]) );
  DRNQHSV2 \pe19/delaycell5/q_reg[4]  ( .D(n15217), .CK(clk), .RDN(n14816), 
        .Q(\pe19/pvq [4]) );
  DRNQHSV1 \pe17/delaycell22/q_reg[3]  ( .D(n5973), .CK(clk), .RDN(n14747), 
        .Q(ao17[6]) );
  DRNQHSV1 \pe16/delaycell4/q_reg  ( .D(po15), .CK(clk), .RDN(n14797), .Q(
        \pe16/pq ) );
  DRNQHSV1 \pe17/delaycell24/q_reg[7]  ( .D(\pe17/poht [7]), .CK(clk), .RDN(
        n14767), .Q(poh17[7]) );
  DRNQHSV2 \pe20/delaycell24/q_reg[2]  ( .D(\pe20/poht [2]), .CK(clk), .RDN(
        n14755), .Q(poh20[2]) );
  DRNQHSV2 \pe20/delaycell21/q_reg[6]  ( .D(n6731), .CK(clk), .RDN(n14803), 
        .Q(\pe20/ti_7t [6]) );
  DRNQHSV2 \pe6/delaycell24/q_reg[7]  ( .D(\pe6/poht [7]), .CK(clk), .RDN(
        n14768), .Q(poh6[7]) );
  DRNQHSV1 \pe11/delaycell5/q_reg[6]  ( .D(n15261), .CK(clk), .RDN(n14753), 
        .Q(\pe11/pvq [6]) );
  DRNQHSV2 \pe9/delaycell21/q_reg[5]  ( .D(n14963), .CK(clk), .RDN(n14721), 
        .Q(\pe9/ti_7t [5]) );
  DRNQHSV2 \pe16/delaycell5/q_reg[5]  ( .D(n15232), .CK(clk), .RDN(n14763), 
        .Q(\pe16/pvq [5]) );
  DRNQHSV1 \pe9/delaycell24/q_reg[6]  ( .D(\pe9/poht [6]), .CK(clk), .RDN(
        n14788), .Q(poh9[6]) );
  DRNQHSV2 \pe1/delaycell1/q_reg[3]  ( .D(ai[6]), .CK(clk), .RDN(n14797), .Q(
        \pe1/aot [6]) );
  DRNQHSV4 \pe8/delaycell5/q_reg[5]  ( .D(\pov7[5] ), .CK(clk), .RDN(n14720), 
        .Q(\pe8/pvq [5]) );
  DRNQHSV2 \pe19/delaycell21/q_reg[6]  ( .D(n14867), .CK(clk), .RDN(n14816), 
        .Q(\pe19/ti_7t [6]) );
  DRNQHSV2 \pe20/delaycell24/q_reg[5]  ( .D(\pe20/poht [5]), .CK(clk), .RDN(
        n14728), .Q(poh20[5]) );
  DRNQHSV2 \pe17/delaycell24/q_reg[5]  ( .D(\pe17/poht [5]), .CK(clk), .RDN(
        n14770), .Q(poh17[5]) );
  DRNQHSV2 \pe9/delaycell24/q_reg[3]  ( .D(\pe9/poht [3]), .CK(clk), .RDN(
        n15094), .Q(poh9[3]) );
  DRNQHSV2 \pe18/delaycell4/q_reg  ( .D(po17), .CK(clk), .RDN(n14814), .Q(
        \pe18/pq ) );
  DRNQHSV2 \pe14/delaycell4/q_reg  ( .D(po13), .CK(clk), .RDN(n14760), .Q(
        \pe14/pq ) );
  DRNQHSV4 \pe2/delaycell24/q_reg[5]  ( .D(\pe2/poht [5]), .CK(clk), .RDN(
        n14778), .Q(poh2[5]) );
  DRNQHSV2 \pe9/delaycell24/q_reg[5]  ( .D(\pe9/poht [5]), .CK(clk), .RDN(rst), 
        .Q(poh9[5]) );
  DRNQHSV2 \pe9/delaycell24/q_reg[2]  ( .D(\pe9/poht [2]), .CK(clk), .RDN(rst), 
        .Q(poh9[2]) );
  DRNQHSV2 \pe9/delaycell24/q_reg[4]  ( .D(\pe9/poht [4]), .CK(clk), .RDN(
        n14729), .Q(poh9[4]) );
  DRNQHSV2 \pe14/delaycell24/q_reg[2]  ( .D(\pe14/poht [2]), .CK(clk), .RDN(
        n14832), .Q(poh14[2]) );
  DRNQHSV2 \pe6/delaycell24/q_reg[6]  ( .D(\pe6/poht [6]), .CK(clk), .RDN(
        n14807), .Q(poh6[6]) );
  DRNQHSV1 \pe7/delaycell24/q_reg[4]  ( .D(\pe7/poht [4]), .CK(clk), .RDN(
        n14816), .Q(poh7[4]) );
  DRNQHSV1 \pe13/delaycell24/q_reg[5]  ( .D(\pe13/poht [5]), .CK(clk), .RDN(
        n14808), .Q(poh13[5]) );
  DRNQHSV2 \pe17/delaycell4/q_reg  ( .D(po16), .CK(clk), .RDN(n14774), .Q(
        \pe17/pq ) );
  DRNQHSV2 \pe2/delaycell24/q_reg[2]  ( .D(\pe2/poht [2]), .CK(clk), .RDN(
        n14722), .Q(poh2[2]) );
  DRNQHSV4 \pe1/delaycell1/q_reg[1]  ( .D(ai[8]), .CK(clk), .RDN(n14793), .Q(
        \pe1/aot [8]) );
  DRNQHSV4 \pe6/delaycell24/q_reg[4]  ( .D(\pe6/poht [4]), .CK(clk), .RDN(
        n14783), .Q(poh6[4]) );
  DRNQHSV2 \pe20/delaycell24/q_reg[6]  ( .D(\pe20/poht [6]), .CK(clk), .RDN(
        n14755), .Q(poh20[6]) );
  DRNQHSV2 \pe20/delaycell24/q_reg[7]  ( .D(\pe20/poht [7]), .CK(clk), .RDN(
        n14782), .Q(poh20[7]) );
  DRNQHSV2 \pe16/delaycell24/q_reg[5]  ( .D(\pe16/poht [5]), .CK(clk), .RDN(
        n14727), .Q(poh16[5]) );
  DRNQHSV4 \pe2/delaycell5/q_reg[3]  ( .D(pov1[3]), .CK(clk), .RDN(n14817), 
        .Q(\pe2/pvq [3]) );
  DRNQHSV2 \pe13/delaycell24/q_reg[4]  ( .D(\pe13/poht [4]), .CK(clk), .RDN(
        n14815), .Q(poh13[4]) );
  DRNQHSV4 \pe6/delaycell5/q_reg[6]  ( .D(n15205), .CK(clk), .RDN(n14759), .Q(
        \pe6/pvq [6]) );
  DRNQHSV2 \pe3/delaycell24/q_reg[3]  ( .D(\pe3/poht [3]), .CK(clk), .RDN(
        n14815), .Q(poh3[3]) );
  DRNQHSV4 \pe14/delaycell24/q_reg[4]  ( .D(\pe14/poht [4]), .CK(clk), .RDN(
        n14809), .Q(poh14[4]) );
  DRNQHSV2 \pe20/delaycell5/q_reg[3]  ( .D(n15212), .CK(clk), .RDN(n14789), 
        .Q(\pe20/pvq [3]) );
  DRNQHSV4 \pe20/delaycell24/q_reg[4]  ( .D(\pe20/poht [4]), .CK(clk), .RDN(
        n14718), .Q(poh20[4]) );
  DRNQHSV2 \pe14/delaycell24/q_reg[5]  ( .D(\pe14/poht [5]), .CK(clk), .RDN(
        n14714), .Q(poh14[5]) );
  DRNQHSV2 \pe14/delaycell5/q_reg[1]  ( .D(n15246), .CK(clk), .RDN(n14770), 
        .Q(\pe14/pvq [1]) );
  DRNQHSV2 \pe17/delaycell24/q_reg[3]  ( .D(\pe17/poht [3]), .CK(clk), .RDN(
        n14799), .Q(poh17[3]) );
  DRNQHSV4 \pe17/delaycell24/q_reg[1]  ( .D(\pe17/poht [1]), .CK(clk), .RDN(
        n14768), .Q(poh17[1]) );
  DRNQHSV2 \pe13/delaycell5/q_reg[1]  ( .D(n15253), .CK(clk), .RDN(n14752), 
        .Q(\pe13/pvq [1]) );
  NAND2HSV4 U6566 ( .A1(n6933), .A2(n6932), .ZN(n14707) );
  CLKNAND2HSV2 U6567 ( .A1(\pe7/got [5]), .A2(n14449), .ZN(n8696) );
  XNOR2HSV4 U6568 ( .A1(n9377), .A2(n5915), .ZN(n6474) );
  XOR2HSV2 U6569 ( .A1(n9376), .A2(n9375), .Z(n5915) );
  INHSV8 U6570 ( .I(ctro14), .ZN(n11156) );
  XOR2HSV2 U6571 ( .A1(n6715), .A2(n5916), .Z(\pe3/poht [1]) );
  CLKNAND2HSV2 U6572 ( .A1(n12973), .A2(n14931), .ZN(n5916) );
  NAND2HSV4 U6573 ( .A1(n15243), .A2(n9881), .ZN(n7471) );
  NAND2HSV4 U6574 ( .A1(n6150), .A2(n5917), .ZN(n9931) );
  INHSV4 U6575 ( .I(n5918), .ZN(n5917) );
  CLKNAND2HSV4 U6576 ( .A1(n9947), .A2(n7565), .ZN(n5918) );
  NAND2HSV2 U6577 ( .A1(n11973), .A2(\pe18/got [7]), .ZN(n11974) );
  CLKNAND2HSV0 U6578 ( .A1(n8418), .A2(n8417), .ZN(n8419) );
  CLKNHSV2 U6579 ( .I(n8964), .ZN(n8961) );
  XNOR2HSV4 U6580 ( .A1(n5920), .A2(n5919), .ZN(n12559) );
  CLKNAND2HSV2 U6581 ( .A1(n7519), .A2(\pe21/got [4]), .ZN(n5919) );
  XOR2HSV2 U6582 ( .A1(n12557), .A2(n5921), .Z(n5920) );
  CLKNHSV2 U6583 ( .I(n12558), .ZN(n5921) );
  NAND2HSV4 U6584 ( .A1(\pe17/aot [8]), .A2(\pe17/bq[8] ), .ZN(n6148) );
  CLKNAND2HSV4 U6585 ( .A1(n10046), .A2(n10045), .ZN(n7238) );
  INHSV4 U6586 ( .I(n13342), .ZN(n13343) );
  NAND2HSV4 U6587 ( .A1(n6583), .A2(n6584), .ZN(n10514) );
  XOR2HSV2 U6588 ( .A1(n12974), .A2(n5922), .Z(\pe3/poht [5]) );
  CLKNAND2HSV2 U6589 ( .A1(n12973), .A2(\pe3/got [3]), .ZN(n5922) );
  INHSV2 U6590 ( .I(n7756), .ZN(n7755) );
  INHSV4 U6591 ( .I(n6534), .ZN(n6535) );
  OAI21HSV2 U6592 ( .A1(n8237), .A2(n8238), .B(n8239), .ZN(\pe13/poht [4]) );
  NAND2HSV4 U6593 ( .A1(\pe2/pvq [3]), .A2(\pe2/ctrq ), .ZN(n6089) );
  MUX2NHSV4 U6594 ( .I0(n7954), .I1(n6090), .S(n6089), .ZN(n6088) );
  CLKXOR2HSV4 U6595 ( .A1(n10365), .A2(n10364), .Z(n10368) );
  INHSV4 U6596 ( .I(n11002), .ZN(n5970) );
  CLKNAND2HSV4 U6597 ( .A1(n7604), .A2(n9886), .ZN(n9903) );
  INHSV4 U6598 ( .I(n9903), .ZN(n6151) );
  NOR2HSV4 U6599 ( .A1(n11467), .A2(n11466), .ZN(n13890) );
  OAI21HSV4 U6600 ( .A1(n11453), .A2(n7157), .B(n11452), .ZN(n11466) );
  XOR3HSV2 U6601 ( .A1(n13675), .A2(n6850), .A3(n13678), .Z(n6055) );
  CLKNHSV4 U6602 ( .I(n9383), .ZN(n13795) );
  NAND2HSV2 U6603 ( .A1(n13749), .A2(\pe20/got [3]), .ZN(n6850) );
  CLKNAND2HSV4 U6604 ( .A1(n13236), .A2(n14864), .ZN(n12539) );
  CLKNAND2HSV2 U6605 ( .A1(n8498), .A2(n8497), .ZN(n8499) );
  NAND2HSV2 U6606 ( .A1(n14709), .A2(\pe20/got [2]), .ZN(n14178) );
  NAND2HSV4 U6607 ( .A1(n13681), .A2(n13682), .ZN(n14709) );
  CLKNAND2HSV4 U6608 ( .A1(n9007), .A2(n9006), .ZN(n9783) );
  CLKNAND2HSV2 U6609 ( .A1(n9783), .A2(n9420), .ZN(n8508) );
  CLKXOR2HSV4 U6610 ( .A1(n13579), .A2(n13578), .Z(n6712) );
  XOR2HSV0 U6611 ( .A1(n6712), .A2(n13586), .Z(n15199) );
  CLKNAND2HSV2 U6612 ( .A1(n6009), .A2(n8413), .ZN(n6008) );
  CLKNAND2HSV2 U6613 ( .A1(n12957), .A2(\pe3/got [6]), .ZN(n5984) );
  INHSV2 U6614 ( .I(n6085), .ZN(n5996) );
  BUFHSV6 U6615 ( .I(\pe10/bq[8] ), .Z(n12272) );
  CLKNAND2HSV4 U6616 ( .A1(\pe20/aot [8]), .A2(\pe20/bq[8] ), .ZN(n8204) );
  CLKNAND2HSV2 U6617 ( .A1(n8205), .A2(n8204), .ZN(n8206) );
  INHSV4 U6618 ( .I(n12538), .ZN(n6561) );
  CLKNHSV1 U6619 ( .I(n9398), .ZN(n10403) );
  CLKNAND2HSV4 U6620 ( .A1(n9735), .A2(n9420), .ZN(n9421) );
  CLKNHSV16 U6621 ( .I(n11093), .ZN(n8948) );
  CLKBUFHSV4 U6622 ( .I(\pe18/got [6]), .Z(n6039) );
  INHSV3 U6623 ( .I(n9056), .ZN(n9054) );
  NAND2HSV2 U6624 ( .A1(n7052), .A2(n10808), .ZN(n7051) );
  CLKNHSV6 U6625 ( .I(ctro11), .ZN(n11943) );
  CLKNHSV4 U6626 ( .I(ctro12), .ZN(n10747) );
  INHSV16 U6627 ( .I(ctro6), .ZN(n9832) );
  CLKNAND2HSV4 U6628 ( .A1(n8935), .A2(\pe6/pvq [6]), .ZN(n7863) );
  OAI21HSV2 U6629 ( .A1(n15237), .A2(n7119), .B(n7116), .ZN(n7855) );
  NAND2HSV2 U6630 ( .A1(n14179), .A2(\pe6/got [3]), .ZN(n12990) );
  INHSV2 U6631 ( .I(n13237), .ZN(n6440) );
  NAND2HSV4 U6632 ( .A1(n12512), .A2(n12511), .ZN(n14061) );
  NAND2HSV2 U6633 ( .A1(n14061), .A2(n14822), .ZN(n8426) );
  CLKNAND2HSV4 U6634 ( .A1(n5923), .A2(n6487), .ZN(n12271) );
  NAND2HSV4 U6635 ( .A1(n9641), .A2(n9640), .ZN(n5923) );
  INHSV4 U6636 ( .I(n8213), .ZN(n7859) );
  XNOR2HSV4 U6637 ( .A1(n5924), .A2(n6919), .ZN(po19) );
  XOR2HSV2 U6638 ( .A1(n6918), .A2(n6916), .Z(n5924) );
  NAND2HSV4 U6639 ( .A1(n15222), .A2(n5925), .ZN(n6441) );
  INHSV4 U6640 ( .I(n6597), .ZN(n5925) );
  CLKNAND2HSV4 U6641 ( .A1(n9359), .A2(n14818), .ZN(n8984) );
  CLKNAND2HSV3 U6642 ( .A1(n6169), .A2(\pe9/phq [3]), .ZN(n6307) );
  NAND2HSV8 U6643 ( .A1(n6489), .A2(n11036), .ZN(n11116) );
  NAND2HSV2 U6644 ( .A1(n7334), .A2(\pe18/got [8]), .ZN(n6835) );
  BUFHSV2 U6645 ( .I(n10836), .Z(n6207) );
  XNOR2HSV4 U6646 ( .A1(n5926), .A2(n7221), .ZN(n7720) );
  XNOR2HSV4 U6647 ( .A1(n7223), .A2(n10991), .ZN(n5926) );
  INHSV4 U6648 ( .I(n13237), .ZN(n6063) );
  OAI21HSV2 U6649 ( .A1(n8413), .A2(n6009), .B(n6008), .ZN(n8414) );
  NAND2HSV4 U6650 ( .A1(n10825), .A2(\pe21/got [7]), .ZN(n6992) );
  XNOR2HSV1 U6651 ( .A1(n14615), .A2(n14614), .ZN(n14616) );
  AOI21HSV2 U6652 ( .A1(n5927), .A2(n13348), .B(n13350), .ZN(n13349) );
  NOR2HSV4 U6653 ( .A1(n13347), .A2(n8913), .ZN(n5927) );
  OAI21HSV2 U6654 ( .A1(n10105), .A2(n8602), .B(n8603), .ZN(n8604) );
  INHSV2 U6655 ( .I(n15183), .ZN(n14465) );
  XNOR2HSV4 U6656 ( .A1(n5928), .A2(\pe18/phq [3]), .ZN(n6891) );
  CLKNAND2HSV2 U6657 ( .A1(\pe18/bq[6] ), .A2(\pe18/aot [8]), .ZN(n5928) );
  NAND2HSV2 U6658 ( .A1(n5929), .A2(n6400), .ZN(\pe17/poht [1]) );
  CLKNAND2HSV2 U6659 ( .A1(n6399), .A2(n6406), .ZN(n5929) );
  NAND2HSV2 U6660 ( .A1(n12997), .A2(\pe13/got [3]), .ZN(n7597) );
  CLKNAND2HSV2 U6661 ( .A1(\pe21/bq[7] ), .A2(\pe21/aot [8]), .ZN(n10364) );
  NAND2HSV2 U6662 ( .A1(n6440), .A2(\pe17/got [6]), .ZN(n6405) );
  NAND2HSV4 U6663 ( .A1(n10836), .A2(n5930), .ZN(n7721) );
  INHSV4 U6664 ( .I(n7729), .ZN(n5930) );
  MUX2NHSV4 U6665 ( .I0(n7273), .I1(n7272), .S(n13886), .ZN(n12512) );
  CLKNAND2HSV4 U6666 ( .A1(\pe18/aot [8]), .A2(\pe18/bq[8] ), .ZN(n9131) );
  INHSV4 U6667 ( .I(n7446), .ZN(n6286) );
  NAND2HSV4 U6668 ( .A1(\pe19/got [6]), .A2(\pe19/ti_1 ), .ZN(n9491) );
  NOR2HSV2 U6669 ( .A1(n13806), .A2(n13552), .ZN(n13553) );
  CLKNAND2HSV4 U6670 ( .A1(\pe21/aot [8]), .A2(\pe21/bq[6] ), .ZN(n7658) );
  CLKNAND2HSV8 U6671 ( .A1(n14572), .A2(\pe8/pvq [3]), .ZN(n10498) );
  AOI21HSV0 U6672 ( .A1(\pe7/got [5]), .A2(n15081), .B(n8591), .ZN(n8592) );
  NAND2HSV2 U6673 ( .A1(n8590), .A2(n5931), .ZN(n8591) );
  NAND2HSV2 U6674 ( .A1(n5933), .A2(n5932), .ZN(n5931) );
  INHSV2 U6675 ( .I(n8589), .ZN(n5932) );
  NOR2HSV0 U6676 ( .A1(n14465), .A2(n14464), .ZN(n5933) );
  NAND2HSV4 U6677 ( .A1(\pe10/bq[5] ), .A2(\pe10/aot [6]), .ZN(n10135) );
  CLKBUFHSV12 U6678 ( .I(n13910), .Z(n6209) );
  NAND2HSV2 U6679 ( .A1(n6209), .A2(\pe9/got [5]), .ZN(n8163) );
  OAI21HSV2 U6680 ( .A1(\pe7/phq [6]), .A2(n8843), .B(n8844), .ZN(n8845) );
  AOI21HSV4 U6681 ( .A1(n15195), .A2(n11117), .B(n7987), .ZN(n11118) );
  CLKNAND2HSV3 U6682 ( .A1(n5934), .A2(n8948), .ZN(n6982) );
  NAND2HSV2 U6683 ( .A1(n15078), .A2(n8955), .ZN(n5934) );
  XNOR2HSV4 U6684 ( .A1(n11119), .A2(n11118), .ZN(n15078) );
  OAI21HSV4 U6685 ( .A1(n7906), .A2(n7874), .B(n7907), .ZN(n11119) );
  NOR2HSV4 U6686 ( .A1(n15288), .A2(n10942), .ZN(n10948) );
  CLKNAND2HSV0 U6687 ( .A1(n15288), .A2(n10789), .ZN(n10972) );
  XNOR2HSV4 U6688 ( .A1(n6333), .A2(n10203), .ZN(n15288) );
  CLKNHSV3 U6689 ( .I(n12253), .ZN(n13624) );
  CLKNAND2HSV4 U6690 ( .A1(n5936), .A2(n5935), .ZN(n12253) );
  CLKNAND2HSV2 U6691 ( .A1(n5941), .A2(n5940), .ZN(n5935) );
  CLKNAND2HSV3 U6692 ( .A1(n5939), .A2(n5938), .ZN(n5936) );
  XNOR2HSV4 U6693 ( .A1(n12244), .A2(n12245), .ZN(n5940) );
  NAND3HSV4 U6694 ( .A1(n12204), .A2(n12308), .A3(n12205), .ZN(n12246) );
  INHSV2 U6695 ( .I(n12246), .ZN(n5937) );
  NOR2HSV4 U6696 ( .A1(n12231), .A2(n5937), .ZN(n5941) );
  INHSV2 U6697 ( .I(n5940), .ZN(n5938) );
  INHSV2 U6698 ( .I(n5941), .ZN(n5939) );
  CLKNAND2HSV3 U6699 ( .A1(n5942), .A2(\pe21/got [6]), .ZN(n10658) );
  INHSV2 U6700 ( .I(n10826), .ZN(n5942) );
  NOR2HSV0 U6701 ( .A1(n10826), .A2(n5943), .ZN(n10827) );
  INHSV2 U6702 ( .I(\pe21/got [5]), .ZN(n5943) );
  CLKNAND2HSV2 U6703 ( .A1(n10876), .A2(\pe21/got [3]), .ZN(n13119) );
  CLKNAND2HSV2 U6704 ( .A1(n10876), .A2(\pe21/got [1]), .ZN(n8384) );
  CLKNAND2HSV2 U6705 ( .A1(n10876), .A2(\pe21/got [2]), .ZN(n8058) );
  CLKNHSV2 U6706 ( .I(n10826), .ZN(n10876) );
  INHSV2 U6707 ( .I(n10825), .ZN(n10826) );
  CLKNAND2HSV4 U6708 ( .A1(\pe20/ti_1 ), .A2(\pe20/got [7]), .ZN(n9023) );
  NAND2HSV4 U6709 ( .A1(n9023), .A2(n9024), .ZN(n9022) );
  NAND2HSV4 U6710 ( .A1(\pe21/got [7]), .A2(n10396), .ZN(n8455) );
  INHSV4 U6711 ( .I(n10064), .ZN(n7024) );
  NAND2HSV2 U6712 ( .A1(n15075), .A2(n10148), .ZN(n10123) );
  CLKNHSV0 U6713 ( .I(n11002), .ZN(n11003) );
  CLKNAND2HSV4 U6714 ( .A1(n6841), .A2(n6840), .ZN(n6839) );
  INHSV6 U6715 ( .I(n10408), .ZN(n7324) );
  INHSV2 U6716 ( .I(n10853), .ZN(n7777) );
  CLKNAND2HSV3 U6717 ( .A1(n12134), .A2(n6398), .ZN(n6387) );
  OR2HSV2 U6718 ( .A1(n13872), .A2(n13269), .Z(n12012) );
  CLKNAND2HSV4 U6719 ( .A1(n6716), .A2(n8010), .ZN(n12059) );
  INHSV3 U6720 ( .I(n10069), .ZN(n10066) );
  CLKNAND2HSV2 U6721 ( .A1(n11880), .A2(n9465), .ZN(n9036) );
  CLKNAND2HSV0 U6722 ( .A1(n14061), .A2(n6721), .ZN(n8710) );
  INHSV6 U6723 ( .I(n10522), .ZN(n12337) );
  OAI21HSV4 U6724 ( .A1(n7203), .A2(n7204), .B(n7115), .ZN(n8430) );
  NAND2HSV2 U6725 ( .A1(n12811), .A2(\pe5/got [7]), .ZN(n10332) );
  CLKNAND2HSV2 U6726 ( .A1(n10145), .A2(\pe10/got [6]), .ZN(n10086) );
  CLKNHSV2 U6727 ( .I(n13882), .ZN(n7456) );
  XNOR2HSV4 U6728 ( .A1(n7462), .A2(n7461), .ZN(n13882) );
  INHSV4 U6729 ( .I(n9882), .ZN(n7602) );
  NAND2HSV4 U6730 ( .A1(n14708), .A2(\pe15/got [4]), .ZN(n12532) );
  XOR2HSV4 U6731 ( .A1(n11456), .A2(n11455), .Z(n11459) );
  INHSV24 U6732 ( .I(\pe8/phq [1]), .ZN(n5944) );
  INHSV2 U6733 ( .I(\pe8/pvq [1]), .ZN(n5945) );
  NOR2HSV4 U6734 ( .A1(n5945), .A2(n5944), .ZN(n10486) );
  NAND2HSV4 U6735 ( .A1(n11492), .A2(n13861), .ZN(n7626) );
  CLKBUFHSV12 U6736 ( .I(n14735), .Z(n5946) );
  CLKNAND2HSV2 U6737 ( .A1(n10052), .A2(n10051), .ZN(n10055) );
  NAND2HSV4 U6738 ( .A1(n10055), .A2(n10054), .ZN(n6225) );
  NAND2HSV4 U6739 ( .A1(n13759), .A2(\pe2/got [7]), .ZN(n7325) );
  NAND2HSV2 U6740 ( .A1(\pe5/got [8]), .A2(\pe5/ti_1 ), .ZN(n10289) );
  CLKNAND2HSV2 U6741 ( .A1(n8952), .A2(\pe10/got [2]), .ZN(n14108) );
  INHSV2 U6742 ( .I(n10933), .ZN(n10936) );
  CLKNAND2HSV2 U6743 ( .A1(n10936), .A2(n10935), .ZN(n10937) );
  NOR2HSV8 U6744 ( .A1(n6144), .A2(n6312), .ZN(n10052) );
  INHSV4 U6745 ( .I(n10368), .ZN(n10366) );
  INHSV4 U6746 ( .I(n8462), .ZN(n6109) );
  CLKNAND2HSV4 U6747 ( .A1(n6109), .A2(n6108), .ZN(n7476) );
  CLKNAND2HSV2 U6748 ( .A1(n6874), .A2(n5977), .ZN(n7608) );
  INHSV4 U6749 ( .I(n11786), .ZN(n14537) );
  AOI21HSV0 U6750 ( .A1(n11002), .A2(n12501), .B(n10996), .ZN(n8007) );
  CLKNAND2HSV4 U6751 ( .A1(\pe21/pvq [2]), .A2(\pe21/ctrq ), .ZN(n10360) );
  DELHS1 U6752 ( .I(\pe16/bq[8] ), .Z(n5947) );
  NAND2HSV2 U6753 ( .A1(n12230), .A2(n12229), .ZN(n12231) );
  CLKNAND2HSV2 U6754 ( .A1(n12957), .A2(n10995), .ZN(n6061) );
  NAND2HSV2 U6755 ( .A1(\pe11/got [5]), .A2(\pe11/ti_7[1] ), .ZN(n7920) );
  NOR2HSV4 U6756 ( .A1(n9135), .A2(n9134), .ZN(n9136) );
  INHSV2 U6757 ( .I(n13603), .ZN(n12991) );
  NOR2HSV8 U6758 ( .A1(n12991), .A2(n11964), .ZN(n11966) );
  CLKNAND2HSV2 U6759 ( .A1(n8183), .A2(n8184), .ZN(n8185) );
  CLKNAND2HSV2 U6760 ( .A1(n6030), .A2(n8182), .ZN(n8183) );
  CLKNAND2HSV2 U6761 ( .A1(\pe10/bq[6] ), .A2(\pe10/aot [8]), .ZN(n10053) );
  CLKXOR2HSV4 U6762 ( .A1(n12087), .A2(n12086), .Z(n7876) );
  DELHS1 U6763 ( .I(\pe8/aot [5]), .Z(n5948) );
  CLKNAND2HSV4 U6764 ( .A1(n10946), .A2(n14931), .ZN(n10204) );
  BUFHSV4 U6765 ( .I(\pe3/ti_7[1] ), .Z(n5949) );
  XOR2HSV2 U6766 ( .A1(n12964), .A2(n12963), .Z(\pe3/poht [4]) );
  NAND2HSV2 U6767 ( .A1(n6168), .A2(n5950), .ZN(n6977) );
  NAND3HSV2 U6768 ( .A1(n5951), .A2(\pe17/bq[7] ), .A3(\pe17/aot [7]), .ZN(
        n5950) );
  INHSV4 U6769 ( .I(\pe17/phq [3]), .ZN(n5951) );
  NAND2HSV4 U6770 ( .A1(\pe21/ctrq ), .A2(\pe21/pvq [1]), .ZN(n9393) );
  XNOR2HSV4 U6771 ( .A1(n6979), .A2(n5952), .ZN(n6978) );
  CLKNAND2HSV4 U6772 ( .A1(\pe17/bq[8] ), .A2(\pe17/aot [6]), .ZN(n5952) );
  NAND2HSV8 U6773 ( .A1(n10825), .A2(n10415), .ZN(n10810) );
  NAND2HSV4 U6774 ( .A1(n5953), .A2(n7872), .ZN(n6511) );
  CLKNAND2HSV4 U6775 ( .A1(n6110), .A2(n8464), .ZN(n5953) );
  NAND2HSV3 U6776 ( .A1(n10396), .A2(\pe21/got [6]), .ZN(n10397) );
  XNOR2HSV4 U6777 ( .A1(n7802), .A2(n13448), .ZN(\pe10/poht [4]) );
  XNOR2HSV4 U6778 ( .A1(n7812), .A2(n7811), .ZN(\pe10/poht [3]) );
  CLKNAND2HSV4 U6779 ( .A1(n15085), .A2(n13107), .ZN(n12100) );
  NOR2HSV3 U6780 ( .A1(n13759), .A2(n9358), .ZN(n7273) );
  NAND2HSV4 U6781 ( .A1(n9920), .A2(n14750), .ZN(n9906) );
  XNOR2HSV4 U6782 ( .A1(n6012), .A2(n5954), .ZN(n10384) );
  OAI21HSV4 U6783 ( .A1(n7656), .A2(n5956), .B(n5955), .ZN(n5954) );
  CLKNAND2HSV2 U6784 ( .A1(n7656), .A2(n8040), .ZN(n5955) );
  CLKNHSV2 U6785 ( .I(\pe21/phq [3]), .ZN(n5956) );
  NAND2HSV4 U6786 ( .A1(n13177), .A2(n13343), .ZN(n11972) );
  CLKNAND2HSV4 U6787 ( .A1(n6063), .A2(\pe17/got [4]), .ZN(n13249) );
  INHSV2 U6788 ( .I(n9947), .ZN(n6467) );
  CLKNAND2HSV4 U6789 ( .A1(n9847), .A2(n9846), .ZN(n6874) );
  NAND2HSV4 U6790 ( .A1(n6874), .A2(\pe6/got [3]), .ZN(n13008) );
  AND2HSV4 U6791 ( .A1(n12257), .A2(n12308), .Z(n12255) );
  INHSV2 U6792 ( .I(n8506), .ZN(n7677) );
  NAND2HSV2 U6793 ( .A1(n6613), .A2(n6611), .ZN(n6620) );
  XNOR2HSV4 U6794 ( .A1(n6446), .A2(n5957), .ZN(n9263) );
  CLKNAND2HSV2 U6795 ( .A1(n9823), .A2(\pe6/got [6]), .ZN(n5957) );
  NAND2HSV4 U6796 ( .A1(\pe5/bq[8] ), .A2(\pe5/aot [8]), .ZN(n10287) );
  CLKNAND2HSV2 U6797 ( .A1(n8710), .A2(n8709), .ZN(n8711) );
  CLKNHSV6 U6798 ( .I(n10404), .ZN(n7871) );
  AOI31HSV2 U6799 ( .A1(n10705), .A2(n13219), .A3(n14064), .B(n7522), .ZN(
        n6214) );
  XNOR2HSV4 U6800 ( .A1(n10675), .A2(n10674), .ZN(n10705) );
  NAND2HSV2 U6801 ( .A1(n10459), .A2(n14852), .ZN(n8600) );
  DELHS1 U6802 ( .I(\pe12/got [8]), .Z(n5958) );
  NAND2HSV2 U6803 ( .A1(n8371), .A2(n8370), .ZN(n8372) );
  CLKNAND2HSV2 U6804 ( .A1(n8369), .A2(n5959), .ZN(n8370) );
  CLKNAND2HSV2 U6805 ( .A1(n5961), .A2(n5960), .ZN(n5959) );
  CLKNHSV2 U6806 ( .I(n8368), .ZN(n5960) );
  CLKNHSV2 U6807 ( .I(n8367), .ZN(n5961) );
  INHSV2 U6808 ( .I(n6519), .ZN(n5975) );
  CLKNAND2HSV4 U6809 ( .A1(n15282), .A2(n14955), .ZN(n12603) );
  NAND2HSV2 U6810 ( .A1(\pe17/aot [8]), .A2(\pe17/bq[7] ), .ZN(n6501) );
  XOR2HSV4 U6811 ( .A1(n12026), .A2(n6664), .Z(n6663) );
  XNOR2HSV2 U6812 ( .A1(n9771), .A2(n9770), .ZN(n9781) );
  NOR2HSV3 U6813 ( .A1(n10191), .A2(n10169), .ZN(n6331) );
  NAND2HSV2 U6814 ( .A1(n14846), .A2(\pe5/got [3]), .ZN(n8537) );
  CLKNAND2HSV3 U6815 ( .A1(n10867), .A2(n7785), .ZN(n7784) );
  CLKNAND2HSV4 U6816 ( .A1(n7053), .A2(n7052), .ZN(n11774) );
  NAND2HSV4 U6817 ( .A1(n6989), .A2(n5962), .ZN(n7053) );
  NAND2HSV2 U6818 ( .A1(n10394), .A2(n10393), .ZN(n5962) );
  CLKNAND2HSV4 U6819 ( .A1(n7424), .A2(n7423), .ZN(n5998) );
  INHSV2 U6820 ( .I(n10589), .ZN(n8643) );
  NAND2HSV4 U6821 ( .A1(n7030), .A2(n7029), .ZN(n10589) );
  NAND2HSV2 U6822 ( .A1(n13811), .A2(\pe11/got [4]), .ZN(n11715) );
  INHSV4 U6823 ( .I(n10873), .ZN(n10874) );
  NAND2HSV2 U6824 ( .A1(n8463), .A2(n8462), .ZN(n7475) );
  CLKNAND2HSV4 U6825 ( .A1(n10644), .A2(n13107), .ZN(n10645) );
  CLKNAND2HSV3 U6826 ( .A1(n11270), .A2(n11271), .ZN(n7747) );
  CLKNAND2HSV3 U6827 ( .A1(n7874), .A2(n7906), .ZN(n7907) );
  XNOR2HSV4 U6828 ( .A1(n7851), .A2(n7854), .ZN(n6329) );
  CLKXOR2HSV4 U6829 ( .A1(n6369), .A2(n6368), .Z(n6105) );
  NAND2HSV4 U6830 ( .A1(n7858), .A2(n7859), .ZN(n7424) );
  OAI21HSV4 U6831 ( .A1(n7529), .A2(n12110), .B(n8213), .ZN(n7423) );
  CLKNHSV6 U6832 ( .I(n13190), .ZN(n14069) );
  NAND2HSV4 U6833 ( .A1(n14069), .A2(\pe16/got [3]), .ZN(n13200) );
  INHSV2 U6834 ( .I(n10470), .ZN(n13841) );
  AOI22HSV4 U6835 ( .A1(n13677), .A2(\pe20/ti_7t [7]), .B1(n11887), .B2(n13794), .ZN(n13682) );
  INHSV2 U6836 ( .I(n7010), .ZN(n7009) );
  CLKNAND2HSV4 U6837 ( .A1(n7490), .A2(n6134), .ZN(n6133) );
  NAND2HSV4 U6838 ( .A1(n6133), .A2(n11468), .ZN(n6132) );
  XNOR2HSV4 U6839 ( .A1(n6822), .A2(n6820), .ZN(\pe10/poht [5]) );
  INHSV4 U6840 ( .I(n8975), .ZN(n6064) );
  INHSV2 U6841 ( .I(n7797), .ZN(n6138) );
  AOI21HSV2 U6842 ( .A1(n6944), .A2(n6941), .B(n6939), .ZN(n9454) );
  XNOR2HSV4 U6843 ( .A1(n7248), .A2(n7251), .ZN(n6701) );
  XNOR2HSV4 U6844 ( .A1(n7923), .A2(n5963), .ZN(n7929) );
  XNOR2HSV4 U6845 ( .A1(n7928), .A2(n7927), .ZN(n5963) );
  NAND2HSV2 U6846 ( .A1(n6181), .A2(\pe4/got [2]), .ZN(n12086) );
  NAND2HSV2 U6847 ( .A1(n10733), .A2(n10734), .ZN(n10732) );
  AOI21HSV0 U6848 ( .A1(n6810), .A2(n5964), .B(n11693), .ZN(n11694) );
  NOR2HSV2 U6849 ( .A1(n11692), .A2(n9794), .ZN(n5964) );
  CLKNHSV0 U6850 ( .I(n12250), .ZN(n12251) );
  NAND2HSV4 U6851 ( .A1(n13857), .A2(n11296), .ZN(n7304) );
  NAND2HSV4 U6852 ( .A1(n9382), .A2(n13796), .ZN(n11238) );
  XOR3HSV2 U6853 ( .A1(n8268), .A2(n7614), .A3(n5965), .Z(n8270) );
  CLKNHSV2 U6854 ( .I(n7613), .ZN(n5965) );
  INHSV2 U6855 ( .I(n7051), .ZN(n7050) );
  XNOR2HSV4 U6856 ( .A1(n12423), .A2(n7760), .ZN(n7759) );
  INHSV4 U6857 ( .I(n11091), .ZN(n11036) );
  CLKNAND2HSV1 U6858 ( .A1(\pe21/got [5]), .A2(n10840), .ZN(n7970) );
  CLKNAND2HSV2 U6859 ( .A1(n13759), .A2(\pe2/got [3]), .ZN(n12917) );
  XNOR2HSV4 U6860 ( .A1(n6046), .A2(n11143), .ZN(\pe14/poht [4]) );
  DELHS1 U6861 ( .I(\pe10/got [6]), .Z(n5966) );
  INHSV4 U6862 ( .I(n13190), .ZN(n14348) );
  CLKNAND2HSV4 U6863 ( .A1(n14348), .A2(\pe16/got [2]), .ZN(n11222) );
  CLKNAND2HSV2 U6864 ( .A1(n13831), .A2(n14822), .ZN(n7101) );
  CLKXOR2HSV2 U6865 ( .A1(n7101), .A2(n12881), .Z(n6086) );
  CLKNAND2HSV4 U6866 ( .A1(n7805), .A2(n7870), .ZN(n10945) );
  NAND2HSV4 U6867 ( .A1(n7871), .A2(n10408), .ZN(n7870) );
  NAND2HSV2 U6868 ( .A1(n14012), .A2(n14011), .ZN(n12134) );
  DELHS1 U6869 ( .I(\pe7/got [8]), .Z(n5967) );
  DELHS1 U6870 ( .I(\pe14/ti_1 ), .Z(n5968) );
  XNOR2HSV4 U6871 ( .A1(n10196), .A2(n10197), .ZN(n7174) );
  NAND2HSV4 U6872 ( .A1(n15086), .A2(\pe4/got [5]), .ZN(n10579) );
  NAND3HSV4 U6873 ( .A1(n8972), .A2(n8973), .A3(n8974), .ZN(n8971) );
  INHSV4 U6874 ( .I(n8971), .ZN(n8977) );
  CLKNAND2HSV2 U6875 ( .A1(\pe2/ti_1 ), .A2(\pe2/got [4]), .ZN(n6505) );
  NOR2HSV4 U6876 ( .A1(n10716), .A2(n14397), .ZN(n12015) );
  NAND2HSV4 U6877 ( .A1(n15242), .A2(n9881), .ZN(n9923) );
  XNOR2HSV4 U6878 ( .A1(n7248), .A2(n7251), .ZN(n10124) );
  CLKNAND2HSV1 U6879 ( .A1(n13089), .A2(\pe14/got [6]), .ZN(n8418) );
  INHSV2 U6880 ( .I(n6560), .ZN(n6559) );
  CLKBUFHSV12 U6881 ( .I(\pe14/ti_7[3] ), .Z(n5969) );
  NAND2HSV2 U6882 ( .A1(\pe15/got [3]), .A2(\pe15/ti_1 ), .ZN(n11381) );
  XNOR2HSV4 U6883 ( .A1(n14613), .A2(n14612), .ZN(n14615) );
  XNOR2HSV4 U6884 ( .A1(n11751), .A2(n11750), .ZN(n11759) );
  NAND2HSV4 U6885 ( .A1(\pe15/bq[5] ), .A2(\pe15/aot [6]), .ZN(n7463) );
  NOR2HSV4 U6886 ( .A1(n5970), .A2(n10994), .ZN(n11001) );
  MUX2NHSV4 U6887 ( .I0(\pe20/phq [1]), .I1(n9010), .S(n5971), .ZN(n9031) );
  NAND2HSV4 U6888 ( .A1(\pe20/ctrq ), .A2(\pe20/pvq [1]), .ZN(n5971) );
  CLKNHSV2 U6889 ( .I(n6213), .ZN(n6211) );
  CLKNAND2HSV2 U6890 ( .A1(n6215), .A2(n6214), .ZN(n6213) );
  CLKNAND2HSV2 U6891 ( .A1(n10595), .A2(n13645), .ZN(n10597) );
  INHSV8 U6892 ( .I(n6241), .ZN(n5972) );
  IOA21HSV4 U6893 ( .A1(n6243), .A2(n8554), .B(n5972), .ZN(n6240) );
  NAND2HSV4 U6894 ( .A1(n6026), .A2(\pe20/got [5]), .ZN(n9482) );
  NAND2HSV4 U6895 ( .A1(n11092), .A2(\pe14/got [7]), .ZN(n7853) );
  BUFHSV2 U6896 ( .I(\pe17/aot [6]), .Z(n5973) );
  NAND2HSV4 U6897 ( .A1(n7360), .A2(n10406), .ZN(n10404) );
  NAND2HSV4 U6898 ( .A1(n8908), .A2(n7828), .ZN(n6885) );
  CLKNHSV8 U6899 ( .I(n10873), .ZN(n10865) );
  NOR2HSV2 U6900 ( .A1(n13749), .A2(n15177), .ZN(n11887) );
  NOR2HSV8 U6901 ( .A1(n11114), .A2(n13852), .ZN(n7986) );
  XNOR3HSV2 U6902 ( .A1(n13228), .A2(n13227), .A3(n13226), .ZN(n13231) );
  XOR3HSV2 U6903 ( .A1(n14296), .A2(n14295), .A3(n14294), .Z(n14300) );
  NAND2HSV4 U6904 ( .A1(n12537), .A2(n6561), .ZN(n14853) );
  XNOR2HSV4 U6905 ( .A1(n6523), .A2(n5974), .ZN(n6518) );
  XNOR2HSV4 U6906 ( .A1(n6522), .A2(n5975), .ZN(n5974) );
  NAND3HSV3 U6907 ( .A1(n13841), .A2(n10439), .A3(n14429), .ZN(n6463) );
  NOR2HSV2 U6908 ( .A1(n6383), .A2(n6572), .ZN(n6382) );
  NAND2HSV4 U6909 ( .A1(n6556), .A2(n6555), .ZN(n6554) );
  NAND2HSV4 U6910 ( .A1(n7500), .A2(n11943), .ZN(n5990) );
  NAND2HSV4 U6911 ( .A1(n5990), .A2(n11714), .ZN(n7502) );
  NAND2HSV4 U6912 ( .A1(\pe10/bq[7] ), .A2(\pe10/aot [6]), .ZN(n6070) );
  AOI21HSV2 U6913 ( .A1(n11978), .A2(n13138), .B(n7009), .ZN(n11979) );
  CLKNAND2HSV4 U6914 ( .A1(n6298), .A2(n6297), .ZN(n6099) );
  NAND2HSV4 U6915 ( .A1(n6099), .A2(n6098), .ZN(n6097) );
  NAND2HSV4 U6916 ( .A1(n6514), .A2(n10690), .ZN(\pe16/ti_7[1] ) );
  CLKBUFHSV12 U6917 ( .I(n13911), .Z(n5976) );
  NAND2HSV4 U6918 ( .A1(n12387), .A2(n14841), .ZN(n6918) );
  NAND3HSV3 U6919 ( .A1(n10677), .A2(n14292), .A3(n10796), .ZN(n10679) );
  DELHS1 U6920 ( .I(\pe6/got [7]), .Z(n5977) );
  NAND2HSV0 U6921 ( .A1(n8467), .A2(n8466), .ZN(n8468) );
  CLKNAND2HSV2 U6922 ( .A1(\pe14/got [7]), .A2(\pe14/ti_1 ), .ZN(n8466) );
  CLKXOR2HSV4 U6923 ( .A1(n10696), .A2(n10695), .Z(n10703) );
  CLKNAND2HSV4 U6924 ( .A1(n14450), .A2(\pe7/got [2]), .ZN(n8687) );
  INHSV2 U6925 ( .I(n14489), .ZN(n6010) );
  NAND2HSV2 U6926 ( .A1(n6126), .A2(n6124), .ZN(n6130) );
  NAND2HSV4 U6927 ( .A1(n15235), .A2(n10521), .ZN(n10790) );
  CLKNAND2HSV2 U6928 ( .A1(n8309), .A2(n7139), .ZN(n7133) );
  INHSV4 U6929 ( .I(n7133), .ZN(n7132) );
  AOI21HSV4 U6930 ( .A1(n9351), .A2(n9364), .B(n9355), .ZN(n9352) );
  XNOR2HSV4 U6931 ( .A1(n11737), .A2(n5978), .ZN(n11741) );
  CLKNAND2HSV2 U6932 ( .A1(n14381), .A2(\pe11/got [7]), .ZN(n5978) );
  NAND2HSV4 U6933 ( .A1(\pe16/bq[8] ), .A2(\pe16/aot [6]), .ZN(n10664) );
  NAND3HSV4 U6934 ( .A1(n11002), .A2(n11773), .A3(n10188), .ZN(n11707) );
  CLKNAND2HSV2 U6935 ( .A1(n11707), .A2(n10188), .ZN(n10940) );
  CLKXOR2HSV4 U6936 ( .A1(n11187), .A2(n11186), .Z(n11188) );
  NAND2HSV4 U6937 ( .A1(n5982), .A2(n5979), .ZN(n10346) );
  CLKNAND2HSV2 U6938 ( .A1(n5981), .A2(n5980), .ZN(n5979) );
  CLKNHSV2 U6939 ( .I(n10320), .ZN(n5980) );
  CLKNHSV2 U6940 ( .I(n10307), .ZN(n5981) );
  CLKNAND2HSV2 U6941 ( .A1(n10527), .A2(n10307), .ZN(n5982) );
  XNOR2HSV4 U6942 ( .A1(n5983), .A2(n6062), .ZN(n6715) );
  XNOR2HSV4 U6943 ( .A1(n5984), .A2(n12767), .ZN(n5983) );
  INHSV3 U6944 ( .I(n10170), .ZN(n10185) );
  CLKNAND2HSV2 U6945 ( .A1(n8573), .A2(n8572), .ZN(n8574) );
  CLKNAND2HSV2 U6946 ( .A1(n15168), .A2(\pe18/got [2]), .ZN(n14698) );
  XNOR2HSV4 U6947 ( .A1(n13187), .A2(n5985), .ZN(po18) );
  CLKNAND2HSV2 U6948 ( .A1(n14695), .A2(n5997), .ZN(n5985) );
  NAND3HSV2 U6949 ( .A1(n10583), .A2(n9713), .A3(n9712), .ZN(n9715) );
  XNOR2HSV4 U6950 ( .A1(n9667), .A2(n9666), .ZN(n10583) );
  CLKNAND2HSV4 U6951 ( .A1(n15241), .A2(n9881), .ZN(n9991) );
  CLKNAND2HSV4 U6952 ( .A1(n9991), .A2(n9990), .ZN(n12997) );
  CLKNHSV0 U6953 ( .I(n11444), .ZN(n7206) );
  NAND2HSV3 U6954 ( .A1(n12940), .A2(n12941), .ZN(n14449) );
  NAND2HSV3 U6955 ( .A1(n8952), .A2(n5966), .ZN(n6024) );
  CLKXOR2HSV4 U6956 ( .A1(n11279), .A2(n11278), .Z(n11281) );
  CLKNAND2HSV1 U6957 ( .A1(n12253), .A2(n12251), .ZN(n12257) );
  CLKNAND2HSV2 U6958 ( .A1(n15168), .A2(n6039), .ZN(n14648) );
  NAND2HSV4 U6959 ( .A1(\pe2/aot [6]), .A2(\pe2/bq[8] ), .ZN(n6085) );
  INHSV2 U6960 ( .I(n15241), .ZN(n8309) );
  INHSV4 U6961 ( .I(n10766), .ZN(n7155) );
  AOI21HSV4 U6962 ( .A1(n5988), .A2(n5987), .B(n5986), .ZN(n6016) );
  INHSV2 U6963 ( .I(n6017), .ZN(n5986) );
  INHSV2 U6964 ( .I(n9713), .ZN(n5987) );
  INHSV4 U6965 ( .I(n10583), .ZN(n5988) );
  XOR2HSV2 U6966 ( .A1(n10890), .A2(n5989), .Z(\pe21/poht [4]) );
  XNOR2HSV4 U6967 ( .A1(n10889), .A2(n10888), .ZN(n5989) );
  NAND2HSV1 U6968 ( .A1(\pe9/got [5]), .A2(\pe9/ti_1 ), .ZN(n9424) );
  CLKNHSV6 U6969 ( .I(n14854), .ZN(n11924) );
  XNOR2HSV4 U6970 ( .A1(n7685), .A2(n11767), .ZN(n7500) );
  INHSV4 U6971 ( .I(n9328), .ZN(n14858) );
  CLKNAND2HSV2 U6972 ( .A1(n14858), .A2(\pe2/bq[3] ), .ZN(n9329) );
  IOA21HSV4 U6973 ( .A1(n14707), .A2(n9378), .B(n9338), .ZN(\pe2/ti_7[1] ) );
  CLKNAND2HSV0 U6974 ( .A1(\pe3/got [4]), .A2(n14819), .ZN(n12963) );
  NAND2HSV4 U6975 ( .A1(n8970), .A2(n8969), .ZN(n8974) );
  NAND3HSV3 U6976 ( .A1(\pe2/phq [2]), .A2(\pe2/bq[7] ), .A3(\pe2/aot [8]), 
        .ZN(n8973) );
  XNOR2HSV4 U6977 ( .A1(n5992), .A2(n5991), .ZN(n12499) );
  CLKNHSV2 U6978 ( .I(n12496), .ZN(n5991) );
  CLKNAND2HSV2 U6979 ( .A1(n12957), .A2(n14931), .ZN(n5992) );
  NAND2HSV2 U6980 ( .A1(n15190), .A2(\pe12/got [2]), .ZN(n14443) );
  XNOR2HSV4 U6981 ( .A1(n5993), .A2(n12220), .ZN(n8902) );
  XNOR2HSV4 U6982 ( .A1(n12221), .A2(n5994), .ZN(n5993) );
  CLKNHSV2 U6983 ( .I(n12222), .ZN(n5994) );
  CLKNAND2HSV4 U6984 ( .A1(n6548), .A2(n6547), .ZN(n12195) );
  INHSV4 U6985 ( .I(n12195), .ZN(n10682) );
  CLKNAND2HSV4 U6986 ( .A1(\pe16/aot [6]), .A2(\pe16/bq[7] ), .ZN(n8548) );
  NAND3HSV2 U6987 ( .A1(n7384), .A2(n7385), .A3(n10307), .ZN(n7380) );
  NAND2HSV2 U6988 ( .A1(n7380), .A2(n11472), .ZN(n6953) );
  NAND2HSV2 U6989 ( .A1(n12957), .A2(\pe3/got [3]), .ZN(n12961) );
  NAND2HSV4 U6990 ( .A1(\pe20/aot [6]), .A2(\pe20/bq[8] ), .ZN(n9016) );
  CLKNAND2HSV4 U6991 ( .A1(n11116), .A2(\pe14/got [7]), .ZN(n7874) );
  NAND2HSV2 U6992 ( .A1(\pe2/bq[7] ), .A2(\pe2/aot [8]), .ZN(n8970) );
  INHSV2 U6993 ( .I(n6725), .ZN(n6116) );
  CLKNAND2HSV4 U6994 ( .A1(\pe2/aot [5]), .A2(\pe2/bq[7] ), .ZN(n9367) );
  CLKXOR2HSV2 U6995 ( .A1(n9368), .A2(n9367), .Z(n9369) );
  BUFHSV6 U6996 ( .I(\pe17/ti_1 ), .Z(n14415) );
  CLKNAND2HSV2 U6997 ( .A1(n5996), .A2(n5995), .ZN(n6083) );
  CLKNAND2HSV2 U6998 ( .A1(\pe2/bq[6] ), .A2(\pe2/aot [8]), .ZN(n5995) );
  CLKNAND2HSV4 U6999 ( .A1(n9133), .A2(\pe18/ti_7t [6]), .ZN(n13176) );
  AND2HSV4 U7000 ( .A1(\pe2/ctrq ), .A2(\pe2/pvq [2]), .Z(n8972) );
  INHSV4 U7001 ( .I(n8463), .ZN(n6108) );
  NAND2HSV4 U7002 ( .A1(n10202), .A2(n15180), .ZN(n6330) );
  CLKNAND2HSV4 U7003 ( .A1(n6569), .A2(\pe17/got [6]), .ZN(n6517) );
  NAND3HSV4 U7004 ( .A1(n10438), .A2(n10470), .A3(n13252), .ZN(n10713) );
  INHSV4 U7005 ( .I(n7736), .ZN(n7361) );
  NAND2HSV2 U7006 ( .A1(\pe19/ctrq ), .A2(\pe19/pvq [3]), .ZN(n9493) );
  CLKXOR2HSV4 U7007 ( .A1(n13509), .A2(n13508), .Z(n13510) );
  CLKNAND2HSV2 U7008 ( .A1(\pe13/ti_7[1] ), .A2(\pe13/got [5]), .ZN(n9918) );
  CLKNAND2HSV2 U7009 ( .A1(n12246), .A2(n12208), .ZN(n12223) );
  DELHS1 U7010 ( .I(\pe18/got [8]), .Z(n5997) );
  NAND2HSV0 U7011 ( .A1(n14179), .A2(\pe6/got [5]), .ZN(n8229) );
  INHSV2 U7012 ( .I(n6428), .ZN(n6427) );
  NAND2HSV4 U7013 ( .A1(n9957), .A2(\pe13/got [6]), .ZN(n6472) );
  CLKNAND2HSV4 U7014 ( .A1(n7693), .A2(n7696), .ZN(n7692) );
  INHSV6 U7015 ( .I(n9977), .ZN(n15087) );
  INHSV4 U7016 ( .I(n6329), .ZN(n6983) );
  CLKNHSV4 U7017 ( .I(\pe17/pvq [1]), .ZN(n9135) );
  CLKNAND2HSV2 U7018 ( .A1(n12973), .A2(n15180), .ZN(n12504) );
  CLKNAND2HSV2 U7019 ( .A1(n12503), .A2(n12502), .ZN(n12973) );
  CLKBUFHSV6 U7020 ( .I(n8942), .Z(n13677) );
  CLKNHSV8 U7021 ( .I(n10058), .ZN(n10599) );
  XNOR2HSV4 U7022 ( .A1(n12005), .A2(n12004), .ZN(n6204) );
  CLKNAND2HSV2 U7023 ( .A1(n11979), .A2(n11975), .ZN(n12005) );
  NAND2HSV4 U7024 ( .A1(n10145), .A2(\pe10/got [7]), .ZN(n7251) );
  NAND2HSV4 U7025 ( .A1(n15078), .A2(n11156), .ZN(n11227) );
  INHSV2 U7026 ( .I(n6433), .ZN(n6432) );
  XOR2HSV4 U7027 ( .A1(n9762), .A2(n9761), .Z(n9796) );
  INHSV4 U7028 ( .I(n10594), .ZN(n10596) );
  NAND2HSV2 U7029 ( .A1(\pe6/ti_1 ), .A2(\pe6/got [6]), .ZN(n9221) );
  XNOR2HSV4 U7030 ( .A1(n11697), .A2(n11696), .ZN(\pe9/poht [3]) );
  CLKNAND2HSV2 U7031 ( .A1(\pe16/aot [7]), .A2(\pe16/bq[7] ), .ZN(n10662) );
  INHSV4 U7032 ( .I(\pe10/bq[7] ), .ZN(n6312) );
  NAND2HSV4 U7033 ( .A1(n7632), .A2(n9799), .ZN(\pe6/ti_7[5] ) );
  INHSV2 U7034 ( .I(n6295), .ZN(n6096) );
  XNOR2HSV4 U7035 ( .A1(n5998), .A2(n8214), .ZN(n7422) );
  CLKXOR2HSV2 U7036 ( .A1(n9930), .A2(n9929), .Z(n8475) );
  INHSV2 U7037 ( .I(n10355), .ZN(n14219) );
  OAI21HSV2 U7038 ( .A1(n8425), .A2(n8426), .B(n8427), .ZN(\pe2/poht [2]) );
  CLKNAND2HSV2 U7039 ( .A1(n13759), .A2(\pe2/got [2]), .ZN(n11240) );
  NAND2HSV1 U7040 ( .A1(\pe13/got [1]), .A2(n14961), .ZN(n8859) );
  CLKNAND2HSV4 U7041 ( .A1(\pe7/ctrq ), .A2(\pe7/pvq [1]), .ZN(n7619) );
  INHSV6 U7042 ( .I(n12629), .ZN(n13089) );
  NAND2HSV4 U7043 ( .A1(n5999), .A2(n10713), .ZN(n6569) );
  INHSV2 U7044 ( .I(n6284), .ZN(n5999) );
  NOR2HSV4 U7045 ( .A1(n7140), .A2(n10403), .ZN(n10859) );
  XNOR2HSV4 U7046 ( .A1(n6000), .A2(n10727), .ZN(n6292) );
  XNOR2HSV4 U7047 ( .A1(n6293), .A2(n6001), .ZN(n6000) );
  XOR2HSV2 U7048 ( .A1(n10722), .A2(\pe12/phq [3]), .Z(n6001) );
  AOI21HSV4 U7049 ( .A1(n11330), .A2(n12317), .B(n10522), .ZN(n11329) );
  CLKNAND2HSV4 U7050 ( .A1(n6282), .A2(n10869), .ZN(n6281) );
  INHSV2 U7051 ( .I(n7913), .ZN(n7829) );
  CLKNAND2HSV4 U7052 ( .A1(n7366), .A2(n6002), .ZN(n7875) );
  NAND2HSV4 U7053 ( .A1(n7792), .A2(n6003), .ZN(n6002) );
  INHSV2 U7054 ( .I(n11692), .ZN(n6003) );
  NAND2HSV4 U7055 ( .A1(n13604), .A2(\pe13/got [2]), .ZN(n6052) );
  CLKNAND2HSV4 U7056 ( .A1(n13752), .A2(n13718), .ZN(n13719) );
  CLKNAND2HSV4 U7057 ( .A1(n10524), .A2(n12194), .ZN(n10677) );
  NAND2HSV4 U7058 ( .A1(n15188), .A2(\pe13/got [6]), .ZN(n10028) );
  BUFHSV4 U7059 ( .I(n14582), .Z(n6810) );
  NAND2HSV4 U7060 ( .A1(n6771), .A2(n6981), .ZN(n13581) );
  NAND2HSV4 U7061 ( .A1(n9847), .A2(n7437), .ZN(n6840) );
  XNOR2HSV1 U7062 ( .A1(n14048), .A2(n14047), .ZN(n14060) );
  CLKBUFHSV12 U7063 ( .I(\pe16/bq[7] ), .Z(n6004) );
  NAND2HSV4 U7064 ( .A1(n7025), .A2(n6005), .ZN(n10062) );
  INHSV2 U7065 ( .I(n6006), .ZN(n6005) );
  NAND2HSV2 U7066 ( .A1(n15264), .A2(n10148), .ZN(n6006) );
  CLKNAND2HSV4 U7067 ( .A1(n7027), .A2(n7026), .ZN(n7025) );
  XNOR2HSV4 U7068 ( .A1(n9892), .A2(n6007), .ZN(n9897) );
  XOR2HSV2 U7069 ( .A1(n9891), .A2(n9890), .Z(n6007) );
  CLKNAND2HSV4 U7070 ( .A1(n12336), .A2(n15235), .ZN(n10523) );
  OAI21HSV2 U7071 ( .A1(n9269), .A2(n9306), .B(n9268), .ZN(n6139) );
  CLKXOR2HSV2 U7072 ( .A1(n12429), .A2(n11925), .Z(n11926) );
  CLKXOR2HSV4 U7073 ( .A1(n11927), .A2(n11926), .Z(n11935) );
  NAND2HSV2 U7074 ( .A1(\pe21/bq[3] ), .A2(\pe21/aot [8]), .ZN(n10817) );
  NAND2HSV2 U7075 ( .A1(n14948), .A2(\pe12/bq[4] ), .ZN(n11423) );
  INHSV4 U7076 ( .I(n10385), .ZN(n10386) );
  CLKNHSV24 U7077 ( .I(n9381), .ZN(n9358) );
  CLKNAND2HSV8 U7078 ( .A1(n15215), .A2(n11976), .ZN(n13177) );
  INAND2HSV4 U7079 ( .A1(n11144), .B1(n6010), .ZN(n6009) );
  INHSV4 U7080 ( .I(n10216), .ZN(n14872) );
  INHSV4 U7081 ( .I(n11743), .ZN(n7499) );
  INHSV2 U7082 ( .I(n10202), .ZN(n10216) );
  XOR2HSV4 U7083 ( .A1(n13200), .A2(n13199), .Z(n13202) );
  CLKNAND2HSV2 U7084 ( .A1(n12347), .A2(n6011), .ZN(n7674) );
  CLKNHSV2 U7085 ( .I(n11948), .ZN(n6011) );
  XNOR2HSV4 U7086 ( .A1(n7502), .A2(n7503), .ZN(n12347) );
  CLKNAND2HSV4 U7087 ( .A1(n6204), .A2(n12006), .ZN(n12009) );
  CLKNAND2HSV4 U7088 ( .A1(n6612), .A2(n7331), .ZN(n6623) );
  NAND2HSV2 U7089 ( .A1(n6623), .A2(n6614), .ZN(n6611) );
  CLKXOR2HSV2 U7090 ( .A1(n13553), .A2(n13577), .Z(n13578) );
  INHSV4 U7091 ( .I(n10682), .ZN(n6965) );
  CLKNAND2HSV4 U7092 ( .A1(n6965), .A2(n6969), .ZN(n6964) );
  CLKNAND2HSV2 U7093 ( .A1(n12264), .A2(n12263), .ZN(n12270) );
  NAND3HSV3 U7094 ( .A1(n9672), .A2(n9671), .A3(n9670), .ZN(n15282) );
  INHSV2 U7095 ( .I(n8180), .ZN(n6032) );
  CLKNAND2HSV4 U7096 ( .A1(n13898), .A2(n9841), .ZN(n7440) );
  XNOR2HSV4 U7097 ( .A1(n7657), .A2(n7658), .ZN(n6012) );
  NAND2HSV4 U7098 ( .A1(n13762), .A2(n6721), .ZN(n9343) );
  CLKNAND2HSV4 U7099 ( .A1(n10050), .A2(n10062), .ZN(n10145) );
  XNOR2HSV4 U7100 ( .A1(n6013), .A2(n10103), .ZN(n10105) );
  XNOR2HSV4 U7101 ( .A1(n10102), .A2(n10104), .ZN(n6013) );
  NAND2HSV2 U7102 ( .A1(n14791), .A2(\pe11/pvq [5]), .ZN(n11716) );
  NAND2HSV4 U7103 ( .A1(n7015), .A2(n9400), .ZN(\pe9/ti_7[1] ) );
  NAND2HSV4 U7104 ( .A1(\pe9/ti_7[1] ), .A2(\pe9/got [5]), .ZN(n7014) );
  XNOR2HSV4 U7105 ( .A1(n12887), .A2(n12886), .ZN(n12889) );
  NOR2HSV4 U7106 ( .A1(n11203), .A2(n8726), .ZN(n11170) );
  XNOR2HSV4 U7107 ( .A1(n6913), .A2(n6915), .ZN(\pe6/poht [6]) );
  INHSV2 U7108 ( .I(n5970), .ZN(n7718) );
  CLKNAND2HSV3 U7109 ( .A1(n7105), .A2(n7103), .ZN(n10721) );
  CLKNAND2HSV4 U7110 ( .A1(\pe18/aot [8]), .A2(\pe18/bq[7] ), .ZN(n9142) );
  NAND2HSV2 U7111 ( .A1(n13752), .A2(\pe20/got [3]), .ZN(n8371) );
  NAND3HSV3 U7112 ( .A1(n6759), .A2(n6758), .A3(n6757), .ZN(n15181) );
  CLKNAND2HSV2 U7113 ( .A1(n14930), .A2(\pe14/got [1]), .ZN(n14436) );
  INOR2HSV4 U7114 ( .A1(\pe21/pvq [5]), .B1(n14537), .ZN(n10648) );
  DELHS1 U7115 ( .I(n15092), .Z(n6014) );
  AOI21HSV4 U7116 ( .A1(n10044), .A2(n10041), .B(n10043), .ZN(n10047) );
  CLKNAND2HSV2 U7117 ( .A1(n6015), .A2(n6544), .ZN(n6498) );
  CLKNAND2HSV2 U7118 ( .A1(n6541), .A2(n6542), .ZN(n6015) );
  CLKNAND2HSV2 U7119 ( .A1(n6540), .A2(\pe17/phq [2]), .ZN(n6541) );
  NAND2HSV4 U7120 ( .A1(\pe18/ti_1 ), .A2(\pe18/got [6]), .ZN(n6893) );
  XOR2HSV4 U7121 ( .A1(n6894), .A2(n6893), .Z(n6892) );
  CLKNAND2HSV4 U7122 ( .A1(\pe10/ti_1 ), .A2(\pe10/got [6]), .ZN(n10056) );
  CLKNAND2HSV4 U7123 ( .A1(n6016), .A2(n9715), .ZN(n13881) );
  CLKNHSV6 U7124 ( .I(n13881), .ZN(n6722) );
  INHSV2 U7125 ( .I(n9711), .ZN(n6017) );
  NAND2HSV4 U7126 ( .A1(n6100), .A2(n11175), .ZN(n11211) );
  NAND2HSV4 U7127 ( .A1(n7155), .A2(n7442), .ZN(n7159) );
  NAND2HSV4 U7128 ( .A1(n7037), .A2(n10217), .ZN(\pe3/ti_7[5] ) );
  INAND2HSV4 U7129 ( .A1(n11612), .B1(n11611), .ZN(n14963) );
  NAND2HSV2 U7130 ( .A1(n14963), .A2(\pe9/got [4]), .ZN(n11662) );
  NAND2HSV4 U7131 ( .A1(n7483), .A2(n8923), .ZN(n11612) );
  CLKNAND2HSV4 U7132 ( .A1(n6287), .A2(n6018), .ZN(n6654) );
  NAND2HSV4 U7133 ( .A1(n11177), .A2(n11178), .ZN(n6018) );
  BUFHSV6 U7134 ( .I(\pe20/ti_1 ), .Z(n13738) );
  NAND2HSV2 U7135 ( .A1(n9763), .A2(n9434), .ZN(n9448) );
  XNOR2HSV4 U7136 ( .A1(n6761), .A2(n6764), .ZN(n8607) );
  NAND2HSV4 U7137 ( .A1(n14872), .A2(\pe3/got [5]), .ZN(n6948) );
  AOI21HSV4 U7138 ( .A1(n9136), .A2(\pe17/ctrq ), .B(n6019), .ZN(n10416) );
  AOI21HSV4 U7139 ( .A1(\pe17/pvq [1]), .A2(\pe17/ctrq ), .B(\pe17/phq [1]), 
        .ZN(n6019) );
  CLKXOR2HSV4 U7140 ( .A1(n11767), .A2(n14381), .Z(n11720) );
  NAND2HSV4 U7141 ( .A1(n14709), .A2(\pe20/got [4]), .ZN(n6851) );
  XOR2HSV0 U7142 ( .A1(n7388), .A2(n6020), .Z(\pe13/poht [1]) );
  XOR2HSV2 U7143 ( .A1(n7386), .A2(n10028), .Z(n6020) );
  INHSV2 U7144 ( .I(n7410), .ZN(n6556) );
  NAND2HSV4 U7145 ( .A1(n7482), .A2(n11611), .ZN(n9754) );
  XNOR2HSV4 U7146 ( .A1(n6530), .A2(n6021), .ZN(n10356) );
  XOR3HSV2 U7147 ( .A1(n6529), .A2(n6528), .A3(n9557), .Z(n6021) );
  NAND3HSV3 U7148 ( .A1(n9167), .A2(n9166), .A3(\pe18/got [6]), .ZN(n9168) );
  OAI21HSV2 U7149 ( .A1(n8323), .A2(n8322), .B(n8324), .ZN(n8325) );
  NAND2HSV2 U7150 ( .A1(n8326), .A2(n8325), .ZN(n8327) );
  CLKXOR2HSV4 U7151 ( .A1(n9330), .A2(n9329), .Z(n9334) );
  CLKNAND2HSV2 U7152 ( .A1(\pe12/pvq [3]), .A2(\pe12/ctrq ), .ZN(n10724) );
  CLKNAND2HSV4 U7153 ( .A1(n14196), .A2(\pe8/got [3]), .ZN(n13532) );
  INOR2HSV4 U7154 ( .A1(n10583), .B1(n15083), .ZN(n6707) );
  XNOR2HSV1 U7155 ( .A1(n6024), .A2(n6022), .ZN(\pe10/poht [2]) );
  XNOR2HSV2 U7156 ( .A1(n7161), .A2(n6023), .ZN(n6022) );
  XNOR2HSV2 U7157 ( .A1(n7163), .A2(n7164), .ZN(n6023) );
  XNOR2HSV4 U7158 ( .A1(n12241), .A2(n6025), .ZN(n12243) );
  CLKNHSV2 U7159 ( .I(n12240), .ZN(n6025) );
  NAND2HSV4 U7160 ( .A1(\pe21/got [8]), .A2(\pe21/ti_1 ), .ZN(n9394) );
  CLKBUFHSV12 U7161 ( .I(n14960), .Z(n6026) );
  INHSV2 U7162 ( .I(n13775), .ZN(n13831) );
  NAND2HSV2 U7163 ( .A1(n11063), .A2(n8948), .ZN(n11065) );
  CLKNAND2HSV2 U7164 ( .A1(n8656), .A2(n8657), .ZN(n8658) );
  DELHS1 U7165 ( .I(\pe1/ti_7[2] ), .Z(n6027) );
  NAND2HSV2 U7166 ( .A1(n11772), .A2(n8505), .ZN(n8506) );
  CLKXOR2HSV2 U7167 ( .A1(n9691), .A2(n9690), .Z(n9695) );
  XNOR2HSV4 U7168 ( .A1(n12847), .A2(n12846), .ZN(n12848) );
  CLKXOR2HSV4 U7169 ( .A1(n11078), .A2(n11077), .Z(n11080) );
  XOR3HSV2 U7170 ( .A1(n6028), .A2(n12746), .A3(n12745), .Z(\pe12/poht [2]) );
  CLKNAND2HSV2 U7171 ( .A1(n15190), .A2(\pe12/got [5]), .ZN(n6028) );
  AOI21HSV4 U7172 ( .A1(n9992), .A2(n9955), .B(n6029), .ZN(n7470) );
  OAI21HSV4 U7173 ( .A1(n9992), .A2(n7471), .B(n7864), .ZN(n6029) );
  CLKNAND2HSV2 U7174 ( .A1(\pe2/aot [8]), .A2(\pe2/bq[4] ), .ZN(n9371) );
  XNOR2HSV2 U7175 ( .A1(n9371), .A2(n6505), .ZN(n9374) );
  NAND3HSV2 U7176 ( .A1(n6085), .A2(\pe2/aot [8]), .A3(\pe2/bq[6] ), .ZN(n6084) );
  AOI21HSV2 U7177 ( .A1(n14707), .A2(n14818), .B(ctro2), .ZN(n7309) );
  NAND2HSV4 U7178 ( .A1(n9925), .A2(n9924), .ZN(n9957) );
  CLKNAND2HSV2 U7179 ( .A1(n12512), .A2(n12511), .ZN(n14957) );
  CLKNAND2HSV4 U7180 ( .A1(\pe18/ti_1 ), .A2(\pe18/got [8]), .ZN(n9132) );
  NAND2HSV4 U7181 ( .A1(n7154), .A2(n8642), .ZN(n7157) );
  NOR2HSV8 U7182 ( .A1(n10040), .A2(n10112), .ZN(n14122) );
  NAND2HSV2 U7183 ( .A1(n10276), .A2(n10263), .ZN(n10268) );
  CLKNAND2HSV4 U7184 ( .A1(n15237), .A2(n8948), .ZN(n6489) );
  NAND2HSV4 U7185 ( .A1(n6489), .A2(n11113), .ZN(n15195) );
  CLKNAND2HSV8 U7186 ( .A1(n6158), .A2(n6157), .ZN(n15217) );
  OAI21HSV4 U7187 ( .A1(n15217), .A2(n13140), .B(n9174), .ZN(n9199) );
  CLKNAND2HSV2 U7188 ( .A1(n6032), .A2(n6031), .ZN(n6030) );
  CLKNHSV2 U7189 ( .I(n8181), .ZN(n6031) );
  NAND2HSV2 U7190 ( .A1(n15068), .A2(\pe9/got [3]), .ZN(n9762) );
  INHSV4 U7191 ( .I(n11122), .ZN(n8085) );
  CLKNAND2HSV8 U7192 ( .A1(n9923), .A2(n9922), .ZN(n13603) );
  CLKNAND2HSV2 U7193 ( .A1(n13603), .A2(\pe13/got [4]), .ZN(n7590) );
  INHSV6 U7194 ( .I(n14856), .ZN(n6763) );
  CLKNAND2HSV2 U7195 ( .A1(n14961), .A2(\pe13/got [3]), .ZN(n11970) );
  XNOR2HSV1 U7196 ( .A1(n11971), .A2(n11970), .ZN(\pe13/poht [5]) );
  NAND2HSV2 U7197 ( .A1(\pe7/bq[6] ), .A2(\pe7/aot [8]), .ZN(n6832) );
  CLKBUFHSV12 U7198 ( .I(n14874), .Z(n6033) );
  NAND2HSV4 U7199 ( .A1(n6141), .A2(n9455), .ZN(n15194) );
  BUFHSV6 U7200 ( .I(\pe11/ti_1 ), .Z(n13811) );
  CLKNAND2HSV4 U7201 ( .A1(n14546), .A2(\pe18/pvq [6]), .ZN(n9185) );
  XNOR2HSV4 U7202 ( .A1(n12306), .A2(n6034), .ZN(n12310) );
  XNOR2HSV4 U7203 ( .A1(n12304), .A2(n12305), .ZN(n6034) );
  CLKNAND2HSV2 U7204 ( .A1(n10187), .A2(n10186), .ZN(n7167) );
  CLKNAND2HSV8 U7205 ( .A1(n7642), .A2(n7641), .ZN(n15185) );
  CLKNAND2HSV4 U7206 ( .A1(n15185), .A2(n14066), .ZN(n11158) );
  INAND2HSV2 U7207 ( .A1(n14396), .B1(\pe11/got [3]), .ZN(n12467) );
  INAND2HSV2 U7208 ( .A1(n14396), .B1(\pe11/got [4]), .ZN(n12569) );
  XNOR2HSV4 U7209 ( .A1(n6035), .A2(n10657), .ZN(n10659) );
  XNOR2HSV4 U7210 ( .A1(n6036), .A2(n10654), .ZN(n6035) );
  XNOR2HSV4 U7211 ( .A1(n10655), .A2(n10656), .ZN(n6036) );
  NAND2HSV4 U7212 ( .A1(n7292), .A2(n7293), .ZN(n6797) );
  INHSV4 U7213 ( .I(\pe10/bq[5] ), .ZN(n10029) );
  CLKNHSV0 U7214 ( .I(n10029), .ZN(n8456) );
  XNOR2HSV4 U7215 ( .A1(n10749), .A2(n10748), .ZN(n10753) );
  XNOR2HSV4 U7216 ( .A1(n6037), .A2(n9428), .ZN(n9433) );
  XOR2HSV2 U7217 ( .A1(n9426), .A2(n9427), .Z(n6037) );
  NAND2HSV4 U7218 ( .A1(n12453), .A2(n12452), .ZN(n14965) );
  DELHS1 U7219 ( .I(\pe7/got [4]), .Z(n6038) );
  XNOR2HSV4 U7220 ( .A1(n9002), .A2(n9001), .ZN(n7880) );
  INAND2HSV2 U7221 ( .A1(n6041), .B1(n6040), .ZN(n7030) );
  CLKNHSV2 U7222 ( .I(n10581), .ZN(n6040) );
  CLKNAND2HSV2 U7223 ( .A1(n14933), .A2(n6042), .ZN(n6041) );
  CLKNHSV2 U7224 ( .I(n12596), .ZN(n6042) );
  CLKNAND2HSV2 U7225 ( .A1(n11306), .A2(n11305), .ZN(n11311) );
  OAI21HSV2 U7226 ( .A1(n8665), .A2(n8666), .B(n8667), .ZN(n8668) );
  CLKNAND2HSV2 U7227 ( .A1(n8669), .A2(n8668), .ZN(n8670) );
  NOR2HSV4 U7228 ( .A1(n9431), .A2(n9430), .ZN(n9432) );
  INAND3HSV4 U7229 ( .A1(n6045), .B1(n6044), .B2(n6043), .ZN(n14846) );
  CLKNHSV2 U7230 ( .I(n7182), .ZN(n6043) );
  CLKNAND2HSV2 U7231 ( .A1(n7183), .A2(n10307), .ZN(n6044) );
  NOR2HSV4 U7232 ( .A1(n7186), .A2(n7184), .ZN(n6045) );
  CLKNAND2HSV2 U7233 ( .A1(n13089), .A2(n6047), .ZN(n6046) );
  CLKNHSV2 U7234 ( .I(n11144), .ZN(n6047) );
  CLKNAND2HSV4 U7235 ( .A1(\pe4/got [6]), .A2(\pe4/ti_1 ), .ZN(n9616) );
  XNOR2HSV4 U7236 ( .A1(n9485), .A2(n6048), .ZN(n9486) );
  OAI21HSV4 U7237 ( .A1(n10409), .A2(n15177), .B(n9467), .ZN(n6048) );
  CLKNAND2HSV2 U7238 ( .A1(n6545), .A2(n7321), .ZN(n6547) );
  NOR2HSV4 U7239 ( .A1(n6147), .A2(n10397), .ZN(n10398) );
  INHSV4 U7240 ( .I(n14011), .ZN(n6386) );
  NAND2HSV4 U7241 ( .A1(n6719), .A2(n6386), .ZN(n12133) );
  CLKNAND2HSV2 U7242 ( .A1(\pe4/got [6]), .A2(\pe4/ti_1 ), .ZN(n9619) );
  NAND2HSV2 U7243 ( .A1(n14930), .A2(\pe14/got [5]), .ZN(n8774) );
  NAND2HSV2 U7244 ( .A1(n8774), .A2(n8773), .ZN(n8775) );
  NAND2HSV2 U7245 ( .A1(\pe12/aot [8]), .A2(\pe12/bq[5] ), .ZN(n10750) );
  CLKNAND2HSV2 U7246 ( .A1(n14948), .A2(\pe12/bq[3] ), .ZN(n11455) );
  NAND2HSV2 U7247 ( .A1(n11580), .A2(\pe8/got [8]), .ZN(n8337) );
  CLKNAND2HSV2 U7248 ( .A1(\pe16/aot [7]), .A2(\pe16/bq[4] ), .ZN(n11185) );
  CLKNAND2HSV8 U7249 ( .A1(n14702), .A2(\pe14/ti_7t [6]), .ZN(n11226) );
  CLKNAND2HSV4 U7250 ( .A1(\pe16/ti_7[1] ), .A2(\pe16/got [5]), .ZN(n6677) );
  NAND2HSV4 U7251 ( .A1(\pe12/bq[8] ), .A2(\pe12/aot [7]), .ZN(n10733) );
  OAI21HSV1 U7252 ( .A1(n8593), .A2(n8594), .B(n8595), .ZN(n8596) );
  INHSV4 U7253 ( .I(n6463), .ZN(n6462) );
  XNOR2HSV4 U7254 ( .A1(n7763), .A2(n7758), .ZN(\pe6/poht [1]) );
  OR2HSV4 U7255 ( .A1(n14396), .A2(n15146), .Z(n12449) );
  CLKXOR2HSV2 U7256 ( .A1(n12449), .A2(n6711), .Z(n12451) );
  CLKNAND2HSV4 U7257 ( .A1(n9324), .A2(\pe2/pvq [6]), .ZN(n9325) );
  CLKNAND2HSV2 U7258 ( .A1(n13738), .A2(\pe20/got [6]), .ZN(n9021) );
  CLKNHSV0 U7259 ( .I(n9021), .ZN(n7414) );
  CLKNAND2HSV4 U7260 ( .A1(\pe8/bq[7] ), .A2(\pe8/aot [8]), .ZN(n10475) );
  XNOR2HSV4 U7261 ( .A1(n10095), .A2(n10094), .ZN(n10103) );
  CLKNAND2HSV2 U7262 ( .A1(\pe3/ti_7[5] ), .A2(\pe3/got [1]), .ZN(n12969) );
  INHSV2 U7263 ( .I(n14396), .ZN(n6049) );
  CLKNAND2HSV2 U7264 ( .A1(n6049), .A2(\pe11/got [5]), .ZN(n14390) );
  AOI21HSV4 U7265 ( .A1(n9603), .A2(\pe11/ctrq ), .B(n9602), .ZN(n6957) );
  MOAI22HSV4 U7266 ( .A1(n13848), .A2(n9033), .B1(ctro20), .B2(\pe20/ti_7t [2]), .ZN(n9071) );
  AOI21HSV4 U7267 ( .A1(n13881), .A2(n13879), .B(n9714), .ZN(n9718) );
  NAND2HSV4 U7268 ( .A1(n14874), .A2(\pe10/got [5]), .ZN(n10084) );
  NAND2HSV2 U7269 ( .A1(n14963), .A2(\pe9/got [3]), .ZN(n11688) );
  CLKNAND2HSV4 U7270 ( .A1(n14348), .A2(\pe16/got [6]), .ZN(n13227) );
  CLKXOR2HSV4 U7271 ( .A1(n10147), .A2(n10146), .Z(n8334) );
  CLKNAND2HSV2 U7272 ( .A1(\pe20/got [5]), .A2(n13738), .ZN(n9048) );
  CLKXOR2HSV2 U7273 ( .A1(n9048), .A2(n9047), .Z(n7455) );
  XOR3HSV2 U7274 ( .A1(n11058), .A2(n11056), .A3(n11057), .Z(n8083) );
  OAI21HSV4 U7275 ( .A1(n9725), .A2(n9724), .B(n9723), .ZN(n9726) );
  CLKNAND2HSV4 U7276 ( .A1(n9170), .A2(n9171), .ZN(n11996) );
  NAND2HSV2 U7277 ( .A1(\pe18/got [4]), .A2(n11996), .ZN(n7898) );
  INHSV8 U7278 ( .I(\pe10/aot [8]), .ZN(n6144) );
  BUFHSV4 U7279 ( .I(\pe17/bq[8] ), .Z(n6456) );
  XNOR2HSV4 U7280 ( .A1(n13720), .A2(n13719), .ZN(\pe20/poht [1]) );
  NOR3HSV4 U7281 ( .A1(n6050), .A2(n13347), .A3(n8913), .ZN(n13351) );
  CLKNHSV2 U7282 ( .I(n13348), .ZN(n6050) );
  NAND3HSV4 U7283 ( .A1(n13344), .A2(n13804), .A3(n13343), .ZN(n13348) );
  XOR2HSV2 U7284 ( .A1(n6051), .A2(n14389), .Z(n14393) );
  XOR2HSV2 U7285 ( .A1(n14390), .A2(n14391), .Z(n6051) );
  OAI21HSV4 U7286 ( .A1(n11116), .A2(n11115), .B(n7986), .ZN(n7987) );
  XOR2HSV2 U7287 ( .A1(n10534), .A2(n6052), .Z(\pe13/poht [6]) );
  NAND2HSV4 U7288 ( .A1(n7066), .A2(n9459), .ZN(n10593) );
  OAI21HSV2 U7289 ( .A1(n8221), .A2(n8222), .B(n8223), .ZN(n8224) );
  NAND2HSV2 U7290 ( .A1(n8225), .A2(n8224), .ZN(n8226) );
  CLKNAND2HSV2 U7291 ( .A1(n13089), .A2(\pe14/got [2]), .ZN(n11232) );
  NAND2HSV2 U7292 ( .A1(n13604), .A2(n14750), .ZN(n8184) );
  NOR2HSV2 U7293 ( .A1(n10940), .A2(n10941), .ZN(n10966) );
  XNOR2HSV4 U7294 ( .A1(n11874), .A2(n11873), .ZN(n11875) );
  CLKXOR2HSV4 U7295 ( .A1(n7157), .A2(n11444), .Z(n15249) );
  NAND2HSV4 U7296 ( .A1(\pe7/ti_1 ), .A2(\pe7/got [8]), .ZN(n7620) );
  INHSV4 U7297 ( .I(n14701), .ZN(n14442) );
  CLKNAND2HSV2 U7298 ( .A1(n11924), .A2(\pe11/aot [4]), .ZN(n7924) );
  XOR2HSV0 U7299 ( .A1(n11716), .A2(n7924), .Z(n7928) );
  NAND2HSV4 U7300 ( .A1(n7147), .A2(n12280), .ZN(n15183) );
  INHSV4 U7301 ( .I(n11005), .ZN(n7038) );
  NAND2HSV4 U7302 ( .A1(n7538), .A2(n6053), .ZN(n11005) );
  INHSV2 U7303 ( .I(n7539), .ZN(n6053) );
  INHSV2 U7304 ( .I(n6054), .ZN(n7786) );
  CLKNAND2HSV2 U7305 ( .A1(n10868), .A2(n13801), .ZN(n6054) );
  XNOR2HSV4 U7306 ( .A1(n6851), .A2(n6055), .ZN(\pe20/poht [4]) );
  INHSV4 U7307 ( .I(n6056), .ZN(n6764) );
  NAND2HSV4 U7308 ( .A1(n8606), .A2(n6057), .ZN(n6056) );
  CLKNAND2HSV4 U7309 ( .A1(n6059), .A2(n6058), .ZN(n6057) );
  INHSV2 U7310 ( .I(n8605), .ZN(n6058) );
  INHSV2 U7311 ( .I(n8604), .ZN(n6059) );
  NAND2HSV4 U7312 ( .A1(n6621), .A2(n6620), .ZN(n7124) );
  INHSV4 U7313 ( .I(n11085), .ZN(n11086) );
  MUX2NHSV4 U7314 ( .I0(n6060), .I1(n12501), .S(n12500), .ZN(n12503) );
  INHSV2 U7315 ( .I(n6061), .ZN(n6060) );
  CLKNHSV2 U7316 ( .I(n12768), .ZN(n6062) );
  INHSV4 U7317 ( .I(n10178), .ZN(n10173) );
  NAND2HSV4 U7318 ( .A1(n6440), .A2(\pe17/got [3]), .ZN(n14329) );
  NAND2HSV4 U7319 ( .A1(n6063), .A2(\pe17/got [2]), .ZN(n14315) );
  NAND2HSV4 U7320 ( .A1(n6063), .A2(n14429), .ZN(n14431) );
  CLKNAND2HSV2 U7321 ( .A1(n13823), .A2(\pe4/aot [3]), .ZN(n9692) );
  XOR2HSV2 U7322 ( .A1(n6069), .A2(n6070), .Z(n10033) );
  NAND3HSV4 U7323 ( .A1(n8965), .A2(n8964), .A3(n8963), .ZN(n6932) );
  CLKNAND2HSV3 U7324 ( .A1(n8962), .A2(n8961), .ZN(n6933) );
  INHSV2 U7325 ( .I(n14707), .ZN(n6065) );
  NOR2HSV4 U7326 ( .A1(n6065), .A2(n6066), .ZN(n7307) );
  CLKNAND2HSV3 U7327 ( .A1(n8982), .A2(n7308), .ZN(n6066) );
  NAND3HSV4 U7328 ( .A1(n6067), .A2(n6064), .A3(n6068), .ZN(n8982) );
  INHSV2 U7329 ( .I(n8976), .ZN(n6067) );
  INHSV2 U7330 ( .I(n8977), .ZN(n6068) );
  NAND2HSV4 U7331 ( .A1(\pe10/got [5]), .A2(\pe10/ti_1 ), .ZN(n6069) );
  CLKNAND2HSV4 U7332 ( .A1(n6071), .A2(n6073), .ZN(n9459) );
  NAND3HSV4 U7333 ( .A1(n6072), .A2(n9456), .A3(n6075), .ZN(n6071) );
  CLKNHSV2 U7334 ( .I(n9060), .ZN(n6072) );
  OAI21HSV4 U7335 ( .A1(n9060), .A2(n9059), .B(n6074), .ZN(n6073) );
  CLKNHSV2 U7336 ( .I(n9456), .ZN(n6074) );
  CLKNHSV2 U7337 ( .I(n9059), .ZN(n6075) );
  INHSV2 U7338 ( .I(n6076), .ZN(n6512) );
  CLKNAND2HSV2 U7339 ( .A1(n12260), .A2(n11691), .ZN(n6076) );
  XNOR2HSV4 U7340 ( .A1(n6078), .A2(n6077), .ZN(n12260) );
  XNOR2HSV4 U7341 ( .A1(n8997), .A2(\pe9/phq [1]), .ZN(n6077) );
  XNOR2HSV4 U7342 ( .A1(n8996), .A2(n8995), .ZN(n6078) );
  CLKNAND2HSV3 U7343 ( .A1(\pe11/ti_1 ), .A2(\pe11/got [6]), .ZN(n6415) );
  CLKNHSV2 U7344 ( .I(n9364), .ZN(n9348) );
  INAND2HSV4 U7345 ( .A1(n10798), .B1(n6079), .ZN(n9364) );
  NOR2HSV4 U7346 ( .A1(n6080), .A2(n9358), .ZN(n6079) );
  CLKNHSV2 U7347 ( .I(n10797), .ZN(n6080) );
  CLKNAND2HSV2 U7348 ( .A1(n9345), .A2(n14818), .ZN(n10798) );
  INAND2HSV4 U7349 ( .A1(n10035), .B1(\pe10/pvq [7]), .ZN(n10093) );
  INAND2HSV4 U7350 ( .A1(n10035), .B1(\pe10/pvq [4]), .ZN(n10036) );
  INAND2HSV4 U7351 ( .A1(n10035), .B1(\pe10/pvq [3]), .ZN(n6222) );
  CLKNAND2HSV2 U7352 ( .A1(n6081), .A2(n7233), .ZN(n7230) );
  NOR2HSV2 U7353 ( .A1(n6081), .A2(n7233), .ZN(n7232) );
  NOR2HSV3 U7354 ( .A1(n10035), .A2(n6082), .ZN(n6081) );
  CLKNHSV4 U7355 ( .I(\pe10/pvq [2]), .ZN(n6082) );
  NAND2HSV2 U7356 ( .A1(n6084), .A2(n6083), .ZN(n6091) );
  XNOR2HSV4 U7357 ( .A1(n9347), .A2(n9346), .ZN(n8983) );
  XNOR2HSV4 U7358 ( .A1(n6087), .A2(n6086), .ZN(n9346) );
  XNOR2HSV4 U7359 ( .A1(n6091), .A2(n6088), .ZN(n6087) );
  CLKNHSV2 U7360 ( .I(n7100), .ZN(n6090) );
  NOR2HSV4 U7361 ( .A1(n8986), .A2(n8968), .ZN(n9347) );
  NOR2HSV4 U7362 ( .A1(n6093), .A2(n6092), .ZN(n8986) );
  CLKNAND2HSV2 U7363 ( .A1(n6932), .A2(n6931), .ZN(n6092) );
  CLKNHSV2 U7364 ( .I(n6933), .ZN(n6093) );
  CLKNAND2HSV2 U7365 ( .A1(n15264), .A2(n10924), .ZN(n7229) );
  XNOR2HSV4 U7366 ( .A1(n6097), .A2(n6094), .ZN(n15264) );
  AOI21HSV4 U7367 ( .A1(n6096), .A2(n6294), .B(n6095), .ZN(n6094) );
  AOI21HSV2 U7368 ( .A1(\pe10/ctrq ), .A2(\pe10/pvq [1]), .B(\pe10/phq [1]), 
        .ZN(n6095) );
  CLKNAND2HSV2 U7369 ( .A1(n6296), .A2(n7102), .ZN(n6098) );
  CLKNAND2HSV4 U7370 ( .A1(n6212), .A2(n6211), .ZN(n6100) );
  NAND3HSV4 U7371 ( .A1(n6100), .A2(n11175), .A3(n11220), .ZN(n6210) );
  CLKNAND2HSV2 U7372 ( .A1(\pe3/pvq [2]), .A2(\pe3/ctrq ), .ZN(n10181) );
  XNOR2HSV4 U7373 ( .A1(n11042), .A2(n6101), .ZN(n9074) );
  CLKNAND2HSV2 U7374 ( .A1(\pe14/aot [8]), .A2(\pe14/bq[6] ), .ZN(n6101) );
  CLKNAND2HSV2 U7375 ( .A1(\pe14/aot [6]), .A2(\pe14/bq[8] ), .ZN(n11042) );
  CLKNAND2HSV4 U7376 ( .A1(n10704), .A2(n7845), .ZN(n14080) );
  CLKNAND2HSV4 U7377 ( .A1(n12195), .A2(n7844), .ZN(n7845) );
  NOR2HSV8 U7378 ( .A1(n7409), .A2(n7846), .ZN(n10704) );
  NOR2HSV8 U7379 ( .A1(n10688), .A2(n7900), .ZN(n10674) );
  CLKNHSV2 U7380 ( .I(n11204), .ZN(n6383) );
  NAND3HSV4 U7381 ( .A1(n10705), .A2(n14080), .A3(n11207), .ZN(n11204) );
  XNOR2HSV4 U7382 ( .A1(n10670), .A2(n10669), .ZN(n10675) );
  CLKNAND2HSV3 U7383 ( .A1(\pe11/bq[6] ), .A2(\pe11/aot [8]), .ZN(n6102) );
  XNOR2HSV4 U7384 ( .A1(n6103), .A2(n6102), .ZN(n6411) );
  CLKNAND2HSV2 U7385 ( .A1(\pe11/bq[7] ), .A2(\pe11/aot [7]), .ZN(n6103) );
  OAI21HSV4 U7386 ( .A1(n7644), .A2(n6106), .B(n6104), .ZN(n6380) );
  NOR2HSV4 U7387 ( .A1(n11210), .A2(n7628), .ZN(n6104) );
  XNOR2HSV4 U7388 ( .A1(n6105), .A2(n6573), .ZN(n11210) );
  CLKNHSV2 U7389 ( .I(n11209), .ZN(n6106) );
  INAND2HSV4 U7390 ( .A1(n10794), .B1(n6107), .ZN(n11209) );
  NOR2HSV4 U7391 ( .A1(n14080), .A2(n8957), .ZN(n6107) );
  NAND2HSV2 U7392 ( .A1(n7476), .A2(n7475), .ZN(n6110) );
  NAND2HSV3 U7393 ( .A1(\pe14/got [6]), .A2(\pe14/ti_1 ), .ZN(n6111) );
  XNOR2HSV4 U7394 ( .A1(n6111), .A2(\pe14/phq [3]), .ZN(n9073) );
  XNOR2HSV4 U7395 ( .A1(n6112), .A2(n13717), .ZN(n13720) );
  XNOR2HSV4 U7396 ( .A1(n6113), .A2(n13716), .ZN(n6112) );
  CLKNAND2HSV2 U7397 ( .A1(n6731), .A2(\pe20/got [6]), .ZN(n6113) );
  CLKNAND2HSV2 U7398 ( .A1(n6795), .A2(n6794), .ZN(n6731) );
  CLKNAND2HSV2 U7399 ( .A1(n15208), .A2(n10412), .ZN(n10150) );
  OAI22HSV4 U7400 ( .A1(n15208), .A2(n13677), .B1(\pe20/ti_7t [5]), .B2(n8939), 
        .ZN(n13751) );
  XNOR2HSV4 U7401 ( .A1(n6775), .A2(n9459), .ZN(n15208) );
  CLKNAND2HSV2 U7402 ( .A1(n6117), .A2(n6114), .ZN(n9262) );
  CLKNAND2HSV2 U7403 ( .A1(n6119), .A2(n6115), .ZN(n6114) );
  CLKNHSV2 U7404 ( .I(n6118), .ZN(n6115) );
  NOR2HSV4 U7405 ( .A1(n6116), .A2(n6120), .ZN(n6119) );
  AOI21HSV4 U7406 ( .A1(n9265), .A2(n6118), .B(n9261), .ZN(n6117) );
  NOR2HSV4 U7407 ( .A1(n6773), .A2(n15095), .ZN(n6118) );
  NOR2HSV4 U7408 ( .A1(n6724), .A2(n9802), .ZN(n9265) );
  MUX2NHSV2 U7409 ( .I0(n8912), .I1(n9241), .S(n9240), .ZN(n6724) );
  AOI21HSV2 U7410 ( .A1(n9306), .A2(n6119), .B(n9267), .ZN(n9268) );
  CLKNHSV2 U7411 ( .I(n10799), .ZN(n6120) );
  CLKNHSV2 U7412 ( .I(n6121), .ZN(n13851) );
  XNOR2HSV4 U7413 ( .A1(n9127), .A2(n9126), .ZN(n6121) );
  AOI22HSV4 U7414 ( .A1(n9680), .A2(\pe4/ti_7t [2]), .B1(n9128), .B2(n6121), 
        .ZN(n6903) );
  CLKNAND2HSV0 U7415 ( .A1(\pe20/bq[7] ), .A2(\pe20/aot [6]), .ZN(n9045) );
  MUX2NHSV2 U7416 ( .I0(n13891), .I1(n6123), .S(n6122), .ZN(n6131) );
  CLKNHSV2 U7417 ( .I(n13893), .ZN(n6122) );
  CLKNHSV2 U7418 ( .I(n13890), .ZN(n6123) );
  CLKNHSV2 U7419 ( .I(n6125), .ZN(n6124) );
  NOR2HSV4 U7420 ( .A1(n13890), .A2(n13893), .ZN(n6125) );
  CLKNAND2HSV2 U7421 ( .A1(n13891), .A2(n13893), .ZN(n6126) );
  XNOR2HSV4 U7422 ( .A1(n6831), .A2(n8080), .ZN(n13893) );
  CLKNAND2HSV2 U7423 ( .A1(n12679), .A2(n12680), .ZN(n14446) );
  AOI22HSV4 U7424 ( .A1(\pe12/ti_7t [7]), .A2(n11471), .B1(n6130), .B2(n6127), 
        .ZN(n12680) );
  CLKNHSV2 U7425 ( .I(n6128), .ZN(n6127) );
  CLKNAND2HSV2 U7426 ( .A1(n15248), .A2(n6129), .ZN(n6128) );
  CLKNHSV2 U7427 ( .I(n11470), .ZN(n6129) );
  CLKNAND2HSV2 U7428 ( .A1(n6132), .A2(n6131), .ZN(n12679) );
  CLKNHSV2 U7429 ( .I(n6135), .ZN(n6134) );
  NOR2HSV4 U7430 ( .A1(n7494), .A2(n7492), .ZN(n6135) );
  CLKNHSV2 U7431 ( .I(n9535), .ZN(n8035) );
  XNOR2HSV4 U7432 ( .A1(n9535), .A2(n6136), .ZN(n9287) );
  XOR2HSV2 U7433 ( .A1(n9534), .A2(n6137), .Z(n6136) );
  CLKNAND2HSV2 U7434 ( .A1(n11951), .A2(n7801), .ZN(n6137) );
  NOR2HSV4 U7435 ( .A1(n6138), .A2(n7798), .ZN(n11951) );
  XNOR2HSV4 U7436 ( .A1(n6140), .A2(n6139), .ZN(n9534) );
  XNOR2HSV4 U7437 ( .A1(n9283), .A2(n9282), .ZN(n6140) );
  AOI21HSV4 U7438 ( .A1(n7468), .A2(n9308), .B(n7466), .ZN(n9535) );
  CLKNAND2HSV2 U7439 ( .A1(n15194), .A2(\pe18/got [5]), .ZN(n12000) );
  CLKNAND2HSV2 U7440 ( .A1(n15194), .A2(\pe18/got [4]), .ZN(n13171) );
  CLKNAND2HSV2 U7441 ( .A1(n15194), .A2(\pe18/got [1]), .ZN(n14659) );
  CLKNAND2HSV2 U7442 ( .A1(n15194), .A2(\pe18/got [3]), .ZN(n14641) );
  CLKNAND2HSV0 U7443 ( .A1(n15194), .A2(\pe18/got [2]), .ZN(n13365) );
  CLKNAND2HSV2 U7444 ( .A1(n15218), .A2(n13145), .ZN(n6141) );
  NOR2HSV3 U7445 ( .A1(n6143), .A2(n6142), .ZN(n8958) );
  CLKNHSV4 U7446 ( .I(\pe2/pvq [1]), .ZN(n6142) );
  CLKNAND2HSV3 U7447 ( .A1(\pe2/got [8]), .A2(\pe2/ti_1 ), .ZN(n6143) );
  NOR2HSV8 U7448 ( .A1(n6145), .A2(n6144), .ZN(n6298) );
  CLKNHSV4 U7449 ( .I(\pe10/bq[8] ), .ZN(n6145) );
  CLKNAND2HSV2 U7450 ( .A1(n15068), .A2(\pe9/got [5]), .ZN(n11665) );
  CLKNAND2HSV2 U7451 ( .A1(n15068), .A2(\pe9/got [2]), .ZN(n11643) );
  CLKNAND2HSV2 U7452 ( .A1(n15068), .A2(\pe9/got [4]), .ZN(n11689) );
  CLKNAND2HSV2 U7453 ( .A1(n15068), .A2(n9420), .ZN(n14583) );
  CLKNAND2HSV2 U7454 ( .A1(n15068), .A2(n9449), .ZN(n7367) );
  NOR2HSV8 U7455 ( .A1(n11692), .A2(n11668), .ZN(n15068) );
  CLKNAND2HSV2 U7456 ( .A1(\pe21/ti_7[1] ), .A2(\pe21/got [5]), .ZN(n10657) );
  CLKNAND2HSV2 U7457 ( .A1(n6146), .A2(n10385), .ZN(\pe21/ti_7[1] ) );
  CLKNAND2HSV2 U7458 ( .A1(n11781), .A2(n9398), .ZN(n6146) );
  XNOR2HSV4 U7459 ( .A1(n10371), .A2(n10370), .ZN(n11781) );
  CLKNAND2HSV2 U7460 ( .A1(\pe20/bq[6] ), .A2(\pe20/aot [7]), .ZN(n9043) );
  NOR2HSV8 U7461 ( .A1(n6147), .A2(n8455), .ZN(n10413) );
  NOR2HSV8 U7462 ( .A1(n11781), .A2(n10386), .ZN(n6147) );
  XNOR2HSV4 U7463 ( .A1(n6149), .A2(n6148), .ZN(n10417) );
  CLKNAND2HSV2 U7464 ( .A1(\pe17/got [8]), .A2(\pe17/ti_1 ), .ZN(n6149) );
  CLKNAND2HSV2 U7465 ( .A1(n9947), .A2(n6150), .ZN(n7599) );
  NOR2HSV8 U7466 ( .A1(n6150), .A2(n9947), .ZN(n9952) );
  NOR2HSV8 U7467 ( .A1(n9946), .A2(n6151), .ZN(n6150) );
  CLKXOR2HSV4 U7468 ( .A1(n6152), .A2(\pe2/phq [1]), .Z(n8964) );
  CLKNAND2HSV3 U7469 ( .A1(\pe2/aot [8]), .A2(\pe2/bq[8] ), .ZN(n6152) );
  CLKNAND2HSV3 U7470 ( .A1(n6153), .A2(n6154), .ZN(n6155) );
  CLKNAND2HSV3 U7471 ( .A1(n9154), .A2(n9217), .ZN(n6153) );
  CLKNHSV2 U7472 ( .I(n6156), .ZN(n6154) );
  CLKNAND2HSV2 U7473 ( .A1(n9154), .A2(n9217), .ZN(n6164) );
  INAND2HSV4 U7474 ( .A1(n6159), .B1(n6155), .ZN(n6158) );
  CLKNHSV2 U7475 ( .I(n6163), .ZN(n6156) );
  XNOR2HSV4 U7476 ( .A1(n9173), .A2(n9172), .ZN(n6159) );
  NAND3HSV4 U7477 ( .A1(n6164), .A2(n6159), .A3(n6163), .ZN(n6157) );
  NAND2HSV8 U7478 ( .A1(n15217), .A2(n13343), .ZN(n11977) );
  OAI21HSV4 U7479 ( .A1(n11977), .A2(n13139), .B(n6160), .ZN(n9219) );
  AOI21HSV4 U7480 ( .A1(n6162), .A2(n13139), .B(n6161), .ZN(n6160) );
  CLKNHSV2 U7481 ( .I(n9218), .ZN(n6161) );
  NOR2HSV4 U7482 ( .A1(n15217), .A2(n13342), .ZN(n6162) );
  CLKNHSV2 U7483 ( .I(n9153), .ZN(n6163) );
  XNOR2HSV4 U7484 ( .A1(n6166), .A2(n6165), .ZN(n13139) );
  XNOR2HSV4 U7485 ( .A1(n9216), .A2(n9215), .ZN(n6165) );
  OAI21HSV4 U7486 ( .A1(n15218), .A2(n13342), .B(n7833), .ZN(n6166) );
  XNOR2HSV4 U7487 ( .A1(n6835), .A2(n9193), .ZN(n15218) );
  NAND2HSV2 U7488 ( .A1(\pe17/aot [7]), .A2(\pe17/bq[7] ), .ZN(n6167) );
  CLKNAND2HSV2 U7489 ( .A1(n6167), .A2(\pe17/phq [3]), .ZN(n6168) );
  CLKNAND2HSV4 U7490 ( .A1(\pe17/got [5]), .A2(\pe17/ti_1 ), .ZN(n8462) );
  CLKNAND2HSV2 U7491 ( .A1(\pe9/ti_1 ), .A2(\pe9/got [6]), .ZN(n6169) );
  CLKBUFHSV2 U7492 ( .I(n6171), .Z(n6170) );
  BUFHSV8 U7493 ( .I(n7160), .Z(n6171) );
  NAND2HSV3 U7494 ( .A1(n7160), .A2(n11242), .ZN(n7749) );
  CLKNAND2HSV4 U7495 ( .A1(n11238), .A2(n11237), .ZN(n7160) );
  CLKNAND2HSV2 U7496 ( .A1(n7160), .A2(n8954), .ZN(n12903) );
  CLKNAND2HSV2 U7497 ( .A1(n6171), .A2(n6172), .ZN(n6318) );
  CLKNHSV2 U7498 ( .I(n6774), .ZN(n6172) );
  CLKNAND2HSV2 U7499 ( .A1(n6170), .A2(n14818), .ZN(n13887) );
  NAND2HSV3 U7500 ( .A1(n6174), .A2(n12340), .ZN(n12387) );
  CLKNAND2HSV2 U7501 ( .A1(n6174), .A2(n6695), .ZN(n13316) );
  CLKNAND2HSV2 U7502 ( .A1(n6174), .A2(n6173), .ZN(n14867) );
  CLKNHSV2 U7503 ( .I(n6359), .ZN(n6173) );
  CLKNAND2HSV4 U7504 ( .A1(n15073), .A2(n9541), .ZN(n6174) );
  XNOR2HSV4 U7505 ( .A1(n6176), .A2(n6175), .ZN(n9986) );
  CLKNAND2HSV2 U7506 ( .A1(\pe13/ti_7[4] ), .A2(\pe13/got [6]), .ZN(n6175) );
  CLKNAND2HSV3 U7507 ( .A1(n9932), .A2(n9931), .ZN(\pe13/ti_7[4] ) );
  AOI21HSV4 U7508 ( .A1(n9952), .A2(n9881), .B(n9951), .ZN(n9932) );
  XNOR2HSV4 U7509 ( .A1(n9976), .A2(n6177), .ZN(n6176) );
  XNOR2HSV4 U7510 ( .A1(n6178), .A2(n9975), .ZN(n6177) );
  XNOR2HSV4 U7511 ( .A1(n9959), .A2(n6179), .ZN(n6178) );
  CLKNHSV2 U7512 ( .I(n9958), .ZN(n6179) );
  CLKNHSV2 U7513 ( .I(\pe17/ti_7[1] ), .ZN(n14401) );
  CLKNAND2HSV2 U7514 ( .A1(\pe17/ti_7[1] ), .A2(\pe17/got [5]), .ZN(n6523) );
  CLKNAND2HSV0 U7515 ( .A1(\pe17/ti_7[1] ), .A2(\pe17/got [4]), .ZN(n12027) );
  CLKNAND2HSV2 U7516 ( .A1(\pe17/ti_7[1] ), .A2(\pe17/got [1]), .ZN(n14343) );
  XOR2HSV2 U7517 ( .A1(n6180), .A2(n13841), .Z(n15224) );
  CLKNAND2HSV2 U7518 ( .A1(\pe17/ti_7[1] ), .A2(\pe17/got [8]), .ZN(n6180) );
  CLKNAND2HSV4 U7519 ( .A1(n6444), .A2(n10526), .ZN(\pe17/ti_7[1] ) );
  BUFHSV8 U7520 ( .I(n12602), .Z(n6181) );
  CLKNAND2HSV4 U7521 ( .A1(n12590), .A2(n9719), .ZN(n12602) );
  CLKNAND2HSV3 U7522 ( .A1(n9718), .A2(n9717), .ZN(n12590) );
  CLKNAND2HSV0 U7523 ( .A1(n6181), .A2(\pe4/got [1]), .ZN(n8152) );
  NOR2HSV4 U7524 ( .A1(n10875), .A2(n10874), .ZN(n6182) );
  XNOR2HSV4 U7525 ( .A1(n7140), .A2(n10858), .ZN(n10875) );
  NOR2HSV8 U7526 ( .A1(n6182), .A2(n6443), .ZN(\pe21/ti_7[5] ) );
  CLKNAND2HSV0 U7527 ( .A1(\pe21/ti_7[5] ), .A2(\pe21/got [5]), .ZN(n8067) );
  CLKNAND2HSV2 U7528 ( .A1(n6183), .A2(n9013), .ZN(n9015) );
  CLKNAND2HSV1 U7529 ( .A1(\pe20/bq[7] ), .A2(\pe20/aot [7]), .ZN(n6183) );
  NAND3HSV4 U7530 ( .A1(n6187), .A2(n6186), .A3(n6184), .ZN(n6594) );
  INAND2HSV4 U7531 ( .A1(n6185), .B1(n6587), .ZN(n6184) );
  CLKNHSV2 U7532 ( .I(n6189), .ZN(n6185) );
  CLKNAND2HSV2 U7533 ( .A1(n6192), .A2(n6587), .ZN(n6186) );
  CLKNAND2HSV2 U7534 ( .A1(n6191), .A2(n6188), .ZN(n6187) );
  NOR2HSV4 U7535 ( .A1(n6190), .A2(n6189), .ZN(n6188) );
  AOI21HSV4 U7536 ( .A1(n14219), .A2(\pe19/got [3]), .B(n14220), .ZN(n6189) );
  CLKNHSV2 U7537 ( .I(n8513), .ZN(n6190) );
  CLKNHSV2 U7538 ( .I(n6192), .ZN(n6191) );
  NOR2HSV4 U7539 ( .A1(n14222), .A2(n6193), .ZN(n6192) );
  CLKNHSV2 U7540 ( .I(n6588), .ZN(n6193) );
  NAND3HSV4 U7541 ( .A1(n6197), .A2(n6195), .A3(n6194), .ZN(n6201) );
  CLKNAND2HSV2 U7542 ( .A1(n6199), .A2(n6202), .ZN(n6194) );
  CLKNAND2HSV2 U7543 ( .A1(n6196), .A2(n8247), .ZN(n6195) );
  NOR2HSV4 U7544 ( .A1(n6199), .A2(n6202), .ZN(n6196) );
  CLKNAND2HSV2 U7545 ( .A1(n6198), .A2(n6202), .ZN(n6197) );
  CLKNHSV2 U7546 ( .I(n8247), .ZN(n6198) );
  NOR2HSV4 U7547 ( .A1(n8245), .A2(n8246), .ZN(n6199) );
  CLKNAND2HSV3 U7548 ( .A1(n13535), .A2(n13533), .ZN(n15182) );
  CLKNAND2HSV2 U7549 ( .A1(n8249), .A2(n8248), .ZN(n8250) );
  XNOR2HSV4 U7550 ( .A1(n6201), .A2(n6200), .ZN(n8248) );
  CLKNAND2HSV2 U7551 ( .A1(n15182), .A2(\pe8/got [5]), .ZN(n6200) );
  CLKNHSV2 U7552 ( .I(n14212), .ZN(n6202) );
  OAI21HSV4 U7553 ( .A1(n15076), .A2(n14190), .B(n8242), .ZN(n8249) );
  XNOR2HSV4 U7554 ( .A1(n6203), .A2(n7175), .ZN(n15076) );
  CLKNHSV2 U7555 ( .I(n7177), .ZN(n6203) );
  CLKNAND2HSV2 U7556 ( .A1(\pe12/ctrq ), .A2(\pe12/pvq [2]), .ZN(n10738) );
  CLKNAND2HSV2 U7557 ( .A1(\pe2/ti_7[1] ), .A2(n6721), .ZN(n9377) );
  NAND2HSV4 U7558 ( .A1(n14736), .A2(n14066), .ZN(n6514) );
  CLKXOR2HSV2 U7559 ( .A1(n9334), .A2(n9333), .Z(n9335) );
  NAND2HSV4 U7560 ( .A1(\pe6/got [8]), .A2(\pe6/ti_1 ), .ZN(n9231) );
  MUX2NHSV4 U7561 ( .I0(\pe15/phq [6]), .I1(n8725), .S(n7463), .ZN(n11383) );
  NAND2HSV2 U7562 ( .A1(n14826), .A2(n9149), .ZN(n9150) );
  CLKNAND2HSV4 U7563 ( .A1(n14511), .A2(\pe18/aot [7]), .ZN(n9143) );
  XNOR2HSV4 U7564 ( .A1(n7406), .A2(n8122), .ZN(n10888) );
  NAND2HSV2 U7565 ( .A1(n14965), .A2(\pe11/got [4]), .ZN(n8225) );
  NAND2HSV2 U7566 ( .A1(n10868), .A2(n10864), .ZN(n10867) );
  NAND2HSV2 U7567 ( .A1(\pe15/aot [3]), .A2(\pe15/bq[8] ), .ZN(n11380) );
  NAND2HSV4 U7568 ( .A1(n9057), .A2(n11880), .ZN(n7417) );
  CLKNAND2HSV2 U7569 ( .A1(\pe2/got [8]), .A2(\pe2/ti_1 ), .ZN(n8960) );
  INHSV8 U7570 ( .I(\pe2/ctrq ), .ZN(n13766) );
  CLKXOR2HSV4 U7571 ( .A1(n10724), .A2(n10723), .Z(n6293) );
  CLKNAND2HSV2 U7572 ( .A1(n8952), .A2(\pe10/got [3]), .ZN(n6822) );
  NAND2HSV4 U7573 ( .A1(\pe14/ti_1 ), .A2(\pe14/got [8]), .ZN(n6742) );
  NAND2HSV4 U7574 ( .A1(n14348), .A2(n14292), .ZN(n14295) );
  NAND2HSV2 U7575 ( .A1(\pe11/got [3]), .A2(n14965), .ZN(n8669) );
  INAND2HSV4 U7576 ( .A1(n12538), .B1(n12537), .ZN(n13236) );
  NAND2HSV2 U7577 ( .A1(n13236), .A2(\pe15/got [3]), .ZN(n8585) );
  NAND2HSV4 U7578 ( .A1(n12386), .A2(n12385), .ZN(n13315) );
  NAND2HSV4 U7579 ( .A1(\pe19/got [8]), .A2(\pe19/ti_1 ), .ZN(n7896) );
  XNOR2HSV2 U7580 ( .A1(n11665), .A2(n11664), .ZN(n7879) );
  NAND2HSV2 U7581 ( .A1(\pe3/bq[7] ), .A2(\pe3/aot [8]), .ZN(n10182) );
  CLKNAND2HSV4 U7582 ( .A1(n13587), .A2(n14750), .ZN(n9999) );
  CLKNAND2HSV2 U7583 ( .A1(\pe18/got [7]), .A2(\pe18/ti_1 ), .ZN(n9145) );
  CLKNAND2HSV4 U7584 ( .A1(n11969), .A2(n11968), .ZN(n14961) );
  OAI21HSV2 U7585 ( .A1(n9533), .A2(n9797), .B(n8036), .ZN(n8037) );
  NAND2HSV4 U7586 ( .A1(n7079), .A2(n10422), .ZN(n6364) );
  INHSV2 U7587 ( .I(n7674), .ZN(n11899) );
  OA22HSV4 U7588 ( .A1(n11705), .A2(n10865), .B1(n7778), .B2(n7777), .Z(n6736)
         );
  INHSV2 U7589 ( .I(n9165), .ZN(n9167) );
  INHSV4 U7590 ( .I(n7500), .ZN(n15258) );
  CLKNAND2HSV2 U7591 ( .A1(n13089), .A2(\pe14/got [3]), .ZN(n11282) );
  CLKNAND2HSV8 U7592 ( .A1(n10401), .A2(n10400), .ZN(n10825) );
  CLKXOR2HSV4 U7593 ( .A1(n11998), .A2(n11997), .Z(n11999) );
  CLKNAND2HSV2 U7594 ( .A1(n8426), .A2(n8425), .ZN(n8427) );
  NAND2HSV2 U7595 ( .A1(n14855), .A2(\pe14/got [4]), .ZN(n8771) );
  XOR2HSV4 U7596 ( .A1(n7174), .A2(n7172), .Z(n7171) );
  CLKNAND2HSV4 U7597 ( .A1(\pe3/aot [8]), .A2(\pe3/bq[8] ), .ZN(n10163) );
  CLKNAND2HSV2 U7598 ( .A1(\pe12/bq[7] ), .A2(\pe12/aot [7]), .ZN(n10722) );
  NAND2HSV2 U7599 ( .A1(n14951), .A2(\pe10/bq[2] ), .ZN(n10092) );
  NAND2HSV4 U7600 ( .A1(\pe3/bq[6] ), .A2(\pe3/aot [8]), .ZN(n10151) );
  NAND2HSV4 U7601 ( .A1(n11398), .A2(n11397), .ZN(n11404) );
  CLKNAND2HSV2 U7602 ( .A1(n6004), .A2(\pe16/aot [8]), .ZN(n7982) );
  NAND2HSV4 U7603 ( .A1(n6498), .A2(n6496), .ZN(n6500) );
  CLKNAND2HSV4 U7604 ( .A1(n7362), .A2(n11782), .ZN(n12248) );
  INHSV4 U7605 ( .I(n6926), .ZN(n6925) );
  NAND2HSV4 U7606 ( .A1(n7795), .A2(n6925), .ZN(n10122) );
  XNOR2HSV4 U7607 ( .A1(n11273), .A2(n11272), .ZN(\pe2/poht [5]) );
  INHSV4 U7608 ( .I(n9828), .ZN(n13057) );
  XNOR2HSV4 U7609 ( .A1(n9468), .A2(\pe20/phq [6]), .ZN(n9470) );
  MAOI22HSV2 U7610 ( .A1(n8265), .A2(n12146), .B1(n7580), .B2(n7579), .ZN(
        n7578) );
  XOR2HSV4 U7611 ( .A1(n7719), .A2(n7715), .Z(n10997) );
  INHSV4 U7612 ( .I(n10997), .ZN(n12500) );
  CLKNAND2HSV2 U7613 ( .A1(n11854), .A2(\pe20/got [5]), .ZN(n11874) );
  INHSV4 U7614 ( .I(n6330), .ZN(n6333) );
  NAND2HSV4 U7615 ( .A1(\pe17/bq[7] ), .A2(\pe17/aot [6]), .ZN(n8463) );
  CLKXOR2HSV4 U7616 ( .A1(n12123), .A2(n12122), .Z(n12124) );
  NAND2HSV2 U7617 ( .A1(n14061), .A2(\pe2/got [4]), .ZN(n12919) );
  NAND2HSV2 U7618 ( .A1(\pe10/phq [1]), .A2(\pe10/ctrq ), .ZN(n6295) );
  CLKNAND2HSV2 U7619 ( .A1(n6874), .A2(\pe6/got [4]), .ZN(n7074) );
  NOR2HSV2 U7620 ( .A1(n7683), .A2(ctro11), .ZN(n11766) );
  CLKNAND2HSV4 U7621 ( .A1(\pe7/got [7]), .A2(\pe7/ti_1 ), .ZN(n10447) );
  NAND2HSV2 U7622 ( .A1(\pe3/aot [6]), .A2(\pe3/bq[8] ), .ZN(n8108) );
  MUX2NHSV2 U7623 ( .I0(\pe3/phq [3]), .I1(n8107), .S(n8108), .ZN(n10154) );
  CLKNAND2HSV2 U7624 ( .A1(n14949), .A2(\pe17/bq[2] ), .ZN(n12114) );
  CLKNAND2HSV4 U7625 ( .A1(n14708), .A2(\pe15/got [5]), .ZN(n14613) );
  NAND2HSV2 U7626 ( .A1(n6706), .A2(\pe4/got [1]), .ZN(n6756) );
  NAND2HSV4 U7627 ( .A1(n13186), .A2(n14681), .ZN(n14695) );
  CLKNAND2HSV4 U7628 ( .A1(n9386), .A2(n9385), .ZN(n9390) );
  XNOR2HSV4 U7629 ( .A1(n13371), .A2(n13370), .ZN(\pe18/poht [2]) );
  INHSV4 U7630 ( .I(n11838), .ZN(n14791) );
  NOR2HSV4 U7631 ( .A1(n6204), .A2(n12010), .ZN(n8408) );
  CLKNAND2HSV4 U7632 ( .A1(n6869), .A2(n6205), .ZN(n9171) );
  CLKNHSV3 U7633 ( .I(n9152), .ZN(n6205) );
  XNOR2HSV1 U7634 ( .A1(n6206), .A2(n9152), .ZN(n15219) );
  CLKNHSV2 U7635 ( .I(n8712), .ZN(n6206) );
  CLKNAND2HSV4 U7636 ( .A1(n11774), .A2(n10402), .ZN(n10836) );
  CLKBUFHSV2 U7637 ( .I(n11774), .Z(n6208) );
  CLKNAND2HSV0 U7638 ( .A1(n11774), .A2(n10641), .ZN(n10643) );
  CLKNAND2HSV3 U7639 ( .A1(n6209), .A2(\pe9/got [1]), .ZN(n9758) );
  CLKNAND2HSV4 U7640 ( .A1(n9748), .A2(n9747), .ZN(n13910) );
  INHSV2 U7641 ( .I(n13910), .ZN(n11674) );
  INHSV2 U7642 ( .I(n6210), .ZN(n11180) );
  CLKNHSV2 U7643 ( .I(n6216), .ZN(n6212) );
  XNOR2HSV4 U7644 ( .A1(n6217), .A2(n6218), .ZN(n6216) );
  CLKNAND2HSV2 U7645 ( .A1(n6216), .A2(n6213), .ZN(n11175) );
  CLKNAND2HSV2 U7646 ( .A1(n7523), .A2(n10795), .ZN(n6215) );
  CLKNAND2HSV2 U7647 ( .A1(n14958), .A2(\pe16/got [6]), .ZN(n6217) );
  XNOR2HSV4 U7648 ( .A1(n6678), .A2(n6677), .ZN(n6218) );
  XNOR2HSV4 U7649 ( .A1(n6220), .A2(n6219), .ZN(n10069) );
  OAI21HSV4 U7650 ( .A1(n15264), .A2(n10073), .B(n10059), .ZN(n6219) );
  XNOR2HSV4 U7651 ( .A1(n6223), .A2(n6221), .ZN(n6220) );
  XNOR2HSV4 U7652 ( .A1(n6222), .A2(n10057), .ZN(n6221) );
  XNOR2HSV4 U7653 ( .A1(n6225), .A2(n6224), .ZN(n6223) );
  XNOR2HSV4 U7654 ( .A1(n10056), .A2(\pe10/phq [3]), .ZN(n6224) );
  CLKNAND2HSV3 U7655 ( .A1(n6227), .A2(n6226), .ZN(n6234) );
  NAND3HSV3 U7656 ( .A1(\pe9/phq [2]), .A2(\pe9/got [7]), .A3(\pe9/ti_1 ), 
        .ZN(n6226) );
  CLKNAND2HSV3 U7657 ( .A1(n8999), .A2(n8998), .ZN(n6227) );
  NAND2HSV2 U7658 ( .A1(\pe9/bq[7] ), .A2(\pe9/aot [8]), .ZN(n6230) );
  XNOR2HSV4 U7659 ( .A1(n9002), .A2(n9000), .ZN(n6513) );
  XNOR2HSV4 U7660 ( .A1(n6229), .A2(n6228), .ZN(n9000) );
  CLKNAND2HSV2 U7661 ( .A1(\pe9/pvq [2]), .A2(\pe9/ctrq ), .ZN(n6228) );
  CLKNHSV2 U7662 ( .I(n6230), .ZN(n6229) );
  XNOR2HSV4 U7663 ( .A1(n6234), .A2(n6231), .ZN(n9002) );
  NOR2HSV4 U7664 ( .A1(n6233), .A2(n6232), .ZN(n6231) );
  CLKNHSV2 U7665 ( .I(\pe9/bq[8] ), .ZN(n6232) );
  CLKNHSV2 U7666 ( .I(\pe9/aot [7]), .ZN(n6233) );
  XNOR2HSV4 U7667 ( .A1(n6235), .A2(n6246), .ZN(n8992) );
  XNOR2HSV4 U7668 ( .A1(n6237), .A2(n6236), .ZN(n6235) );
  XNOR2HSV4 U7669 ( .A1(n6238), .A2(n8988), .ZN(n6236) );
  CLKNAND2HSV2 U7670 ( .A1(n6240), .A2(n6239), .ZN(n6237) );
  XNOR2HSV4 U7671 ( .A1(n6300), .A2(n8989), .ZN(n6238) );
  NAND3HSV4 U7672 ( .A1(n6241), .A2(n8554), .A3(n6243), .ZN(n6239) );
  XNOR2HSV4 U7673 ( .A1(n6242), .A2(n6299), .ZN(n6241) );
  CLKNHSV2 U7674 ( .I(n8555), .ZN(n6242) );
  CLKNAND2HSV2 U7675 ( .A1(n6245), .A2(n6244), .ZN(n6243) );
  CLKNHSV2 U7676 ( .I(\pe2/phq [4]), .ZN(n6244) );
  CLKNHSV2 U7677 ( .I(n8553), .ZN(n6245) );
  NOR2HSV4 U7678 ( .A1(n8986), .A2(n6247), .ZN(n6246) );
  CLKNAND2HSV2 U7679 ( .A1(n8987), .A2(n8954), .ZN(n6247) );
  OAI21HSV4 U7680 ( .A1(n7175), .A2(n6252), .B(n6248), .ZN(n15091) );
  AOI21HSV4 U7681 ( .A1(n6250), .A2(n7175), .B(n6249), .ZN(n6248) );
  CLKNHSV2 U7682 ( .I(n12371), .ZN(n6249) );
  NOR2HSV4 U7683 ( .A1(n7177), .A2(n6251), .ZN(n6250) );
  CLKNHSV2 U7684 ( .I(n6253), .ZN(n6251) );
  CLKNAND2HSV2 U7685 ( .A1(n7180), .A2(n6253), .ZN(n6252) );
  XNOR2HSV4 U7686 ( .A1(n7179), .A2(n7178), .ZN(n7175) );
  CLKNHSV2 U7687 ( .I(n7176), .ZN(n6253) );
  NOR2HSV4 U7688 ( .A1(n6863), .A2(n7181), .ZN(n7177) );
  NAND2HSV2 U7689 ( .A1(n11408), .A2(n6254), .ZN(n7370) );
  XNOR2HSV4 U7690 ( .A1(n11359), .A2(n11360), .ZN(n6254) );
  INHSV2 U7691 ( .I(n6254), .ZN(n7369) );
  XNOR2HSV4 U7692 ( .A1(n11408), .A2(n6254), .ZN(n11410) );
  XNOR2HSV4 U7693 ( .A1(n9915), .A2(n6255), .ZN(n9919) );
  XNOR2HSV4 U7694 ( .A1(n6258), .A2(n6256), .ZN(n6255) );
  XNOR2HSV4 U7695 ( .A1(n6257), .A2(\pe13/phq [5]), .ZN(n6256) );
  CLKNAND2HSV2 U7696 ( .A1(n14552), .A2(\pe13/pvq [5]), .ZN(n6257) );
  XNOR2HSV4 U7697 ( .A1(n6260), .A2(n6259), .ZN(n6258) );
  CLKNAND2HSV2 U7698 ( .A1(n7583), .A2(\pe13/aot [4]), .ZN(n6259) );
  CLKNAND2HSV2 U7699 ( .A1(n14939), .A2(\pe13/bq[4] ), .ZN(n6260) );
  AOI22HSV4 U7700 ( .A1(n14010), .A2(\pe17/ti_7t [7]), .B1(n15220), .B2(n13252), .ZN(n13261) );
  CLKNAND2HSV2 U7701 ( .A1(n12134), .A2(n12133), .ZN(n15220) );
  CLKNHSV2 U7702 ( .I(n12942), .ZN(n14450) );
  CLKNHSV0 U7703 ( .I(n14043), .ZN(n14044) );
  XNOR2HSV4 U7704 ( .A1(n6263), .A2(n6261), .ZN(n14043) );
  CLKXOR2HSV4 U7705 ( .A1(n6262), .A2(n14042), .Z(n6261) );
  NOR2HSV2 U7706 ( .A1(n14465), .A2(n14029), .ZN(n6262) );
  NOR2HSV3 U7707 ( .A1(n12942), .A2(n6264), .ZN(n6263) );
  CLKNHSV4 U7708 ( .I(\pe7/got [3]), .ZN(n6264) );
  CLKNHSV3 U7709 ( .I(\pe3/ctrq ), .ZN(n6266) );
  CLKNHSV2 U7710 ( .I(\pe3/phq [1]), .ZN(n6269) );
  CLKNAND2HSV2 U7711 ( .A1(\pe3/ctrq ), .A2(\pe3/pvq [1]), .ZN(n6268) );
  NOR2HSV4 U7712 ( .A1(n6266), .A2(n6265), .ZN(n6267) );
  CLKNAND2HSV2 U7713 ( .A1(\pe3/phq [1]), .A2(\pe3/pvq [1]), .ZN(n6265) );
  AOI21HSV4 U7714 ( .A1(n6269), .A2(n6268), .B(n6267), .ZN(n10165) );
  CLKNHSV0 U7715 ( .I(n6270), .ZN(n10712) );
  CLKNAND2HSV3 U7716 ( .A1(n6672), .A2(n6671), .ZN(n6270) );
  CLKNAND2HSV4 U7717 ( .A1(n6272), .A2(n6271), .ZN(n6672) );
  CLKNHSV4 U7718 ( .I(n10470), .ZN(n6271) );
  CLKNHSV4 U7719 ( .I(n10471), .ZN(n6272) );
  XNOR2HSV4 U7720 ( .A1(n6277), .A2(n6273), .ZN(n11259) );
  NOR2HSV4 U7721 ( .A1(n12879), .A2(n12878), .ZN(n6273) );
  AOI21HSV4 U7722 ( .A1(n15293), .A2(n6276), .B(n6274), .ZN(n12879) );
  CLKNHSV2 U7723 ( .I(n6275), .ZN(n6274) );
  CLKNAND2HSV2 U7724 ( .A1(n9358), .A2(\pe2/ti_7t [3]), .ZN(n6275) );
  CLKNHSV2 U7725 ( .I(n9358), .ZN(n6276) );
  XNOR2HSV1 U7726 ( .A1(n10798), .A2(n10797), .ZN(n15293) );
  XNOR2HSV4 U7727 ( .A1(n6279), .A2(n6278), .ZN(n6277) );
  CLKNHSV2 U7728 ( .I(n11258), .ZN(n6278) );
  XNOR2HSV4 U7729 ( .A1(n6280), .A2(n11243), .ZN(n6279) );
  CLKNAND2HSV2 U7730 ( .A1(n13762), .A2(\pe2/got [4]), .ZN(n6280) );
  XNOR2HSV4 U7731 ( .A1(n10371), .A2(n10370), .ZN(n6282) );
  CLKNHSV3 U7732 ( .I(n6281), .ZN(n10372) );
  OAI21HSV4 U7733 ( .A1(n6282), .A2(n10863), .B(n10374), .ZN(n10379) );
  CLKNAND2HSV3 U7734 ( .A1(n15225), .A2(n6283), .ZN(n10471) );
  INHSV2 U7735 ( .I(n7659), .ZN(n6283) );
  OAI21HSV4 U7736 ( .A1(n10471), .A2(n10470), .B(n10469), .ZN(n6284) );
  XNOR2HSV4 U7737 ( .A1(n6500), .A2(n6499), .ZN(n10470) );
  CLKNAND2HSV2 U7738 ( .A1(n10421), .A2(n12103), .ZN(n10438) );
  NAND2HSV2 U7739 ( .A1(n6285), .A2(\pe18/got [4]), .ZN(n14684) );
  CLKNAND2HSV2 U7740 ( .A1(n6285), .A2(n6039), .ZN(n13371) );
  CLKNAND2HSV3 U7741 ( .A1(n14682), .A2(n14681), .ZN(n6285) );
  OAI21HSV2 U7742 ( .A1(n10071), .A2(n10119), .B(n10118), .ZN(n14856) );
  AOI21HSV4 U7743 ( .A1(n6286), .A2(n7447), .B(n7449), .ZN(n10118) );
  NAND3HSV3 U7744 ( .A1(n7510), .A2(n7514), .A3(n7513), .ZN(n6287) );
  CLKNHSV2 U7745 ( .I(n9419), .ZN(n8507) );
  XNOR2HSV4 U7746 ( .A1(n6290), .A2(n6288), .ZN(n9419) );
  XNOR2HSV4 U7747 ( .A1(n6289), .A2(n6309), .ZN(n6288) );
  XNOR2HSV4 U7748 ( .A1(n6302), .A2(n6301), .ZN(n6289) );
  NOR2HSV4 U7749 ( .A1(n9430), .A2(n9009), .ZN(n6290) );
  NOR2HSV4 U7750 ( .A1(n12260), .A2(n9008), .ZN(n9430) );
  XNOR2HSV4 U7751 ( .A1(n6292), .A2(n6291), .ZN(n11434) );
  NOR2HSV4 U7752 ( .A1(n10759), .A2(n10730), .ZN(n6291) );
  NOR2HSV4 U7753 ( .A1(n15253), .A2(n7332), .ZN(n10759) );
  XNOR2HSV4 U7754 ( .A1(n6353), .A2(n6351), .ZN(n15253) );
  CLKNAND2HSV2 U7755 ( .A1(n15264), .A2(\pe10/got [8]), .ZN(n10064) );
  CLKNHSV2 U7756 ( .I(n14929), .ZN(n6294) );
  CLKNAND2HSV1 U7757 ( .A1(\pe10/aot [8]), .A2(\pe10/bq[8] ), .ZN(n6296) );
  CLKNHSV2 U7758 ( .I(n7102), .ZN(n6297) );
  CLKNAND2HSV2 U7759 ( .A1(\pe2/got [5]), .A2(\pe2/ti_1 ), .ZN(n6299) );
  CLKNAND2HSV2 U7760 ( .A1(\pe2/bq[7] ), .A2(\pe2/aot [6]), .ZN(n6300) );
  CLKNAND2HSV2 U7761 ( .A1(n13910), .A2(\pe9/got [6]), .ZN(n6815) );
  CLKNAND2HSV4 U7762 ( .A1(\pe9/aot [8]), .A2(\pe9/bq[6] ), .ZN(n6306) );
  OAI21HSV4 U7763 ( .A1(n6308), .A2(\pe9/phq [3]), .B(n6307), .ZN(n6301) );
  INAND2HSV4 U7764 ( .A1(n6304), .B1(n6305), .ZN(n6302) );
  BUFHSV8 U7765 ( .I(\pe9/aot [7]), .Z(n6303) );
  AOI21HSV4 U7766 ( .A1(\pe9/aot [7]), .A2(\pe9/bq[7] ), .B(n6306), .ZN(n6304)
         );
  NAND3HSV4 U7767 ( .A1(n6306), .A2(n6303), .A3(n13911), .ZN(n6305) );
  CLKNAND2HSV2 U7768 ( .A1(\pe9/got [6]), .A2(\pe9/ti_1 ), .ZN(n6308) );
  XOR2HSV2 U7769 ( .A1(n6311), .A2(n6310), .Z(n6309) );
  CLKNAND2HSV2 U7770 ( .A1(\pe9/pvq [3]), .A2(\pe9/ctrq ), .ZN(n6310) );
  NOR2HSV4 U7771 ( .A1(n9773), .A2(n15093), .ZN(n6311) );
  CLKNHSV2 U7772 ( .I(\pe9/aot [6]), .ZN(n9773) );
  NAND2HSV2 U7773 ( .A1(n15225), .A2(n8928), .ZN(n6444) );
  XNOR2HSV4 U7774 ( .A1(n10417), .A2(n10416), .ZN(n15225) );
  INAND2HSV1 U7775 ( .A1(n6313), .B1(n6563), .ZN(n15223) );
  NOR2HSV4 U7776 ( .A1(n6314), .A2(n6313), .ZN(n12111) );
  NOR2HSV3 U7777 ( .A1(n10714), .A2(n10715), .ZN(n6313) );
  CLKNAND2HSV2 U7778 ( .A1(n6563), .A2(n6315), .ZN(n6314) );
  CLKNHSV2 U7779 ( .I(n12020), .ZN(n6315) );
  AOI22HSV4 U7780 ( .A1(\pe19/ti_7t [2]), .A2(n9721), .B1(n9514), .B2(n6316), 
        .ZN(n9516) );
  NOR2HSV4 U7781 ( .A1(n9555), .A2(n9513), .ZN(n6316) );
  CLKNAND2HSV3 U7782 ( .A1(n9581), .A2(\pe19/got [6]), .ZN(n6528) );
  CLKNAND2HSV4 U7783 ( .A1(n9517), .A2(n9516), .ZN(n9581) );
  CLKNAND2HSV3 U7784 ( .A1(n13845), .A2(n6317), .ZN(n9517) );
  AOI21HSV4 U7785 ( .A1(n9500), .A2(n13844), .B(n9721), .ZN(n6317) );
  CLKNHSV2 U7786 ( .I(n9514), .ZN(n13845) );
  XOR3HSV0 U7787 ( .A1(n6320), .A2(n6319), .A3(n6318), .Z(n8709) );
  NOR2HSV3 U7788 ( .A1(n13102), .A2(n13101), .ZN(n6319) );
  MUX2NHSV1 U7789 ( .I0(n6324), .I1(n6323), .S(n6321), .ZN(n6320) );
  XNOR2HSV1 U7790 ( .A1(n13099), .A2(n6322), .ZN(n6321) );
  XNOR2HSV1 U7791 ( .A1(n8707), .A2(n13096), .ZN(n6322) );
  CLKNAND2HSV3 U7792 ( .A1(n14935), .A2(\pe2/got [2]), .ZN(n6323) );
  CLKNHSV3 U7793 ( .I(n6325), .ZN(n6324) );
  CLKNAND2HSV4 U7794 ( .A1(n14935), .A2(n8708), .ZN(n6325) );
  CLKBUFHSV2 U7795 ( .I(n14840), .Z(n6326) );
  CLKNHSV2 U7796 ( .I(n14840), .ZN(n7042) );
  CLKNAND2HSV2 U7797 ( .A1(n14840), .A2(\pe3/got [3]), .ZN(n11017) );
  CLKNAND2HSV2 U7798 ( .A1(n6326), .A2(\pe3/got [1]), .ZN(n12956) );
  CLKNAND2HSV2 U7799 ( .A1(n6326), .A2(\pe3/got [5]), .ZN(n12495) );
  CLKNAND2HSV2 U7800 ( .A1(n6326), .A2(\pe3/got [4]), .ZN(n12766) );
  XNOR2HSV4 U7801 ( .A1(n6328), .A2(n6327), .ZN(n8566) );
  CLKNAND2HSV2 U7802 ( .A1(n6326), .A2(\pe3/got [2]), .ZN(n6327) );
  OAI21HSV4 U7803 ( .A1(n10168), .A2(n10993), .B(n10992), .ZN(n14840) );
  CLKNHSV2 U7804 ( .I(n8565), .ZN(n6328) );
  OAI21HSV4 U7805 ( .A1(n13581), .A2(n6329), .B(n13582), .ZN(n6980) );
  CLKNAND2HSV2 U7806 ( .A1(n6329), .A2(n13582), .ZN(n13584) );
  XOR2HSV2 U7807 ( .A1(n8850), .A2(n6983), .Z(\pov14[7] ) );
  XNOR2HSV4 U7808 ( .A1(n6332), .A2(n6331), .ZN(n10203) );
  XNOR2HSV4 U7809 ( .A1(n10162), .A2(n10161), .ZN(n6332) );
  NOR2HSV8 U7810 ( .A1(n10433), .A2(n10419), .ZN(n10473) );
  NOR2HSV4 U7811 ( .A1(n10421), .A2(n10418), .ZN(n10433) );
  XNOR2HSV4 U7812 ( .A1(n10417), .A2(n10416), .ZN(n10421) );
  MUX2NHSV4 U7813 ( .I0(n9303), .I1(n9302), .S(n6341), .ZN(n6340) );
  XNOR2HSV4 U7814 ( .A1(n6334), .A2(n9299), .ZN(n6341) );
  XNOR2HSV4 U7815 ( .A1(n9300), .A2(n6335), .ZN(n6334) );
  CLKNHSV2 U7816 ( .I(n6341), .ZN(n6343) );
  CLKNHSV2 U7817 ( .I(n6344), .ZN(n6335) );
  CLKNHSV2 U7818 ( .I(n9829), .ZN(n9828) );
  XNOR2HSV4 U7819 ( .A1(n6338), .A2(n6336), .ZN(n9317) );
  CLKNAND2HSV2 U7820 ( .A1(n9829), .A2(n6337), .ZN(n6336) );
  CLKNHSV2 U7821 ( .I(n12410), .ZN(n6337) );
  CLKNAND2HSV2 U7822 ( .A1(n7813), .A2(n9533), .ZN(n9829) );
  NAND3HSV4 U7823 ( .A1(n6340), .A2(n6342), .A3(n6339), .ZN(n6338) );
  NAND3HSV4 U7824 ( .A1(n6341), .A2(n15071), .A3(n9536), .ZN(n6339) );
  CLKNAND2HSV2 U7825 ( .A1(n8910), .A2(n6343), .ZN(n6342) );
  CLKNHSV2 U7826 ( .I(n9301), .ZN(n6344) );
  CLKNAND2HSV3 U7827 ( .A1(n15246), .A2(n9978), .ZN(n7373) );
  XNOR2HSV4 U7828 ( .A1(n6346), .A2(n6345), .ZN(n15246) );
  OAI21HSV4 U7829 ( .A1(n6348), .A2(\pe13/phq [1]), .B(n6347), .ZN(n6345) );
  XNOR2HSV4 U7830 ( .A1(n6350), .A2(n6349), .ZN(n6346) );
  IOA21HSV4 U7831 ( .A1(\pe13/bq[8] ), .A2(\pe13/aot [8]), .B(\pe13/phq [1]), 
        .ZN(n6347) );
  CLKNAND2HSV2 U7832 ( .A1(\pe13/aot [8]), .A2(\pe13/bq[8] ), .ZN(n6348) );
  NAND2HSV3 U7833 ( .A1(\pe13/ti_1 ), .A2(\pe13/got [8]), .ZN(n6349) );
  CLKNAND2HSV2 U7834 ( .A1(\pe13/pvq [1]), .A2(\pe13/ctrq ), .ZN(n6350) );
  CLKNAND2HSV3 U7835 ( .A1(\pe12/bq[8] ), .A2(\pe12/aot [8]), .ZN(n6352) );
  CLKNAND2HSV3 U7836 ( .A1(\pe12/got [8]), .A2(\pe12/ti_1 ), .ZN(n6354) );
  XNOR2HSV4 U7837 ( .A1(n6352), .A2(\pe12/phq [1]), .ZN(n6351) );
  XNOR2HSV4 U7838 ( .A1(n6355), .A2(n6354), .ZN(n6353) );
  CLKNAND2HSV2 U7839 ( .A1(\pe12/pvq [1]), .A2(\pe12/ctrq ), .ZN(n6355) );
  NOR2HSV4 U7840 ( .A1(n13808), .A2(n13807), .ZN(n14650) );
  NOR2HSV4 U7841 ( .A1(n13803), .A2(n13143), .ZN(n13808) );
  CLKNAND2HSV2 U7842 ( .A1(n6356), .A2(n13804), .ZN(n13803) );
  CLKNAND2HSV2 U7843 ( .A1(n13138), .A2(n5997), .ZN(n6356) );
  CLKNHSV2 U7844 ( .I(n12183), .ZN(n12182) );
  OAI21HSV4 U7845 ( .A1(n6361), .A2(n6360), .B(n6357), .ZN(n12183) );
  CLKNAND2HSV2 U7846 ( .A1(n6358), .A2(n6361), .ZN(n6357) );
  CLKNAND2HSV2 U7847 ( .A1(n14867), .A2(\pe19/got [3]), .ZN(n6358) );
  CLKNHSV2 U7848 ( .I(n12340), .ZN(n6359) );
  CLKNAND2HSV2 U7849 ( .A1(n13316), .A2(\pe19/got [3]), .ZN(n6360) );
  XNOR2HSV4 U7850 ( .A1(n6363), .A2(n6362), .ZN(n6361) );
  CLKNAND2HSV2 U7851 ( .A1(n15084), .A2(\pe19/got [2]), .ZN(n6362) );
  XOR2HSV2 U7852 ( .A1(n12180), .A2(n12179), .Z(n6363) );
  CLKNAND2HSV2 U7853 ( .A1(\pe21/got [3]), .A2(\pe21/ti_1 ), .ZN(n10811) );
  NAND3HSV4 U7854 ( .A1(n6364), .A2(n12017), .A3(n12015), .ZN(n12013) );
  CLKNAND2HSV0 U7855 ( .A1(n6364), .A2(n12019), .ZN(n6428) );
  NOR2HSV8 U7856 ( .A1(n14736), .A2(n10673), .ZN(n10688) );
  XNOR2HSV4 U7857 ( .A1(n10672), .A2(n10671), .ZN(n14736) );
  XNOR2HSV4 U7858 ( .A1(n6365), .A2(n6370), .ZN(n6369) );
  XNOR2HSV4 U7859 ( .A1(n6367), .A2(n6366), .ZN(n6365) );
  XOR2HSV2 U7860 ( .A1(n8548), .A2(n7782), .Z(n6366) );
  XNOR2HSV4 U7861 ( .A1(n6372), .A2(n8549), .ZN(n6367) );
  NOR2HSV4 U7862 ( .A1(n10688), .A2(n10687), .ZN(n6368) );
  XOR2HSV2 U7863 ( .A1(n6371), .A2(n10684), .Z(n6370) );
  XNOR2HSV4 U7864 ( .A1(n7783), .A2(n10685), .ZN(n6371) );
  NOR2HSV4 U7865 ( .A1(n11827), .A2(n10683), .ZN(n6372) );
  CLKNAND2HSV3 U7866 ( .A1(n6374), .A2(n6375), .ZN(n6373) );
  CLKNHSV8 U7867 ( .I(\pe13/phq [2]), .ZN(n6375) );
  CLKNAND2HSV4 U7868 ( .A1(\pe13/bq[7] ), .A2(\pe13/aot [8]), .ZN(n6374) );
  OAI21HSV4 U7869 ( .A1(n6375), .A2(n6374), .B(n6373), .ZN(n9871) );
  CLKNHSV2 U7870 ( .I(n6376), .ZN(n6477) );
  CLKNAND2HSV2 U7871 ( .A1(n9363), .A2(n6377), .ZN(n6376) );
  CLKNHSV2 U7872 ( .I(n6478), .ZN(n6377) );
  CLKNAND2HSV2 U7873 ( .A1(n6378), .A2(n10798), .ZN(n9363) );
  NOR2HSV2 U7874 ( .A1(n10797), .A2(n6379), .ZN(n6378) );
  CLKNHSV2 U7875 ( .I(n9378), .ZN(n6379) );
  CLKNAND2HSV2 U7876 ( .A1(n6381), .A2(n6380), .ZN(n7123) );
  AOI31HSV2 U7877 ( .A1(n11210), .A2(n6382), .A3(n11209), .B(n11208), .ZN(
        n6381) );
  CLKNHSV1 U7878 ( .I(n12907), .ZN(n9388) );
  CLKNAND2HSV4 U7879 ( .A1(n9380), .A2(n10709), .ZN(n12907) );
  NAND3HSV4 U7880 ( .A1(n6385), .A2(n6384), .A3(n9386), .ZN(n13796) );
  INAND2HSV4 U7881 ( .A1(n9380), .B1(n11267), .ZN(n9386) );
  CLKNHSV2 U7882 ( .I(n9379), .ZN(n6384) );
  INAND2HSV4 U7883 ( .A1(n12907), .B1(n11264), .ZN(n6385) );
  NOR2HSV4 U7884 ( .A1(n11267), .A2(n9358), .ZN(n11264) );
  INHSV2 U7885 ( .I(n12133), .ZN(n6388) );
  NOR2HSV3 U7886 ( .A1(n14310), .A2(n14319), .ZN(n13271) );
  OAI22HSV4 U7887 ( .A1(n6387), .A2(n6388), .B1(n6407), .B2(n6409), .ZN(n14310) );
  CLKNAND2HSV2 U7888 ( .A1(n7887), .A2(n7886), .ZN(n7888) );
  XNOR2HSV4 U7889 ( .A1(n6390), .A2(n6389), .ZN(n7886) );
  NOR2HSV4 U7890 ( .A1(n11161), .A2(n14096), .ZN(n6389) );
  XOR2HSV2 U7891 ( .A1(n6392), .A2(n6391), .Z(n6390) );
  MUX2NHSV2 U7892 ( .I0(n7884), .I1(n13211), .S(n7822), .ZN(n6391) );
  XNOR2HSV4 U7893 ( .A1(n7820), .A2(n7819), .ZN(n6392) );
  CLKNHSV2 U7894 ( .I(n15086), .ZN(n12645) );
  CLKNAND2HSV2 U7895 ( .A1(n6395), .A2(n6393), .ZN(n12653) );
  CLKNAND2HSV2 U7896 ( .A1(n15086), .A2(n6394), .ZN(n6393) );
  CLKNHSV2 U7897 ( .I(n12644), .ZN(n6394) );
  CLKNAND2HSV2 U7898 ( .A1(n6396), .A2(n12643), .ZN(n6395) );
  CLKNAND2HSV2 U7899 ( .A1(n15086), .A2(n6397), .ZN(n6396) );
  CLKNHSV2 U7900 ( .I(n8009), .ZN(n6397) );
  CLKNAND2HSV2 U7901 ( .A1(n10512), .A2(n10511), .ZN(n15086) );
  CLKNHSV2 U7902 ( .I(n6407), .ZN(n6398) );
  CLKNHSV2 U7903 ( .I(n6401), .ZN(n6399) );
  INAND2HSV4 U7904 ( .A1(n6406), .B1(n6401), .ZN(n6400) );
  XNOR2HSV4 U7905 ( .A1(n6404), .A2(n6402), .ZN(n6401) );
  NAND2HSV2 U7906 ( .A1(n14824), .A2(\pe17/got [5]), .ZN(n6402) );
  INAND2HSV4 U7907 ( .A1(n6403), .B1(n6441), .ZN(n14824) );
  CLKNHSV2 U7908 ( .I(n6596), .ZN(n6403) );
  MUX2NHSV2 U7909 ( .I0(n7630), .I1(n7629), .S(n6405), .ZN(n6404) );
  NOR2HSV4 U7910 ( .A1(n14310), .A2(n14333), .ZN(n6406) );
  CLKNHSV2 U7911 ( .I(n6408), .ZN(n6407) );
  CLKNAND2HSV2 U7912 ( .A1(n13269), .A2(\pe17/ti_7t [7]), .ZN(n6408) );
  CLKNHSV2 U7913 ( .I(n13269), .ZN(n6409) );
  XNOR2HSV4 U7914 ( .A1(n6418), .A2(n6410), .ZN(n11767) );
  XOR4HSV2 U7915 ( .A1(n6416), .A2(n6414), .A3(n6412), .A4(n6411), .Z(n6410)
         );
  NOR2HSV4 U7916 ( .A1(n14854), .A2(n6413), .ZN(n6412) );
  CLKNHSV2 U7917 ( .I(\pe11/aot [6]), .ZN(n6413) );
  XOR2HSV2 U7918 ( .A1(n6415), .A2(\pe11/phq [3]), .Z(n6414) );
  NOR2HSV4 U7919 ( .A1(n11838), .A2(n6417), .ZN(n6416) );
  CLKNHSV2 U7920 ( .I(\pe11/pvq [3]), .ZN(n6417) );
  NOR2HSV4 U7921 ( .A1(n11734), .A2(n9610), .ZN(n6418) );
  NOR2HSV4 U7922 ( .A1(n15260), .A2(n11914), .ZN(n11734) );
  XNOR2HSV4 U7923 ( .A1(n6958), .A2(n6957), .ZN(n15260) );
  XNOR2HSV1 U7924 ( .A1(n6420), .A2(n6419), .ZN(n12935) );
  CLKNAND2HSV3 U7925 ( .A1(n15188), .A2(\pe13/got [4]), .ZN(n6419) );
  CLKNAND2HSV4 U7926 ( .A1(n9991), .A2(n9990), .ZN(n15188) );
  XNOR2HSV2 U7927 ( .A1(n6422), .A2(n6421), .ZN(n6420) );
  AOI31HSV1 U7928 ( .A1(\pe13/got [2]), .A2(n12933), .A3(n13587), .B(n12932), 
        .ZN(n6421) );
  CLKNAND2HSV3 U7929 ( .A1(n13603), .A2(n6423), .ZN(n6422) );
  INHSV2 U7930 ( .I(n12921), .ZN(n6423) );
  NOR2HSV4 U7931 ( .A1(n15167), .A2(n14400), .ZN(n13246) );
  NOR2HSV4 U7932 ( .A1(n15167), .A2(n14398), .ZN(n14428) );
  NOR2HSV4 U7933 ( .A1(n15167), .A2(n14319), .ZN(n14327) );
  CLKNHSV2 U7934 ( .I(ctro16), .ZN(n10796) );
  CLKNHSV2 U7935 ( .I(n10690), .ZN(n10673) );
  CLKNAND2HSV2 U7936 ( .A1(n10690), .A2(ctro16), .ZN(n10686) );
  CLKNAND2HSV2 U7937 ( .A1(\pe16/ti_7t [1]), .A2(ctro16), .ZN(n10690) );
  CLKNAND2HSV2 U7938 ( .A1(n6429), .A2(n12037), .ZN(n12040) );
  AOI21HSV4 U7939 ( .A1(n8911), .A2(n6427), .B(n6424), .ZN(n12037) );
  OAI21HSV2 U7940 ( .A1(n6426), .A2(n12019), .B(n6425), .ZN(n6424) );
  CLKNHSV2 U7941 ( .I(n12018), .ZN(n6425) );
  CLKNAND2HSV0 U7942 ( .A1(n12013), .A2(n13252), .ZN(n6426) );
  CLKNAND2HSV2 U7943 ( .A1(n12033), .A2(n12036), .ZN(n6429) );
  OAI21HSV4 U7944 ( .A1(n12111), .A2(n12032), .B(n6433), .ZN(n12036) );
  CLKNAND2HSV2 U7945 ( .A1(n6432), .A2(n6430), .ZN(n12033) );
  NOR2HSV4 U7946 ( .A1(n12111), .A2(n6431), .ZN(n6430) );
  CLKNHSV2 U7947 ( .I(n12035), .ZN(n6431) );
  XNOR2HSV4 U7948 ( .A1(n12030), .A2(n6434), .ZN(n6433) );
  CLKNHSV2 U7949 ( .I(n12029), .ZN(n6434) );
  BUFHSV8 U7950 ( .I(n6459), .Z(n6435) );
  NOR2HSV4 U7951 ( .A1(n6435), .A2(n13801), .ZN(n13802) );
  AOI21HSV4 U7952 ( .A1(n6459), .A2(n9398), .B(n10645), .ZN(n10661) );
  AOI21HSV4 U7953 ( .A1(n6435), .A2(n10841), .B(n7970), .ZN(n7532) );
  XNOR2HSV4 U7954 ( .A1(n10809), .A2(n10810), .ZN(n6459) );
  XNOR2HSV4 U7955 ( .A1(n12624), .A2(n6436), .ZN(n12626) );
  XNOR2HSV4 U7956 ( .A1(n6438), .A2(n6437), .ZN(n6436) );
  CLKNAND2HSV2 U7957 ( .A1(n7127), .A2(\pe15/got [2]), .ZN(n6437) );
  XNOR2HSV4 U7958 ( .A1(n6439), .A2(n12622), .ZN(n6438) );
  CLKNHSV2 U7959 ( .I(n12623), .ZN(n6439) );
  XNOR2HSV4 U7960 ( .A1(n6442), .A2(n12108), .ZN(n15222) );
  NOR2HSV4 U7961 ( .A1(n15167), .A2(n14397), .ZN(n6442) );
  CLKNAND2HSV0 U7962 ( .A1(\pe21/ti_7[5] ), .A2(\pe21/got [3]), .ZN(n12557) );
  CLKNHSV2 U7963 ( .I(n7405), .ZN(n6443) );
  CLKNHSV2 U7964 ( .I(\pe2/aot [8]), .ZN(n9328) );
  CLKBUFHSV2 U7965 ( .I(n9823), .Z(n6445) );
  CLKNAND2HSV4 U7966 ( .A1(n6773), .A2(n6772), .ZN(n9823) );
  XNOR2HSV4 U7967 ( .A1(n9263), .A2(n9262), .ZN(n9834) );
  XNOR2HSV4 U7968 ( .A1(n6447), .A2(n9260), .ZN(n6446) );
  XNOR2HSV4 U7969 ( .A1(n9256), .A2(n9255), .ZN(n6447) );
  CLKNHSV2 U7970 ( .I(\pe2/got [8]), .ZN(n10708) );
  CLKNAND2HSV2 U7971 ( .A1(n6448), .A2(\pe21/phq [1]), .ZN(n9396) );
  NAND2HSV2 U7972 ( .A1(\pe21/aot [8]), .A2(\pe21/bq[8] ), .ZN(n6448) );
  AOI21HSV4 U7973 ( .A1(n6454), .A2(n6453), .B(n6449), .ZN(n7681) );
  NAND3HSV4 U7974 ( .A1(n6452), .A2(n7682), .A3(n6450), .ZN(n6449) );
  CLKNAND2HSV2 U7975 ( .A1(n6451), .A2(n7321), .ZN(n6450) );
  CLKNHSV2 U7976 ( .I(n6554), .ZN(n6451) );
  INAND2HSV4 U7977 ( .A1(n7321), .B1(n7842), .ZN(n6452) );
  CLKNAND2HSV2 U7978 ( .A1(n7321), .A2(n6555), .ZN(n6453) );
  NOR2HSV4 U7979 ( .A1(n6455), .A2(n6551), .ZN(n6454) );
  NOR2HSV4 U7980 ( .A1(n7321), .A2(n6552), .ZN(n6455) );
  CLKNAND2HSV2 U7981 ( .A1(n6456), .A2(\pe17/aot [3]), .ZN(n6665) );
  CLKNAND2HSV2 U7982 ( .A1(n6456), .A2(\pe17/aot [2]), .ZN(n12119) );
  CLKNAND2HSV2 U7983 ( .A1(n6456), .A2(\pe17/aot [1]), .ZN(n14413) );
  MUX2NHSV2 U7984 ( .I0(n6458), .I1(n6457), .S(n14571), .ZN(n15057) );
  CLKNHSV2 U7985 ( .I(n6456), .ZN(n6457) );
  CLKNHSV2 U7986 ( .I(bo17[8]), .ZN(n6458) );
  CLKNAND2HSV4 U7987 ( .A1(n14740), .A2(n6817), .ZN(n6760) );
  XNOR2HSV4 U7988 ( .A1(n12019), .A2(n12013), .ZN(n14740) );
  XNOR2HSV4 U7989 ( .A1(n6461), .A2(n6460), .ZN(n12019) );
  NAND3HSV4 U7990 ( .A1(n10423), .A2(n13252), .A3(n6569), .ZN(n12017) );
  NOR2HSV4 U7991 ( .A1(n6462), .A2(n6536), .ZN(n6460) );
  XNOR2HSV4 U7992 ( .A1(n6539), .A2(n10434), .ZN(n6461) );
  XNOR2HSV4 U7993 ( .A1(n6468), .A2(n6464), .ZN(n7472) );
  CLKNAND2HSV2 U7994 ( .A1(n6465), .A2(n9950), .ZN(n6464) );
  OAI211HSV2 U7995 ( .A1(n7624), .A2(n8027), .B(n6466), .C(n7623), .ZN(n6465)
         );
  CLKNAND2HSV2 U7996 ( .A1(n7624), .A2(n6467), .ZN(n6466) );
  XNOR2HSV4 U7997 ( .A1(n6472), .A2(n6469), .ZN(n6468) );
  XOR3HSV2 U7998 ( .A1(n9945), .A2(n9944), .A3(n6470), .Z(n6469) );
  XNOR2HSV4 U7999 ( .A1(n6752), .A2(n6471), .ZN(n6470) );
  CLKNHSV2 U8000 ( .I(n9942), .ZN(n6471) );
  XNOR2HSV4 U8001 ( .A1(n6476), .A2(n6473), .ZN(n11267) );
  XNOR2HSV4 U8002 ( .A1(n6475), .A2(n6474), .ZN(n6473) );
  CLKNAND2HSV2 U8003 ( .A1(n13762), .A2(n14822), .ZN(n6475) );
  CLKNAND2HSV2 U8004 ( .A1(n9364), .A2(n6477), .ZN(n6476) );
  CLKNHSV2 U8005 ( .I(n9362), .ZN(n6478) );
  XNOR2HSV4 U8006 ( .A1(n6486), .A2(n6479), .ZN(n13879) );
  OAI21HSV4 U8007 ( .A1(n6483), .A2(n9709), .B(n6480), .ZN(n6479) );
  NAND3HSV4 U8008 ( .A1(n9709), .A2(n6482), .A3(n6481), .ZN(n6480) );
  NOR2HSV4 U8009 ( .A1(n9708), .A2(n9706), .ZN(n6481) );
  CLKNHSV2 U8010 ( .I(n9707), .ZN(n6482) );
  NOR2HSV4 U8011 ( .A1(n6485), .A2(n6484), .ZN(n6483) );
  CLKNAND2HSV2 U8012 ( .A1(n9703), .A2(n9705), .ZN(n6484) );
  CLKNHSV2 U8013 ( .I(n9704), .ZN(n6485) );
  OAI21HSV4 U8014 ( .A1(n12271), .A2(n9676), .B(n9675), .ZN(n6486) );
  CLKNAND2HSV2 U8015 ( .A1(n9638), .A2(n9639), .ZN(n6487) );
  XNOR2HSV4 U8016 ( .A1(n8033), .A2(n6849), .ZN(n15073) );
  INHSV6 U8017 ( .I(n6488), .ZN(n10373) );
  CLKNAND2HSV3 U8018 ( .A1(n10377), .A2(n10376), .ZN(n6488) );
  XNOR2HSV4 U8019 ( .A1(n13798), .A2(n10373), .ZN(n13799) );
  AOI22HSV4 U8020 ( .A1(n9746), .A2(n9449), .B1(n9744), .B2(n9435), .ZN(n7315)
         );
  XNOR2HSV4 U8021 ( .A1(n6494), .A2(n6490), .ZN(n9744) );
  XNOR2HSV4 U8022 ( .A1(n6492), .A2(n6491), .ZN(n6490) );
  CLKNAND2HSV2 U8023 ( .A1(n9783), .A2(n9434), .ZN(n6491) );
  XNOR2HSV4 U8024 ( .A1(n9433), .A2(n6493), .ZN(n6492) );
  CLKNHSV2 U8025 ( .I(n9432), .ZN(n6493) );
  AOI21HSV4 U8026 ( .A1(n6495), .A2(n9739), .B(n9421), .ZN(n6494) );
  XNOR2HSV4 U8027 ( .A1(n9419), .A2(n9783), .ZN(n6495) );
  NAND3HSV4 U8028 ( .A1(n6541), .A2(n6497), .A3(n6542), .ZN(n6496) );
  CLKNHSV2 U8029 ( .I(n6544), .ZN(n6497) );
  XNOR2HSV4 U8030 ( .A1(n6502), .A2(n6501), .ZN(n6499) );
  CLKNAND2HSV2 U8031 ( .A1(\pe17/bq[8] ), .A2(\pe17/aot [7]), .ZN(n6502) );
  XNOR2HSV4 U8032 ( .A1(n6504), .A2(n6503), .ZN(n7905) );
  CLKNAND2HSV2 U8033 ( .A1(n14944), .A2(\pe14/got [5]), .ZN(n6503) );
  XNOR2HSV4 U8034 ( .A1(n11112), .A2(n11111), .ZN(n6504) );
  CLKNHSV2 U8035 ( .I(\pe2/got [4]), .ZN(n13760) );
  CLKNHSV2 U8036 ( .I(\pe2/ti_1 ), .ZN(n13775) );
  XNOR2HSV4 U8037 ( .A1(n12507), .A2(n12506), .ZN(n15231) );
  XNOR2HSV4 U8038 ( .A1(n6507), .A2(n6506), .ZN(n12506) );
  OAI21HSV4 U8039 ( .A1(n15232), .A2(n12320), .B(n12319), .ZN(n6506) );
  XOR3HSV2 U8040 ( .A1(n6733), .A2(n6937), .A3(n6508), .Z(n6507) );
  NOR2HSV4 U8041 ( .A1(n11407), .A2(n6936), .ZN(n6508) );
  CLKNAND2HSV2 U8042 ( .A1(n14914), .A2(n15178), .ZN(n12507) );
  NAND2HSV2 U8043 ( .A1(n11084), .A2(n11085), .ZN(n6509) );
  OAI21HSV4 U8044 ( .A1(n11088), .A2(n11087), .B(n11086), .ZN(n6510) );
  CLKNAND2HSV4 U8045 ( .A1(n6510), .A2(n6509), .ZN(n11094) );
  INHSV2 U8046 ( .I(n11094), .ZN(n11121) );
  XNOR2HSV4 U8047 ( .A1(n6511), .A2(n8465), .ZN(n10430) );
  INHSV1 U8048 ( .I(n9000), .ZN(n9001) );
  AOI21HSV4 U8049 ( .A1(n6513), .A2(n6512), .B(n9004), .ZN(n9007) );
  XNOR2HSV4 U8050 ( .A1(n7245), .A2(\pe16/phq [1]), .ZN(n10671) );
  XNOR2HSV4 U8051 ( .A1(n7247), .A2(n7246), .ZN(n10672) );
  CLKNAND2HSV2 U8052 ( .A1(\pe6/bq[5] ), .A2(\pe6/aot [6]), .ZN(n9298) );
  XNOR2HSV4 U8053 ( .A1(n6516), .A2(n6515), .ZN(n6522) );
  XNOR2HSV4 U8054 ( .A1(n6660), .A2(n6659), .ZN(n6515) );
  XNOR2HSV4 U8055 ( .A1(n10719), .A2(n10718), .ZN(n6516) );
  XNOR2HSV4 U8056 ( .A1(n6518), .A2(n6517), .ZN(n10720) );
  XNOR2HSV4 U8057 ( .A1(n6521), .A2(n6520), .ZN(n6519) );
  XOR2HSV2 U8058 ( .A1(n6662), .A2(\pe17/phq [5]), .Z(n6520) );
  XNOR2HSV4 U8059 ( .A1(n14335), .A2(n6661), .ZN(n6521) );
  AOI21HSV2 U8060 ( .A1(n15073), .A2(n13844), .B(n6524), .ZN(n6954) );
  CLKNHSV2 U8061 ( .I(n9541), .ZN(n6524) );
  XNOR2HSV4 U8062 ( .A1(n6525), .A2(n6663), .ZN(n12028) );
  XOR4HSV2 U8063 ( .A1(n12024), .A2(n14408), .A3(n6527), .A4(n6526), .Z(n6525)
         );
  XNOR2HSV4 U8064 ( .A1(n6669), .A2(n6668), .ZN(n6526) );
  CLKNAND2HSV2 U8065 ( .A1(n14415), .A2(\pe17/got [3]), .ZN(n6527) );
  NOR2HSV4 U8066 ( .A1(n6667), .A2(n6666), .ZN(n14408) );
  XOR2HSV2 U8067 ( .A1(n9553), .A2(n9554), .Z(n6529) );
  OAI21HSV4 U8068 ( .A1(n15212), .A2(n10357), .B(n9543), .ZN(n6530) );
  XNOR2HSV4 U8069 ( .A1(n7377), .A2(n9540), .ZN(n15212) );
  CLKNAND2HSV2 U8070 ( .A1(n10356), .A2(n9541), .ZN(n9558) );
  CLKNAND2HSV4 U8071 ( .A1(n6532), .A2(n6531), .ZN(n7331) );
  CLKNHSV2 U8072 ( .I(n10794), .ZN(n6531) );
  XNOR2HSV4 U8073 ( .A1(n10675), .A2(n10674), .ZN(n10794) );
  CLKAND2HSV4 U8074 ( .A1(n7850), .A2(n6533), .Z(n6532) );
  CLKNHSV2 U8075 ( .I(n7849), .ZN(n6533) );
  CLKNHSV2 U8076 ( .I(n14914), .ZN(n6534) );
  NAND2HSV4 U8077 ( .A1(n6676), .A2(n6570), .ZN(n14914) );
  XNOR2HSV2 U8078 ( .A1(n12019), .A2(n12013), .ZN(n12107) );
  CLKNAND2HSV2 U8079 ( .A1(n6538), .A2(n6537), .ZN(n6536) );
  CLKNHSV2 U8080 ( .I(n10436), .ZN(n6537) );
  NAND3HSV2 U8081 ( .A1(n10438), .A2(n10470), .A3(n10437), .ZN(n6538) );
  XNOR2HSV4 U8082 ( .A1(n10430), .A2(n10429), .ZN(n6539) );
  CLKNAND2HSV3 U8083 ( .A1(\pe17/ti_1 ), .A2(\pe17/got [7]), .ZN(n6540) );
  NAND3HSV4 U8084 ( .A1(n6543), .A2(\pe17/ti_1 ), .A3(\pe17/got [7]), .ZN(
        n6542) );
  CLKNHSV2 U8085 ( .I(\pe17/phq [2]), .ZN(n6543) );
  CLKNAND2HSV2 U8086 ( .A1(\pe17/pvq [2]), .A2(\pe17/ctrq ), .ZN(n6544) );
  CLKNAND2HSV2 U8087 ( .A1(n6554), .A2(n6546), .ZN(n6545) );
  CLKNAND2HSV2 U8088 ( .A1(n7196), .A2(n7197), .ZN(n6546) );
  CLKNHSV4 U8089 ( .I(n7197), .ZN(n6555) );
  CLKNAND2HSV2 U8090 ( .A1(n6550), .A2(n6549), .ZN(n6548) );
  CLKNHSV2 U8091 ( .I(n7321), .ZN(n6549) );
  CLKNAND2HSV2 U8092 ( .A1(n6553), .A2(n7843), .ZN(n6550) );
  CLKNHSV2 U8093 ( .I(n7196), .ZN(n6551) );
  CLKNHSV2 U8094 ( .I(n7847), .ZN(n6552) );
  INAND2HSV4 U8095 ( .A1(n7847), .B1(n7196), .ZN(n6553) );
  INHSV24 U8096 ( .I(n7698), .ZN(n6557) );
  INHSV24 U8097 ( .I(n7697), .ZN(n6558) );
  CLKNAND2HSV3 U8098 ( .A1(n6559), .A2(n12507), .ZN(n12537) );
  CLKNAND2HSV2 U8099 ( .A1(n12506), .A2(n12337), .ZN(n6560) );
  IOA22HSV4 U8100 ( .B1(n12506), .B2(n6562), .A1(n6558), .A2(n6557), .ZN(
        n12538) );
  CLKNAND2HSV2 U8101 ( .A1(n14914), .A2(n12336), .ZN(n6562) );
  CLKNAND2HSV2 U8102 ( .A1(n6565), .A2(n10714), .ZN(n6563) );
  XNOR2HSV4 U8103 ( .A1(n10473), .A2(n10472), .ZN(n10714) );
  INAND2HSV4 U8104 ( .A1(n6564), .B1(n14962), .ZN(n10715) );
  CLKNHSV2 U8105 ( .I(n6568), .ZN(n6564) );
  CLKNAND2HSV2 U8106 ( .A1(n14962), .A2(n6566), .ZN(n6565) );
  CLKNHSV2 U8107 ( .I(n6567), .ZN(n6566) );
  NAND3HSV4 U8108 ( .A1(n10713), .A2(n6672), .A3(n6671), .ZN(n14962) );
  INHSV8 U8109 ( .I(n12103), .ZN(n6567) );
  XNOR2HSV4 U8110 ( .A1(n6976), .A2(n6974), .ZN(n10472) );
  CLKNHSV2 U8111 ( .I(n6670), .ZN(n6568) );
  NOR2HSV4 U8112 ( .A1(n6569), .A2(n12021), .ZN(n10422) );
  NAND2HSV2 U8113 ( .A1(n6842), .A2(n6995), .ZN(n6570) );
  CLKNAND2HSV2 U8114 ( .A1(n8581), .A2(n8582), .ZN(n8583) );
  XNOR2HSV4 U8115 ( .A1(n6571), .A2(n8580), .ZN(n8581) );
  CLKNAND2HSV2 U8116 ( .A1(n14914), .A2(\pe15/got [2]), .ZN(n6571) );
  NAND2HSV2 U8117 ( .A1(n14962), .A2(\pe17/got [5]), .ZN(n12029) );
  CLKNHSV2 U8118 ( .I(n7627), .ZN(n6572) );
  CLKNAND2HSV2 U8119 ( .A1(n6964), .A2(n7544), .ZN(n6573) );
  CLKNAND2HSV2 U8120 ( .A1(\pe21/ti_7[5] ), .A2(\pe21/got [4]), .ZN(n8393) );
  CLKNHSV2 U8121 ( .I(n6579), .ZN(n8901) );
  MUX2NHSV2 U8122 ( .I0(n6576), .I1(n6575), .S(n6574), .ZN(n7731) );
  XOR2HSV2 U8123 ( .A1(n10828), .A2(n10827), .Z(n6574) );
  CLKNHSV2 U8124 ( .I(n10834), .ZN(n6575) );
  NOR2HSV4 U8125 ( .A1(n10829), .A2(n6577), .ZN(n6576) );
  CLKNAND2HSV2 U8126 ( .A1(n6579), .A2(n6578), .ZN(n6577) );
  CLKNHSV2 U8127 ( .I(n10830), .ZN(n6578) );
  CLKNAND2HSV2 U8128 ( .A1(n10387), .A2(n6580), .ZN(n6579) );
  NOR2HSV4 U8129 ( .A1(n10810), .A2(n6581), .ZN(n6580) );
  CLKNHSV2 U8130 ( .I(n10841), .ZN(n6581) );
  NAND2HSV3 U8131 ( .A1(\pe15/bq[8] ), .A2(\pe15/aot [7]), .ZN(n6582) );
  CLKNAND2HSV2 U8132 ( .A1(n6582), .A2(\pe15/phq [2]), .ZN(n6583) );
  NAND3HSV4 U8133 ( .A1(n6585), .A2(\pe15/bq[8] ), .A3(\pe15/aot [7]), .ZN(
        n6584) );
  CLKNHSV2 U8134 ( .I(\pe15/phq [2]), .ZN(n6585) );
  NOR2HSV4 U8135 ( .A1(n6586), .A2(n13144), .ZN(n13344) );
  NOR2HSV4 U8136 ( .A1(n15217), .A2(n13140), .ZN(n6586) );
  CLKNHSV4 U8137 ( .I(n8513), .ZN(n6587) );
  CLKNHSV2 U8138 ( .I(n6589), .ZN(n6588) );
  CLKNHSV2 U8139 ( .I(n6590), .ZN(n6589) );
  INHSV24 U8140 ( .I(n14221), .ZN(n6590) );
  CLKNAND2HSV3 U8141 ( .A1(n7581), .A2(n7578), .ZN(n15084) );
  XNOR2HSV4 U8142 ( .A1(n6592), .A2(n6591), .ZN(n8514) );
  CLKNAND2HSV2 U8143 ( .A1(n12387), .A2(\pe19/got [5]), .ZN(n6591) );
  XOR2HSV2 U8144 ( .A1(n6594), .A2(n6593), .Z(n6592) );
  CLKNAND2HSV2 U8145 ( .A1(n15084), .A2(\pe19/got [4]), .ZN(n6593) );
  CLKNAND2HSV2 U8146 ( .A1(n6595), .A2(\pe15/phq [1]), .ZN(n6826) );
  CLKNAND2HSV2 U8147 ( .A1(\pe15/bq[8] ), .A2(\pe15/aot [8]), .ZN(n6595) );
  CLKNAND2HSV2 U8148 ( .A1(n14824), .A2(\pe17/got [4]), .ZN(n6628) );
  INAND2HSV4 U8149 ( .A1(n8928), .B1(\pe17/ti_7t [5]), .ZN(n6596) );
  CLKNHSV2 U8150 ( .I(n8928), .ZN(n6597) );
  CLKNHSV4 U8151 ( .I(n11827), .ZN(n6599) );
  CLKBUFHSV2 U8152 ( .I(n11827), .Z(n6598) );
  CLKNAND2HSV2 U8153 ( .A1(n6599), .A2(\pe16/pvq [7]), .ZN(n11164) );
  CLKNAND2HSV2 U8154 ( .A1(n6599), .A2(\pe16/pvq [6]), .ZN(n11187) );
  MUX2NHSV2 U8155 ( .I0(n6601), .I1(n6600), .S(n6598), .ZN(n14992) );
  CLKNHSV2 U8156 ( .I(bo16[2]), .ZN(n6600) );
  CLKNHSV2 U8157 ( .I(\pe16/bq[2] ), .ZN(n6601) );
  MUX2NHSV2 U8158 ( .I0(n6603), .I1(n6602), .S(n6598), .ZN(n15001) );
  CLKNHSV2 U8159 ( .I(bo16[6]), .ZN(n6602) );
  CLKNHSV2 U8160 ( .I(n14527), .ZN(n6603) );
  CLKNAND2HSV0 U8161 ( .A1(n8679), .A2(n6604), .ZN(n8680) );
  INAND2HSV1 U8162 ( .A1(n8678), .B1(n6605), .ZN(n6604) );
  NOR2HSV0 U8163 ( .A1(n15167), .A2(n14347), .ZN(n6605) );
  XNOR2HSV2 U8164 ( .A1(n6608), .A2(n6606), .ZN(n8678) );
  XOR3HSV1 U8165 ( .A1(n14344), .A2(n6607), .A3(n8676), .Z(n6606) );
  INHSV2 U8166 ( .I(n14346), .ZN(n6607) );
  INHSV2 U8167 ( .I(n8677), .ZN(n6608) );
  INHSV2 U8168 ( .I(n6622), .ZN(n6613) );
  XNOR2HSV4 U8169 ( .A1(n6610), .A2(n6609), .ZN(n6622) );
  CLKNAND2HSV2 U8170 ( .A1(n14958), .A2(\pe16/got [5]), .ZN(n6609) );
  XNOR2HSV4 U8171 ( .A1(n11199), .A2(n11198), .ZN(n6610) );
  AOI21HSV4 U8172 ( .A1(n6615), .A2(n10794), .B(n6618), .ZN(n6612) );
  INHSV24 U8173 ( .I(n11202), .ZN(n6614) );
  CLKNHSV2 U8174 ( .I(n6623), .ZN(n11203) );
  CLKNAND2HSV2 U8175 ( .A1(n7850), .A2(n6616), .ZN(n6615) );
  CLKNHSV2 U8176 ( .I(n6619), .ZN(n6616) );
  CLKNAND2HSV2 U8177 ( .A1(n6617), .A2(n10794), .ZN(n7848) );
  CLKNAND2HSV2 U8178 ( .A1(n7850), .A2(n12194), .ZN(n6617) );
  CLKNHSV2 U8179 ( .I(n6895), .ZN(n6618) );
  CLKNHSV2 U8180 ( .I(n12194), .ZN(n6619) );
  NAND3HSV4 U8181 ( .A1(n6623), .A2(n6622), .A3(n11201), .ZN(n6621) );
  CLKNAND2HSV0 U8182 ( .A1(n6626), .A2(n6624), .ZN(\pe17/poht [2]) );
  NAND3HSV2 U8183 ( .A1(n6633), .A2(n6630), .A3(n6625), .ZN(n6624) );
  CLKNHSV3 U8184 ( .I(n6627), .ZN(n6625) );
  CLKNAND2HSV3 U8185 ( .A1(n6629), .A2(n6627), .ZN(n6626) );
  XNOR2HSV2 U8186 ( .A1(n6628), .A2(n8188), .ZN(n6627) );
  CLKNAND2HSV3 U8187 ( .A1(n6633), .A2(n6630), .ZN(n6629) );
  CLKNAND2HSV3 U8188 ( .A1(n6632), .A2(n6631), .ZN(n6630) );
  CLKNHSV4 U8189 ( .I(n6643), .ZN(n6631) );
  INHSV2 U8190 ( .I(n6644), .ZN(n6632) );
  CLKNAND2HSV3 U8191 ( .A1(n6636), .A2(n6634), .ZN(n6633) );
  CLKNAND2HSV3 U8192 ( .A1(n6643), .A2(n6635), .ZN(n6634) );
  CLKNHSV3 U8193 ( .I(n6637), .ZN(n6635) );
  NAND2HSV2 U8194 ( .A1(n6642), .A2(n6637), .ZN(n6636) );
  CLKNAND2HSV3 U8195 ( .A1(n6641), .A2(n6638), .ZN(n6637) );
  INHSV2 U8196 ( .I(n6639), .ZN(n6638) );
  NAND2HSV2 U8197 ( .A1(n14012), .A2(n8928), .ZN(n6639) );
  INAND2HSV2 U8198 ( .A1(n6640), .B1(n7631), .ZN(n14012) );
  CLKNHSV3 U8199 ( .I(n12103), .ZN(n6640) );
  INHSV2 U8200 ( .I(n14011), .ZN(n6641) );
  CLKNAND2HSV1 U8201 ( .A1(n6644), .A2(n6643), .ZN(n6642) );
  CLKNAND2HSV4 U8202 ( .A1(n7039), .A2(\pe17/got [5]), .ZN(n6643) );
  AOI21HSV2 U8203 ( .A1(n6646), .A2(n7039), .B(n6645), .ZN(n6644) );
  INHSV1 U8204 ( .I(n14014), .ZN(n6645) );
  INHSV2 U8205 ( .I(n6647), .ZN(n6646) );
  CLKNAND2HSV3 U8206 ( .A1(n14011), .A2(n14007), .ZN(n6647) );
  INHSV2 U8207 ( .I(n6732), .ZN(n14708) );
  XNOR2HSV4 U8208 ( .A1(n6652), .A2(n6648), .ZN(n12847) );
  XOR3HSV2 U8209 ( .A1(n12843), .A2(n6650), .A3(n6649), .Z(n6648) );
  CLKNHSV2 U8210 ( .I(n12845), .ZN(n6649) );
  NOR2HSV4 U8211 ( .A1(n6732), .A2(n6651), .ZN(n6650) );
  CLKNHSV2 U8212 ( .I(\pe15/got [3]), .ZN(n6651) );
  CLKNAND2HSV2 U8213 ( .A1(n12614), .A2(n6653), .ZN(n6652) );
  CLKNHSV2 U8214 ( .I(n12844), .ZN(n6653) );
  CLKNAND2HSV2 U8215 ( .A1(n7436), .A2(n7435), .ZN(n12614) );
  CLKNAND2HSV3 U8216 ( .A1(n6654), .A2(n14065), .ZN(n6655) );
  CLKNAND2HSV3 U8217 ( .A1(n15186), .A2(n7647), .ZN(n14065) );
  OAI21HSV4 U8218 ( .A1(n15226), .A2(n8956), .B(n13188), .ZN(n14364) );
  OAI21HSV4 U8219 ( .A1(n14065), .A2(n6654), .B(n6655), .ZN(n15226) );
  NOR2HSV4 U8220 ( .A1(n14364), .A2(n14349), .ZN(n13377) );
  CLKNAND2HSV2 U8221 ( .A1(n8625), .A2(n8624), .ZN(n8626) );
  XNOR2HSV4 U8222 ( .A1(n6658), .A2(n6656), .ZN(n8624) );
  CLKNHSV2 U8223 ( .I(n6657), .ZN(n6656) );
  CLKNAND2HSV2 U8224 ( .A1(n15084), .A2(\pe19/got [3]), .ZN(n6657) );
  CLKNHSV2 U8225 ( .I(n8623), .ZN(n6658) );
  CLKNAND2HSV2 U8226 ( .A1(n13316), .A2(\pe19/got [4]), .ZN(n8625) );
  CLKNAND2HSV2 U8227 ( .A1(\pe17/bq[5] ), .A2(\pe17/aot [7]), .ZN(n6659) );
  CLKNAND2HSV2 U8228 ( .A1(\pe17/aot [5]), .A2(\pe17/bq[7] ), .ZN(n14335) );
  CLKNAND2HSV2 U8229 ( .A1(\pe17/pvq [5]), .A2(\pe17/ctrq ), .ZN(n6660) );
  CLKNAND2HSV2 U8230 ( .A1(\pe17/bq[6] ), .A2(\pe17/aot [6]), .ZN(n6661) );
  CLKNAND2HSV2 U8231 ( .A1(\pe17/bq[8] ), .A2(\pe17/aot [4]), .ZN(n6662) );
  XOR2HSV2 U8232 ( .A1(n12025), .A2(n6665), .Z(n6664) );
  CLKNHSV2 U8233 ( .I(\pe17/bq[3] ), .ZN(n6666) );
  CLKNHSV2 U8234 ( .I(n14949), .ZN(n6667) );
  CLKNAND2HSV2 U8235 ( .A1(\pe17/aot [5]), .A2(\pe17/bq[6] ), .ZN(n6668) );
  CLKNAND2HSV2 U8236 ( .A1(\pe17/aot [4]), .A2(\pe17/bq[7] ), .ZN(n6669) );
  CLKNAND2HSV2 U8237 ( .A1(n10714), .A2(n10715), .ZN(n7097) );
  CLKNHSV2 U8238 ( .I(n12103), .ZN(n6670) );
  CLKNHSV2 U8239 ( .I(n7691), .ZN(n6671) );
  CLKNAND2HSV2 U8240 ( .A1(n11404), .A2(n11403), .ZN(n11701) );
  NAND3HSV4 U8241 ( .A1(n6673), .A2(n11700), .A3(n11699), .ZN(n6676) );
  NOR2HSV4 U8242 ( .A1(n6675), .A2(n6674), .ZN(n6673) );
  CLKNAND2HSV2 U8243 ( .A1(n11403), .A2(n6848), .ZN(n6674) );
  CLKNHSV2 U8244 ( .I(n11404), .ZN(n6675) );
  CLKNAND2HSV4 U8245 ( .A1(n10704), .A2(n7845), .ZN(n14958) );
  XNOR2HSV4 U8246 ( .A1(n10703), .A2(n10702), .ZN(n6678) );
  CLKNHSV2 U8247 ( .I(n6732), .ZN(n7127) );
  CLKNAND2HSV2 U8248 ( .A1(n7371), .A2(n6679), .ZN(n11700) );
  CLKNHSV2 U8249 ( .I(n6680), .ZN(n6679) );
  CLKNAND2HSV2 U8250 ( .A1(n6732), .A2(n7372), .ZN(n6680) );
  CLKNAND2HSV2 U8251 ( .A1(n7336), .A2(n11702), .ZN(n11699) );
  CLKNHSV2 U8252 ( .I(n6681), .ZN(n7737) );
  CLKNAND2HSV2 U8253 ( .A1(\pe13/ti_7[4] ), .A2(\pe13/got [3]), .ZN(n6681) );
  CLKNAND2HSV4 U8254 ( .A1(n11323), .A2(n11324), .ZN(n11390) );
  CLKNAND2HSV3 U8255 ( .A1(n7305), .A2(n13857), .ZN(n11324) );
  CLKNAND2HSV4 U8256 ( .A1(n7304), .A2(n7303), .ZN(n11323) );
  CLKNAND2HSV2 U8257 ( .A1(n15232), .A2(n12337), .ZN(n7436) );
  OAI21HSV4 U8258 ( .A1(n6934), .A2(n6732), .B(n6682), .ZN(n15232) );
  OAI21HSV4 U8259 ( .A1(n6732), .A2(n8744), .B(n11702), .ZN(n6682) );
  CLKNAND2HSV2 U8260 ( .A1(n7370), .A2(n7368), .ZN(n11702) );
  XNOR2HSV4 U8261 ( .A1(n6687), .A2(n6683), .ZN(n13260) );
  XNOR2HSV4 U8262 ( .A1(n6686), .A2(n6684), .ZN(n6683) );
  NOR2HSV4 U8263 ( .A1(n10355), .A2(n6685), .ZN(n6684) );
  CLKNHSV2 U8264 ( .I(\pe19/got [6]), .ZN(n6685) );
  XOR2HSV2 U8265 ( .A1(n12169), .A2(n12168), .Z(n6686) );
  CLKNAND2HSV2 U8266 ( .A1(n12147), .A2(n6688), .ZN(n6687) );
  AOI31HSV2 U8267 ( .A1(n14219), .A2(n12146), .A3(n12145), .B(n12144), .ZN(
        n6688) );
  NOR2HSV4 U8268 ( .A1(n10356), .A2(n12135), .ZN(n12146) );
  XNOR2HSV4 U8269 ( .A1(n6697), .A2(n6689), .ZN(\pe19/poht [5]) );
  MUX2NHSV2 U8270 ( .I0(n6696), .I1(n6693), .S(n6690), .ZN(n6689) );
  XNOR2HSV4 U8271 ( .A1(n6692), .A2(n6691), .ZN(n6690) );
  CLKNHSV2 U8272 ( .I(n8675), .ZN(n6691) );
  CLKNAND2HSV2 U8273 ( .A1(n15084), .A2(\pe19/got [1]), .ZN(n6692) );
  CLKNHSV2 U8274 ( .I(n6694), .ZN(n6693) );
  CLKNAND2HSV2 U8275 ( .A1(n13316), .A2(\pe19/got [2]), .ZN(n6694) );
  CLKNHSV2 U8276 ( .I(n6785), .ZN(n6695) );
  CLKNAND2HSV2 U8277 ( .A1(n12387), .A2(\pe19/got [2]), .ZN(n6696) );
  CLKNAND2HSV2 U8278 ( .A1(n13315), .A2(\pe19/got [3]), .ZN(n6697) );
  CLKXOR2HSV4 U8279 ( .A1(n9552), .A2(n9551), .Z(n9553) );
  AOI21HSV0 U8280 ( .A1(n10281), .A2(n12866), .B(n7901), .ZN(n10282) );
  AND2HSV4 U8281 ( .A1(n10281), .A2(n10601), .Z(n10232) );
  AOI22HSV4 U8282 ( .A1(n10225), .A2(n10224), .B1(n10281), .B2(n10223), .ZN(
        n10226) );
  INAND2HSV2 U8283 ( .A1(n7398), .B1(n9727), .ZN(n9537) );
  NAND3HSV2 U8284 ( .A1(n9560), .A2(n9541), .A3(n9730), .ZN(n9562) );
  NOR2HSV2 U8285 ( .A1(n10222), .A2(n8931), .ZN(n10281) );
  INHSV4 U8286 ( .I(\pe1/aot [8]), .ZN(n10222) );
  CLKNAND2HSV2 U8287 ( .A1(n10230), .A2(n10229), .ZN(n10231) );
  NAND2HSV2 U8288 ( .A1(n14867), .A2(n8435), .ZN(n7637) );
  NAND2HSV2 U8289 ( .A1(n14867), .A2(\pe19/got [6]), .ZN(n7639) );
  NAND2HSV4 U8290 ( .A1(n10271), .A2(n10270), .ZN(n10272) );
  CLKNAND2HSV2 U8291 ( .A1(n10273), .A2(n10269), .ZN(n10271) );
  INHSV4 U8292 ( .I(n10272), .ZN(n10627) );
  CLKXOR2HSV4 U8293 ( .A1(n11706), .A2(poh21[6]), .Z(po[7]) );
  CLKNAND2HSV2 U8294 ( .A1(\pe1/aot [8]), .A2(\pe1/bq[7] ), .ZN(n10225) );
  NOR2HSV4 U8295 ( .A1(n10268), .A2(n10267), .ZN(n10269) );
  CLKXOR2HSV4 U8296 ( .A1(n10253), .A2(n10252), .Z(n10254) );
  XNOR2HSV4 U8297 ( .A1(n6698), .A2(n10254), .ZN(n10258) );
  XNOR2HSV4 U8298 ( .A1(n10251), .A2(n10250), .ZN(n6698) );
  BUFHSV8 U8299 ( .I(n13879), .Z(n13880) );
  NOR2HSV4 U8300 ( .A1(n12658), .A2(n10587), .ZN(n8644) );
  CLKNAND2HSV4 U8301 ( .A1(n7551), .A2(n7550), .ZN(\pe8/ti_7[1] ) );
  CLKNAND2HSV4 U8302 ( .A1(n7774), .A2(n7775), .ZN(n6750) );
  NAND2HSV2 U8303 ( .A1(\pe8/ti_7[1] ), .A2(n13488), .ZN(n7282) );
  XNOR2HSV4 U8304 ( .A1(n11562), .A2(n6699), .ZN(n7178) );
  CLKXOR2HSV4 U8305 ( .A1(n11559), .A2(n11558), .Z(n6699) );
  NAND2HSV4 U8306 ( .A1(n7771), .A2(n7772), .ZN(n7181) );
  NAND3HSV3 U8307 ( .A1(n12769), .A2(n11602), .A3(n7773), .ZN(n7772) );
  NAND2HSV2 U8308 ( .A1(n12787), .A2(n12775), .ZN(n6923) );
  CLKNAND2HSV8 U8309 ( .A1(n6751), .A2(n6750), .ZN(n11607) );
  OAI21HSV2 U8310 ( .A1(n6863), .A2(n6866), .B(n6864), .ZN(n13538) );
  NOR2HSV2 U8311 ( .A1(n7181), .A2(n6863), .ZN(n7180) );
  CLKNAND2HSV4 U8312 ( .A1(n8965), .A2(n8963), .ZN(n8962) );
  CLKXOR2HSV4 U8313 ( .A1(n11489), .A2(n11488), .Z(n11491) );
  NAND2HSV4 U8314 ( .A1(n9342), .A2(n9341), .ZN(n9345) );
  NAND2HSV2 U8315 ( .A1(n9342), .A2(n9341), .ZN(n8990) );
  NAND2HSV4 U8316 ( .A1(n7141), .A2(n14247), .ZN(\pe12/ti_7[3] ) );
  NAND2HSV2 U8317 ( .A1(n15251), .A2(n11446), .ZN(n7141) );
  INHSV2 U8318 ( .I(n7391), .ZN(n8903) );
  NAND2HSV2 U8319 ( .A1(n11444), .A2(n11448), .ZN(n7391) );
  NAND2HSV4 U8320 ( .A1(n7113), .A2(n7114), .ZN(n7508) );
  OAI21HSV0 U8321 ( .A1(n6700), .A2(n8833), .B(n8834), .ZN(n15268) );
  NOR2HSV4 U8322 ( .A1(n10496), .A2(n13516), .ZN(n10480) );
  CLKXOR2HSV2 U8323 ( .A1(n10482), .A2(n10481), .Z(n6700) );
  INHSV4 U8324 ( .I(n7274), .ZN(n11519) );
  BUFHSV8 U8325 ( .I(n11606), .Z(n6863) );
  BUFHSV4 U8326 ( .I(n12981), .Z(n14941) );
  NAND2HSV2 U8327 ( .A1(\pe15/pvq [1]), .A2(\pe15/ctrq ), .ZN(n6824) );
  XOR2HSV4 U8328 ( .A1(n10087), .A2(n10086), .Z(n10111) );
  XNOR2HSV4 U8329 ( .A1(n13787), .A2(n13786), .ZN(n15269) );
  CLKNHSV0 U8330 ( .I(n13257), .ZN(n8612) );
  CLKNAND2HSV2 U8331 ( .A1(n7965), .A2(n7964), .ZN(n7966) );
  CLKNAND2HSV2 U8332 ( .A1(\pov7[5] ), .A2(n12308), .ZN(n7374) );
  NAND2HSV2 U8333 ( .A1(n7962), .A2(n7961), .ZN(n7963) );
  NAND2HSV0 U8334 ( .A1(\pe1/aot [6]), .A2(\pe1/bq[7] ), .ZN(n10252) );
  NAND2HSV0 U8335 ( .A1(\pe1/aot [6]), .A2(n14502), .ZN(n10218) );
  CLKNAND2HSV2 U8336 ( .A1(\pe1/aot [6]), .A2(\pe1/bq[3] ), .ZN(n13965) );
  NAND2HSV2 U8337 ( .A1(n8819), .A2(n8818), .ZN(n8820) );
  CLKNAND2HSV2 U8338 ( .A1(n8822), .A2(n8821), .ZN(n8823) );
  NAND2HSV4 U8339 ( .A1(n10640), .A2(n10638), .ZN(n7710) );
  INHSV4 U8340 ( .I(n7710), .ZN(n7709) );
  BUFHSV2 U8341 ( .I(n13859), .Z(n6702) );
  CLKXOR2HSV4 U8342 ( .A1(n10247), .A2(n10246), .Z(n10248) );
  AOI21HSV0 U8343 ( .A1(n14000), .A2(n10238), .B(n10237), .ZN(n10239) );
  NOR2HSV0 U8344 ( .A1(n10255), .A2(n10633), .ZN(n10256) );
  INAND2HSV4 U8345 ( .A1(n10266), .B1(n10265), .ZN(n10275) );
  INHSV4 U8346 ( .I(n10264), .ZN(n10265) );
  NOR2HSV2 U8347 ( .A1(n13258), .A2(n10634), .ZN(n8028) );
  OAI21HSV2 U8348 ( .A1(n13256), .A2(\pe1/ti_7[5] ), .B(n7713), .ZN(n7712) );
  INHSV2 U8349 ( .I(n10275), .ZN(n10267) );
  XOR2HSV0 U8350 ( .A1(n7152), .A2(n7150), .Z(\pe8/poht [6]) );
  NAND2HSV4 U8351 ( .A1(n11563), .A2(n7289), .ZN(n14857) );
  INHSV4 U8352 ( .I(n9638), .ZN(n9641) );
  XNOR2HSV1 U8353 ( .A1(n6756), .A2(n6755), .ZN(\pe4/poht [7]) );
  NAND2HSV2 U8354 ( .A1(\pe1/ti_7[7] ), .A2(\pe1/got [4]), .ZN(n12860) );
  NAND2HSV2 U8355 ( .A1(n14703), .A2(\pe1/ti_7[7] ), .ZN(n8825) );
  NAND2HSV4 U8356 ( .A1(n7709), .A2(n10639), .ZN(\pe1/ti_7[7] ) );
  NAND2HSV4 U8357 ( .A1(n11587), .A2(n11585), .ZN(n11589) );
  NAND2HSV4 U8358 ( .A1(n6747), .A2(n6746), .ZN(n7776) );
  NAND2HSV4 U8359 ( .A1(\pe4/bq[6] ), .A2(\pe4/aot [8]), .ZN(n9614) );
  NAND2HSV4 U8360 ( .A1(n9621), .A2(n9620), .ZN(n9622) );
  NAND2HSV4 U8361 ( .A1(n13315), .A2(\pe19/got [2]), .ZN(n6790) );
  CLKNAND2HSV2 U8362 ( .A1(n12603), .A2(n11284), .ZN(n14850) );
  CLKNHSV0 U8363 ( .I(n12791), .ZN(n12816) );
  XOR2HSV4 U8364 ( .A1(n11536), .A2(n7281), .Z(n6703) );
  CLKAND2HSV4 U8365 ( .A1(n7280), .A2(n15267), .Z(n11588) );
  OAI21HSV2 U8366 ( .A1(n8165), .A2(n8166), .B(n8167), .ZN(n8168) );
  OAI21HSV2 U8367 ( .A1(n8169), .A2(n8170), .B(n8171), .ZN(po9) );
  CLKNAND2HSV2 U8368 ( .A1(n8169), .A2(n8170), .ZN(n8171) );
  XNOR2HSV4 U8369 ( .A1(n8168), .A2(n7367), .ZN(n8169) );
  XNOR2HSV4 U8370 ( .A1(n10299), .A2(n10298), .ZN(n10304) );
  XNOR2HSV4 U8371 ( .A1(n10304), .A2(n10303), .ZN(n10305) );
  OAI21HSV2 U8372 ( .A1(n8821), .A2(n8822), .B(n8823), .ZN(n8824) );
  XNOR2HSV2 U8373 ( .A1(n12813), .A2(n12812), .ZN(n12814) );
  XOR2HSV4 U8374 ( .A1(n10315), .A2(n10314), .Z(n6704) );
  AOI21HSV2 U8375 ( .A1(n11592), .A2(n11775), .B(n7770), .ZN(n6745) );
  NAND2HSV0 U8376 ( .A1(n8166), .A2(n8165), .ZN(n8167) );
  AND2HSV4 U8377 ( .A1(n7157), .A2(n8903), .Z(n11467) );
  BUFHSV6 U8378 ( .I(n11492), .Z(n14952) );
  NAND2HSV0 U8379 ( .A1(n11492), .A2(n11473), .ZN(n7383) );
  NAND2HSV4 U8380 ( .A1(n7385), .A2(n7384), .ZN(n11492) );
  XOR2HSV0 U8381 ( .A1(n13638), .A2(n6705), .Z(\pe7/poht [1]) );
  XOR2HSV0 U8382 ( .A1(n6860), .A2(n6857), .Z(n6705) );
  CLKNAND2HSV2 U8383 ( .A1(n13605), .A2(n14829), .ZN(n13638) );
  AOI21HSV2 U8384 ( .A1(n6953), .A2(n10331), .B(n6952), .ZN(n7107) );
  CLKNAND2HSV4 U8385 ( .A1(n11520), .A2(n11519), .ZN(n11596) );
  CLKNAND2HSV2 U8386 ( .A1(n11711), .A2(n11710), .ZN(n11539) );
  INHSV4 U8387 ( .I(n10353), .ZN(n10351) );
  XNOR2HSV4 U8388 ( .A1(n10350), .A2(n10349), .ZN(n10353) );
  XNOR2HSV4 U8389 ( .A1(n13311), .A2(n13310), .ZN(\pe5/poht [2]) );
  XOR2HSV4 U8390 ( .A1(n13309), .A2(n13308), .Z(n13310) );
  XNOR2HSV4 U8391 ( .A1(n9540), .A2(n11777), .ZN(n9515) );
  NAND2HSV2 U8392 ( .A1(n13236), .A2(\pe15/got [4]), .ZN(n8657) );
  XNOR2HSV2 U8393 ( .A1(n13433), .A2(n13432), .ZN(n13434) );
  NAND2HSV2 U8394 ( .A1(n14179), .A2(\pe6/got [1]), .ZN(n7007) );
  NAND2HSV2 U8395 ( .A1(n7107), .A2(n7381), .ZN(n12811) );
  NAND2HSV2 U8396 ( .A1(n12786), .A2(n12774), .ZN(n7244) );
  NAND3HSV2 U8397 ( .A1(n12787), .A2(n12786), .A3(n12785), .ZN(n12788) );
  NAND3HSV4 U8398 ( .A1(n6759), .A2(n6758), .A3(n6757), .ZN(n6706) );
  INHSV4 U8399 ( .I(n6765), .ZN(n6757) );
  NAND2HSV2 U8400 ( .A1(\pe5/bq[7] ), .A2(\pe5/aot [7]), .ZN(n7085) );
  NAND2HSV4 U8401 ( .A1(n13840), .A2(n6987), .ZN(n10067) );
  INHSV4 U8402 ( .I(n7025), .ZN(n13840) );
  NAND2HSV4 U8403 ( .A1(n10068), .A2(n10067), .ZN(n10065) );
  CLKNAND2HSV2 U8404 ( .A1(n13855), .A2(n10313), .ZN(n7384) );
  XOR2HSV0 U8405 ( .A1(n7640), .A2(n7633), .Z(\pe19/poht [1]) );
  NAND3HSV4 U8406 ( .A1(n12601), .A2(n12600), .A3(n12599), .ZN(n12612) );
  XNOR2HSV4 U8407 ( .A1(n7557), .A2(n7556), .ZN(n7555) );
  CLKNAND2HSV2 U8408 ( .A1(n7555), .A2(n7558), .ZN(n7554) );
  NAND2HSV0 U8409 ( .A1(n13406), .A2(\pe5/got [2]), .ZN(n7257) );
  NAND2HSV2 U8410 ( .A1(n8755), .A2(n8754), .ZN(n8756) );
  NAND2HSV2 U8411 ( .A1(n15181), .A2(\pe4/got [7]), .ZN(n7835) );
  NAND2HSV2 U8412 ( .A1(n14132), .A2(\pe10/got [1]), .ZN(n7704) );
  XOR2HSV0 U8413 ( .A1(n7740), .A2(n6708), .Z(\pe21/poht [6]) );
  CLKXOR2HSV2 U8414 ( .A1(n7739), .A2(n10872), .Z(n6708) );
  NAND2HSV2 U8415 ( .A1(n6731), .A2(n13718), .ZN(n7557) );
  OAI21HSV0 U8416 ( .A1(n14827), .A2(n11176), .B(n7515), .ZN(n6709) );
  OAI21HSV2 U8417 ( .A1(n14827), .A2(n11176), .B(n7515), .ZN(n7517) );
  NAND2HSV4 U8418 ( .A1(n14068), .A2(n14067), .ZN(n14072) );
  OAI21HSV2 U8419 ( .A1(n8866), .A2(n8867), .B(n8868), .ZN(n8869) );
  OAI21HSV2 U8420 ( .A1(n8869), .A2(n8870), .B(n8871), .ZN(n8872) );
  CLKNAND2HSV2 U8421 ( .A1(n8869), .A2(n8870), .ZN(n8871) );
  INHSV2 U8422 ( .I(n15081), .ZN(n12942) );
  NAND2HSV2 U8423 ( .A1(n7394), .A2(n12277), .ZN(n15081) );
  CLKNAND2HSV2 U8424 ( .A1(n7107), .A2(n7381), .ZN(n6710) );
  INHSV4 U8425 ( .I(n7185), .ZN(n7183) );
  NAND3HSV3 U8426 ( .A1(n10640), .A2(n10639), .A3(n10638), .ZN(n8947) );
  XNOR2HSV1 U8427 ( .A1(n12663), .A2(n7835), .ZN(\pe4/poht [1]) );
  NAND2HSV4 U8428 ( .A1(n13257), .A2(n7711), .ZN(n10640) );
  XNOR2HSV2 U8429 ( .A1(n9448), .A2(n9741), .ZN(n7312) );
  XNOR2HSV4 U8430 ( .A1(n10306), .A2(n10305), .ZN(n10315) );
  AOI21HSV2 U8431 ( .A1(n10328), .A2(n6704), .B(n10327), .ZN(n10329) );
  NAND2HSV4 U8432 ( .A1(n7824), .A2(n7823), .ZN(\pe10/ti_7[6] ) );
  NAND2HSV4 U8433 ( .A1(n7431), .A2(n10729), .ZN(\pe12/ti_7[1] ) );
  AND3HSV2 U8434 ( .A1(n12787), .A2(n12773), .A3(n12786), .Z(n13014) );
  CLKNAND2HSV2 U8435 ( .A1(n8857), .A2(n8856), .ZN(n8858) );
  CLKNAND2HSV2 U8436 ( .A1(n12824), .A2(n12823), .ZN(n12825) );
  NAND2HSV2 U8437 ( .A1(n10227), .A2(n10226), .ZN(n10230) );
  XNOR2HSV4 U8438 ( .A1(n10241), .A2(n10240), .ZN(n10247) );
  XOR2HSV0 U8439 ( .A1(n12448), .A2(n12447), .Z(n6711) );
  NAND3HSV2 U8440 ( .A1(n7243), .A2(n7242), .A3(n12776), .ZN(n7241) );
  NAND2HSV2 U8441 ( .A1(n12776), .A2(n12787), .ZN(n13305) );
  CLKNAND2HSV2 U8442 ( .A1(n12776), .A2(n12775), .ZN(n13012) );
  NAND2HSV0 U8443 ( .A1(n12777), .A2(n10307), .ZN(n12782) );
  CLKNAND2HSV4 U8444 ( .A1(n9457), .A2(n9462), .ZN(n15184) );
  NAND2HSV2 U8445 ( .A1(n14709), .A2(\pe20/got [6]), .ZN(n8755) );
  NAND2HSV2 U8446 ( .A1(n14709), .A2(\pe20/got [1]), .ZN(n7496) );
  NAND2HSV4 U8447 ( .A1(n12041), .A2(n12040), .ZN(n13875) );
  XOR2HSV1 U8448 ( .A1(poh21[7]), .A2(n8474), .Z(po[8]) );
  NAND2HSV2 U8449 ( .A1(\pe5/pvq [3]), .A2(\pe5/ctrq ), .ZN(n7088) );
  NAND3HSV2 U8450 ( .A1(n7241), .A2(n13304), .A3(n7240), .ZN(n7239) );
  MAOI22HSV2 U8451 ( .A1(n14131), .A2(n14130), .B1(n14129), .B2(n14128), .ZN(
        n14153) );
  XNOR2HSV2 U8452 ( .A1(n14155), .A2(n14154), .ZN(n14156) );
  CLKNHSV0 U8453 ( .I(n14924), .ZN(n6713) );
  INHSV2 U8454 ( .I(n11441), .ZN(n7572) );
  INHSV4 U8455 ( .I(n7338), .ZN(n7129) );
  NAND2HSV2 U8456 ( .A1(n10401), .A2(n9398), .ZN(n10388) );
  NAND2HSV2 U8457 ( .A1(n15192), .A2(\pe12/got [7]), .ZN(n7443) );
  AOI21HSV2 U8458 ( .A1(n11906), .A2(n7335), .B(n11905), .ZN(n11907) );
  XOR2HSV4 U8459 ( .A1(n10857), .A2(n7531), .Z(n7530) );
  AOI21HSV2 U8460 ( .A1(n7050), .A2(n7053), .B(n7047), .ZN(n7732) );
  AOI21HSV2 U8461 ( .A1(n11010), .A2(n11016), .B(n7003), .ZN(n7002) );
  NOR2HSV2 U8462 ( .A1(n11016), .A2(n11017), .ZN(n7005) );
  NAND2HSV2 U8463 ( .A1(\pe21/ti_7[5] ), .A2(\pe21/got [2]), .ZN(n7406) );
  NAND2HSV2 U8464 ( .A1(n10764), .A2(n10765), .ZN(n14255) );
  NAND2HSV4 U8465 ( .A1(n11711), .A2(n11710), .ZN(n14196) );
  NAND2HSV2 U8466 ( .A1(n11539), .A2(\pe8/got [7]), .ZN(n7179) );
  OAI22HSV4 U8467 ( .A1(n14074), .A2(n14073), .B1(n14075), .B2(n14072), .ZN(
        n14079) );
  INHSV2 U8468 ( .I(n7456), .ZN(n6714) );
  CLKNAND2HSV2 U8469 ( .A1(n7302), .A2(\pe6/got [1]), .ZN(n6914) );
  NAND2HSV4 U8470 ( .A1(n7302), .A2(n7762), .ZN(n7761) );
  NAND2HSV4 U8471 ( .A1(n9847), .A2(n7764), .ZN(n7302) );
  XNOR2HSV4 U8472 ( .A1(n6914), .A2(n13934), .ZN(n6913) );
  NAND2HSV2 U8473 ( .A1(n8150), .A2(n8149), .ZN(n8151) );
  XNOR2HSV4 U8474 ( .A1(n10219), .A2(n10218), .ZN(n10220) );
  NAND2HSV4 U8475 ( .A1(n7154), .A2(n11416), .ZN(n7204) );
  NAND2HSV0 U8476 ( .A1(n14546), .A2(\pe18/pvq [7]), .ZN(n11983) );
  NAND2HSV0 U8477 ( .A1(n14546), .A2(\pe18/pq ), .ZN(n13153) );
  CKMUX2HSV2 U8478 ( .I0(bo18[6]), .I1(\pe18/bq[6] ), .S(n14546), .Z(n15017)
         );
  INHSV4 U8479 ( .I(n10802), .ZN(n14546) );
  XNOR2HSV4 U8480 ( .A1(n9189), .A2(n9188), .ZN(n9191) );
  INHSV4 U8481 ( .I(n7054), .ZN(n6989) );
  INHSV2 U8482 ( .I(n9946), .ZN(n7622) );
  MUX2NHSV2 U8483 ( .I0(n12224), .I1(n12223), .S(n8902), .ZN(n12227) );
  CLKNAND2HSV4 U8484 ( .A1(n7187), .A2(n7189), .ZN(n7186) );
  NAND2HSV2 U8485 ( .A1(n9129), .A2(n10586), .ZN(n9118) );
  XNOR2HSV4 U8486 ( .A1(n6905), .A2(n6902), .ZN(n9639) );
  CLKNAND2HSV4 U8487 ( .A1(n12271), .A2(n9712), .ZN(n9713) );
  XOR2HSV0 U8488 ( .A1(n10455), .A2(n10454), .Z(n6716) );
  CLKXOR2HSV4 U8489 ( .A1(n10453), .A2(n10452), .Z(n10454) );
  OAI21HSV2 U8490 ( .A1(n8256), .A2(n8257), .B(n8258), .ZN(n8259) );
  OAI21HSV2 U8491 ( .A1(n8259), .A2(n8260), .B(n8261), .ZN(n8262) );
  CLKAND2HSV4 U8492 ( .A1(n8430), .A2(n7507), .Z(n6717) );
  NAND3HSV3 U8493 ( .A1(n11589), .A2(n11594), .A3(n11595), .ZN(n11775) );
  CLKXOR2HSV4 U8494 ( .A1(n10895), .A2(n10894), .Z(n10896) );
  XNOR2HSV4 U8495 ( .A1(n10897), .A2(n10896), .ZN(n10898) );
  AOI21HSV0 U8496 ( .A1(n8925), .A2(\pe6/pvq [5]), .B(\pe6/phq [5]), .ZN(n8727) );
  CLKXOR2HSV2 U8497 ( .A1(n12469), .A2(n12468), .Z(n12471) );
  CLKXOR2HSV2 U8498 ( .A1(n12571), .A2(n12570), .Z(n12573) );
  OAI21HSV2 U8499 ( .A1(n9454), .A2(n9748), .B(n9453), .ZN(n7311) );
  CLKXOR2HSV2 U8500 ( .A1(n12451), .A2(n12450), .Z(n12455) );
  NOR2HSV8 U8501 ( .A1(n11336), .A2(n11337), .ZN(n6732) );
  XOR2HSV2 U8502 ( .A1(n7597), .A2(n6718), .Z(n8237) );
  AND2HSV4 U8503 ( .A1(n7595), .A2(n7593), .Z(n6718) );
  CLKAND2HSV2 U8504 ( .A1(n7631), .A2(n12103), .Z(n6719) );
  CLKNHSV0 U8505 ( .I(n14397), .ZN(n12103) );
  NAND2HSV2 U8506 ( .A1(n6710), .A2(\pe5/got [6]), .ZN(n7111) );
  AND2HSV4 U8507 ( .A1(n10527), .A2(n11473), .Z(n8904) );
  NAND2HSV2 U8508 ( .A1(n8501), .A2(n8500), .ZN(n8502) );
  CLKNAND2HSV4 U8509 ( .A1(n7411), .A2(n9070), .ZN(n9057) );
  CLKXOR2HSV4 U8510 ( .A1(n10480), .A2(n10479), .Z(n10481) );
  NAND2HSV4 U8511 ( .A1(n11588), .A2(n13862), .ZN(n11594) );
  OAI21HSV2 U8512 ( .A1(n8352), .A2(n8353), .B(n8354), .ZN(n8355) );
  OAI21HSV2 U8513 ( .A1(n8355), .A2(n8356), .B(n8357), .ZN(n8358) );
  NAND2HSV2 U8514 ( .A1(n9982), .A2(n9977), .ZN(n10000) );
  NAND2HSV2 U8515 ( .A1(n15262), .A2(n10070), .ZN(n6927) );
  OAI21HSV2 U8516 ( .A1(n8581), .A2(n8582), .B(n8583), .ZN(n8584) );
  INHSV4 U8517 ( .I(n7365), .ZN(n7362) );
  CLKNAND2HSV2 U8518 ( .A1(n6795), .A2(n6794), .ZN(n13749) );
  NAND2HSV2 U8519 ( .A1(n14077), .A2(n14072), .ZN(n14074) );
  NOR2HSV4 U8520 ( .A1(n14079), .A2(n14078), .ZN(n14102) );
  NAND2HSV2 U8521 ( .A1(n7186), .A2(n7185), .ZN(n15276) );
  OAI21HSV2 U8522 ( .A1(n8566), .A2(n8567), .B(n8568), .ZN(n8569) );
  NAND2HSV2 U8523 ( .A1(\pe3/ti_7[5] ), .A2(\pe3/got [3]), .ZN(n8567) );
  NAND2HSV2 U8524 ( .A1(n8567), .A2(n8566), .ZN(n8568) );
  NAND2HSV0 U8525 ( .A1(n8570), .A2(n8569), .ZN(n8571) );
  NAND2HSV4 U8526 ( .A1(n7493), .A2(n7494), .ZN(n15248) );
  XNOR2HSV4 U8527 ( .A1(n9164), .A2(n9163), .ZN(n9169) );
  NAND2HSV2 U8528 ( .A1(\pe7/ti_1 ), .A2(\pe7/got [4]), .ZN(n7961) );
  NAND2HSV2 U8529 ( .A1(n7937), .A2(n10121), .ZN(n6884) );
  AND2HSV4 U8530 ( .A1(n10121), .A2(n10924), .Z(n8908) );
  NAND3HSV2 U8531 ( .A1(n9763), .A2(n9434), .A3(n9741), .ZN(n6940) );
  CLKNAND2HSV2 U8532 ( .A1(n10047), .A2(n10052), .ZN(n7237) );
  NAND2HSV0 U8533 ( .A1(n11777), .A2(\pe19/got [4]), .ZN(n12166) );
  INHSV4 U8534 ( .I(n7491), .ZN(n7490) );
  XNOR2HSV1 U8535 ( .A1(n11643), .A2(n11642), .ZN(n7882) );
  AOI21HSV2 U8536 ( .A1(n11342), .A2(n11341), .B(n11340), .ZN(n11373) );
  CLKXOR2HSV2 U8537 ( .A1(n12653), .A2(n12652), .Z(n12654) );
  IAO21HSV4 U8538 ( .A1(n15233), .A2(n12829), .B(n6720), .ZN(n6733) );
  OR2HSV2 U8539 ( .A1(n12335), .A2(n12513), .Z(n6720) );
  INHSV4 U8540 ( .I(n12878), .ZN(n6721) );
  XNOR2HSV4 U8541 ( .A1(n7074), .A2(n7069), .ZN(n8228) );
  NAND2HSV2 U8542 ( .A1(n9083), .A2(n9082), .ZN(n6729) );
  AOI21HSV2 U8543 ( .A1(n7357), .A2(n7355), .B(n7354), .ZN(n7686) );
  XNOR2HSV1 U8544 ( .A1(n11327), .A2(n13864), .ZN(n13867) );
  NOR2HSV2 U8545 ( .A1(n13864), .A2(n11317), .ZN(n11361) );
  NOR2HSV2 U8546 ( .A1(n13864), .A2(n11327), .ZN(n11331) );
  CLKNAND2HSV8 U8547 ( .A1(n11610), .A2(n7506), .ZN(n15190) );
  NOR2HSV0 U8548 ( .A1(n14492), .A2(n11042), .ZN(n11044) );
  XOR2HSV4 U8549 ( .A1(n13136), .A2(n13137), .Z(n8856) );
  CLKXOR2HSV4 U8550 ( .A1(n13135), .A2(n13134), .Z(n13136) );
  AOI21HSV4 U8551 ( .A1(n10839), .A2(n7724), .B(n7723), .ZN(n7728) );
  OAI21HSV4 U8552 ( .A1(n7721), .A2(n10839), .B(n10838), .ZN(n7723) );
  CLKNHSV0 U8553 ( .I(n11791), .ZN(n6723) );
  NAND2HSV2 U8554 ( .A1(\pe21/aot [6]), .A2(\pe21/bq[7] ), .ZN(n7671) );
  NAND2HSV2 U8555 ( .A1(\pe21/aot [7]), .A2(\pe21/bq[7] ), .ZN(n7657) );
  INHSV4 U8556 ( .I(n10174), .ZN(n10177) );
  CLKNAND2HSV4 U8557 ( .A1(n11238), .A2(n11237), .ZN(n13759) );
  NAND2HSV2 U8558 ( .A1(\pe10/bq[4] ), .A2(\pe10/aot [8]), .ZN(n6963) );
  MUX2NHSV1 U8559 ( .I0(n8912), .I1(n9241), .S(n9240), .ZN(n6725) );
  NOR2HSV4 U8560 ( .A1(n9246), .A2(n9247), .ZN(n6726) );
  MUX2NHSV1 U8561 ( .I0(n8912), .I1(n9241), .S(n9240), .ZN(n9304) );
  OAI21HSV4 U8562 ( .A1(n9304), .A2(n6773), .B(n9243), .ZN(n9247) );
  NOR2HSV0 U8563 ( .A1(n11902), .A2(n11901), .ZN(n11906) );
  BUFHSV4 U8564 ( .I(n9783), .Z(n14896) );
  MUX2NHSV4 U8565 ( .I0(n11892), .I1(n11893), .S(n6727), .ZN(n13681) );
  CLKXOR2HSV4 U8566 ( .A1(n11891), .A2(n11890), .Z(n6727) );
  CLKNHSV0 U8567 ( .I(n8508), .ZN(n7390) );
  CLKNAND2HSV2 U8568 ( .A1(n6943), .A2(n6942), .ZN(n10442) );
  CLKNHSV0 U8569 ( .I(n12253), .ZN(n7458) );
  OAI31HSV0 U8570 ( .A1(n13401), .A2(n8701), .A3(n8698), .B(n8702), .ZN(n8703)
         );
  OAI21HSV0 U8571 ( .A1(n13401), .A2(n8698), .B(n8701), .ZN(n8702) );
  XNOR2HSV4 U8572 ( .A1(n13403), .A2(n13402), .ZN(n13404) );
  MUX2NHSV1 U8573 ( .I0(n13648), .I1(n13647), .S(n6775), .ZN(n13650) );
  NAND2HSV4 U8574 ( .A1(n15184), .A2(n11880), .ZN(n6775) );
  OAI21HSV2 U8575 ( .A1(n8749), .A2(n8748), .B(n8750), .ZN(n8751) );
  CLKNHSV0 U8576 ( .I(n9265), .ZN(n9269) );
  INHSV2 U8577 ( .I(\pe10/got [7]), .ZN(n7653) );
  NAND2HSV2 U8578 ( .A1(n14125), .A2(\pe10/got [7]), .ZN(n7714) );
  INHSV4 U8579 ( .I(n10598), .ZN(n6793) );
  AOI21HSV2 U8580 ( .A1(n6760), .A2(n7425), .B(n12106), .ZN(n7421) );
  NAND2HSV2 U8581 ( .A1(\pe13/bq[6] ), .A2(\pe13/aot [8]), .ZN(n7585) );
  INAND2HSV2 U8582 ( .A1(n10944), .B1(n7870), .ZN(n7541) );
  AO22HSV2 U8583 ( .A1(n12146), .A2(n11713), .B1(n12141), .B2(n11712), .Z(
        n15210) );
  OAI21HSV0 U8584 ( .A1(n8625), .A2(n8624), .B(n8626), .ZN(n8627) );
  MUX2NHSV1 U8585 ( .I0(n12234), .I1(n8842), .S(n8845), .ZN(n12218) );
  OAI21HSV2 U8586 ( .A1(n8085), .A2(n11115), .B(n7852), .ZN(n7851) );
  XNOR2HSV4 U8587 ( .A1(n11421), .A2(n14243), .ZN(n11429) );
  NAND2HSV2 U8588 ( .A1(\pe15/aot [7]), .A2(\pe15/bq[7] ), .ZN(n7347) );
  XOR2HSV0 U8589 ( .A1(n12990), .A2(n6728), .Z(\pe6/poht [5]) );
  CLKXOR2HSV2 U8590 ( .A1(n12989), .A2(n12988), .Z(n6728) );
  NAND2HSV2 U8591 ( .A1(n6830), .A2(\pe12/got [4]), .ZN(n7319) );
  NAND2HSV2 U8592 ( .A1(n11390), .A2(n10521), .ZN(n11291) );
  MUX2NHSV2 U8593 ( .I0(n8643), .I1(n10589), .S(n8644), .ZN(n10585) );
  OAI21HSV2 U8594 ( .A1(n8342), .A2(n8343), .B(n8344), .ZN(n8345) );
  NAND2HSV2 U8595 ( .A1(n8343), .A2(n8342), .ZN(n8344) );
  NAND2HSV2 U8596 ( .A1(n8346), .A2(n8345), .ZN(n8347) );
  CLKNAND2HSV4 U8597 ( .A1(n9103), .A2(n9080), .ZN(n9083) );
  XNOR2HSV4 U8598 ( .A1(n13549), .A2(n13548), .ZN(n13550) );
  CLKNAND2HSV2 U8599 ( .A1(n13874), .A2(n12042), .ZN(n12044) );
  OAI21HSV2 U8600 ( .A1(n14740), .A2(n12132), .B(n8212), .ZN(n8214) );
  XNOR2HSV4 U8601 ( .A1(n10952), .A2(n10951), .ZN(n10960) );
  XNOR2HSV4 U8602 ( .A1(n13369), .A2(n13368), .ZN(n13370) );
  NAND2HSV0 U8603 ( .A1(n12260), .A2(n9450), .ZN(n7015) );
  CLKNAND2HSV2 U8604 ( .A1(n14805), .A2(\pe2/pvq [4]), .ZN(n8553) );
  CLKNHSV0 U8605 ( .I(n13881), .ZN(n6730) );
  NAND2HSV2 U8606 ( .A1(n7360), .A2(n10407), .ZN(n7359) );
  NAND2HSV4 U8607 ( .A1(n10404), .A2(n7324), .ZN(n7805) );
  OAI21HSV2 U8608 ( .A1(n8802), .A2(n8803), .B(n8804), .ZN(n8805) );
  NAND2HSV2 U8609 ( .A1(n7302), .A2(\pe6/got [5]), .ZN(n8803) );
  XNOR2HSV4 U8610 ( .A1(n7608), .A2(n7609), .ZN(n8331) );
  AOI21HSV2 U8611 ( .A1(n12078), .A2(n12077), .B(n8737), .ZN(n8738) );
  IOA22HSV1 U8612 ( .B1(n12078), .B2(n12077), .A1(n12267), .A2(n8905), .ZN(
        n8737) );
  NAND2HSV4 U8613 ( .A1(n8738), .A2(n7363), .ZN(n12265) );
  NAND2HSV0 U8614 ( .A1(n8637), .A2(n8636), .ZN(n8638) );
  CLKNHSV0 U8615 ( .I(n12264), .ZN(n12199) );
  CLKNAND2HSV2 U8616 ( .A1(n12060), .A2(n12059), .ZN(n12232) );
  NAND2HSV4 U8617 ( .A1(n12680), .A2(n12679), .ZN(n14959) );
  NAND3HSV2 U8618 ( .A1(n9727), .A2(n9725), .A3(n9722), .ZN(n7401) );
  NOR2HSV2 U8619 ( .A1(n9727), .A2(n9725), .ZN(n7402) );
  NOR2HSV2 U8620 ( .A1(n9725), .A2(n9722), .ZN(n7400) );
  INAND2HSV2 U8621 ( .A1(n8231), .B1(n13603), .ZN(n7594) );
  NAND2HSV2 U8622 ( .A1(n15182), .A2(\pe8/got [1]), .ZN(n7151) );
  CLKNAND2HSV2 U8623 ( .A1(n14381), .A2(n15179), .ZN(n7685) );
  NAND2HSV4 U8624 ( .A1(n9608), .A2(n9607), .ZN(n14381) );
  NOR2HSV4 U8625 ( .A1(n7498), .A2(n7499), .ZN(n11902) );
  NAND2HSV2 U8626 ( .A1(n11742), .A2(n7501), .ZN(n7498) );
  OAI21HSV2 U8627 ( .A1(n6771), .A2(n11136), .B(n11135), .ZN(n11139) );
  INHSV2 U8628 ( .I(n11139), .ZN(n11137) );
  CLKNAND2HSV4 U8629 ( .A1(n12259), .A2(n12258), .ZN(n15189) );
  AOI21HSV2 U8630 ( .A1(n12102), .A2(n12107), .B(n13872), .ZN(n12042) );
  NAND2HSV4 U8631 ( .A1(n15255), .A2(n11943), .ZN(n12193) );
  INHSV8 U8632 ( .I(n13832), .ZN(n14570) );
  NAND2HSV4 U8633 ( .A1(n11215), .A2(n11214), .ZN(n15186) );
  NAND2HSV0 U8634 ( .A1(n8881), .A2(n13871), .ZN(n8882) );
  NAND3HSV2 U8635 ( .A1(n11213), .A2(n13871), .A3(n14066), .ZN(n11214) );
  OAI21HSV2 U8636 ( .A1(n7673), .A2(n12347), .B(n11744), .ZN(n7672) );
  INAND2HSV2 U8637 ( .A1(n7722), .B1(n6207), .ZN(n12542) );
  AOI21HSV2 U8638 ( .A1(n10836), .A2(n7725), .B(n10403), .ZN(n7724) );
  NAND2HSV0 U8639 ( .A1(\pe5/ti_7[7] ), .A2(\pe5/got [4]), .ZN(n8637) );
  NAND3HSV2 U8640 ( .A1(n7212), .A2(\pe5/ctrq ), .A3(\pe5/pvq [2]), .ZN(n7211)
         );
  NAND2HSV4 U8641 ( .A1(\pe5/pvq [2]), .A2(\pe5/ctrq ), .ZN(n7208) );
  INAND2HSV2 U8642 ( .A1(n13012), .B1(n13014), .ZN(n7065) );
  NAND3HSV4 U8643 ( .A1(n10377), .A2(n10376), .A3(n10375), .ZN(n10378) );
  CLKNAND2HSV4 U8644 ( .A1(n10367), .A2(n10366), .ZN(n10377) );
  CLKNAND2HSV2 U8645 ( .A1(n7390), .A2(n9419), .ZN(n6942) );
  NAND3HSV2 U8646 ( .A1(n11770), .A2(n11769), .A3(n11768), .ZN(n8505) );
  NAND2HSV2 U8647 ( .A1(n15085), .A2(n13797), .ZN(n8857) );
  NAND2HSV2 U8648 ( .A1(n7513), .A2(n7512), .ZN(n11178) );
  NAND2HSV2 U8649 ( .A1(n7512), .A2(n7516), .ZN(n7511) );
  NAND2HSV4 U8650 ( .A1(n6856), .A2(n6855), .ZN(n14365) );
  NAND2HSV0 U8651 ( .A1(n14365), .A2(\pe11/got [5]), .ZN(n12448) );
  NAND2HSV2 U8652 ( .A1(n14365), .A2(\pe11/got [6]), .ZN(n6854) );
  XOR2HSV0 U8653 ( .A1(n9158), .A2(n9157), .Z(n9159) );
  NAND2HSV2 U8654 ( .A1(\pe18/ti_7[1] ), .A2(\pe18/got [5]), .ZN(n7542) );
  NAND2HSV4 U8655 ( .A1(n6791), .A2(n10598), .ZN(n6794) );
  CLKNHSV0 U8656 ( .I(n12036), .ZN(n12031) );
  NAND2HSV2 U8657 ( .A1(n7104), .A2(n10715), .ZN(n7103) );
  NAND2HSV2 U8658 ( .A1(\pe17/pvq [3]), .A2(\pe17/ctrq ), .ZN(n6975) );
  NAND2HSV4 U8659 ( .A1(n10071), .A2(n7446), .ZN(n15075) );
  NAND2HSV4 U8660 ( .A1(n9932), .A2(n9931), .ZN(n13587) );
  NOR2HSV0 U8661 ( .A1(n7813), .A2(n7356), .ZN(n7355) );
  CLKNAND2HSV2 U8662 ( .A1(n7813), .A2(n9832), .ZN(n7467) );
  NOR2HSV2 U8663 ( .A1(n12602), .A2(n7841), .ZN(n7840) );
  OAI21HSV2 U8664 ( .A1(n12276), .A2(n7397), .B(n7395), .ZN(n12305) );
  CLKAND2HSV2 U8665 ( .A1(n12276), .A2(n12252), .Z(n7459) );
  NOR2HSV4 U8666 ( .A1(n13695), .A2(n11877), .ZN(n11886) );
  NAND3HSV2 U8667 ( .A1(n7368), .A2(n7370), .A3(n6935), .ZN(n6934) );
  NAND2HSV0 U8668 ( .A1(n14914), .A2(\pe15/got [3]), .ZN(n7695) );
  NOR2HSV2 U8669 ( .A1(n11336), .A2(n11337), .ZN(n11407) );
  NOR2HSV0 U8670 ( .A1(n6732), .A2(n7337), .ZN(n7336) );
  XNOR2HSV4 U8671 ( .A1(n13088), .A2(n13087), .ZN(n13091) );
  INAND2HSV2 U8672 ( .A1(n7598), .B1(n14961), .ZN(n8238) );
  NAND2HSV4 U8673 ( .A1(n11969), .A2(n11968), .ZN(n13604) );
  CLKNAND2HSV2 U8674 ( .A1(n13406), .A2(\pe5/got [6]), .ZN(n7994) );
  CLKXOR2HSV4 U8675 ( .A1(n13303), .A2(n13302), .Z(n13309) );
  INHSV2 U8676 ( .I(n10585), .ZN(n12595) );
  NAND2HSV2 U8677 ( .A1(n15212), .A2(n9541), .ZN(n7376) );
  MUX2NHSV4 U8678 ( .I0(\pe19/phq [1]), .I1(n7895), .S(n7896), .ZN(n9511) );
  AOI21HSV2 U8679 ( .A1(n10859), .A2(n10858), .B(n7779), .ZN(n8207) );
  NOR2HSV2 U8680 ( .A1(n10858), .A2(n7537), .ZN(n7536) );
  NAND2HSV2 U8681 ( .A1(n7875), .A2(\pe9/got [8]), .ZN(n8170) );
  NAND2HSV2 U8682 ( .A1(n7875), .A2(\pe9/got [2]), .ZN(n11673) );
  NAND2HSV2 U8683 ( .A1(n7875), .A2(\pe9/got [1]), .ZN(n13909) );
  CLKXOR2HSV4 U8684 ( .A1(n11689), .A2(n6734), .Z(n11697) );
  XNOR2HSV4 U8685 ( .A1(n11688), .A2(n11687), .ZN(n6734) );
  XOR2HSV0 U8686 ( .A1(n12005), .A2(n12004), .Z(n6735) );
  OAI31HSV2 U8687 ( .A1(n13809), .A2(n7996), .A3(n13429), .B(n7997), .ZN(n7998) );
  CLKNAND2HSV2 U8688 ( .A1(n7241), .A2(n13304), .ZN(n13809) );
  NAND2HSV2 U8689 ( .A1(n8608), .A2(n8607), .ZN(n8609) );
  BUFHSV6 U8690 ( .I(n7631), .Z(n7039) );
  INHSV2 U8691 ( .I(n6776), .ZN(n7825) );
  NOR2HSV2 U8692 ( .A1(n15261), .A2(n10930), .ZN(n13468) );
  OAI21HSV2 U8693 ( .A1(n15075), .A2(n10784), .B(n10128), .ZN(n6776) );
  NAND2HSV4 U8694 ( .A1(n15075), .A2(n10925), .ZN(n10116) );
  CLKNHSV0 U8695 ( .I(n10123), .ZN(n7661) );
  AOI21HSV0 U8696 ( .A1(n14132), .A2(n10124), .B(n10120), .ZN(n7937) );
  AOI21HSV2 U8697 ( .A1(n7661), .A2(n6701), .B(n7660), .ZN(n7827) );
  NOR2HSV2 U8698 ( .A1(n10124), .A2(ctro10), .ZN(n10107) );
  NAND2HSV2 U8699 ( .A1(n10124), .A2(n10925), .ZN(n6926) );
  NAND2HSV0 U8700 ( .A1(n12387), .A2(n6787), .ZN(n6786) );
  NAND2HSV4 U8701 ( .A1(n12386), .A2(n12385), .ZN(n14862) );
  NAND2HSV4 U8702 ( .A1(n15070), .A2(n11266), .ZN(n9380) );
  INHSV4 U8703 ( .I(n11972), .ZN(n13185) );
  INHSV4 U8704 ( .I(n7749), .ZN(n7272) );
  OAI21HSV2 U8705 ( .A1(n8037), .A2(n9534), .B(n8038), .ZN(n8039) );
  OAI21HSV0 U8706 ( .A1(n13476), .A2(n7700), .B(n7699), .ZN(n7810) );
  OAI21HSV0 U8707 ( .A1(n13476), .A2(n8776), .B(n7702), .ZN(n7699) );
  CLKXOR2HSV4 U8708 ( .A1(n13443), .A2(n13442), .Z(n13445) );
  NAND2HSV2 U8709 ( .A1(n11081), .A2(\pe14/got [7]), .ZN(n9114) );
  NAND2HSV4 U8710 ( .A1(n9744), .A2(n7083), .ZN(n9748) );
  OAI21HSV2 U8711 ( .A1(n9744), .A2(n9790), .B(n9743), .ZN(n7484) );
  AOI31HSV2 U8712 ( .A1(n11523), .A2(n11515), .A3(n11514), .B(n11513), .ZN(
        n7275) );
  IAO22HSV4 U8713 ( .B1(\pe8/ti_7t [5]), .B2(n7934), .A1(n11596), .A2(n11560), 
        .ZN(n11710) );
  CLKNAND2HSV2 U8714 ( .A1(n9537), .A2(n9728), .ZN(n9560) );
  CLKNAND2HSV8 U8715 ( .A1(n6904), .A2(n6903), .ZN(n14733) );
  CLKNAND2HSV4 U8716 ( .A1(n13851), .A2(n9130), .ZN(n6904) );
  MUX2NHSV4 U8717 ( .I0(n8002), .I1(n12416), .S(n7547), .ZN(n7546) );
  NAND2HSV2 U8718 ( .A1(n14061), .A2(\pe2/got [1]), .ZN(n14063) );
  CLKNAND2HSV4 U8719 ( .A1(n11720), .A2(n11944), .ZN(n11740) );
  NAND2HSV2 U8720 ( .A1(n12997), .A2(\pe13/got [5]), .ZN(n7588) );
  NOR2HSV2 U8721 ( .A1(n13401), .A2(n13307), .ZN(n13308) );
  INHSV4 U8722 ( .I(n9071), .ZN(n7411) );
  CLKXOR2HSV4 U8723 ( .A1(n14327), .A2(n14326), .Z(n14330) );
  NAND3HSV3 U8724 ( .A1(n13870), .A2(n13869), .A3(n11183), .ZN(n7125) );
  CLKNAND2HSV4 U8725 ( .A1(n11180), .A2(n7126), .ZN(n13870) );
  NOR2HSV2 U8726 ( .A1(n11606), .A2(n6868), .ZN(n13535) );
  CLKNAND2HSV8 U8727 ( .A1(n7742), .A2(n7741), .ZN(n15085) );
  NAND2HSV4 U8728 ( .A1(n10442), .A2(n10441), .ZN(n9763) );
  NOR2HSV4 U8729 ( .A1(n15262), .A2(n14122), .ZN(n14129) );
  XNOR2HSV4 U8730 ( .A1(n7314), .A2(n7310), .ZN(n6737) );
  MUX2NHSV4 U8731 ( .I0(n14273), .I1(n7885), .S(n7877), .ZN(n7822) );
  XNOR2HSV4 U8732 ( .A1(n9094), .A2(n9093), .ZN(n15176) );
  OAI21HSV4 U8733 ( .A1(n6740), .A2(n6739), .B(n6738), .ZN(n9093) );
  CLKNAND2HSV2 U8734 ( .A1(n9079), .A2(\pe14/phq [1]), .ZN(n6738) );
  CLKNHSV2 U8735 ( .I(\pe14/pvq [1]), .ZN(n6739) );
  CLKNAND2HSV2 U8736 ( .A1(n6741), .A2(\pe14/ctrq ), .ZN(n6740) );
  CLKNHSV2 U8737 ( .I(\pe14/phq [1]), .ZN(n6741) );
  XNOR2HSV4 U8738 ( .A1(n6743), .A2(n6742), .ZN(n9094) );
  CLKNAND2HSV2 U8739 ( .A1(\pe14/aot [8]), .A2(\pe14/bq[8] ), .ZN(n6743) );
  NOR2HSV4 U8740 ( .A1(n7773), .A2(n6744), .ZN(n11606) );
  CLKNAND2HSV2 U8741 ( .A1(n7776), .A2(n6745), .ZN(n6744) );
  CLKNHSV2 U8742 ( .I(n11593), .ZN(n6746) );
  CLKNHSV2 U8743 ( .I(n13878), .ZN(n6747) );
  XNOR2HSV4 U8744 ( .A1(n11607), .A2(n11608), .ZN(n7773) );
  XNOR2HSV4 U8745 ( .A1(n6749), .A2(n6748), .ZN(n11608) );
  XOR3HSV2 U8746 ( .A1(n11584), .A2(n11583), .A3(n11582), .Z(n6748) );
  CLKNAND2HSV2 U8747 ( .A1(n14857), .A2(\pe8/got [6]), .ZN(n6749) );
  AOI21HSV4 U8748 ( .A1(n8008), .A2(n6703), .B(n11513), .ZN(n6751) );
  XOR3HSV2 U8749 ( .A1(n9935), .A2(n9943), .A3(n6753), .Z(n6752) );
  OAI21HSV4 U8750 ( .A1(n8469), .A2(\pe13/phq [6]), .B(n8470), .ZN(n6753) );
  CLKBUFHSV2 U8751 ( .I(n10071), .Z(n6754) );
  OAI21HSV4 U8752 ( .A1(n10119), .A2(n6754), .B(n10118), .ZN(n14132) );
  CLKNHSV2 U8753 ( .I(n13907), .ZN(n6755) );
  CLKNAND2HSV2 U8754 ( .A1(n6766), .A2(n12602), .ZN(n6758) );
  CLKNAND2HSV2 U8755 ( .A1(n7840), .A2(n12595), .ZN(n6759) );
  NAND2HSV4 U8756 ( .A1(n6760), .A2(n6818), .ZN(n6816) );
  NOR2HSV4 U8757 ( .A1(n6763), .A2(n6762), .ZN(n6761) );
  CLKNHSV2 U8758 ( .I(\pe10/got [5]), .ZN(n6762) );
  CLKNAND2HSV3 U8759 ( .A1(n7836), .A2(n6770), .ZN(n6765) );
  INHSV2 U8760 ( .I(n6767), .ZN(n6766) );
  CLKNAND2HSV1 U8761 ( .A1(n10585), .A2(n6768), .ZN(n6767) );
  INHSV2 U8762 ( .I(n6769), .ZN(n6768) );
  INHSV2 U8763 ( .I(n10586), .ZN(n6769) );
  CLKNAND2HSV0 U8764 ( .A1(n15181), .A2(\pe4/got [3]), .ZN(n12088) );
  INHSV2 U8765 ( .I(n12591), .ZN(n6770) );
  XNOR2HSV4 U8766 ( .A1(n11119), .A2(n11118), .ZN(n6771) );
  CLKNAND2HSV4 U8767 ( .A1(n9242), .A2(n9285), .ZN(n6773) );
  CLKNAND2HSV3 U8768 ( .A1(n9802), .A2(\pe6/ti_7t [1]), .ZN(n6772) );
  CLKNHSV4 U8769 ( .I(\pe2/got [4]), .ZN(n6774) );
  NAND3HSV4 U8770 ( .A1(n10069), .A2(n6985), .A3(n10067), .ZN(n7446) );
  CLKNAND2HSV4 U8771 ( .A1(n10066), .A2(n10065), .ZN(n10071) );
  CLKNAND2HSV1 U8772 ( .A1(\pe2/ti_1 ), .A2(\pe2/got [7]), .ZN(n6778) );
  CLKNHSV2 U8773 ( .I(\pe2/got [7]), .ZN(n9360) );
  OAI21HSV4 U8774 ( .A1(n6779), .A2(n6778), .B(n6777), .ZN(n8975) );
  CLKNAND2HSV2 U8775 ( .A1(n6779), .A2(n6778), .ZN(n6777) );
  NOR2HSV4 U8776 ( .A1(n6781), .A2(n6780), .ZN(n6779) );
  CLKNHSV2 U8777 ( .I(\pe2/bq[8] ), .ZN(n6780) );
  CLKNHSV2 U8778 ( .I(\pe2/aot [7]), .ZN(n6781) );
  XNOR2HSV4 U8779 ( .A1(n6790), .A2(n6782), .ZN(\pe19/poht [6]) );
  CLKNAND2HSV2 U8780 ( .A1(n6786), .A2(n6783), .ZN(n6782) );
  CLKNAND2HSV2 U8781 ( .A1(n6784), .A2(n6789), .ZN(n6783) );
  CLKNAND2HSV2 U8782 ( .A1(n13316), .A2(\pe19/got [1]), .ZN(n6784) );
  CLKNHSV2 U8783 ( .I(n12340), .ZN(n6785) );
  NOR2HSV4 U8784 ( .A1(n6789), .A2(n6788), .ZN(n6787) );
  CLKNHSV2 U8785 ( .I(\pe19/got [1]), .ZN(n6788) );
  CLKNHSV2 U8786 ( .I(n8760), .ZN(n6789) );
  CLKNAND2HSV2 U8787 ( .A1(n10597), .A2(n10596), .ZN(n6791) );
  AOI21HSV4 U8788 ( .A1(n6793), .A2(n6792), .B(n8915), .ZN(n6795) );
  NOR2HSV4 U8789 ( .A1(n7322), .A2(n10594), .ZN(n6792) );
  CLKNAND2HSV0 U8790 ( .A1(n13749), .A2(\pe20/got [2]), .ZN(n8365) );
  CLKNAND2HSV3 U8791 ( .A1(n6796), .A2(\pe16/phq [2]), .ZN(n7292) );
  CLKNAND2HSV3 U8792 ( .A1(\pe16/got [7]), .A2(\pe16/ti_1 ), .ZN(n6796) );
  CLKNHSV3 U8793 ( .I(\pe16/phq [2]), .ZN(n6798) );
  CLKNAND2HSV3 U8794 ( .A1(n6797), .A2(n7980), .ZN(n7981) );
  NAND3HSV4 U8795 ( .A1(n6798), .A2(\pe16/ti_1 ), .A3(\pe16/got [7]), .ZN(
        n7293) );
  CLKNAND2HSV4 U8796 ( .A1(n9391), .A2(n9392), .ZN(n11237) );
  XNOR2HSV4 U8797 ( .A1(n6806), .A2(n6799), .ZN(n8422) );
  OAI21HSV4 U8798 ( .A1(n6802), .A2(n6801), .B(n6800), .ZN(n6799) );
  CLKNAND2HSV2 U8799 ( .A1(n6801), .A2(n6802), .ZN(n6800) );
  CLKNAND2HSV2 U8800 ( .A1(n14935), .A2(\pe2/got [3]), .ZN(n6801) );
  AOI21HSV4 U8801 ( .A1(n6805), .A2(n6804), .B(n6803), .ZN(n6802) );
  CLKNHSV2 U8802 ( .I(n8421), .ZN(n6803) );
  CLKNHSV2 U8803 ( .I(n13761), .ZN(n6804) );
  NOR2HSV4 U8804 ( .A1(n8420), .A2(n13100), .ZN(n6805) );
  CLKNAND2HSV2 U8805 ( .A1(n13759), .A2(n6721), .ZN(n6806) );
  NOR2HSV4 U8806 ( .A1(n14582), .A2(n9794), .ZN(n7792) );
  XNOR2HSV4 U8807 ( .A1(n6809), .A2(n6807), .ZN(n14582) );
  AOI21HSV4 U8808 ( .A1(n11612), .A2(n9434), .B(n6808), .ZN(n6807) );
  NOR2HSV4 U8809 ( .A1(n11674), .A2(n6811), .ZN(n6808) );
  XNOR2HSV4 U8810 ( .A1(n6815), .A2(n6813), .ZN(n6809) );
  CLKNAND2HSV2 U8811 ( .A1(n9789), .A2(n6812), .ZN(n6811) );
  CLKNHSV2 U8812 ( .I(n8922), .ZN(n6812) );
  XNOR2HSV4 U8813 ( .A1(n6814), .A2(n9787), .ZN(n6813) );
  CLKNHSV2 U8814 ( .I(n9788), .ZN(n6814) );
  INHSV6 U8815 ( .I(n6816), .ZN(n15167) );
  CLKNHSV3 U8816 ( .I(n6819), .ZN(n6817) );
  INHSV2 U8817 ( .I(n10440), .ZN(n6818) );
  CLKNHSV2 U8818 ( .I(n8928), .ZN(n6819) );
  NAND2HSV4 U8819 ( .A1(n10591), .A2(n10590), .ZN(n8952) );
  CLKNAND2HSV4 U8820 ( .A1(n15201), .A2(n10599), .ZN(n10591) );
  XNOR2HSV2 U8821 ( .A1(n14115), .A2(n6821), .ZN(n6820) );
  CLKNAND2HSV3 U8822 ( .A1(\pe10/ti_7[6] ), .A2(\pe10/got [2]), .ZN(n6821) );
  CLKNAND2HSV3 U8823 ( .A1(n6825), .A2(n6823), .ZN(n6829) );
  CLKNAND2HSV2 U8824 ( .A1(n6824), .A2(n7082), .ZN(n6823) );
  CLKNAND2HSV2 U8825 ( .A1(n7080), .A2(\pe15/pvq [1]), .ZN(n6825) );
  OAI21HSV4 U8826 ( .A1(\pe15/phq [1]), .A2(n6827), .B(n6826), .ZN(n6828) );
  CLKNAND2HSV2 U8827 ( .A1(\pe15/bq[8] ), .A2(\pe15/aot [8]), .ZN(n6827) );
  XNOR2HSV4 U8828 ( .A1(n6829), .A2(n6828), .ZN(n15235) );
  CLKBUFHSV2 U8829 ( .I(n14943), .Z(n6830) );
  CLKNAND2HSV3 U8830 ( .A1(n14943), .A2(\pe12/got [6]), .ZN(n6831) );
  CLKNAND2HSV4 U8831 ( .A1(n11445), .A2(n11415), .ZN(n14943) );
  CLKNAND2HSV3 U8832 ( .A1(n15250), .A2(n11448), .ZN(n11445) );
  XNOR2HSV4 U8833 ( .A1(n6833), .A2(n6832), .ZN(n10464) );
  CLKNAND2HSV2 U8834 ( .A1(\pe7/aot [7]), .A2(\pe7/bq[7] ), .ZN(n6833) );
  OAI21HSV4 U8835 ( .A1(n6726), .A2(n9284), .B(n6834), .ZN(n7813) );
  AOI21HSV4 U8836 ( .A1(n7755), .A2(n7814), .B(n7815), .ZN(n6834) );
  XNOR2HSV4 U8837 ( .A1(n7757), .A2(n9248), .ZN(n9284) );
  NOR2HSV4 U8838 ( .A1(n9246), .A2(n9247), .ZN(n7814) );
  XNOR2HSV4 U8839 ( .A1(n6871), .A2(n6873), .ZN(n9193) );
  CLKNAND2HSV4 U8840 ( .A1(n6839), .A2(n6836), .ZN(n14179) );
  CLKNAND2HSV1 U8841 ( .A1(n6838), .A2(n6837), .ZN(n6836) );
  OAI21HSV2 U8842 ( .A1(n12369), .A2(n7228), .B(n7225), .ZN(n6837) );
  CLKNHSV3 U8843 ( .I(n13898), .ZN(n6838) );
  CLKNAND2HSV3 U8844 ( .A1(n7440), .A2(n7439), .ZN(n6841) );
  AOI31HSV2 U8845 ( .A1(n6847), .A2(n11412), .A3(n6998), .B(n6843), .ZN(n6842)
         );
  OAI31HSV2 U8846 ( .A1(n11410), .A2(n6732), .A3(n6845), .B(n6844), .ZN(n6843)
         );
  CLKNHSV2 U8847 ( .I(n6996), .ZN(n6844) );
  CLKNAND2HSV2 U8848 ( .A1(n6846), .A2(n6998), .ZN(n6845) );
  CLKNHSV2 U8849 ( .I(n11409), .ZN(n6846) );
  CLKNAND2HSV2 U8850 ( .A1(n7127), .A2(n12337), .ZN(n6847) );
  CLKNHSV2 U8851 ( .I(n11406), .ZN(n6848) );
  AOI21HSV4 U8852 ( .A1(n9559), .A2(n8034), .B(n9563), .ZN(n6849) );
  XNOR2HSV4 U8853 ( .A1(n6854), .A2(n6852), .ZN(n11940) );
  XNOR2HSV4 U8854 ( .A1(n11939), .A2(n6853), .ZN(n6852) );
  XOR3HSV2 U8855 ( .A1(n11937), .A2(n11936), .A3(n11938), .Z(n6853) );
  AOI31HSV2 U8856 ( .A1(n11741), .A2(n11740), .A3(n7793), .B(n11895), .ZN(
        n6855) );
  CLKNAND2HSV2 U8857 ( .A1(n11738), .A2(n11765), .ZN(n6856) );
  MUX2NHSV2 U8858 ( .I0(n13636), .I1(n13635), .S(n6858), .ZN(n6857) );
  XNOR2HSV4 U8859 ( .A1(n6859), .A2(n13619), .ZN(n6858) );
  CLKNAND2HSV2 U8860 ( .A1(n14450), .A2(\pe7/got [4]), .ZN(n6859) );
  CLKNHSV2 U8861 ( .I(n13637), .ZN(n6860) );
  XNOR2HSV4 U8862 ( .A1(n9953), .A2(n9954), .ZN(n9982) );
  OAI21HSV4 U8863 ( .A1(n15244), .A2(n9988), .B(n9909), .ZN(n9954) );
  XNOR2HSV4 U8864 ( .A1(n9907), .A2(n9906), .ZN(n15244) );
  XNOR2HSV4 U8865 ( .A1(n6862), .A2(n6861), .ZN(n9953) );
  CLKNAND2HSV2 U8866 ( .A1(n9882), .A2(\pe13/got [6]), .ZN(n6861) );
  XNOR2HSV4 U8867 ( .A1(n9919), .A2(n9918), .ZN(n6862) );
  CLKNHSV2 U8868 ( .I(n6865), .ZN(n6864) );
  CLKNAND2HSV2 U8869 ( .A1(n13532), .A2(\pe8/got [4]), .ZN(n6865) );
  CLKNAND2HSV2 U8870 ( .A1(n13533), .A2(n6867), .ZN(n6866) );
  CLKNHSV2 U8871 ( .I(n6868), .ZN(n6867) );
  NAND3HSV4 U8872 ( .A1(n12770), .A2(n12769), .A3(n11591), .ZN(n13533) );
  XNOR2HSV4 U8873 ( .A1(n11607), .A2(n11608), .ZN(n12770) );
  CLKNAND2HSV4 U8874 ( .A1(n7776), .A2(n11601), .ZN(n12769) );
  INHSV2 U8875 ( .I(n11605), .ZN(n6868) );
  AOI21HSV2 U8876 ( .A1(n7199), .A2(\pe18/got [8]), .B(n9133), .ZN(n6869) );
  AOI21HSV4 U8877 ( .A1(n9152), .A2(n6870), .B(n9151), .ZN(n9170) );
  CLKNHSV2 U8878 ( .I(n9150), .ZN(n6870) );
  XNOR2HSV4 U8879 ( .A1(n9193), .A2(n11996), .ZN(n9154) );
  XNOR2HSV4 U8880 ( .A1(n6872), .A2(n6887), .ZN(n6871) );
  XNOR2HSV4 U8881 ( .A1(n6892), .A2(n6891), .ZN(n6872) );
  NOR2HSV4 U8882 ( .A1(n9165), .A2(n9140), .ZN(n6873) );
  NOR2HSV4 U8883 ( .A1(n7199), .A2(n7198), .ZN(n9165) );
  CLKNAND2HSV3 U8884 ( .A1(n6874), .A2(\pe6/got [2]), .ZN(n12989) );
  XNOR2HSV4 U8885 ( .A1(n6878), .A2(n6875), .ZN(n15261) );
  XNOR2HSV4 U8886 ( .A1(n6877), .A2(n6876), .ZN(n6875) );
  CLKNAND2HSV2 U8887 ( .A1(n7827), .A2(n7826), .ZN(n6876) );
  XNOR2HSV4 U8888 ( .A1(n7825), .A2(n8334), .ZN(n6877) );
  OAI21HSV4 U8889 ( .A1(n6886), .A2(n6885), .B(n6879), .ZN(n6878) );
  CLKNAND2HSV2 U8890 ( .A1(n6884), .A2(n6880), .ZN(n6879) );
  NAND3HSV4 U8891 ( .A1(n10115), .A2(n10114), .A3(n6881), .ZN(n6880) );
  CLKNAND2HSV2 U8892 ( .A1(n6883), .A2(n6882), .ZN(n6881) );
  CLKNHSV2 U8893 ( .I(n10116), .ZN(n6882) );
  CLKNHSV2 U8894 ( .I(n10117), .ZN(n6883) );
  CLKNHSV2 U8895 ( .I(n7829), .ZN(n6886) );
  XOR2HSV2 U8896 ( .A1(n6889), .A2(n6888), .Z(n6887) );
  CLKNAND2HSV2 U8897 ( .A1(\pe18/aot [6]), .A2(\pe18/bq[8] ), .ZN(n6888) );
  NOR2HSV4 U8898 ( .A1(n10802), .A2(n6890), .ZN(n6889) );
  CLKNHSV2 U8899 ( .I(\pe18/pvq [3]), .ZN(n6890) );
  CLKNAND2HSV2 U8900 ( .A1(\pe18/bq[7] ), .A2(\pe18/aot [7]), .ZN(n6894) );
  CLKNAND2HSV2 U8901 ( .A1(n12272), .A2(\pe10/aot [6]), .ZN(n10057) );
  CLKNAND2HSV2 U8902 ( .A1(n7848), .A2(n7331), .ZN(n15229) );
  CLKNHSV2 U8903 ( .I(n11159), .ZN(n6895) );
  CLKNAND2HSV2 U8904 ( .A1(n15229), .A2(n11207), .ZN(n7330) );
  MUX2NHSV2 U8905 ( .I0(n13014), .I1(n13013), .S(n13012), .ZN(n15205) );
  XNOR2HSV4 U8906 ( .A1(n6897), .A2(n6896), .ZN(n6900) );
  XOR2HSV2 U8907 ( .A1(n9633), .A2(\pe4/phq [4]), .Z(n6896) );
  XOR2HSV2 U8908 ( .A1(n9634), .A2(n8281), .Z(n6897) );
  XNOR2HSV4 U8909 ( .A1(n6898), .A2(n6909), .ZN(n6905) );
  XOR2HSV2 U8910 ( .A1(n6900), .A2(n6899), .Z(n6898) );
  XOR2HSV2 U8911 ( .A1(n6901), .A2(n9632), .Z(n6899) );
  CLKNAND2HSV2 U8912 ( .A1(n6906), .A2(n8280), .ZN(n6901) );
  CLKNAND2HSV3 U8913 ( .A1(n14733), .A2(\pe4/got [7]), .ZN(n6902) );
  CLKNAND2HSV1 U8914 ( .A1(n6908), .A2(n6907), .ZN(n6906) );
  CLKNHSV1 U8915 ( .I(n8279), .ZN(n6907) );
  CLKNHSV1 U8916 ( .I(n8278), .ZN(n6908) );
  NOR2HSV3 U8917 ( .A1(n9635), .A2(n6910), .ZN(n6909) );
  INHSV2 U8918 ( .I(n9637), .ZN(n6910) );
  CLKNAND2HSV4 U8919 ( .A1(n15248), .A2(n7495), .ZN(n11610) );
  CLKNAND2HSV4 U8920 ( .A1(n6912), .A2(n6911), .ZN(n7494) );
  CLKNAND2HSV4 U8921 ( .A1(n6717), .A2(n7508), .ZN(n7493) );
  INHSV2 U8922 ( .I(n8430), .ZN(n6911) );
  CLKNAND2HSV3 U8923 ( .A1(n7508), .A2(n7507), .ZN(n6912) );
  CLKNAND2HSV4 U8924 ( .A1(n14179), .A2(\pe6/got [2]), .ZN(n6915) );
  XNOR2HSV4 U8925 ( .A1(n7959), .A2(n6917), .ZN(n6916) );
  CLKNAND2HSV2 U8926 ( .A1(n15084), .A2(\pe19/got [6]), .ZN(n6917) );
  CLKNAND2HSV2 U8927 ( .A1(n13315), .A2(n13844), .ZN(n6919) );
  CLKNAND2HSV2 U8928 ( .A1(n6954), .A2(n13260), .ZN(n12385) );
  NOR2HSV4 U8929 ( .A1(n6955), .A2(n12171), .ZN(n12386) );
  CLKNAND2HSV2 U8930 ( .A1(n8174), .A2(n8175), .ZN(n8176) );
  XNOR2HSV4 U8931 ( .A1(n8173), .A2(n6920), .ZN(n8174) );
  XNOR2HSV4 U8932 ( .A1(n13602), .A2(n6921), .ZN(n6920) );
  XNOR2HSV4 U8933 ( .A1(n8172), .A2(n13599), .ZN(n6921) );
  INHSV2 U8934 ( .I(n12791), .ZN(n6922) );
  NOR2HSV4 U8935 ( .A1(n11494), .A2(n13429), .ZN(n12779) );
  INHSV2 U8936 ( .I(n6923), .ZN(n7242) );
  CLKBUFHSV2 U8937 ( .I(n12791), .Z(n6924) );
  CLKNHSV2 U8938 ( .I(n7075), .ZN(n12819) );
  INHSV2 U8939 ( .I(n12791), .ZN(n12780) );
  CLKNAND2HSV2 U8940 ( .A1(n12780), .A2(n12779), .ZN(n12775) );
  INAND2HSV4 U8941 ( .A1(n7075), .B1(n6924), .ZN(n12787) );
  CLKNAND2HSV3 U8942 ( .A1(n6927), .A2(n10926), .ZN(\pe10/ti_7[5] ) );
  XNOR2HSV4 U8943 ( .A1(n6930), .A2(n6928), .ZN(n15262) );
  CLKNAND2HSV3 U8944 ( .A1(n10107), .A2(n10116), .ZN(n10121) );
  XNOR2HSV4 U8945 ( .A1(n6929), .A2(n10111), .ZN(n6928) );
  CLKNAND2HSV2 U8946 ( .A1(n10075), .A2(n10074), .ZN(n6929) );
  NAND3HSV4 U8947 ( .A1(n10122), .A2(n10121), .A3(n10072), .ZN(n6930) );
  CLKNHSV2 U8948 ( .I(n8967), .ZN(n6931) );
  CLKNHSV2 U8949 ( .I(n8744), .ZN(n6935) );
  CLKNHSV2 U8950 ( .I(\pe15/got [6]), .ZN(n6936) );
  XNOR2HSV4 U8951 ( .A1(n6938), .A2(n12332), .ZN(n6937) );
  XNOR2HSV4 U8952 ( .A1(n12333), .A2(n12334), .ZN(n6938) );
  INHSV2 U8953 ( .I(n6940), .ZN(n6939) );
  CLKNAND2HSV1 U8954 ( .A1(n9763), .A2(n9449), .ZN(n6941) );
  AOI21HSV2 U8955 ( .A1(n8507), .A2(n8508), .B(n7389), .ZN(n6943) );
  CLKNHSV2 U8956 ( .I(n9741), .ZN(n6944) );
  XNOR2HSV4 U8957 ( .A1(n6945), .A2(n9447), .ZN(n9741) );
  XNOR2HSV4 U8958 ( .A1(n6946), .A2(n7014), .ZN(n6945) );
  XNOR2HSV4 U8959 ( .A1(n7018), .A2(n7016), .ZN(n6946) );
  XNOR2HSV4 U8960 ( .A1(n10968), .A2(n10967), .ZN(n11709) );
  XNOR2HSV4 U8961 ( .A1(n10963), .A2(n6947), .ZN(n10967) );
  XOR3HSV2 U8962 ( .A1(n10962), .A2(n6949), .A3(n6948), .Z(n6947) );
  XNOR2HSV4 U8963 ( .A1(n6950), .A2(n10959), .ZN(n6949) );
  XNOR2HSV4 U8964 ( .A1(n10960), .A2(n6951), .ZN(n6950) );
  CLKNHSV2 U8965 ( .I(n10961), .ZN(n6951) );
  OAI21HSV4 U8966 ( .A1(n10945), .A2(n10944), .B(n7868), .ZN(n10968) );
  CLKNHSV2 U8967 ( .I(n7379), .ZN(n6952) );
  XNOR2HSV4 U8968 ( .A1(n7382), .A2(n10323), .ZN(n10331) );
  NOR2HSV4 U8969 ( .A1(n13260), .A2(n6956), .ZN(n6955) );
  CLKNAND2HSV2 U8970 ( .A1(n15073), .A2(n12137), .ZN(n6956) );
  CLKNAND2HSV4 U8971 ( .A1(n15260), .A2(n12353), .ZN(n11921) );
  XNOR2HSV4 U8972 ( .A1(n9601), .A2(n9600), .ZN(n6958) );
  CLKNAND2HSV3 U8973 ( .A1(n11921), .A2(n11916), .ZN(\pe11/ti_7[1] ) );
  XOR3HSV2 U8974 ( .A1(n6963), .A2(n6961), .A3(n6959), .Z(n10082) );
  XNOR2HSV4 U8975 ( .A1(n6960), .A2(\pe10/phq [5]), .ZN(n6959) );
  CLKNAND2HSV2 U8976 ( .A1(\pe10/aot [4]), .A2(\pe10/bq[8] ), .ZN(n6960) );
  NOR2HSV4 U8977 ( .A1(n10035), .A2(n6962), .ZN(n6961) );
  CLKNHSV2 U8978 ( .I(\pe10/pvq [5]), .ZN(n6962) );
  CLKNAND2HSV4 U8979 ( .A1(n6967), .A2(n6966), .ZN(n7641) );
  CLKNHSV2 U8980 ( .I(n11210), .ZN(n6966) );
  NOR2HSV3 U8981 ( .A1(n6968), .A2(n7644), .ZN(n6967) );
  CLKNHSV4 U8982 ( .I(n11209), .ZN(n6968) );
  CLKNAND2HSV4 U8983 ( .A1(n11204), .A2(n11205), .ZN(n7644) );
  INHSV2 U8984 ( .I(n10679), .ZN(n6969) );
  XOR3HSV2 U8985 ( .A1(n14362), .A2(n6971), .A3(n6970), .Z(\pe16/poht [3]) );
  NOR2HSV4 U8986 ( .A1(n14364), .A2(n14363), .ZN(n6970) );
  XNOR2HSV4 U8987 ( .A1(n6973), .A2(n6972), .ZN(n6971) );
  XOR2HSV2 U8988 ( .A1(n14361), .A2(n14360), .Z(n6972) );
  CLKNAND2HSV2 U8989 ( .A1(n14348), .A2(\pe16/got [4]), .ZN(n6973) );
  XOR2HSV2 U8990 ( .A1(n10420), .A2(n6975), .Z(n6974) );
  XNOR2HSV4 U8991 ( .A1(n6978), .A2(n6977), .ZN(n6976) );
  CLKNAND2HSV2 U8992 ( .A1(\pe17/aot [8]), .A2(\pe17/bq[6] ), .ZN(n6979) );
  NOR2HSV4 U8993 ( .A1(n13583), .A2(n6980), .ZN(n12629) );
  CLKNHSV2 U8994 ( .I(n7473), .ZN(n6981) );
  NOR2HSV4 U8995 ( .A1(n6982), .A2(n6983), .ZN(n13583) );
  CLKNAND2HSV1 U8996 ( .A1(n15257), .A2(n11765), .ZN(n7673) );
  OAI21HSV4 U8997 ( .A1(n15257), .A2(n11895), .B(n8504), .ZN(n7678) );
  CLKNAND2HSV4 U8998 ( .A1(n11743), .A2(n11742), .ZN(n15257) );
  NOR2HSV4 U8999 ( .A1(n6286), .A2(n6984), .ZN(n7448) );
  CLKNHSV2 U9000 ( .I(n6986), .ZN(n6984) );
  CLKNHSV2 U9001 ( .I(n10063), .ZN(n6985) );
  CLKNHSV2 U9002 ( .I(n10063), .ZN(n10068) );
  CLKNHSV2 U9003 ( .I(n7449), .ZN(n6986) );
  CLKNHSV2 U9004 ( .I(n6988), .ZN(n6987) );
  CLKNAND2HSV2 U9005 ( .A1(n10064), .A2(n10148), .ZN(n6988) );
  XOR2HSV4 U9006 ( .A1(n10399), .A2(n10398), .Z(n6993) );
  AOI21HSV4 U9007 ( .A1(n6991), .A2(n6990), .B(n10403), .ZN(n6994) );
  CLKNHSV2 U9008 ( .I(n10389), .ZN(n6990) );
  CLKNHSV2 U9009 ( .I(n10380), .ZN(n6991) );
  XNOR2HSV4 U9010 ( .A1(n6993), .A2(n6992), .ZN(n7054) );
  CLKNAND2HSV3 U9011 ( .A1(n10387), .A2(n6994), .ZN(n10394) );
  CLKNHSV4 U9012 ( .I(n10392), .ZN(n10387) );
  AOI21HSV4 U9013 ( .A1(n10391), .A2(n10392), .B(n10390), .ZN(n10393) );
  NAND3HSV4 U9014 ( .A1(n11404), .A2(n6998), .A3(n11403), .ZN(n6995) );
  NOR2HSV4 U9015 ( .A1(n6997), .A2(n7680), .ZN(n6996) );
  CLKNHSV2 U9016 ( .I(n6999), .ZN(n6997) );
  CLKNHSV2 U9017 ( .I(n7680), .ZN(n6998) );
  CLKNHSV2 U9018 ( .I(n12337), .ZN(n6999) );
  XOR2HSV2 U9019 ( .A1(n11033), .A2(n7000), .Z(n11034) );
  XNOR2HSV4 U9020 ( .A1(n7002), .A2(n7001), .ZN(n7000) );
  CLKNHSV2 U9021 ( .I(n11032), .ZN(n7001) );
  CLKNAND2HSV2 U9022 ( .A1(n11015), .A2(n7004), .ZN(n7003) );
  CLKNHSV2 U9023 ( .I(n7005), .ZN(n7004) );
  XNOR2HSV1 U9024 ( .A1(n7007), .A2(n7006), .ZN(\pe6/poht [7]) );
  CLKNHSV2 U9025 ( .I(n14180), .ZN(n7006) );
  CLKNAND2HSV2 U9026 ( .A1(n13139), .A2(n7008), .ZN(n13341) );
  CLKNHSV2 U9027 ( .I(n7013), .ZN(n7008) );
  NAND3HSV4 U9028 ( .A1(n13139), .A2(n11977), .A3(n7011), .ZN(n7010) );
  NOR2HSV4 U9029 ( .A1(n7013), .A2(n7012), .ZN(n7011) );
  CLKNAND2HSV4 U9030 ( .A1(n13142), .A2(n11977), .ZN(n13138) );
  CLKNHSV2 U9031 ( .I(n13142), .ZN(n7012) );
  CLKNHSV2 U9032 ( .I(n11976), .ZN(n7013) );
  XNOR2HSV4 U9033 ( .A1(n9446), .A2(n7017), .ZN(n7016) );
  XNOR2HSV4 U9034 ( .A1(n9443), .A2(n9767), .ZN(n7017) );
  XNOR2HSV4 U9035 ( .A1(n7019), .A2(n9442), .ZN(n7018) );
  CLKNAND2HSV2 U9036 ( .A1(n9439), .A2(n7020), .ZN(n7019) );
  CLKNAND2HSV2 U9037 ( .A1(n7022), .A2(n13920), .ZN(n7020) );
  CLKNHSV2 U9038 ( .I(n9441), .ZN(n7021) );
  CLKNHSV2 U9039 ( .I(n9440), .ZN(n7022) );
  CLKNAND2HSV2 U9040 ( .A1(\pe10/aot [5]), .A2(\pe10/bq[8] ), .ZN(n10037) );
  NOR2HSV4 U9041 ( .A1(n7024), .A2(n7023), .ZN(n10049) );
  NAND3HSV4 U9042 ( .A1(n7027), .A2(n7026), .A3(n10040), .ZN(n7023) );
  NAND3HSV4 U9043 ( .A1(n7238), .A2(n7236), .A3(n7237), .ZN(n7026) );
  CLKNAND2HSV3 U9044 ( .A1(n7234), .A2(n7235), .ZN(n7027) );
  XNOR2HSV4 U9045 ( .A1(n7028), .A2(n8069), .ZN(n13785) );
  CLKNAND2HSV2 U9046 ( .A1(n13762), .A2(\pe2/got [3]), .ZN(n7028) );
  CLKNHSV2 U9047 ( .I(n10589), .ZN(n8614) );
  CLKNAND2HSV2 U9048 ( .A1(n10580), .A2(n10581), .ZN(n7029) );
  AOI21HSV1 U9049 ( .A1(n8615), .A2(n8614), .B(n7031), .ZN(n8616) );
  CLKNAND2HSV2 U9050 ( .A1(n7033), .A2(n7032), .ZN(n7031) );
  CLKNHSV0 U9051 ( .I(\pe4/got [8]), .ZN(n7032) );
  CLKNHSV2 U9052 ( .I(n9714), .ZN(n7033) );
  XOR2HSV2 U9053 ( .A1(n7034), .A2(n12493), .Z(n12494) );
  XOR2HSV2 U9054 ( .A1(n12492), .A2(n7035), .Z(n7034) );
  XNOR2HSV4 U9055 ( .A1(n12484), .A2(n7036), .ZN(n7035) );
  XNOR2HSV4 U9056 ( .A1(n12491), .A2(n12483), .ZN(n7036) );
  CLKNAND2HSV2 U9057 ( .A1(n15287), .A2(n10789), .ZN(n7037) );
  XNOR2HSV4 U9058 ( .A1(n7718), .A2(n7038), .ZN(n15287) );
  CLKNHSV4 U9059 ( .I(n7631), .ZN(n13237) );
  NAND3HSV4 U9060 ( .A1(n12047), .A2(n12046), .A3(n12045), .ZN(n7631) );
  CLKNAND2HSV2 U9061 ( .A1(n7039), .A2(\pe17/got [1]), .ZN(n13265) );
  XNOR3HSV2 U9062 ( .A1(n8341), .A2(n7316), .A3(n7040), .ZN(n8342) );
  NOR2HSV4 U9063 ( .A1(n14442), .A2(n8338), .ZN(n7040) );
  CLKNHSV2 U9064 ( .I(n10458), .ZN(n7041) );
  XNOR2HSV4 U9065 ( .A1(n8897), .A2(n7041), .ZN(n15272) );
  CLKNAND2HSV2 U9066 ( .A1(n11001), .A2(n7042), .ZN(n7716) );
  CLKNAND2HSV2 U9067 ( .A1(n7806), .A2(n10404), .ZN(n10993) );
  XNOR2HSV4 U9068 ( .A1(n7808), .A2(n7807), .ZN(n11002) );
  CLKNHSV2 U9069 ( .I(n8328), .ZN(n7612) );
  XNOR2HSV4 U9070 ( .A1(n7044), .A2(n7043), .ZN(n8328) );
  CLKNAND2HSV2 U9071 ( .A1(n15077), .A2(\pe6/got [5]), .ZN(n7043) );
  XNOR2HSV4 U9072 ( .A1(n7045), .A2(n13058), .ZN(n7044) );
  XNOR2HSV4 U9073 ( .A1(n13056), .A2(n7046), .ZN(n7045) );
  CLKNHSV2 U9074 ( .I(n13055), .ZN(n7046) );
  NAND3HSV4 U9075 ( .A1(n7054), .A2(n10393), .A3(n10394), .ZN(n7052) );
  OAI21HSV4 U9076 ( .A1(n7049), .A2(n10402), .B(n7048), .ZN(n7047) );
  CLKNHSV2 U9077 ( .I(n7733), .ZN(n7048) );
  CLKNHSV2 U9078 ( .I(n10808), .ZN(n7049) );
  AOI21HSV4 U9079 ( .A1(n12631), .A2(\pe4/got [5]), .B(n8350), .ZN(n8351) );
  CLKNAND2HSV2 U9080 ( .A1(n8349), .A2(n7055), .ZN(n8350) );
  CLKNAND2HSV2 U9081 ( .A1(n7057), .A2(n7056), .ZN(n7055) );
  NOR2HSV4 U9082 ( .A1(n12645), .A2(n10536), .ZN(n7056) );
  CLKNHSV2 U9083 ( .I(n8348), .ZN(n7057) );
  XNOR2HSV4 U9084 ( .A1(n7058), .A2(n10539), .ZN(n8348) );
  XNOR2HSV4 U9085 ( .A1(n10558), .A2(n7059), .ZN(n7058) );
  CLKNHSV2 U9086 ( .I(n10538), .ZN(n7059) );
  CLKNAND2HSV4 U9087 ( .A1(n10360), .A2(n10359), .ZN(n10358) );
  CLKNHSV8 U9088 ( .I(\pe21/phq [2]), .ZN(n10359) );
  NAND3HSV4 U9089 ( .A1(n7060), .A2(n10599), .A3(n10116), .ZN(n10115) );
  AOI21HSV4 U9090 ( .A1(n7060), .A2(n10113), .B(n10120), .ZN(n10114) );
  CLKNAND2HSV2 U9091 ( .A1(n7912), .A2(n7060), .ZN(n7828) );
  OAI21HSV1 U9092 ( .A1(n7912), .A2(n7060), .B(n10122), .ZN(n7913) );
  CLKNHSV4 U9093 ( .I(n10111), .ZN(n7060) );
  CLKNHSV4 U9094 ( .I(\pe21/bq[8] ), .ZN(n10361) );
  NAND2HSV4 U9095 ( .A1(n7064), .A2(n7061), .ZN(\pe5/ti_7[7] ) );
  CLKNAND2HSV3 U9096 ( .A1(n7063), .A2(n7062), .ZN(n7061) );
  NOR2HSV4 U9097 ( .A1(n13019), .A2(n13018), .ZN(n7062) );
  CLKNAND2HSV3 U9098 ( .A1(n15205), .A2(n11472), .ZN(n7063) );
  AOI31HSV2 U9099 ( .A1(n13019), .A2(n13017), .A3(n7065), .B(n13016), .ZN(
        n7064) );
  XNOR2HSV4 U9100 ( .A1(n12826), .A2(n12825), .ZN(n13019) );
  CLKNHSV3 U9101 ( .I(n9457), .ZN(n7066) );
  CLKNAND2HSV4 U9102 ( .A1(n14821), .A2(n13645), .ZN(n9457) );
  CLKNAND2HSV3 U9103 ( .A1(n10593), .A2(n7067), .ZN(n10595) );
  CLKNHSV2 U9104 ( .I(n10592), .ZN(n7067) );
  XNOR2HSV4 U9105 ( .A1(n7068), .A2(n7294), .ZN(n9456) );
  XNOR2HSV4 U9106 ( .A1(n7295), .A2(n9072), .ZN(n7068) );
  XNOR2HSV2 U9107 ( .A1(n7073), .A2(n7070), .ZN(n7069) );
  OAI21HSV1 U9108 ( .A1(n9860), .A2(n9861), .B(n7071), .ZN(n7070) );
  CLKNAND2HSV3 U9109 ( .A1(n9860), .A2(n7072), .ZN(n7071) );
  NOR2HSV3 U9110 ( .A1(n8227), .A2(n12998), .ZN(n7072) );
  CLKNAND2HSV4 U9111 ( .A1(\pe6/ti_7[5] ), .A2(\pe6/got [3]), .ZN(n7073) );
  CLKNAND2HSV4 U9112 ( .A1(n12369), .A2(n9536), .ZN(n9847) );
  CLKNAND2HSV3 U9113 ( .A1(n11495), .A2(n10307), .ZN(n7075) );
  CLKNAND2HSV4 U9114 ( .A1(n7078), .A2(n7076), .ZN(n11495) );
  CLKNAND2HSV2 U9115 ( .A1(n10353), .A2(n7077), .ZN(n7076) );
  CLKNAND2HSV0 U9116 ( .A1(n12811), .A2(\pe5/got [7]), .ZN(n7077) );
  NAND2HSV2 U9117 ( .A1(n10352), .A2(n10351), .ZN(n7078) );
  INHSV4 U9118 ( .I(n10423), .ZN(n7079) );
  NOR2HSV3 U9119 ( .A1(n7082), .A2(n7081), .ZN(n7080) );
  CLKNHSV4 U9120 ( .I(\pe15/ctrq ), .ZN(n7081) );
  CLKNAND2HSV4 U9121 ( .A1(\pe15/got [8]), .A2(\pe15/ti_1 ), .ZN(n7082) );
  INHSV2 U9122 ( .I(n7375), .ZN(n7083) );
  XNOR2HSV4 U9123 ( .A1(n7086), .A2(n7084), .ZN(n7679) );
  XOR2HSV2 U9124 ( .A1(n7085), .A2(\pe5/phq [3]), .Z(n7084) );
  XNOR2HSV4 U9125 ( .A1(n7088), .A2(n7087), .ZN(n7086) );
  CLKNAND2HSV2 U9126 ( .A1(\pe5/bq[6] ), .A2(\pe5/aot [8]), .ZN(n7087) );
  AOI21HSV4 U9127 ( .A1(n7093), .A2(n7089), .B(n7095), .ZN(n7094) );
  CLKNHSV2 U9128 ( .I(n7090), .ZN(n7089) );
  CLKNAND2HSV2 U9129 ( .A1(n14962), .A2(n7091), .ZN(n7090) );
  NOR2HSV4 U9130 ( .A1(n7096), .A2(n7092), .ZN(n7091) );
  CLKNHSV2 U9131 ( .I(n12103), .ZN(n7092) );
  CLKNHSV2 U9132 ( .I(n10714), .ZN(n7093) );
  OAI21HSV4 U9133 ( .A1(n7097), .A2(n7096), .B(n7094), .ZN(\pe17/ti_7[3] ) );
  CLKNHSV2 U9134 ( .I(n12022), .ZN(n7095) );
  CLKNHSV2 U9135 ( .I(n12043), .ZN(n7096) );
  CLKNAND2HSV4 U9136 ( .A1(n7099), .A2(n7098), .ZN(n14821) );
  CLKNAND2HSV2 U9137 ( .A1(n9056), .A2(n9055), .ZN(n7098) );
  CLKNAND2HSV3 U9138 ( .A1(n9054), .A2(n9053), .ZN(n7099) );
  CLKNAND2HSV4 U9139 ( .A1(n9170), .A2(n9171), .ZN(n7334) );
  CLKNHSV2 U9140 ( .I(n13766), .ZN(n14805) );
  CLKNHSV2 U9141 ( .I(\pe2/phq [3]), .ZN(n7100) );
  CLKNAND2HSV2 U9142 ( .A1(\pe2/aot [7]), .A2(\pe2/bq[7] ), .ZN(n12881) );
  CLKNAND2HSV4 U9143 ( .A1(\pe10/ti_1 ), .A2(\pe10/got [8]), .ZN(n7102) );
  NOR2HSV4 U9144 ( .A1(n10714), .A2(n12130), .ZN(n7104) );
  AOI31HSV2 U9145 ( .A1(n14399), .A2(n10714), .A3(n14007), .B(n7106), .ZN(
        n7105) );
  CLKNHSV2 U9146 ( .I(n10717), .ZN(n7106) );
  XNOR2HSV4 U9147 ( .A1(n7111), .A2(n7108), .ZN(n11494) );
  XNOR2HSV4 U9148 ( .A1(n7110), .A2(n7109), .ZN(n7108) );
  XOR2HSV2 U9149 ( .A1(n11491), .A2(n11490), .Z(n7109) );
  CLKNAND2HSV2 U9150 ( .A1(n14952), .A2(\pe5/got [5]), .ZN(n7110) );
  AOI21HSV4 U9151 ( .A1(n7112), .A2(n11449), .B(n7205), .ZN(n7507) );
  CLKNHSV2 U9152 ( .I(n11445), .ZN(n7112) );
  CLKNHSV4 U9153 ( .I(n14943), .ZN(n7113) );
  INHSV2 U9154 ( .I(n7391), .ZN(n7114) );
  CLKNAND2HSV3 U9155 ( .A1(n7204), .A2(n7128), .ZN(n7115) );
  AOI21HSV2 U9156 ( .A1(n7118), .A2(n11036), .B(n7117), .ZN(n7116) );
  CLKNHSV4 U9157 ( .I(\pe14/got [6]), .ZN(n7117) );
  CLKNHSV4 U9158 ( .I(n8948), .ZN(n7118) );
  INHSV2 U9159 ( .I(n11036), .ZN(n7119) );
  XNOR2HSV4 U9160 ( .A1(n7166), .A2(n7165), .ZN(n15237) );
  INHSV24 U9161 ( .I(n11172), .ZN(n7120) );
  INHSV24 U9162 ( .I(n11173), .ZN(n7121) );
  CLKNHSV2 U9163 ( .I(n11211), .ZN(n11174) );
  OA21HSV4 U9164 ( .A1(n11211), .A2(n7121), .B(n7120), .Z(n7515) );
  AOI21HSV4 U9165 ( .A1(\pe16/ti_7t [6]), .A2(n8956), .B(n7122), .ZN(n11215)
         );
  NOR2HSV4 U9166 ( .A1(n7125), .A2(n13871), .ZN(n7122) );
  XNOR2HSV4 U9167 ( .A1(n7124), .A2(n7123), .ZN(n13871) );
  NAND3HSV4 U9168 ( .A1(n15185), .A2(n11211), .A3(n11220), .ZN(n13869) );
  CLKNHSV2 U9169 ( .I(n15185), .ZN(n7126) );
  CLKNAND2HSV3 U9170 ( .A1(n10766), .A2(n10767), .ZN(n7158) );
  CLKNAND2HSV3 U9171 ( .A1(n7159), .A2(n7158), .ZN(n15250) );
  CLKNAND2HSV3 U9172 ( .A1(n7567), .A2(n7571), .ZN(n7128) );
  CLKNAND2HSV4 U9173 ( .A1(n7568), .A2(n7129), .ZN(n7567) );
  NOR2HSV4 U9174 ( .A1(n9989), .A2(n7138), .ZN(n7137) );
  XNOR2HSV4 U9175 ( .A1(n9986), .A2(n9985), .ZN(n9989) );
  MUX2NHSV4 U9176 ( .I0(n7132), .I1(n7130), .S(n9989), .ZN(n11969) );
  CLKNHSV3 U9177 ( .I(n7131), .ZN(n7130) );
  CLKNAND2HSV3 U9178 ( .A1(n15241), .A2(n9978), .ZN(n7131) );
  NOR2HSV4 U9179 ( .A1(n7137), .A2(n7134), .ZN(n11968) );
  NOR2HSV4 U9180 ( .A1(n7136), .A2(n7135), .ZN(n7134) );
  CLKNHSV2 U9181 ( .I(\pe13/ti_7t [7]), .ZN(n7135) );
  CLKNHSV2 U9182 ( .I(n9988), .ZN(n7136) );
  CLKNHSV2 U9183 ( .I(n9987), .ZN(n7138) );
  CLKNHSV2 U9184 ( .I(n7857), .ZN(n7139) );
  CLKNHSV3 U9185 ( .I(n10839), .ZN(n7140) );
  CLKNAND2HSV3 U9186 ( .A1(n10643), .A2(n10642), .ZN(n10858) );
  CLKNAND2HSV2 U9187 ( .A1(\pe12/ti_7[3] ), .A2(\pe12/got [5]), .ZN(n8078) );
  CLKNAND2HSV2 U9188 ( .A1(\pe12/ti_7[3] ), .A2(\pe12/got [1]), .ZN(n12672) );
  CLKNAND2HSV2 U9189 ( .A1(\pe12/ti_7[3] ), .A2(\pe12/got [4]), .ZN(n12703) );
  CLKNAND2HSV2 U9190 ( .A1(\pe12/ti_7[3] ), .A2(\pe12/got [2]), .ZN(n12740) );
  CLKNAND2HSV2 U9191 ( .A1(n7144), .A2(n7142), .ZN(n8088) );
  CLKNAND2HSV2 U9192 ( .A1(n15183), .A2(n7143), .ZN(n7142) );
  NOR2HSV4 U9193 ( .A1(n8087), .A2(n8086), .ZN(n7143) );
  CLKNAND2HSV2 U9194 ( .A1(n7145), .A2(n8087), .ZN(n7144) );
  CLKNAND2HSV2 U9195 ( .A1(n15183), .A2(n7146), .ZN(n7145) );
  CLKNHSV2 U9196 ( .I(n13617), .ZN(n7146) );
  CLKNAND2HSV2 U9197 ( .A1(n15271), .A2(n12252), .ZN(n7147) );
  CLKNHSV2 U9198 ( .I(n10941), .ZN(n11708) );
  CLKNHSV2 U9199 ( .I(n7148), .ZN(n10965) );
  INAND2HSV4 U9200 ( .A1(n10942), .B1(n10941), .ZN(n7148) );
  OAI21HSV4 U9201 ( .A1(n7149), .A2(n11002), .B(n7803), .ZN(n10941) );
  CLKNAND2HSV2 U9202 ( .A1(n10945), .A2(n10789), .ZN(n7149) );
  XNOR2HSV4 U9203 ( .A1(n7151), .A2(n12377), .ZN(n7150) );
  OAI21HSV4 U9204 ( .A1(n15076), .A2(n12374), .B(n12373), .ZN(n7152) );
  XNOR2HSV4 U9205 ( .A1(n7153), .A2(n7392), .ZN(n11444) );
  OAI21HSV4 U9206 ( .A1(n15251), .A2(n14831), .B(n10769), .ZN(n7153) );
  NAND3HSV4 U9207 ( .A1(n7159), .A2(n7158), .A3(n7156), .ZN(n7154) );
  CLKNHSV2 U9208 ( .I(n11417), .ZN(n7156) );
  CLKNHSV2 U9209 ( .I(n11444), .ZN(n11449) );
  INAND2HSV2 U9210 ( .A1(n13468), .B1(n7162), .ZN(n7161) );
  NOR2HSV2 U9211 ( .A1(n13467), .A2(n13466), .ZN(n7162) );
  XNOR2HSV2 U9212 ( .A1(n13465), .A2(n13464), .ZN(n7163) );
  NAND2HSV2 U9213 ( .A1(\pe10/ti_7[5] ), .A2(\pe10/got [4]), .ZN(n7164) );
  OAI21HSV4 U9214 ( .A1(n15237), .A2(n11091), .B(n7953), .ZN(n11122) );
  XNOR2HSV4 U9215 ( .A1(n9115), .A2(n9114), .ZN(n7165) );
  AOI21HSV4 U9216 ( .A1(n9102), .A2(n8948), .B(n9101), .ZN(n7166) );
  CLKNAND2HSV2 U9217 ( .A1(\pe6/ti_1 ), .A2(\pe6/got [7]), .ZN(n9236) );
  AOI22HSV4 U9218 ( .A1(\pe3/ti_7t [2]), .A2(n10942), .B1(n10185), .B2(n13842), 
        .ZN(n7168) );
  CLKNAND2HSV4 U9219 ( .A1(n7168), .A2(n7167), .ZN(n10202) );
  XNOR2HSV4 U9220 ( .A1(n7170), .A2(n7169), .ZN(n10408) );
  CLKNAND2HSV2 U9221 ( .A1(n10202), .A2(n14931), .ZN(n7169) );
  XNOR2HSV4 U9222 ( .A1(n7171), .A2(n10200), .ZN(n7170) );
  XOR3HSV2 U9223 ( .A1(\pe3/phq [4]), .A2(n7173), .A3(n10198), .Z(n7172) );
  CLKNHSV2 U9224 ( .I(n10199), .ZN(n7173) );
  CLKNHSV2 U9225 ( .I(n12316), .ZN(n7176) );
  INHSV24 U9226 ( .I(n13284), .ZN(n7182) );
  CLKNHSV2 U9227 ( .I(n10307), .ZN(n7184) );
  CLKNAND2HSV2 U9228 ( .A1(n15276), .A2(n10307), .ZN(n13285) );
  CLKNAND2HSV2 U9229 ( .A1(n7188), .A2(n11495), .ZN(n7185) );
  CLKNHSV2 U9230 ( .I(n7188), .ZN(n7187) );
  CLKNAND2HSV2 U9231 ( .A1(n10329), .A2(n10330), .ZN(n7188) );
  CLKNHSV4 U9232 ( .I(n11495), .ZN(n7189) );
  XNOR2HSV4 U9233 ( .A1(n7195), .A2(n7190), .ZN(n10634) );
  XNOR2HSV4 U9234 ( .A1(n7194), .A2(n7191), .ZN(n7190) );
  XNOR2HSV4 U9235 ( .A1(n10623), .A2(n7192), .ZN(n7191) );
  XNOR2HSV4 U9236 ( .A1(n7193), .A2(n10615), .ZN(n7192) );
  CLKNAND2HSV2 U9237 ( .A1(\pe1/ti_7[2] ), .A2(\pe1/got [4]), .ZN(n7193) );
  NOR2HSV4 U9238 ( .A1(n13953), .A2(n10625), .ZN(n7194) );
  AOI21HSV4 U9239 ( .A1(pov1[3]), .A2(n10228), .B(n10624), .ZN(n13953) );
  CLKNAND2HSV2 U9240 ( .A1(n7268), .A2(n8510), .ZN(pov1[3]) );
  CLKNAND2HSV2 U9241 ( .A1(n14847), .A2(\pe1/got [6]), .ZN(n7195) );
  CLKNAND2HSV2 U9242 ( .A1(n10627), .A2(n10626), .ZN(n14847) );
  NAND3HSV4 U9243 ( .A1(n13859), .A2(n10228), .A3(n13860), .ZN(n10626) );
  NOR2HSV4 U9244 ( .A1(n12195), .A2(n10680), .ZN(n7409) );
  CLKNHSV2 U9245 ( .I(n7983), .ZN(n7196) );
  CLKNHSV2 U9246 ( .I(n7982), .ZN(n7197) );
  CLKNAND2HSV4 U9247 ( .A1(\pe14/aot [7]), .A2(\pe14/bq[8] ), .ZN(n9086) );
  CLKNHSV2 U9248 ( .I(n9139), .ZN(n7198) );
  XNOR2HSV4 U9249 ( .A1(n9138), .A2(n9137), .ZN(n7199) );
  CLKNHSV2 U9250 ( .I(n7200), .ZN(n10374) );
  CLKNAND2HSV2 U9251 ( .A1(n10375), .A2(n7201), .ZN(n7200) );
  CLKNAND2HSV2 U9252 ( .A1(n10873), .A2(n10837), .ZN(n7201) );
  INAND2HSV4 U9253 ( .A1(n10873), .B1(\pe21/ti_7t [2]), .ZN(n10375) );
  XNOR2HSV4 U9254 ( .A1(n11855), .A2(n7202), .ZN(n11872) );
  CLKNAND2HSV2 U9255 ( .A1(n14960), .A2(\pe20/got [4]), .ZN(n7202) );
  CLKNAND2HSV2 U9256 ( .A1(n7411), .A2(n9070), .ZN(n14960) );
  CLKNAND2HSV2 U9257 ( .A1(n13848), .A2(n9035), .ZN(n9070) );
  CLKNAND2HSV2 U9258 ( .A1(n7567), .A2(n7571), .ZN(n7203) );
  CLKNHSV2 U9259 ( .I(n11443), .ZN(n7205) );
  NOR2HSV2 U9260 ( .A1(n10705), .A2(n7207), .ZN(n7523) );
  CLKNHSV2 U9261 ( .I(n11207), .ZN(n7207) );
  CLKNAND2HSV3 U9262 ( .A1(n7208), .A2(\pe5/phq [2]), .ZN(n7210) );
  XNOR2HSV4 U9263 ( .A1(n7209), .A2(n7213), .ZN(n10311) );
  CLKNAND2HSV2 U9264 ( .A1(n7211), .A2(n7210), .ZN(n7209) );
  CLKNHSV2 U9265 ( .I(\pe5/phq [2]), .ZN(n7212) );
  CLKNHSV2 U9266 ( .I(n11477), .ZN(n7213) );
  CLKNAND2HSV2 U9267 ( .A1(\pe5/bq[7] ), .A2(\pe5/aot [8]), .ZN(n11477) );
  CLKNAND2HSV2 U9268 ( .A1(n9480), .A2(n9481), .ZN(n9479) );
  XNOR2HSV4 U9269 ( .A1(n9478), .A2(n7214), .ZN(n9481) );
  XNOR2HSV4 U9270 ( .A1(n9477), .A2(n7215), .ZN(n7214) );
  CLKNAND2HSV2 U9271 ( .A1(n13738), .A2(\pe20/got [3]), .ZN(n7215) );
  CLKNAND2HSV2 U9272 ( .A1(n8951), .A2(\pe20/got [4]), .ZN(n9480) );
  CLKNAND2HSV2 U9273 ( .A1(n7216), .A2(n9062), .ZN(n8951) );
  CLKNAND2HSV2 U9274 ( .A1(n9061), .A2(n10412), .ZN(n7216) );
  OAI21HSV4 U9275 ( .A1(n7220), .A2(n7218), .B(n7217), .ZN(n11568) );
  CLKNAND2HSV2 U9276 ( .A1(n7220), .A2(n7218), .ZN(n7217) );
  CLKNHSV2 U9277 ( .I(n7219), .ZN(n7218) );
  CLKNAND2HSV2 U9278 ( .A1(n14950), .A2(\pe8/bq[3] ), .ZN(n7219) );
  NOR2HSV4 U9279 ( .A1(n11567), .A2(n13516), .ZN(n7220) );
  AOI21HSV4 U9280 ( .A1(n10972), .A2(n10971), .B(n7222), .ZN(n7221) );
  CLKNHSV2 U9281 ( .I(\pe3/got [5]), .ZN(n7222) );
  XNOR2HSV4 U9282 ( .A1(n7224), .A2(n10973), .ZN(n7223) );
  CLKNAND2HSV2 U9283 ( .A1(n14872), .A2(\pe3/got [4]), .ZN(n7224) );
  AOI21HSV4 U9284 ( .A1(n7441), .A2(n7227), .B(n7226), .ZN(n7225) );
  CLKNHSV2 U9285 ( .I(n9845), .ZN(n7226) );
  CLKNHSV2 U9286 ( .I(n9536), .ZN(n7227) );
  CLKNHSV2 U9287 ( .I(n7441), .ZN(n7228) );
  MUX2NHSV4 U9288 ( .I0(n9320), .I1(n9319), .S(n9318), .ZN(n12369) );
  CLKNAND2HSV4 U9289 ( .A1(n7229), .A2(n10088), .ZN(n14874) );
  CLKNAND2HSV2 U9290 ( .A1(n7231), .A2(n7230), .ZN(n7236) );
  CLKNHSV2 U9291 ( .I(n7232), .ZN(n7231) );
  CLKNAND2HSV2 U9292 ( .A1(\pe10/bq[8] ), .A2(\pe10/aot [7]), .ZN(n7233) );
  CLKNAND2HSV3 U9293 ( .A1(n7238), .A2(n7237), .ZN(n7234) );
  INHSV2 U9294 ( .I(n7236), .ZN(n7235) );
  XOR2HSV2 U9295 ( .A1(n13019), .A2(n7239), .Z(n15275) );
  CLKNHSV2 U9296 ( .I(n12790), .ZN(n7240) );
  CLKNAND2HSV2 U9297 ( .A1(n7243), .A2(n12775), .ZN(n13306) );
  CLKNAND2HSV3 U9298 ( .A1(n12789), .A2(n12788), .ZN(n13304) );
  CLKNHSV2 U9299 ( .I(n7244), .ZN(n7243) );
  CLKNAND2HSV3 U9300 ( .A1(\pe16/bq[8] ), .A2(\pe16/aot [8]), .ZN(n7246) );
  CLKNAND2HSV3 U9301 ( .A1(\pe16/pvq [1]), .A2(\pe16/ctrq ), .ZN(n7245) );
  CLKNAND2HSV2 U9302 ( .A1(\pe16/got [8]), .A2(\pe16/ti_1 ), .ZN(n7247) );
  CLKNAND2HSV4 U9303 ( .A1(n14874), .A2(\pe10/got [6]), .ZN(n7250) );
  XNOR2HSV4 U9304 ( .A1(n7250), .A2(n7249), .ZN(n7248) );
  XNOR2HSV4 U9305 ( .A1(n10039), .A2(n10038), .ZN(n7249) );
  CLKNHSV4 U9306 ( .I(\pe20/ctrq ), .ZN(n11795) );
  CLKNAND2HSV2 U9307 ( .A1(n8749), .A2(n8748), .ZN(n8750) );
  OAI22HSV4 U9308 ( .A1(n13652), .A2(n13653), .B1(n7253), .B2(n7252), .ZN(
        n8749) );
  CLKNHSV2 U9309 ( .I(n13651), .ZN(n7252) );
  CLKNHSV2 U9310 ( .I(n7254), .ZN(n7253) );
  CLKNAND2HSV2 U9311 ( .A1(n13650), .A2(n13649), .ZN(n7254) );
  OAI21HSV4 U9312 ( .A1(n7259), .A2(n7256), .B(n7255), .ZN(n8636) );
  CLKNAND2HSV2 U9313 ( .A1(n7256), .A2(n7259), .ZN(n7255) );
  XNOR2HSV4 U9314 ( .A1(n7258), .A2(n7257), .ZN(n7256) );
  CLKNHSV2 U9315 ( .I(n8635), .ZN(n7258) );
  NOR2HSV4 U9316 ( .A1(n13809), .A2(n8630), .ZN(n7259) );
  OAI21HSV4 U9317 ( .A1(n7267), .A2(n7261), .B(n7260), .ZN(n8149) );
  CLKNAND2HSV2 U9318 ( .A1(n7261), .A2(n7267), .ZN(n7260) );
  XNOR2HSV4 U9319 ( .A1(n7263), .A2(n7262), .ZN(n7261) );
  CLKNHSV2 U9320 ( .I(n8148), .ZN(n7262) );
  CLKNAND2HSV2 U9321 ( .A1(n8147), .A2(n7264), .ZN(n7263) );
  CLKNAND2HSV2 U9322 ( .A1(n7266), .A2(n7265), .ZN(n7264) );
  CLKNHSV2 U9323 ( .I(n8146), .ZN(n7265) );
  CLKNHSV2 U9324 ( .I(n8145), .ZN(n7266) );
  NOR2HSV4 U9325 ( .A1(n14005), .A2(n8139), .ZN(n7267) );
  AOI21HSV4 U9326 ( .A1(pov1[3]), .A2(n10631), .B(n10624), .ZN(n14005) );
  CLKNAND2HSV2 U9327 ( .A1(n7270), .A2(n7269), .ZN(n7268) );
  CLKNHSV2 U9328 ( .I(n8509), .ZN(n7269) );
  CLKNHSV2 U9329 ( .I(n10264), .ZN(n7270) );
  CLKNAND2HSV2 U9330 ( .A1(\pe8/got [8]), .A2(\pe8/ti_1 ), .ZN(n10484) );
  NOR2HSV4 U9331 ( .A1(n7271), .A2(n7743), .ZN(n12511) );
  NOR2HSV4 U9332 ( .A1(n13886), .A2(n7745), .ZN(n7271) );
  XNOR2HSV4 U9333 ( .A1(n7748), .A2(n7747), .ZN(n13886) );
  NOR2HSV4 U9334 ( .A1(n11517), .A2(n11518), .ZN(n7274) );
  OAI21HSV4 U9335 ( .A1(n11516), .A2(n7276), .B(n7275), .ZN(n11518) );
  CLKNAND2HSV2 U9336 ( .A1(n11511), .A2(n11512), .ZN(n7276) );
  NOR2HSV4 U9337 ( .A1(n15079), .A2(n10509), .ZN(n11516) );
  XNOR2HSV4 U9338 ( .A1(n7277), .A2(n11510), .ZN(n11517) );
  XNOR2HSV4 U9339 ( .A1(n11509), .A2(n11508), .ZN(n7277) );
  CLKNAND2HSV3 U9340 ( .A1(n12193), .A2(n12192), .ZN(n14388) );
  XNOR2HSV4 U9341 ( .A1(n7278), .A2(n7279), .ZN(n15255) );
  XNOR2HSV4 U9342 ( .A1(n7678), .A2(n7675), .ZN(n7278) );
  AOI21HSV4 U9343 ( .A1(n11899), .A2(n11776), .B(n7672), .ZN(n7279) );
  INHSV24 U9344 ( .I(n10509), .ZN(n7280) );
  XNOR2HSV4 U9345 ( .A1(n11536), .A2(n7281), .ZN(n13862) );
  XNOR2HSV4 U9346 ( .A1(n11535), .A2(n7282), .ZN(n7281) );
  MUX2NHSV2 U9347 ( .I0(n11523), .I1(n8336), .S(n8337), .ZN(n15267) );
  NOR2HSV4 U9348 ( .A1(n11343), .A2(n11373), .ZN(n11408) );
  CLKNAND2HSV2 U9349 ( .A1(n7285), .A2(n7283), .ZN(n11342) );
  CLKNHSV2 U9350 ( .I(n7284), .ZN(n7283) );
  CLKNAND2HSV0 U9351 ( .A1(n11324), .A2(n11296), .ZN(n7284) );
  CLKNHSV2 U9352 ( .I(n11297), .ZN(n7285) );
  CLKNAND2HSV2 U9353 ( .A1(n11371), .A2(n11339), .ZN(n11343) );
  CLKNAND2HSV2 U9354 ( .A1(n7286), .A2(n11340), .ZN(n11371) );
  XNOR2HSV4 U9355 ( .A1(n11290), .A2(n11289), .ZN(n11340) );
  CLKNHSV2 U9356 ( .I(n11338), .ZN(n7286) );
  OAI22HSV2 U9357 ( .A1(n8082), .A2(n7287), .B1(n8081), .B2(n11523), .ZN(n7289) );
  CLKNAND2HSV2 U9358 ( .A1(n7288), .A2(n7290), .ZN(n7287) );
  CLKNHSV2 U9359 ( .I(n8081), .ZN(n7288) );
  INHSV2 U9360 ( .I(n11538), .ZN(n7290) );
  NAND3HSV4 U9361 ( .A1(n7292), .A2(n7293), .A3(n7291), .ZN(n7320) );
  CLKNHSV2 U9362 ( .I(n7980), .ZN(n7291) );
  CLKNAND2HSV2 U9363 ( .A1(\pe16/pvq [2]), .A2(\pe16/ctrq ), .ZN(n7980) );
  CLKNAND2HSV2 U9364 ( .A1(n14960), .A2(\pe20/got [6]), .ZN(n7294) );
  XNOR2HSV4 U9365 ( .A1(n7298), .A2(n7296), .ZN(n7295) );
  XNOR2HSV4 U9366 ( .A1(n9067), .A2(n7297), .ZN(n7296) );
  XOR2HSV2 U9367 ( .A1(n9066), .A2(\pe20/phq [5]), .Z(n7297) );
  XNOR2HSV4 U9368 ( .A1(n7300), .A2(n7299), .ZN(n7298) );
  XOR2HSV2 U9369 ( .A1(n9069), .A2(n9068), .Z(n7299) );
  XNOR2HSV4 U9370 ( .A1(n9065), .A2(n7301), .ZN(n7300) );
  CLKNAND2HSV2 U9371 ( .A1(n12362), .A2(\pe20/pvq [5]), .ZN(n7301) );
  CLKNHSV2 U9372 ( .I(n7302), .ZN(n12411) );
  AOI22HSV4 U9373 ( .A1(n10520), .A2(n14704), .B1(n15235), .B2(n10519), .ZN(
        n7303) );
  CLKNHSV1 U9374 ( .I(n10523), .ZN(n7305) );
  AOI21HSV4 U9375 ( .A1(n7307), .A2(n7306), .B(n8981), .ZN(n9341) );
  CLKNHSV2 U9376 ( .I(n8980), .ZN(n7306) );
  CLKNAND2HSV2 U9377 ( .A1(n8990), .A2(\pe2/got [7]), .ZN(n8991) );
  CLKNHSV2 U9378 ( .I(n8979), .ZN(n7308) );
  CLKNAND2HSV2 U9379 ( .A1(n11778), .A2(n7309), .ZN(n9342) );
  CLKNAND2HSV2 U9380 ( .A1(n8978), .A2(n8982), .ZN(n11778) );
  NOR2HSV8 U9381 ( .A1(n15196), .A2(n14866), .ZN(n11692) );
  XNOR2HSV4 U9382 ( .A1(n7314), .A2(n7310), .ZN(n15196) );
  AOI21HSV4 U9383 ( .A1(n7313), .A2(n7312), .B(n7311), .ZN(n7310) );
  NOR2HSV4 U9384 ( .A1(n15069), .A2(n14866), .ZN(n7313) );
  XNOR2HSV4 U9385 ( .A1(n9436), .A2(n7315), .ZN(n7314) );
  CLKNAND2HSV2 U9386 ( .A1(n7318), .A2(n7317), .ZN(n7316) );
  CLKNAND2HSV2 U9387 ( .A1(n7560), .A2(n6830), .ZN(n7317) );
  CLKNAND2HSV2 U9388 ( .A1(n7319), .A2(n7561), .ZN(n7318) );
  CLKNAND2HSV4 U9389 ( .A1(n7320), .A2(n7981), .ZN(n7321) );
  CLKNAND2HSV2 U9390 ( .A1(n10593), .A2(n7892), .ZN(n7322) );
  NAND3HSV4 U9391 ( .A1(n7361), .A2(n7735), .A3(n10188), .ZN(n7360) );
  BUFHSV8 U9392 ( .I(n10408), .Z(n7323) );
  XNOR2HSV4 U9393 ( .A1(n8496), .A2(n7325), .ZN(n8497) );
  XNOR2HSV4 U9394 ( .A1(n7328), .A2(n7326), .ZN(n7807) );
  NOR2HSV2 U9395 ( .A1(n10216), .A2(n7327), .ZN(n7326) );
  CLKNHSV2 U9396 ( .I(\pe3/got [6]), .ZN(n7327) );
  XNOR2HSV4 U9397 ( .A1(n10215), .A2(n7329), .ZN(n7328) );
  CLKNAND2HSV2 U9398 ( .A1(\pe3/ti_7[1] ), .A2(\pe3/got [5]), .ZN(n7329) );
  CLKNAND2HSV2 U9399 ( .A1(n10214), .A2(n10213), .ZN(\pe3/ti_7[1] ) );
  CLKNAND2HSV2 U9400 ( .A1(n7330), .A2(n11160), .ZN(\pe16/ti_7[3] ) );
  CLKNHSV2 U9401 ( .I(n10729), .ZN(n7332) );
  CLKNAND2HSV2 U9402 ( .A1(n15253), .A2(n11469), .ZN(n10731) );
  CLKNAND2HSV2 U9403 ( .A1(n15253), .A2(n10747), .ZN(n7431) );
  AOI21HSV2 U9404 ( .A1(n15253), .A2(\pe12/got [8]), .B(n11471), .ZN(n10744)
         );
  CLKBUFHSV2 U9405 ( .I(n7334), .Z(n7333) );
  CLKNAND2HSV2 U9406 ( .A1(n7334), .A2(\pe18/got [7]), .ZN(n9172) );
  CLKNAND2HSV2 U9407 ( .A1(n7333), .A2(\pe18/got [3]), .ZN(n13149) );
  CLKNAND2HSV2 U9408 ( .A1(n7333), .A2(\pe18/got [2]), .ZN(n14638) );
  CLKNAND2HSV2 U9409 ( .A1(n7333), .A2(\pe18/got [1]), .ZN(n13363) );
  CLKNHSV2 U9410 ( .I(n12347), .ZN(n7335) );
  CLKNHSV2 U9411 ( .I(n12337), .ZN(n7337) );
  CLKNAND2HSV2 U9412 ( .A1(n8393), .A2(n8392), .ZN(n8394) );
  CLKNAND2HSV0 U9413 ( .A1(n7339), .A2(n11440), .ZN(n7573) );
  CLKNAND2HSV2 U9414 ( .A1(n11441), .A2(n7339), .ZN(n7338) );
  CLKNAND2HSV1 U9415 ( .A1(n7341), .A2(n7340), .ZN(n7339) );
  NOR2HSV0 U9416 ( .A1(n11436), .A2(n11447), .ZN(n7340) );
  INHSV2 U9417 ( .I(n11437), .ZN(n7341) );
  CLKNAND2HSV2 U9418 ( .A1(\pe7/ti_7[1] ), .A2(\pe7/got [5]), .ZN(n12242) );
  CLKNAND2HSV2 U9419 ( .A1(n7342), .A2(n11783), .ZN(\pe7/ti_7[1] ) );
  CLKNAND2HSV2 U9420 ( .A1(n15273), .A2(n11782), .ZN(n7342) );
  XNOR2HSV4 U9421 ( .A1(n7344), .A2(n7343), .ZN(n15273) );
  XNOR2HSV4 U9422 ( .A1(n7619), .A2(\pe7/phq [1]), .ZN(n7343) );
  XNOR2HSV4 U9423 ( .A1(n7621), .A2(n7620), .ZN(n7344) );
  XNOR2HSV4 U9424 ( .A1(n7348), .A2(n7345), .ZN(n10793) );
  XNOR2HSV4 U9425 ( .A1(n7347), .A2(n7346), .ZN(n7345) );
  CLKNAND2HSV2 U9426 ( .A1(\pe15/bq[6] ), .A2(\pe15/aot [8]), .ZN(n7346) );
  XNOR2HSV4 U9427 ( .A1(n11304), .A2(n7349), .ZN(n7348) );
  CLKNAND2HSV2 U9428 ( .A1(\pe15/ti_1 ), .A2(\pe15/got [6]), .ZN(n7349) );
  CLKNAND2HSV2 U9429 ( .A1(\pe15/bq[8] ), .A2(\pe15/aot [6]), .ZN(n11304) );
  CLKNAND2HSV2 U9430 ( .A1(n7350), .A2(n8023), .ZN(n8026) );
  CLKNHSV2 U9431 ( .I(n7564), .ZN(n7350) );
  AOI21HSV4 U9432 ( .A1(n7353), .A2(n7352), .B(n7351), .ZN(n7564) );
  CLKNHSV2 U9433 ( .I(n8024), .ZN(n7351) );
  CLKNHSV2 U9434 ( .I(n8025), .ZN(n7352) );
  CLKNHSV2 U9435 ( .I(n15251), .ZN(n7353) );
  CLKNHSV2 U9436 ( .I(n7813), .ZN(n9835) );
  NOR2HSV4 U9437 ( .A1(n7688), .A2(n7687), .ZN(n7354) );
  CLKNHSV2 U9438 ( .I(n7689), .ZN(n7356) );
  CLKNHSV2 U9439 ( .I(n9834), .ZN(n7357) );
  OAI21HSV4 U9440 ( .A1(n10993), .A2(n10939), .B(n10992), .ZN(n8005) );
  AOI21HSV4 U9441 ( .A1(n7323), .A2(n7358), .B(n10944), .ZN(n10992) );
  CLKNHSV2 U9442 ( .I(n7359), .ZN(n7358) );
  CLKNAND2HSV2 U9443 ( .A1(n7365), .A2(n7364), .ZN(n7363) );
  CLKNHSV2 U9444 ( .I(n8736), .ZN(n7364) );
  XNOR2HSV4 U9445 ( .A1(n12202), .A2(n14860), .ZN(n7365) );
  OAI21HSV2 U9446 ( .A1(n14582), .A2(n8428), .B(n7497), .ZN(n7366) );
  OAI21HSV4 U9447 ( .A1(n11343), .A2(n11373), .B(n7369), .ZN(n7368) );
  INHSV2 U9448 ( .I(n11702), .ZN(n7371) );
  CLKNHSV3 U9449 ( .I(n12320), .ZN(n7372) );
  CLKNHSV2 U9450 ( .I(n7373), .ZN(n8907) );
  XNOR2HSV4 U9451 ( .A1(n13621), .A2(n13624), .ZN(\pov7[5] ) );
  CLKNAND2HSV3 U9452 ( .A1(n7374), .A2(n13620), .ZN(\pe7/ti_7[5] ) );
  CLKNAND2HSV0 U9453 ( .A1(\pe7/ti_7[5] ), .A2(\pe7/got [1]), .ZN(n8523) );
  CLKNHSV2 U9454 ( .I(n9450), .ZN(n7375) );
  CLKNAND2HSV2 U9455 ( .A1(n12148), .A2(\pe19/got [5]), .ZN(n12169) );
  CLKNAND2HSV2 U9456 ( .A1(n7376), .A2(n10468), .ZN(n12148) );
  CLKNAND2HSV2 U9457 ( .A1(n9581), .A2(n13844), .ZN(n7377) );
  XNOR2HSV4 U9458 ( .A1(n9499), .A2(n9498), .ZN(n9540) );
  CLKNHSV0 U9459 ( .I(n14821), .ZN(n12048) );
  CLKNAND2HSV2 U9460 ( .A1(\pe6/aot [8]), .A2(\pe6/bq[8] ), .ZN(n8303) );
  AOI22HSV4 U9461 ( .A1(\pe5/ti_7t [2]), .A2(n10322), .B1(n8904), .B2(n10312), 
        .ZN(n7385) );
  INHSV2 U9462 ( .I(n10331), .ZN(n7378) );
  CLKNAND2HSV2 U9463 ( .A1(n13015), .A2(\pe5/ti_7t [3]), .ZN(n7379) );
  INAND2HSV4 U9464 ( .A1(n7383), .B1(n7378), .ZN(n7381) );
  XNOR2HSV4 U9465 ( .A1(n7679), .A2(n10319), .ZN(n7382) );
  XNOR2HSV4 U9466 ( .A1(n7387), .A2(n10027), .ZN(n7386) );
  AOI21HSV4 U9467 ( .A1(n10006), .A2(n10005), .B(n10004), .ZN(n7387) );
  CLKNAND2HSV2 U9468 ( .A1(n13604), .A2(\pe13/got [7]), .ZN(n7388) );
  CLKNAND2HSV0 U9469 ( .A1(n9763), .A2(\pe9/got [6]), .ZN(n9418) );
  INHSV2 U9470 ( .I(n9399), .ZN(n7389) );
  XNOR2HSV4 U9471 ( .A1(n10781), .A2(n7393), .ZN(n7392) );
  CLKNAND2HSV2 U9472 ( .A1(n14255), .A2(\pe12/got [6]), .ZN(n7393) );
  XNOR2HSV4 U9473 ( .A1(n11436), .A2(n11434), .ZN(n15251) );
  CLKNAND2HSV2 U9474 ( .A1(n12276), .A2(n12252), .ZN(n7394) );
  CLKNHSV2 U9475 ( .I(n7396), .ZN(n7395) );
  OAI21HSV4 U9476 ( .A1(n12252), .A2(n7397), .B(\pe7/got [6]), .ZN(n7396) );
  CLKNHSV2 U9477 ( .I(n12277), .ZN(n7397) );
  NAND2HSV3 U9478 ( .A1(n12265), .A2(n12264), .ZN(n12276) );
  CLKNHSV2 U9479 ( .I(n9725), .ZN(n9728) );
  CLKNHSV2 U9480 ( .I(n9722), .ZN(n7398) );
  OAI21HSV4 U9481 ( .A1(n15211), .A2(n9565), .B(n8032), .ZN(n7751) );
  INAND3HSV4 U9482 ( .A1(n7402), .B1(n7401), .B2(n7399), .ZN(n15211) );
  CLKNHSV2 U9483 ( .I(n7400), .ZN(n7399) );
  CLKNAND2HSV4 U9484 ( .A1(n9515), .A2(n9541), .ZN(n9727) );
  XNOR2HSV4 U9485 ( .A1(n9532), .A2(n9531), .ZN(n9725) );
  CLKNAND2HSV2 U9486 ( .A1(n7583), .A2(\pe13/aot [5]), .ZN(n9894) );
  CLKNAND2HSV2 U9487 ( .A1(n7583), .A2(\pe13/aot [2]), .ZN(n9968) );
  MUX2NHSV2 U9488 ( .I0(n7404), .I1(n7403), .S(n13820), .ZN(n15147) );
  CLKNHSV2 U9489 ( .I(n7583), .ZN(n7403) );
  CLKNHSV2 U9490 ( .I(bo13[8]), .ZN(n7404) );
  INHSV24 U9491 ( .I(n7407), .ZN(n7405) );
  NOR2HSV4 U9492 ( .A1(n10873), .A2(\pe21/ti_7t [5]), .ZN(n7407) );
  CLKNAND2HSV2 U9493 ( .A1(\pe7/aot [8]), .A2(\pe7/bq[4] ), .ZN(n7962) );
  XNOR2HSV4 U9494 ( .A1(n7408), .A2(n11295), .ZN(n15233) );
  CLKNAND2HSV2 U9495 ( .A1(n11390), .A2(n15178), .ZN(n7408) );
  CLKNHSV1 U9496 ( .I(n7983), .ZN(n7410) );
  NOR2HSV4 U9497 ( .A1(n10409), .A2(n15177), .ZN(n9060) );
  XOR2HSV4 U9498 ( .A1(n7417), .A2(n9058), .Z(n10409) );
  XNOR2HSV4 U9499 ( .A1(n7412), .A2(n7416), .ZN(n9058) );
  XNOR2HSV4 U9500 ( .A1(n7415), .A2(n7413), .ZN(n7412) );
  XNOR2HSV4 U9501 ( .A1(n7414), .A2(n9019), .ZN(n7413) );
  XNOR2HSV4 U9502 ( .A1(n9018), .A2(n9020), .ZN(n7415) );
  NOR2HSV4 U9503 ( .A1(n9038), .A2(n9012), .ZN(n7416) );
  XNOR2HSV4 U9504 ( .A1(n7422), .A2(n7418), .ZN(n14011) );
  OAI21HSV4 U9505 ( .A1(n7421), .A2(n7420), .B(n7419), .ZN(n7418) );
  NOR2HSV4 U9506 ( .A1(n7427), .A2(n12105), .ZN(n7419) );
  CLKNHSV2 U9507 ( .I(n12108), .ZN(n7420) );
  NOR2HSV4 U9508 ( .A1(n10440), .A2(n7426), .ZN(n7425) );
  CLKNHSV2 U9509 ( .I(n7790), .ZN(n7426) );
  NOR2HSV4 U9510 ( .A1(n12108), .A2(n7428), .ZN(n7427) );
  CLKNAND2HSV2 U9511 ( .A1(n12107), .A2(n7429), .ZN(n7428) );
  CLKNHSV2 U9512 ( .I(n7789), .ZN(n7429) );
  XNOR2HSV4 U9513 ( .A1(n7432), .A2(n7430), .ZN(n10781) );
  CLKNAND2HSV2 U9514 ( .A1(\pe12/ti_7[1] ), .A2(\pe12/got [5]), .ZN(n7430) );
  XNOR2HSV4 U9515 ( .A1(n10780), .A2(n7433), .ZN(n7432) );
  XNOR2HSV4 U9516 ( .A1(n7434), .A2(n10773), .ZN(n7433) );
  XOR2HSV2 U9517 ( .A1(n10772), .A2(\pe12/phq [5]), .Z(n7434) );
  CLKNHSV2 U9518 ( .I(n11704), .ZN(n7435) );
  NOR2HSV4 U9519 ( .A1(n7438), .A2(n7816), .ZN(n7437) );
  CLKNHSV2 U9520 ( .I(n7764), .ZN(n7438) );
  CLKNHSV2 U9521 ( .I(n7816), .ZN(n7439) );
  CLKNHSV3 U9522 ( .I(n7817), .ZN(n7441) );
  CLKNHSV2 U9523 ( .I(n10767), .ZN(n7442) );
  XNOR2HSV4 U9524 ( .A1(n7444), .A2(n7443), .ZN(n10767) );
  XNOR2HSV4 U9525 ( .A1(n10763), .A2(n10762), .ZN(n7444) );
  AOI21HSV4 U9526 ( .A1(n7445), .A2(n10747), .B(n10746), .ZN(n10766) );
  XNOR2HSV4 U9527 ( .A1(n11434), .A2(n15192), .ZN(n7445) );
  CLKNHSV2 U9528 ( .I(n10119), .ZN(n7447) );
  CLKNAND2HSV0 U9529 ( .A1(n7448), .A2(n10071), .ZN(n10075) );
  CLKNHSV2 U9530 ( .I(n10127), .ZN(n7449) );
  XNOR2HSV4 U9531 ( .A1(n7451), .A2(n7450), .ZN(n9055) );
  CLKNAND2HSV2 U9532 ( .A1(n9057), .A2(n13718), .ZN(n7450) );
  XNOR2HSV4 U9533 ( .A1(n9052), .A2(n7452), .ZN(n7451) );
  XNOR2HSV4 U9534 ( .A1(n7454), .A2(n7453), .ZN(n7452) );
  XNOR2HSV4 U9535 ( .A1(n9046), .A2(n9050), .ZN(n7453) );
  XNOR2HSV4 U9536 ( .A1(n7455), .A2(n9051), .ZN(n7454) );
  CLKNAND2HSV2 U9537 ( .A1(n12256), .A2(n12257), .ZN(n13883) );
  AOI21HSV4 U9538 ( .A1(n7459), .A2(n7458), .B(n7457), .ZN(n12256) );
  CLKNHSV2 U9539 ( .I(n7460), .ZN(n7457) );
  NAND3HSV4 U9540 ( .A1(n7456), .A2(n13883), .A3(n12308), .ZN(n12258) );
  CLKNHSV2 U9541 ( .I(n8211), .ZN(n7460) );
  CLKNAND2HSV2 U9542 ( .A1(n12227), .A2(n12226), .ZN(n7461) );
  OAI21HSV4 U9543 ( .A1(n12200), .A2(n12199), .B(n12198), .ZN(n7462) );
  AOI21HSV4 U9544 ( .A1(n7464), .A2(n10412), .B(n10411), .ZN(n11854) );
  CLKNHSV2 U9545 ( .I(n10409), .ZN(n7464) );
  CLKBUFHSV2 U9546 ( .I(n8951), .Z(n7465) );
  CLKNAND2HSV2 U9547 ( .A1(n8951), .A2(\pe20/got [5]), .ZN(n9072) );
  CLKNAND2HSV2 U9548 ( .A1(n7465), .A2(\pe20/got [3]), .ZN(n11855) );
  CLKNAND2HSV2 U9549 ( .A1(n7465), .A2(\pe20/got [1]), .ZN(n13708) );
  CLKNAND2HSV2 U9550 ( .A1(n7465), .A2(\pe20/got [2]), .ZN(n13721) );
  CLKNAND2HSV2 U9551 ( .A1(n7465), .A2(n14865), .ZN(n8876) );
  OAI21HSV2 U9552 ( .A1(n7467), .A2(n9834), .B(n9264), .ZN(n7466) );
  NOR2HSV3 U9553 ( .A1(n7469), .A2(n9842), .ZN(n7468) );
  CLKNHSV3 U9554 ( .I(n9835), .ZN(n7469) );
  XNOR2HSV4 U9555 ( .A1(n7472), .A2(n7470), .ZN(n15241) );
  XNOR2HSV4 U9556 ( .A1(n9953), .A2(n9954), .ZN(n9992) );
  CLKNHSV2 U9557 ( .I(n11120), .ZN(n7473) );
  CLKNAND2HSV2 U9558 ( .A1(n8098), .A2(n8099), .ZN(n8100) );
  CLKNAND2HSV2 U9559 ( .A1(\pe19/aot [8]), .A2(\pe19/bq[8] ), .ZN(n8099) );
  CLKNAND2HSV2 U9560 ( .A1(\pe19/pvq [1]), .A2(\pe19/ctrq ), .ZN(n8098) );
  NAND3HSV2 U9561 ( .A1(n7476), .A2(n7475), .A3(n7474), .ZN(n7872) );
  CLKNHSV2 U9562 ( .I(n8464), .ZN(n7474) );
  CLKNAND2HSV4 U9563 ( .A1(\pe17/bq[6] ), .A2(\pe17/aot [7]), .ZN(n8464) );
  CLKNHSV2 U9564 ( .I(n10978), .ZN(n10805) );
  XNOR2HSV4 U9565 ( .A1(n10205), .A2(n7477), .ZN(n10212) );
  XOR2HSV2 U9566 ( .A1(n7478), .A2(n8841), .Z(n7477) );
  NOR2HSV4 U9567 ( .A1(n10978), .A2(n7479), .ZN(n7478) );
  CLKNHSV2 U9568 ( .I(\pe3/pvq [5]), .ZN(n7479) );
  CLKNHSV2 U9569 ( .I(n9745), .ZN(n9789) );
  CLKNAND2HSV2 U9570 ( .A1(n13910), .A2(n7480), .ZN(n11611) );
  NOR2HSV4 U9571 ( .A1(n9745), .A2(n7481), .ZN(n7480) );
  CLKNHSV2 U9572 ( .I(n11691), .ZN(n7481) );
  CLKNHSV2 U9573 ( .I(n11612), .ZN(n7482) );
  CLKNAND2HSV2 U9574 ( .A1(n9745), .A2(n7484), .ZN(n7483) );
  XNOR2HSV4 U9575 ( .A1(n9742), .A2(n9741), .ZN(n9745) );
  CLKNAND2HSV0 U9576 ( .A1(n7486), .A2(n7485), .ZN(n14293) );
  INAND2HSV2 U9577 ( .A1(n11220), .B1(\pe16/ti_7t [5]), .ZN(n7485) );
  CLKNAND2HSV3 U9578 ( .A1(n15228), .A2(n11220), .ZN(n7486) );
  MUX2NHSV4 U9579 ( .I0(n8503), .I1(n11174), .S(n7487), .ZN(n15228) );
  CLKNAND2HSV4 U9580 ( .A1(n14827), .A2(n11179), .ZN(n7487) );
  CLKNAND2HSV4 U9581 ( .A1(n11158), .A2(n11157), .ZN(n14827) );
  XOR3HSV2 U9582 ( .A1(n13531), .A2(n7489), .A3(n7488), .Z(n8477) );
  CLKNAND2HSV2 U9583 ( .A1(n14191), .A2(\pe8/got [3]), .ZN(n7488) );
  XOR2HSV2 U9584 ( .A1(n8476), .A2(n13529), .Z(n7489) );
  OAI21HSV4 U9585 ( .A1(n7493), .A2(n7492), .B(n10747), .ZN(n7491) );
  CLKNHSV2 U9586 ( .I(n7495), .ZN(n7492) );
  CLKNHSV2 U9587 ( .I(n7509), .ZN(n7495) );
  XOR2HSV0 U9588 ( .A1(n7496), .A2(n14172), .Z(\pe20/poht [7]) );
  OAI21HSV4 U9589 ( .A1(n6737), .A2(n9790), .B(n8429), .ZN(n7497) );
  NOR2HSV4 U9590 ( .A1(n11902), .A2(n11898), .ZN(n12348) );
  CLKNHSV2 U9591 ( .I(n11895), .ZN(n7501) );
  XNOR2HSV4 U9592 ( .A1(n12348), .A2(n12347), .ZN(n15256) );
  XOR3HSV2 U9593 ( .A1(n7920), .A2(n7929), .A3(n7930), .Z(n7503) );
  CLKNHSV2 U9594 ( .I(n13344), .ZN(n13805) );
  NOR2HSV4 U9595 ( .A1(n14650), .A2(n13147), .ZN(n13175) );
  CLKNAND2HSV2 U9596 ( .A1(n7504), .A2(n7933), .ZN(n13807) );
  CLKNAND2HSV2 U9597 ( .A1(n7505), .A2(n13344), .ZN(n7504) );
  NOR2HSV4 U9598 ( .A1(n13804), .A2(n7932), .ZN(n7505) );
  NOR2HSV4 U9599 ( .A1(n9284), .A2(n6726), .ZN(n7798) );
  CLKNAND2HSV2 U9600 ( .A1(n9284), .A2(n6726), .ZN(n7797) );
  CLKNHSV2 U9601 ( .I(n7576), .ZN(n7506) );
  CLKNHSV2 U9602 ( .I(n11446), .ZN(n7509) );
  INAND2HSV4 U9603 ( .A1(n7517), .B1(n7516), .ZN(n11177) );
  CLKNHSV2 U9604 ( .I(n7511), .ZN(n7510) );
  NAND3HSV3 U9605 ( .A1(n11171), .A2(n13191), .A3(\pe16/got [6]), .ZN(n7512)
         );
  CLKNAND2HSV3 U9606 ( .A1(n7577), .A2(n7518), .ZN(n7513) );
  CLKNHSV1 U9607 ( .I(n6709), .ZN(n7514) );
  CLKNAND2HSV3 U9608 ( .A1(n8906), .A2(n14827), .ZN(n7516) );
  INHSV2 U9609 ( .I(n11171), .ZN(n7518) );
  BUFHSV8 U9610 ( .I(n7738), .Z(n7519) );
  CLKNHSV2 U9611 ( .I(n7520), .ZN(n7788) );
  CLKNAND2HSV2 U9612 ( .A1(n7738), .A2(n10869), .ZN(n7520) );
  CLKNAND2HSV2 U9613 ( .A1(n7519), .A2(n13797), .ZN(n8472) );
  CLKNAND2HSV2 U9614 ( .A1(n7519), .A2(\pe21/got [5]), .ZN(n10885) );
  CLKNAND2HSV2 U9615 ( .A1(n7519), .A2(n13107), .ZN(n13137) );
  OAI22HSV4 U9616 ( .A1(n11705), .A2(n10865), .B1(n7778), .B2(n7777), .ZN(
        n7738) );
  CLKBUFHSV2 U9617 ( .I(n13105), .Z(n7521) );
  CLKNHSV2 U9618 ( .I(n13105), .ZN(n9308) );
  XOR2HSV2 U9619 ( .A1(n9263), .A2(n9262), .Z(n13105) );
  CLKNHSV2 U9620 ( .I(n10707), .ZN(n7522) );
  CLKNAND2HSV2 U9621 ( .A1(\pe14/ti_7[3] ), .A2(\pe14/got [5]), .ZN(n8084) );
  CLKNAND2HSV2 U9622 ( .A1(n5969), .A2(\pe14/got [1]), .ZN(n8763) );
  CLKNAND2HSV2 U9623 ( .A1(n5969), .A2(\pe14/got [4]), .ZN(n13080) );
  CLKNAND2HSV2 U9624 ( .A1(n5969), .A2(\pe14/got [3]), .ZN(n13574) );
  XOR2HSV2 U9625 ( .A1(n7524), .A2(n8409), .Z(n8410) );
  CLKNAND2HSV2 U9626 ( .A1(n5969), .A2(\pe14/got [2]), .ZN(n7524) );
  AOI21HSV4 U9627 ( .A1(n12630), .A2(n7527), .B(n7525), .ZN(\pe14/ti_7[3] ) );
  CLKNHSV2 U9628 ( .I(n7526), .ZN(n7525) );
  CLKNAND2HSV2 U9629 ( .A1(n11090), .A2(n11039), .ZN(n7526) );
  CLKNHSV2 U9630 ( .I(n11090), .ZN(n7527) );
  CLKBUFHSV2 U9631 ( .I(n14958), .Z(n7528) );
  CLKNAND2HSV2 U9632 ( .A1(n7528), .A2(\pe16/got [3]), .ZN(n14265) );
  CLKBUFHSV2 U9633 ( .I(n12111), .Z(n7529) );
  XNOR2HSV4 U9634 ( .A1(n7534), .A2(n7530), .ZN(n10868) );
  XOR3HSV2 U9635 ( .A1(n7648), .A2(n7533), .A3(n7532), .Z(n7531) );
  XNOR2HSV4 U9636 ( .A1(n7649), .A2(n7651), .ZN(n7533) );
  CLKNAND2HSV2 U9637 ( .A1(n8207), .A2(n7535), .ZN(n7534) );
  CLKNAND2HSV2 U9638 ( .A1(n7140), .A2(n7536), .ZN(n7535) );
  CLKNHSV2 U9639 ( .I(n10402), .ZN(n7537) );
  CLKNAND2HSV2 U9640 ( .A1(n7540), .A2(n7805), .ZN(n7538) );
  CLKNHSV2 U9641 ( .I(n8304), .ZN(n7539) );
  CLKNHSV2 U9642 ( .I(n7541), .ZN(n7540) );
  XNOR2HSV4 U9643 ( .A1(n9214), .A2(n7542), .ZN(n9216) );
  CLKNAND2HSV2 U9644 ( .A1(n7543), .A2(n9139), .ZN(\pe18/ti_7[1] ) );
  CLKNAND2HSV2 U9645 ( .A1(n14826), .A2(n9217), .ZN(n7543) );
  XNOR2HSV4 U9646 ( .A1(n9138), .A2(n9137), .ZN(n14826) );
  AOI21HSV4 U9647 ( .A1(n7681), .A2(n10681), .B(n7545), .ZN(n7544) );
  NOR2HSV3 U9648 ( .A1(n10678), .A2(n13229), .ZN(n7545) );
  MUX2NHSV2 U9649 ( .I0(n8001), .I1(n9298), .S(n7546), .ZN(n9300) );
  XNOR2HSV4 U9650 ( .A1(n7549), .A2(n7548), .ZN(n7547) );
  CLKNAND2HSV2 U9651 ( .A1(n13824), .A2(\pe6/got [3]), .ZN(n7548) );
  XNOR2HSV4 U9652 ( .A1(n7863), .A2(\pe6/phq [6]), .ZN(n7549) );
  CLKNAND2HSV2 U9653 ( .A1(\pe8/ti_7[1] ), .A2(\pe8/got [5]), .ZN(n11508) );
  CLKNAND2HSV2 U9654 ( .A1(n11521), .A2(\pe8/ti_7t [1]), .ZN(n7550) );
  CLKNAND2HSV2 U9655 ( .A1(n11796), .A2(n12316), .ZN(n7551) );
  XNOR2HSV4 U9656 ( .A1(n7553), .A2(n7552), .ZN(n11796) );
  AOI21HSV4 U9657 ( .A1(n10486), .A2(n11574), .B(n10485), .ZN(n7552) );
  XNOR2HSV4 U9658 ( .A1(n10484), .A2(n10483), .ZN(n7553) );
  CLKNAND2HSV0 U9659 ( .A1(n8194), .A2(n8193), .ZN(n8195) );
  OAI21HSV2 U9660 ( .A1(n7558), .A2(n7555), .B(n7554), .ZN(n8193) );
  INHSV2 U9661 ( .I(n8192), .ZN(n7556) );
  NOR2HSV8 U9662 ( .A1(n13751), .A2(n13750), .ZN(n7558) );
  INAND2HSV2 U9663 ( .A1(n7559), .B1(n13752), .ZN(n8194) );
  CLKNAND2HSV3 U9664 ( .A1(n13681), .A2(n13682), .ZN(n13752) );
  INHSV2 U9665 ( .I(n14865), .ZN(n7559) );
  NOR2HSV4 U9666 ( .A1(n7561), .A2(n14248), .ZN(n7560) );
  CLKNAND2HSV2 U9667 ( .A1(n8026), .A2(n7562), .ZN(n7561) );
  CLKNAND2HSV2 U9668 ( .A1(n7564), .A2(n7563), .ZN(n7562) );
  CLKNHSV2 U9669 ( .I(n8023), .ZN(n7563) );
  CLKNHSV2 U9670 ( .I(n7566), .ZN(n7565) );
  CLKNHSV4 U9671 ( .I(n9881), .ZN(n7566) );
  NOR2HSV4 U9672 ( .A1(n7570), .A2(n7569), .ZN(n7568) );
  CLKNHSV2 U9673 ( .I(n11440), .ZN(n7569) );
  CLKNHSV2 U9674 ( .I(n11435), .ZN(n7570) );
  OAI21HSV4 U9675 ( .A1(n11439), .A2(n7573), .B(n7572), .ZN(n7571) );
  XOR3HSV2 U9676 ( .A1(n7575), .A2(n12722), .A3(n7574), .Z(\pe12/poht [4]) );
  CLKNAND2HSV2 U9677 ( .A1(n14959), .A2(\pe12/got [4]), .ZN(n7574) );
  CLKNAND2HSV2 U9678 ( .A1(n15190), .A2(\pe12/got [3]), .ZN(n7575) );
  CLKNHSV2 U9679 ( .I(n11609), .ZN(n7576) );
  CLKNAND2HSV3 U9680 ( .A1(n13191), .A2(\pe16/got [6]), .ZN(n7577) );
  CLKNAND2HSV3 U9681 ( .A1(n11158), .A2(n11157), .ZN(n13191) );
  CLKNHSV2 U9682 ( .I(n10357), .ZN(n7579) );
  CLKNHSV2 U9683 ( .I(\pe19/ti_7t [5]), .ZN(n7580) );
  NAND3HSV4 U9684 ( .A1(n12141), .A2(n9541), .A3(n11712), .ZN(n7581) );
  NAND2HSV2 U9685 ( .A1(\pe13/bq[8] ), .A2(\pe13/aot [6]), .ZN(n7582) );
  CLKXOR2HSV4 U9686 ( .A1(n9862), .A2(n7582), .Z(n7586) );
  CLKBUFHSV2 U9687 ( .I(\pe13/bq[8] ), .Z(n7583) );
  XNOR2HSV4 U9688 ( .A1(n7586), .A2(n7584), .ZN(n9865) );
  XOR2HSV2 U9689 ( .A1(n7585), .A2(\pe13/phq [3]), .Z(n7584) );
  XOR2HSV0 U9690 ( .A1(n7592), .A2(n7587), .Z(\pe13/poht [2]) );
  XOR2HSV2 U9691 ( .A1(n7589), .A2(n7588), .Z(n7587) );
  XNOR2HSV4 U9692 ( .A1(n7591), .A2(n7590), .ZN(n7589) );
  XOR3HSV2 U9693 ( .A1(n9928), .A2(n7737), .A3(n8475), .Z(n7591) );
  CLKNAND2HSV2 U9694 ( .A1(n13604), .A2(\pe13/got [6]), .ZN(n7592) );
  CLKNAND2HSV2 U9695 ( .A1(n8237), .A2(n8238), .ZN(n8239) );
  CLKNAND2HSV2 U9696 ( .A1(n7594), .A2(n8236), .ZN(n7593) );
  CLKNAND2HSV2 U9697 ( .A1(n7596), .A2(n13603), .ZN(n7595) );
  NOR2HSV4 U9698 ( .A1(n8236), .A2(n8231), .ZN(n7596) );
  CLKNHSV2 U9699 ( .I(\pe13/got [4]), .ZN(n7598) );
  INAND2HSV4 U9700 ( .A1(n9952), .B1(n7599), .ZN(n15243) );
  XNOR2HSV4 U9701 ( .A1(n7601), .A2(n7600), .ZN(n9947) );
  NAND2HSV2 U9702 ( .A1(n9920), .A2(\pe13/got [7]), .ZN(n7600) );
  XNOR2HSV4 U9703 ( .A1(n9902), .A2(n9901), .ZN(n7601) );
  OAI21HSV4 U9704 ( .A1(n7603), .A2(n7602), .B(n9883), .ZN(n9946) );
  CLKNAND2HSV2 U9705 ( .A1(n9885), .A2(n9881), .ZN(n7603) );
  CLKNHSV2 U9706 ( .I(n9887), .ZN(n7604) );
  AOI21HSV4 U9707 ( .A1(n15292), .A2(n7607), .B(n7605), .ZN(n13102) );
  CLKNHSV2 U9708 ( .I(n7606), .ZN(n7605) );
  CLKNAND2HSV2 U9709 ( .A1(n9358), .A2(\pe2/ti_7t [5]), .ZN(n7606) );
  CLKNHSV2 U9710 ( .I(n9358), .ZN(n7607) );
  CLKNAND2HSV0 U9711 ( .A1(n8332), .A2(n8331), .ZN(n8333) );
  NAND2HSV2 U9712 ( .A1(n8330), .A2(n7610), .ZN(n7609) );
  CLKNAND2HSV1 U9713 ( .A1(n7612), .A2(n7611), .ZN(n7610) );
  CLKNHSV1 U9714 ( .I(n8329), .ZN(n7611) );
  CLKNAND2HSV3 U9715 ( .A1(n14179), .A2(\pe6/got [8]), .ZN(n8332) );
  CLKNAND2HSV2 U9716 ( .A1(n8270), .A2(n8271), .ZN(n8272) );
  CLKNAND2HSV2 U9717 ( .A1(n13752), .A2(\pe20/got [5]), .ZN(n8271) );
  CLKNHSV2 U9718 ( .I(n8269), .ZN(n7613) );
  CLKNAND2HSV2 U9719 ( .A1(\pe20/ti_7[5] ), .A2(\pe20/got [3]), .ZN(n7614) );
  XNOR2HSV4 U9720 ( .A1(n7617), .A2(n7615), .ZN(n15201) );
  AOI21HSV4 U9721 ( .A1(n15261), .A2(n10148), .B(n7616), .ZN(n7615) );
  NOR2HSV4 U9722 ( .A1(n7862), .A2(n7861), .ZN(n7616) );
  XNOR2HSV4 U9723 ( .A1(n8610), .A2(n7618), .ZN(n7617) );
  NOR2HSV4 U9724 ( .A1(n14129), .A2(n7714), .ZN(n7618) );
  AOI21HSV4 U9725 ( .A1(n15273), .A2(n10459), .B(n12311), .ZN(n8010) );
  CLKNAND2HSV2 U9726 ( .A1(\pe7/bq[8] ), .A2(\pe7/aot [8]), .ZN(n7621) );
  CLKNAND2HSV2 U9727 ( .A1(n7622), .A2(n9903), .ZN(n7624) );
  CLKNHSV2 U9728 ( .I(n9951), .ZN(n7623) );
  OAI21HSV4 U9729 ( .A1(n11475), .A2(n7625), .B(n11474), .ZN(n7894) );
  CLKNAND2HSV2 U9730 ( .A1(n15278), .A2(n11473), .ZN(n7625) );
  XNOR2HSV4 U9731 ( .A1(n7626), .A2(n10331), .ZN(n15278) );
  CLKNHSV2 U9732 ( .I(n11206), .ZN(n7627) );
  CLKNHSV2 U9733 ( .I(n11220), .ZN(n7628) );
  CLKNHSV2 U9734 ( .I(n8680), .ZN(n7629) );
  CLKNHSV2 U9735 ( .I(n7873), .ZN(n7630) );
  XNOR2HSV4 U9736 ( .A1(n7730), .A2(n7728), .ZN(n11705) );
  CLKNAND2HSV2 U9737 ( .A1(\pe6/ti_7[5] ), .A2(\pe6/got [1]), .ZN(n12987) );
  CLKNAND2HSV2 U9738 ( .A1(n15198), .A2(n9536), .ZN(n7632) );
  MUX2NHSV2 U9739 ( .I0(n8035), .I1(n9535), .S(n8039), .ZN(n15198) );
  MUX2NHSV2 U9740 ( .I0(n7638), .I1(n7637), .S(n7634), .ZN(n7633) );
  XNOR2HSV4 U9741 ( .A1(n7636), .A2(n7635), .ZN(n7634) );
  CLKNAND2HSV2 U9742 ( .A1(n15084), .A2(\pe19/got [5]), .ZN(n7635) );
  CLKNHSV2 U9743 ( .I(n8434), .ZN(n7636) );
  CLKNHSV2 U9744 ( .I(n7639), .ZN(n7638) );
  CLKNAND2HSV2 U9745 ( .A1(n14862), .A2(n14841), .ZN(n7640) );
  OAI21HSV4 U9746 ( .A1(n7643), .A2(n7644), .B(n11210), .ZN(n7642) );
  CLKNHSV2 U9747 ( .I(n11209), .ZN(n7643) );
  NOR2HSV4 U9748 ( .A1(n7646), .A2(n7645), .ZN(n14067) );
  CLKNHSV2 U9749 ( .I(n14066), .ZN(n7645) );
  CLKNHSV2 U9750 ( .I(n14065), .ZN(n7646) );
  CLKNHSV2 U9751 ( .I(n11181), .ZN(n7647) );
  XNOR2HSV1 U9752 ( .A1(n7977), .A2(n7976), .ZN(n7648) );
  NOR2HSV2 U9753 ( .A1(n10826), .A2(n7650), .ZN(n7649) );
  CLKNHSV4 U9754 ( .I(\pe21/got [4]), .ZN(n7650) );
  CLKXOR2HSV2 U9755 ( .A1(n7975), .A2(n10844), .Z(n7651) );
  OAI21HSV1 U9756 ( .A1(n15201), .A2(n7655), .B(n7652), .ZN(n14157) );
  AOI21HSV2 U9757 ( .A1(n10590), .A2(n7654), .B(n7653), .ZN(n7652) );
  INHSV2 U9758 ( .I(n10599), .ZN(n7654) );
  CLKNHSV3 U9759 ( .I(n10590), .ZN(n7655) );
  CLKNAND2HSV2 U9760 ( .A1(n10591), .A2(n10590), .ZN(n15187) );
  CLKNAND2HSV2 U9761 ( .A1(\pe21/got [6]), .A2(\pe21/ti_1 ), .ZN(n7656) );
  CLKNHSV2 U9762 ( .I(n14007), .ZN(n7659) );
  CLKNHSV2 U9763 ( .I(n10126), .ZN(n7660) );
  XNOR2HSV4 U9764 ( .A1(n7666), .A2(n7662), .ZN(n10399) );
  XNOR2HSV4 U9765 ( .A1(n7664), .A2(n7663), .ZN(n7662) );
  CLKNAND2HSV2 U9766 ( .A1(n11786), .A2(\pe21/pvq [4]), .ZN(n7663) );
  XOR2HSV2 U9767 ( .A1(n7665), .A2(\pe21/phq [4]), .Z(n7664) );
  CLKNAND2HSV2 U9768 ( .A1(\pe21/aot [8]), .A2(\pe21/bq[5] ), .ZN(n7665) );
  XNOR2HSV4 U9769 ( .A1(n7670), .A2(n7667), .ZN(n7666) );
  XNOR2HSV4 U9770 ( .A1(n7669), .A2(n7668), .ZN(n7667) );
  CLKNAND2HSV2 U9771 ( .A1(\pe21/aot [7]), .A2(\pe21/bq[6] ), .ZN(n7668) );
  CLKNAND2HSV2 U9772 ( .A1(\pe21/ti_1 ), .A2(\pe21/got [5]), .ZN(n7669) );
  XNOR2HSV4 U9773 ( .A1(n10395), .A2(n7671), .ZN(n7670) );
  NOR2HSV4 U9774 ( .A1(n7677), .A2(n7676), .ZN(n7675) );
  NOR2HSV4 U9775 ( .A1(n11771), .A2(n11772), .ZN(n7676) );
  CLKNHSV2 U9776 ( .I(n11413), .ZN(n7680) );
  INHSV2 U9777 ( .I(n7705), .ZN(n7682) );
  CLKBUFHSV2 U9778 ( .I(n7685), .Z(n7683) );
  CLKBUFHSV2 U9779 ( .I(n11767), .Z(n7684) );
  NAND3HSV4 U9780 ( .A1(n7683), .A2(n11765), .A3(n7684), .ZN(n11770) );
  CLKNAND2HSV2 U9781 ( .A1(n9858), .A2(\pe6/got [6]), .ZN(n9836) );
  OAI21HSV4 U9782 ( .A1(n9833), .A2(n13103), .B(n7686), .ZN(n9858) );
  CLKNHSV2 U9783 ( .I(\pe6/ti_7t [4]), .ZN(n7687) );
  CLKNHSV2 U9784 ( .I(n15088), .ZN(n7688) );
  CLKNHSV2 U9785 ( .I(n9840), .ZN(n7689) );
  CLKNAND2HSV0 U9786 ( .A1(n7994), .A2(n7993), .ZN(n7995) );
  XNOR2HSV2 U9787 ( .A1(n7992), .A2(n7690), .ZN(n7993) );
  CLKNAND2HSV3 U9788 ( .A1(n6922), .A2(\pe5/got [5]), .ZN(n7690) );
  CLKNAND2HSV3 U9789 ( .A1(n13285), .A2(n13284), .ZN(n13406) );
  CLKNHSV2 U9790 ( .I(n10469), .ZN(n7691) );
  OAI21HSV4 U9791 ( .A1(n7696), .A2(n7693), .B(n7692), .ZN(n8656) );
  XNOR2HSV4 U9792 ( .A1(n7695), .A2(n7694), .ZN(n7693) );
  CLKNHSV2 U9793 ( .I(n8655), .ZN(n7694) );
  NOR2HSV4 U9794 ( .A1(n14585), .A2(n8649), .ZN(n7696) );
  CLKNHSV2 U9795 ( .I(\pe15/ti_7t [7]), .ZN(n7697) );
  CLKNHSV2 U9796 ( .I(n12829), .ZN(n7698) );
  INAND2HSV4 U9797 ( .A1(n8776), .B1(n7701), .ZN(n7700) );
  CLKNHSV2 U9798 ( .I(n7702), .ZN(n7701) );
  XNOR2HSV4 U9799 ( .A1(n7704), .A2(n7703), .ZN(n7702) );
  XNOR2HSV4 U9800 ( .A1(n8777), .A2(n13473), .ZN(n7703) );
  CLKNHSV2 U9801 ( .I(n14873), .ZN(n7705) );
  CLKNAND2HSV2 U9802 ( .A1(n15176), .A2(n11120), .ZN(n9084) );
  INAND2HSV4 U9803 ( .A1(n13257), .B1(n7706), .ZN(n10639) );
  CLKNHSV2 U9804 ( .I(n7707), .ZN(n7706) );
  CLKNAND2HSV2 U9805 ( .A1(n10637), .A2(n7708), .ZN(n7707) );
  CLKNHSV2 U9806 ( .I(n10632), .ZN(n7708) );
  NOR2HSV4 U9807 ( .A1(n8028), .A2(n7712), .ZN(n7711) );
  AOI21HSV4 U9808 ( .A1(n10634), .A2(n10633), .B(n14868), .ZN(n7713) );
  NAND3HSV4 U9809 ( .A1(n10604), .A2(n8395), .A3(n8396), .ZN(n13257) );
  OAI211HSV2 U9810 ( .A1(n7718), .A2(n7717), .B(n8007), .C(n7716), .ZN(n7715)
         );
  CLKNAND2HSV2 U9811 ( .A1(n8005), .A2(n10995), .ZN(n7717) );
  XNOR2HSV4 U9812 ( .A1(n8006), .A2(n7720), .ZN(n7719) );
  XNOR2HSV4 U9813 ( .A1(n10660), .A2(n10661), .ZN(n10839) );
  CLKNHSV2 U9814 ( .I(n7725), .ZN(n7722) );
  CLKNAND2HSV2 U9815 ( .A1(n7727), .A2(n7726), .ZN(n7725) );
  CLKNHSV2 U9816 ( .I(n10835), .ZN(n7726) );
  CLKNHSV2 U9817 ( .I(n10402), .ZN(n7727) );
  CLKNHSV2 U9818 ( .I(n10402), .ZN(n7729) );
  XNOR2HSV4 U9819 ( .A1(n7732), .A2(n7731), .ZN(n7730) );
  CLKNHSV2 U9820 ( .I(n13107), .ZN(n7733) );
  CLKNAND2HSV2 U9821 ( .A1(n7734), .A2(\pe10/got [4]), .ZN(n10079) );
  CLKNHSV2 U9822 ( .I(n15139), .ZN(n7734) );
  CLKNAND2HSV2 U9823 ( .A1(n10202), .A2(n10203), .ZN(n7735) );
  NOR2HSV4 U9824 ( .A1(n10203), .A2(n10202), .ZN(n7736) );
  AOI21HSV4 U9825 ( .A1(n7786), .A2(n6736), .B(n7784), .ZN(n7742) );
  CLKNAND2HSV2 U9826 ( .A1(n7519), .A2(\pe21/got [1]), .ZN(n7739) );
  CLKNAND2HSV3 U9827 ( .A1(n15085), .A2(\pe21/got [2]), .ZN(n7740) );
  CLKNAND2HSV3 U9828 ( .A1(n7788), .A2(n13338), .ZN(n7741) );
  CLKNHSV2 U9829 ( .I(n7744), .ZN(n7743) );
  CLKNAND2HSV2 U9830 ( .A1(n9358), .A2(\pe2/ti_7t [7]), .ZN(n7744) );
  CLKNAND2HSV2 U9831 ( .A1(n8310), .A2(n7746), .ZN(n7745) );
  CLKNHSV2 U9832 ( .I(n9358), .ZN(n7746) );
  XNOR2HSV4 U9833 ( .A1(n11260), .A2(n11259), .ZN(n7748) );
  OAI21HSV4 U9834 ( .A1(n7752), .A2(n7751), .B(n7750), .ZN(n8033) );
  CLKNAND2HSV2 U9835 ( .A1(n7751), .A2(n7752), .ZN(n7750) );
  CLKNAND2HSV2 U9836 ( .A1(n7754), .A2(n7753), .ZN(n7752) );
  CLKNHSV2 U9837 ( .I(n8031), .ZN(n7753) );
  CLKNHSV2 U9838 ( .I(n8030), .ZN(n7754) );
  MUX2NHSV2 U9839 ( .I0(n8375), .I1(n9248), .S(n7757), .ZN(n7756) );
  NOR2HSV4 U9840 ( .A1(n9244), .A2(n9232), .ZN(n9248) );
  XNOR2HSV4 U9841 ( .A1(n9229), .A2(n9228), .ZN(n7757) );
  XNOR2HSV2 U9842 ( .A1(n7761), .A2(n7759), .ZN(n7758) );
  CLKNAND2HSV3 U9843 ( .A1(\pe6/ti_7[5] ), .A2(\pe6/got [5]), .ZN(n7760) );
  INHSV2 U9844 ( .I(n12410), .ZN(n7762) );
  CLKNAND2HSV3 U9845 ( .A1(n14179), .A2(n5977), .ZN(n7763) );
  INHSV2 U9846 ( .I(n7818), .ZN(n7764) );
  CLKNAND2HSV2 U9847 ( .A1(n8534), .A2(n8533), .ZN(n8535) );
  XNOR2HSV4 U9848 ( .A1(n7766), .A2(n7765), .ZN(n8533) );
  XNOR2HSV4 U9849 ( .A1(n8532), .A2(n13391), .ZN(n7765) );
  CLKNAND2HSV2 U9850 ( .A1(n14916), .A2(\pe5/got [1]), .ZN(n7766) );
  XNOR2HSV4 U9851 ( .A1(n7769), .A2(n7767), .ZN(n8409) );
  XOR2HSV2 U9852 ( .A1(n11155), .A2(n7768), .Z(n7767) );
  CLKNHSV2 U9853 ( .I(n11154), .ZN(n7768) );
  CLKNAND2HSV2 U9854 ( .A1(n14944), .A2(\pe14/got [1]), .ZN(n7769) );
  CLKNAND2HSV2 U9855 ( .A1(n11597), .A2(n11591), .ZN(n7770) );
  CLKNHSV2 U9856 ( .I(n11604), .ZN(n7771) );
  CLKNHSV2 U9857 ( .I(n11587), .ZN(n7774) );
  CLKNHSV2 U9858 ( .I(n11588), .ZN(n7775) );
  CLKNHSV2 U9859 ( .I(\pe21/ti_7t [6]), .ZN(n7778) );
  CLKNAND2HSV2 U9860 ( .A1(n7781), .A2(n7780), .ZN(n7779) );
  CLKNHSV2 U9861 ( .I(n10860), .ZN(n7780) );
  CLKNHSV2 U9862 ( .I(n10861), .ZN(n7781) );
  CLKNAND2HSV2 U9863 ( .A1(\pe16/aot [5]), .A2(\pe16/bq[8] ), .ZN(n7782) );
  CLKNAND2HSV2 U9864 ( .A1(\pe16/bq[6] ), .A2(\pe16/aot [7]), .ZN(n7783) );
  CLKNHSV2 U9865 ( .I(n7787), .ZN(n7785) );
  CLKNHSV2 U9866 ( .I(n10866), .ZN(n7787) );
  CLKNHSV2 U9867 ( .I(n14007), .ZN(n7789) );
  CLKNHSV2 U9868 ( .I(n14010), .ZN(n7790) );
  XNOR2HSV4 U9869 ( .A1(n7791), .A2(n10721), .ZN(n12108) );
  CLKNHSV2 U9870 ( .I(n10720), .ZN(n7791) );
  XNOR2HSV4 U9871 ( .A1(n10721), .A2(n10720), .ZN(n12102) );
  CLKNHSV2 U9872 ( .I(n7794), .ZN(n7793) );
  CLKNAND2HSV2 U9873 ( .A1(n11739), .A2(n11944), .ZN(n7794) );
  AOI21HSV4 U9874 ( .A1(n11740), .A2(n11739), .B(n11741), .ZN(n11738) );
  CLKNAND2HSV1 U9875 ( .A1(n6754), .A2(n10118), .ZN(n7795) );
  INHSV2 U9876 ( .I(n7798), .ZN(n7796) );
  NAND3HSV4 U9877 ( .A1(n7797), .A2(n7796), .A3(n7799), .ZN(n8036) );
  CLKNHSV2 U9878 ( .I(n7800), .ZN(n7799) );
  CLKNAND2HSV2 U9879 ( .A1(n7801), .A2(n9832), .ZN(n7800) );
  CLKBUFHSV2 U9880 ( .I(n5977), .Z(n7801) );
  CLKNAND2HSV3 U9881 ( .A1(n15187), .A2(\pe10/got [4]), .ZN(n7802) );
  CLKNHSV2 U9882 ( .I(n7804), .ZN(n7803) );
  CLKNAND2HSV2 U9883 ( .A1(n11006), .A2(n15180), .ZN(n7804) );
  CLKNHSV2 U9884 ( .I(n10408), .ZN(n7806) );
  NOR2HSV4 U9885 ( .A1(n10948), .A2(n10204), .ZN(n7808) );
  XOR2HSV2 U9886 ( .A1(n7809), .A2(n8779), .Z(n7811) );
  XOR2HSV2 U9887 ( .A1(n7810), .A2(n8778), .Z(n7809) );
  CLKNAND2HSV3 U9888 ( .A1(n15187), .A2(\pe10/got [5]), .ZN(n7812) );
  CLKNHSV2 U9889 ( .I(n8376), .ZN(n7815) );
  CLKNHSV2 U9890 ( .I(n9844), .ZN(n7816) );
  INAND2HSV4 U9891 ( .A1(n9842), .B1(n9846), .ZN(n7817) );
  CLKNHSV2 U9892 ( .I(n9846), .ZN(n7818) );
  XNOR2HSV4 U9893 ( .A1(n9839), .A2(n9838), .ZN(n13898) );
  CLKNHSV2 U9894 ( .I(n12411), .ZN(n15089) );
  CLKNAND2HSV2 U9895 ( .A1(n14179), .A2(\pe6/got [4]), .ZN(n13010) );
  XNOR2HSV4 U9896 ( .A1(n11167), .A2(n11163), .ZN(n7819) );
  XNOR2HSV4 U9897 ( .A1(n7883), .A2(n7821), .ZN(n7820) );
  XOR2HSV2 U9898 ( .A1(n11168), .A2(n11162), .Z(n7821) );
  CLKNHSV2 U9899 ( .I(n10930), .ZN(n7823) );
  CLKNAND2HSV2 U9900 ( .A1(n15261), .A2(n10599), .ZN(n7824) );
  CLKNAND2HSV2 U9901 ( .A1(n8335), .A2(n10787), .ZN(n7826) );
  XOR3HSV2 U9902 ( .A1(n8072), .A2(n7832), .A3(n7830), .Z(n8074) );
  MUX2NHSV2 U9903 ( .I0(n8070), .I1(n12667), .S(n7831), .ZN(n7830) );
  XNOR2HSV4 U9904 ( .A1(n8071), .A2(n11458), .ZN(n7831) );
  CLKNHSV2 U9905 ( .I(n8073), .ZN(n7832) );
  CLKNHSV2 U9906 ( .I(n7834), .ZN(n7833) );
  CLKNAND2HSV2 U9907 ( .A1(n9200), .A2(n8041), .ZN(n7834) );
  CLKNAND2HSV2 U9908 ( .A1(n8616), .A2(n7837), .ZN(n7836) );
  CLKNAND2HSV2 U9909 ( .A1(n7839), .A2(n7838), .ZN(n7837) );
  CLKNHSV2 U9910 ( .I(n8615), .ZN(n7838) );
  CLKNHSV2 U9911 ( .I(n8614), .ZN(n7839) );
  CLKNHSV2 U9912 ( .I(n10510), .ZN(n7841) );
  INHSV2 U9913 ( .I(n7843), .ZN(n7842) );
  NAND2HSV2 U9914 ( .A1(n7847), .A2(n7983), .ZN(n7843) );
  CLKAND2HSV4 U9915 ( .A1(n10677), .A2(n10796), .Z(n7844) );
  CLKNHSV2 U9916 ( .I(n10678), .ZN(n7846) );
  CLKNAND2HSV2 U9917 ( .A1(n10524), .A2(n14064), .ZN(n10680) );
  XNOR2HSV4 U9918 ( .A1(n10672), .A2(n10671), .ZN(n10524) );
  CLKNHSV2 U9919 ( .I(n7982), .ZN(n7847) );
  CLKNAND2HSV4 U9920 ( .A1(n10704), .A2(n7845), .ZN(n7850) );
  CLKNAND2HSV2 U9921 ( .A1(n7850), .A2(n12194), .ZN(n10795) );
  CLKNHSV2 U9922 ( .I(n12194), .ZN(n7849) );
  AOI21HSV4 U9923 ( .A1(n8085), .A2(n11117), .B(n7853), .ZN(n7852) );
  XNOR2HSV4 U9924 ( .A1(n7856), .A2(n7855), .ZN(n7854) );
  XNOR2HSV4 U9925 ( .A1(n8083), .A2(n8084), .ZN(n7856) );
  CLKNHSV2 U9926 ( .I(n9989), .ZN(n13259) );
  CLKNHSV2 U9927 ( .I(n8308), .ZN(n7857) );
  NOR2HSV4 U9928 ( .A1(n7529), .A2(n12110), .ZN(n7858) );
  XNOR2HSV4 U9929 ( .A1(n7860), .A2(n12129), .ZN(n8213) );
  XOR2HSV2 U9930 ( .A1(n12127), .A2(n12128), .Z(n7860) );
  INHSV2 U9931 ( .I(\pe10/got [8]), .ZN(n7861) );
  INHSV24 U9932 ( .I(n10930), .ZN(n7862) );
  NOR2HSV4 U9933 ( .A1(n9996), .A2(n9956), .ZN(n7864) );
  XNOR2HSV4 U9934 ( .A1(n7905), .A2(n7865), .ZN(n7906) );
  CLKNAND2HSV2 U9935 ( .A1(n7867), .A2(n7866), .ZN(n7865) );
  NOR2HSV4 U9936 ( .A1(n11095), .A2(n13059), .ZN(n7866) );
  CLKNAND2HSV2 U9937 ( .A1(n12630), .A2(n11156), .ZN(n7867) );
  XNOR2HSV4 U9938 ( .A1(n11062), .A2(n11064), .ZN(n12630) );
  CLKNHSV2 U9939 ( .I(n7869), .ZN(n7868) );
  CLKNAND2HSV2 U9940 ( .A1(n8109), .A2(n14931), .ZN(n7869) );
  NAND2HSV0 U9941 ( .A1(n6706), .A2(\pe4/got [5]), .ZN(n8873) );
  CLKNHSV2 U9942 ( .I(n8680), .ZN(n7873) );
  NAND2HSV0 U9943 ( .A1(\pe10/ti_7[6] ), .A2(n5966), .ZN(n14154) );
  NAND2HSV0 U9944 ( .A1(\pe10/ti_7[5] ), .A2(n5966), .ZN(n10927) );
  INOR2HSV2 U9945 ( .A1(n5966), .B1(n10125), .ZN(n10108) );
  CLKNAND2HSV4 U9946 ( .A1(n10999), .A2(n10998), .ZN(n12957) );
  INHSV4 U9947 ( .I(n9982), .ZN(n9979) );
  XNOR2HSV4 U9948 ( .A1(n12499), .A2(n12498), .ZN(n12505) );
  CLKNAND2HSV2 U9949 ( .A1(n10704), .A2(n7845), .ZN(n13219) );
  XOR2HSV0 U9950 ( .A1(n7876), .A2(n12088), .Z(\pe4/poht [5]) );
  XNOR2HSV4 U9951 ( .A1(n11164), .A2(\pe16/phq [7]), .ZN(n7877) );
  XOR2HSV0 U9952 ( .A1(n7878), .A2(n11673), .Z(\pe9/poht [6]) );
  CLKXOR2HSV4 U9953 ( .A1(n11672), .A2(n11671), .Z(n7878) );
  AOI21HSV4 U9954 ( .A1(n11394), .A2(n11393), .B(n11392), .ZN(n11395) );
  CLKXOR2HSV4 U9955 ( .A1(n10081), .A2(n10080), .Z(n10083) );
  OAI21HSV2 U9956 ( .A1(n8607), .A2(n8608), .B(n8609), .ZN(n8610) );
  XOR2HSV0 U9957 ( .A1(n7879), .A2(n11666), .Z(\pe9/poht [2]) );
  INHSV2 U9958 ( .I(n10842), .ZN(n8544) );
  OAI21HSV2 U9959 ( .A1(n8414), .A2(n8415), .B(n8416), .ZN(n8417) );
  XNOR2HSV4 U9960 ( .A1(n10822), .A2(n10821), .ZN(n10823) );
  AOI21HSV4 U9961 ( .A1(n12092), .A2(n8544), .B(n8545), .ZN(n10843) );
  NAND2HSV2 U9962 ( .A1(n15085), .A2(\pe21/got [4]), .ZN(n10890) );
  NAND2HSV2 U9963 ( .A1(n15085), .A2(\pe21/got [5]), .ZN(n12560) );
  MUX2NHSV2 U9964 ( .I0(n7971), .I1(n12089), .S(n7974), .ZN(n7975) );
  MUX2NHSV1 U9965 ( .I0(n9419), .I1(n8507), .S(n8508), .ZN(n7881) );
  XOR2HSV0 U9966 ( .A1(n7882), .A2(n11644), .Z(\pe9/poht [5]) );
  XOR2HSV0 U9967 ( .A1(n10698), .A2(n10697), .Z(n10701) );
  NAND2HSV2 U9968 ( .A1(\pe6/aot [5]), .A2(\pe6/bq[8] ), .ZN(n9257) );
  NAND2HSV4 U9969 ( .A1(n12453), .A2(n12452), .ZN(n14257) );
  NAND2HSV2 U9970 ( .A1(\pe21/bq[7] ), .A2(\pe21/aot [5]), .ZN(n10651) );
  XOR2HSV0 U9971 ( .A1(n9045), .A2(n9044), .Z(n9046) );
  NAND2HSV2 U9972 ( .A1(n9015), .A2(n9014), .ZN(n9020) );
  NAND2HSV2 U9973 ( .A1(\pe18/ctrq ), .A2(\pe18/pvq [5]), .ZN(n9202) );
  XOR2HSV0 U9974 ( .A1(n9625), .A2(n9624), .Z(n9626) );
  OAI21HSV2 U9975 ( .A1(n9481), .A2(n9480), .B(n9479), .ZN(n9483) );
  AOI22HSV2 U9976 ( .A1(n11303), .A2(n11302), .B1(n11301), .B2(n11300), .ZN(
        n11307) );
  NAND2HSV4 U9977 ( .A1(n11334), .A2(n11333), .ZN(n13865) );
  NAND2HSV4 U9978 ( .A1(n11227), .A2(n11226), .ZN(n13086) );
  NAND2HSV2 U9979 ( .A1(n12603), .A2(n11284), .ZN(n12079) );
  NAND2HSV2 U9980 ( .A1(n9061), .A2(n11888), .ZN(n9033) );
  INHSV4 U9981 ( .I(n6735), .ZN(n13255) );
  CLKXOR2HSV4 U9982 ( .A1(n10083), .A2(n10082), .Z(n10085) );
  INHSV2 U9983 ( .I(n10997), .ZN(n13888) );
  NAND2HSV2 U9984 ( .A1(\pe3/got [8]), .A2(\pe3/ti_1 ), .ZN(n10164) );
  NOR2HSV2 U9985 ( .A1(n11946), .A2(n11948), .ZN(n11945) );
  AND2HSV4 U9986 ( .A1(n11946), .A2(n11942), .Z(n8909) );
  IOA22HSV1 U9987 ( .B1(n10014), .B2(n11832), .A1(n13591), .A2(\pe13/aot [1]), 
        .ZN(n10015) );
  XNOR2HSV1 U9988 ( .A1(n12662), .A2(n12661), .ZN(n12663) );
  NAND2HSV2 U9989 ( .A1(\pe20/pvq [3]), .A2(\pe20/ctrq ), .ZN(n9017) );
  NAND2HSV2 U9990 ( .A1(\pe3/pvq [4]), .A2(\pe3/ctrq ), .ZN(n10192) );
  NAND2HSV2 U9991 ( .A1(\pe19/aot [8]), .A2(\pe19/bq[5] ), .ZN(n12152) );
  CLKXOR2HSV2 U9992 ( .A1(n9049), .A2(\pe20/phq [4]), .Z(n9051) );
  NAND2HSV0 U9993 ( .A1(n13824), .A2(\pe6/got [1]), .ZN(n13042) );
  NAND2HSV0 U9994 ( .A1(\pe21/ti_7[1] ), .A2(\pe21/got [1]), .ZN(n12097) );
  NAND2HSV2 U9995 ( .A1(n14505), .A2(\pe14/aot [3]), .ZN(n11105) );
  MUX2NHSV1 U9996 ( .I0(n9440), .I1(n7908), .S(n7911), .ZN(n9428) );
  CLKNAND2HSV2 U9997 ( .A1(n12232), .A2(n10459), .ZN(n12201) );
  AND2HSV2 U9998 ( .A1(n11267), .A2(n11266), .Z(n11268) );
  NAND2HSV4 U9999 ( .A1(n11367), .A2(n11366), .ZN(n11336) );
  OAI21HSV2 U10000 ( .A1(n15198), .A2(n9801), .B(n9800), .ZN(n9839) );
  NOR2HSV2 U10001 ( .A1(n11605), .A2(n11603), .ZN(n11604) );
  NAND2HSV2 U10002 ( .A1(n9729), .A2(n9728), .ZN(n9731) );
  NAND3HSV2 U10003 ( .A1(n10608), .A2(n13884), .A3(n10601), .ZN(n10604) );
  NAND2HSV2 U10004 ( .A1(n14257), .A2(\pe11/got [2]), .ZN(n14263) );
  XOR2HSV0 U10005 ( .A1(n12455), .A2(n12454), .Z(po11) );
  NAND2HSV2 U10006 ( .A1(n14257), .A2(n15179), .ZN(n12454) );
  XOR2HSV0 U10007 ( .A1(n12471), .A2(n12470), .Z(\pe11/poht [3]) );
  NAND2HSV2 U10008 ( .A1(n14257), .A2(\pe11/got [5]), .ZN(n12470) );
  XNOR2HSV1 U10009 ( .A1(n12463), .A2(n12462), .ZN(n12465) );
  XOR2HSV0 U10010 ( .A1(n12573), .A2(n12572), .Z(\pe11/poht [2]) );
  XOR2HSV0 U10011 ( .A1(n9796), .A2(n9795), .Z(\pe9/poht [4]) );
  CLKXOR2HSV2 U10012 ( .A1(n9760), .A2(n9759), .Z(n9761) );
  AOI22HSV2 U10013 ( .A1(n9754), .A2(n9753), .B1(n9752), .B2(n9751), .ZN(n9760) );
  NAND2HSV2 U10014 ( .A1(n13086), .A2(n13085), .ZN(n13087) );
  NAND2HSV2 U10015 ( .A1(n14933), .A2(n6707), .ZN(n9672) );
  CLKNAND2HSV2 U10016 ( .A1(n15283), .A2(n10510), .ZN(n10512) );
  BUFHSV2 U10017 ( .I(n13762), .Z(n14934) );
  NAND2HSV2 U10018 ( .A1(n10150), .A2(n10149), .ZN(\pe20/ti_7[5] ) );
  NOR2HSV2 U10019 ( .A1(n12713), .A2(n14245), .ZN(n12676) );
  NAND2HSV2 U10020 ( .A1(n6171), .A2(\pe2/got [1]), .ZN(n13433) );
  NAND2HSV4 U10021 ( .A1(n9713), .A2(n9674), .ZN(n14933) );
  XOR2HSV0 U10022 ( .A1(n13106), .A2(n13105), .Z(n15197) );
  XOR2HSV0 U10023 ( .A1(n11166), .A2(n11165), .Z(n7883) );
  CLKNHSV0 U10024 ( .I(n13211), .ZN(n7884) );
  CLKNHSV0 U10025 ( .I(n14273), .ZN(n7885) );
  NAND2HSV0 U10026 ( .A1(\pe16/got [4]), .A2(n13219), .ZN(n7887) );
  OAI21HSV0 U10027 ( .A1(n7886), .A2(n7887), .B(n7888), .ZN(n11169) );
  CLKNAND2HSV0 U10028 ( .A1(\pe14/pvq [4]), .A2(\pe14/ctrq ), .ZN(n7889) );
  NAND2HSV0 U10029 ( .A1(\pe14/bq[6] ), .A2(\pe14/aot [7]), .ZN(n7890) );
  NAND2HSV0 U10030 ( .A1(n7890), .A2(n7889), .ZN(n7891) );
  OAI21HSV2 U10031 ( .A1(n7889), .A2(n7890), .B(n7891), .ZN(n9106) );
  NOR2HSV0 U10032 ( .A1(n10592), .A2(ctro20), .ZN(n7892) );
  OAI21HSV2 U10033 ( .A1(n15278), .A2(n13018), .B(n11472), .ZN(n7893) );
  AOI21HSV4 U10034 ( .A1(n11476), .A2(n7893), .B(n7894), .ZN(n12791) );
  CLKNHSV0 U10035 ( .I(\pe19/phq [1]), .ZN(n7895) );
  INAND2HSV2 U10036 ( .A1(\pe21/ti_7t [1]), .B1(n11780), .ZN(n10396) );
  NAND2HSV0 U10037 ( .A1(\pe18/ti_7[1] ), .A2(\pe18/got [3]), .ZN(n7897) );
  NAND2HSV0 U10038 ( .A1(n7898), .A2(n7897), .ZN(n7899) );
  OAI21HSV0 U10039 ( .A1(n7897), .A2(n7898), .B(n7899), .ZN(n11997) );
  INOR2HSV1 U10040 ( .A1(n11512), .B1(n11538), .ZN(n11514) );
  INAND2HSV0 U10041 ( .A1(\pe19/ti_7t [5]), .B1(n10357), .ZN(n12138) );
  NAND2HSV0 U10042 ( .A1(n10686), .A2(\pe16/got [7]), .ZN(n7900) );
  INOR2HSV2 U10043 ( .A1(\pe17/ti_7t [1]), .B1(n12014), .ZN(n10418) );
  AOI22HSV0 U10044 ( .A1(\pe1/bq[8] ), .A2(\pe1/aot [3]), .B1(\pe1/bq[3] ), 
        .B2(\pe1/aot [8]), .ZN(n7901) );
  NAND2HSV0 U10045 ( .A1(\pe13/ti_7[1] ), .A2(\pe13/got [2]), .ZN(n7902) );
  NAND2HSV0 U10046 ( .A1(\pe13/got [3]), .A2(n9882), .ZN(n7903) );
  NAND2HSV2 U10047 ( .A1(n7903), .A2(n7902), .ZN(n7904) );
  OAI21HSV2 U10048 ( .A1(n7902), .A2(n7903), .B(n7904), .ZN(n13602) );
  INAND2HSV0 U10049 ( .A1(\pe21/ti_7t [3]), .B1(n10863), .ZN(n10644) );
  INHSV2 U10050 ( .I(n9440), .ZN(n7908) );
  NAND2HSV0 U10051 ( .A1(\pe9/pvq [4]), .A2(\pe9/ctrq ), .ZN(n7909) );
  NAND2HSV0 U10052 ( .A1(n7909), .A2(\pe9/phq [4]), .ZN(n7910) );
  OAI21HSV2 U10053 ( .A1(\pe9/phq [4]), .A2(n7909), .B(n7910), .ZN(n7911) );
  INAND2HSV0 U10054 ( .A1(\pe17/ti_7t [5]), .B1(n12021), .ZN(n12104) );
  NAND2HSV2 U10055 ( .A1(n9133), .A2(\pe18/ti_7t [1]), .ZN(n9139) );
  NAND2HSV0 U10056 ( .A1(\pe10/got [7]), .A2(n15075), .ZN(n7912) );
  NAND2HSV0 U10057 ( .A1(n14964), .A2(\pe14/got [2]), .ZN(n7914) );
  NAND2HSV0 U10058 ( .A1(\pe14/got [3]), .A2(n14944), .ZN(n7915) );
  NAND2HSV0 U10059 ( .A1(n7915), .A2(n7914), .ZN(n7916) );
  OAI21HSV2 U10060 ( .A1(n7914), .A2(n7915), .B(n7916), .ZN(n13078) );
  NAND2HSV0 U10061 ( .A1(\pe1/bq[2] ), .A2(\pe1/aot [7]), .ZN(n7917) );
  OAI21HSV0 U10062 ( .A1(n13968), .A2(n13969), .B(n7917), .ZN(n7918) );
  OAI31HSV0 U10063 ( .A1(n13968), .A2(n7917), .A3(n13969), .B(n7918), .ZN(
        n13973) );
  NAND2HSV0 U10064 ( .A1(n9898), .A2(\pe13/got [7]), .ZN(n7919) );
  NOR2HSV4 U10065 ( .A1(n9900), .A2(n7919), .ZN(n9904) );
  INAND2HSV0 U10066 ( .A1(\pe3/ti_7t [3]), .B1(n10994), .ZN(n10946) );
  INOR2HSV0 U10067 ( .A1(\pe17/ti_7t [3]), .B1(n12014), .ZN(n12020) );
  XOR2HSV0 U10068 ( .A1(n11717), .A2(n11718), .Z(n7921) );
  XOR2HSV0 U10069 ( .A1(\pe11/phq [5]), .A2(n11719), .Z(n7922) );
  XOR2HSV0 U10070 ( .A1(n7921), .A2(n7922), .Z(n7923) );
  CLKNHSV0 U10071 ( .I(n11715), .ZN(n7925) );
  NAND2HSV0 U10072 ( .A1(n11797), .A2(n14837), .ZN(n7926) );
  MUX2NHSV2 U10073 ( .I0(n7925), .I1(n11715), .S(n7926), .ZN(n7927) );
  NAND2HSV0 U10074 ( .A1(n14381), .A2(\pe11/got [6]), .ZN(n7930) );
  NAND2HSV0 U10075 ( .A1(n9636), .A2(\pe4/got [7]), .ZN(n7931) );
  NOR2HSV4 U10076 ( .A1(n9635), .A2(n7931), .ZN(n9643) );
  CLKNHSV0 U10077 ( .I(n13145), .ZN(n7932) );
  NAND2HSV0 U10078 ( .A1(n13146), .A2(\pe18/ti_7t [5]), .ZN(n7933) );
  CLKNHSV0 U10079 ( .I(n15082), .ZN(n7934) );
  INAND2HSV2 U10080 ( .A1(n10799), .B1(\pe6/ti_7t [6]), .ZN(n9846) );
  NAND2HSV0 U10081 ( .A1(\pe18/pvq [4]), .A2(\pe18/ctrq ), .ZN(n7935) );
  NAND2HSV0 U10082 ( .A1(n7935), .A2(\pe18/phq [4]), .ZN(n7936) );
  OAI21HSV2 U10083 ( .A1(\pe18/phq [4]), .A2(n7935), .B(n7936), .ZN(n9162) );
  NAND2HSV0 U10084 ( .A1(\pe13/bq[6] ), .A2(\pe13/aot [1]), .ZN(n7938) );
  NAND2HSV0 U10085 ( .A1(\pe13/bq[1] ), .A2(\pe13/aot [6]), .ZN(n7939) );
  CLKNAND2HSV0 U10086 ( .A1(n7939), .A2(n7938), .ZN(n7940) );
  OAI21HSV0 U10087 ( .A1(n7938), .A2(n7939), .B(n7940), .ZN(n7941) );
  AOI22HSV0 U10088 ( .A1(\pe13/bq[5] ), .A2(\pe13/aot [2]), .B1(\pe13/aot [5]), 
        .B2(\pe13/bq[2] ), .ZN(n7942) );
  AOI21HSV0 U10089 ( .A1(n13592), .A2(n12922), .B(n7942), .ZN(n7943) );
  NAND2HSV0 U10090 ( .A1(n7943), .A2(n7941), .ZN(n7944) );
  OAI21HSV2 U10091 ( .A1(n7943), .A2(n7941), .B(n7944), .ZN(n7945) );
  NAND2HSV0 U10092 ( .A1(\pe13/aot [3]), .A2(\pe13/bq[4] ), .ZN(n7946) );
  NAND2HSV2 U10093 ( .A1(n7946), .A2(n7945), .ZN(n7947) );
  OAI21HSV2 U10094 ( .A1(n7945), .A2(n7946), .B(n7947), .ZN(n7948) );
  NAND2HSV0 U10095 ( .A1(\pe13/bq[3] ), .A2(\pe13/aot [4]), .ZN(n7949) );
  NAND2HSV2 U10096 ( .A1(n7949), .A2(n7948), .ZN(n7950) );
  OAI21HSV2 U10097 ( .A1(n7948), .A2(n7949), .B(n7950), .ZN(n9928) );
  CLKNHSV0 U10098 ( .I(n13970), .ZN(n7951) );
  AOI22HSV0 U10099 ( .A1(\pe1/aot [1]), .A2(n14502), .B1(\pe1/bq[5] ), .B2(
        \pe1/aot [4]), .ZN(n7952) );
  AOI21HSV0 U10100 ( .A1(n13971), .A2(n7951), .B(n7952), .ZN(n13972) );
  AOI21HSV0 U10101 ( .A1(n11113), .A2(n11093), .B(n11089), .ZN(n7953) );
  CLKNHSV0 U10102 ( .I(\pe2/phq [3]), .ZN(n7954) );
  NAND2HSV0 U10103 ( .A1(\pe19/got [5]), .A2(n14219), .ZN(n7955) );
  XOR2HSV0 U10104 ( .A1(n12409), .A2(n12408), .Z(n7956) );
  NAND2HSV0 U10105 ( .A1(n12148), .A2(\pe19/got [4]), .ZN(n7957) );
  XOR2HSV0 U10106 ( .A1(n7956), .A2(n7957), .Z(n7958) );
  XOR2HSV0 U10107 ( .A1(n7955), .A2(n7958), .Z(n7959) );
  AOI22HSV0 U10108 ( .A1(\pe5/bq[3] ), .A2(\pe5/aot [8]), .B1(\pe5/bq[7] ), 
        .B2(\pe5/aot [4]), .ZN(n7960) );
  IAO21HSV2 U10109 ( .A1(n13290), .A2(n11477), .B(n7960), .ZN(n11481) );
  OAI21HSV2 U10110 ( .A1(n7961), .A2(n7962), .B(n7963), .ZN(n7964) );
  NAND2HSV0 U10111 ( .A1(\pe7/aot [7]), .A2(\pe7/bq[5] ), .ZN(n7965) );
  OAI21HSV2 U10112 ( .A1(n7964), .A2(n7965), .B(n7966), .ZN(n7967) );
  NAND2HSV0 U10113 ( .A1(\pe7/aot [4]), .A2(\pe7/bq[8] ), .ZN(n7968) );
  NAND2HSV2 U10114 ( .A1(n7968), .A2(n7967), .ZN(n7969) );
  OAI21HSV2 U10115 ( .A1(n7967), .A2(n7968), .B(n7969), .ZN(n12241) );
  CLKNHSV0 U10116 ( .I(n12089), .ZN(n7971) );
  INHSV2 U10117 ( .I(n10843), .ZN(n7972) );
  NAND2HSV0 U10118 ( .A1(n15092), .A2(\pe21/pvq [7]), .ZN(n7973) );
  MUX2NHSV2 U10119 ( .I0(n7972), .I1(n10843), .S(n7973), .ZN(n7974) );
  XOR2HSV0 U10120 ( .A1(n10850), .A2(n10851), .Z(n7976) );
  NAND2HSV0 U10121 ( .A1(\pe21/got [3]), .A2(\pe21/ti_7[1] ), .ZN(n7977) );
  NAND2HSV0 U10122 ( .A1(\pe19/pvq [6]), .A2(\pe19/ctrq ), .ZN(n7978) );
  NAND2HSV2 U10123 ( .A1(n7978), .A2(\pe19/phq [6]), .ZN(n7979) );
  OAI21HSV2 U10124 ( .A1(\pe19/phq [6]), .A2(n7978), .B(n7979), .ZN(n9569) );
  NAND2HSV0 U10125 ( .A1(\pe16/aot [7]), .A2(\pe16/bq[8] ), .ZN(n7983) );
  IOA21HSV2 U10126 ( .A1(n10800), .A2(n10799), .B(n10801), .ZN(n13034) );
  CLKNHSV0 U10127 ( .I(\pe18/phq [1]), .ZN(n7984) );
  NAND2HSV2 U10128 ( .A1(\pe18/pvq [1]), .A2(\pe18/ctrq ), .ZN(n7985) );
  MUX2NHSV4 U10129 ( .I0(\pe18/phq [1]), .I1(n7984), .S(n7985), .ZN(n9137) );
  INOR2HSV0 U10130 ( .A1(\pe9/ti_7t [4]), .B1(n15074), .ZN(n9746) );
  INOR2HSV0 U10131 ( .A1(\pe1/aot [4]), .B1(n8931), .ZN(n13971) );
  XOR2HSV0 U10132 ( .A1(n13426), .A2(n13428), .Z(n7988) );
  XOR2HSV0 U10133 ( .A1(n13427), .A2(n7988), .Z(n7989) );
  NAND2HSV0 U10134 ( .A1(\pe5/got [4]), .A2(n14916), .ZN(n7990) );
  CLKNAND2HSV0 U10135 ( .A1(n7990), .A2(n7989), .ZN(n7991) );
  OAI21HSV0 U10136 ( .A1(n7989), .A2(n7990), .B(n7991), .ZN(n7992) );
  OAI21HSV2 U10137 ( .A1(n7993), .A2(n7994), .B(n7995), .ZN(n7996) );
  OAI21HSV0 U10138 ( .A1(n13809), .A2(n13429), .B(n7996), .ZN(n7997) );
  NAND2HSV0 U10139 ( .A1(\pe5/ti_7[7] ), .A2(n13861), .ZN(n7999) );
  NAND2HSV0 U10140 ( .A1(n7999), .A2(n7998), .ZN(n8000) );
  OAI21HSV0 U10141 ( .A1(n7998), .A2(n7999), .B(n8000), .ZN(po5) );
  CLKNHSV0 U10142 ( .I(n9298), .ZN(n8001) );
  CLKNHSV0 U10143 ( .I(n12416), .ZN(n8002) );
  NAND2HSV0 U10144 ( .A1(n12475), .A2(\pe3/got [1]), .ZN(n8003) );
  AOI21HSV2 U10145 ( .A1(\pe3/pq ), .A2(n12474), .B(n8003), .ZN(n8004) );
  AO31HSV0 U10146 ( .A1(\pe3/pq ), .A2(n12474), .A3(n8003), .B(n8004), .Z(
        n12480) );
  NAND2HSV0 U10147 ( .A1(n8005), .A2(\pe3/got [6]), .ZN(n8006) );
  NOR2HSV2 U10148 ( .A1(n11586), .A2(n11585), .ZN(n8008) );
  CLKNHSV0 U10149 ( .I(\pe4/got [3]), .ZN(n8009) );
  CLKNHSV0 U10150 ( .I(n13590), .ZN(n8011) );
  AOI22HSV0 U10151 ( .A1(n13591), .A2(\pe13/aot [2]), .B1(\pe13/aot [7]), .B2(
        \pe13/bq[2] ), .ZN(n8012) );
  AOI21HSV0 U10152 ( .A1(n13592), .A2(n8011), .B(n8012), .ZN(n8013) );
  CLKNAND2HSV0 U10153 ( .A1(\pe13/pq ), .A2(n14795), .ZN(n8014) );
  NAND2HSV0 U10154 ( .A1(\pe13/bq[1] ), .A2(n14939), .ZN(n8015) );
  NAND2HSV0 U10155 ( .A1(n8015), .A2(n8014), .ZN(n8016) );
  OAI21HSV0 U10156 ( .A1(n8014), .A2(n8015), .B(n8016), .ZN(n8017) );
  XOR2HSV0 U10157 ( .A1(n8013), .A2(n8017), .Z(n13600) );
  NAND2HSV0 U10158 ( .A1(\pe11/ti_7[1] ), .A2(\pe11/got [2]), .ZN(n8018) );
  NAND2HSV0 U10159 ( .A1(n12561), .A2(\pe11/got [3]), .ZN(n8019) );
  NAND2HSV2 U10160 ( .A1(n8019), .A2(n8018), .ZN(n8020) );
  OAI21HSV2 U10161 ( .A1(n8018), .A2(n8019), .B(n8020), .ZN(n12444) );
  OAI21HSV0 U10162 ( .A1(n14244), .A2(n14243), .B(n14242), .ZN(n8021) );
  XOR2HSV0 U10163 ( .A1(n14239), .A2(n14238), .Z(n8022) );
  XOR2HSV0 U10164 ( .A1(n8021), .A2(n8022), .Z(n8023) );
  AOI21HSV0 U10165 ( .A1(n14246), .A2(n14247), .B(n14245), .ZN(n8024) );
  CLKNHSV0 U10166 ( .I(n14247), .ZN(n8025) );
  CLKNHSV0 U10167 ( .I(n9947), .ZN(n8027) );
  CLKNHSV0 U10168 ( .I(n9587), .ZN(n8029) );
  AOI21HSV2 U10169 ( .A1(n9584), .A2(n9588), .B(n8029), .ZN(n8030) );
  AOI21HSV2 U10170 ( .A1(n9585), .A2(n9589), .B(n9587), .ZN(n8031) );
  AOI21HSV0 U10171 ( .A1(n9723), .A2(n10357), .B(n12139), .ZN(n8032) );
  NAND2HSV0 U10172 ( .A1(n9730), .A2(n9560), .ZN(n8034) );
  NAND2HSV0 U10173 ( .A1(n8037), .A2(n9534), .ZN(n8038) );
  CLKNHSV0 U10174 ( .I(\pe21/phq [3]), .ZN(n8040) );
  CLKNHSV0 U10175 ( .I(n9201), .ZN(n8041) );
  INAND2HSV0 U10176 ( .A1(\pe3/ti_7t [5]), .B1(n10939), .ZN(n11006) );
  OAI31HSV2 U10177 ( .A1(n10583), .A2(n10584), .A3(n10582), .B(n10588), .ZN(
        n12658) );
  AO22HSV2 U10178 ( .A1(\pe2/aot [1]), .A2(n14510), .B1(\pe2/bq[3] ), .B2(
        \pe2/aot [4]), .Z(n8042) );
  AOI22HSV0 U10179 ( .A1(\pe2/bq[2] ), .A2(\pe2/aot [5]), .B1(\pe2/bq[1] ), 
        .B2(\pe2/aot [6]), .ZN(n8043) );
  IAO21HSV2 U10180 ( .A1(n13098), .A2(n12880), .B(n8043), .ZN(n8044) );
  OAI21HSV2 U10181 ( .A1(n12508), .A2(n13092), .B(n8042), .ZN(n8045) );
  NAND2HSV2 U10182 ( .A1(n8045), .A2(n8044), .ZN(n8046) );
  OAI21HSV2 U10183 ( .A1(n8045), .A2(n8044), .B(n8046), .ZN(n8047) );
  NAND2HSV0 U10184 ( .A1(\pe2/aot [2]), .A2(\pe2/bq[5] ), .ZN(n8048) );
  NAND2HSV2 U10185 ( .A1(n8048), .A2(n8047), .ZN(n8049) );
  OAI21HSV2 U10186 ( .A1(n8047), .A2(n8048), .B(n8049), .ZN(n8050) );
  NAND2HSV0 U10187 ( .A1(\pe2/aot [3]), .A2(\pe2/bq[4] ), .ZN(n8051) );
  CLKNAND2HSV0 U10188 ( .A1(n8051), .A2(n8050), .ZN(n8052) );
  OAI21HSV2 U10189 ( .A1(n8050), .A2(n8051), .B(n8052), .ZN(n12509) );
  CLKNHSV0 U10190 ( .I(n12090), .ZN(n8053) );
  MUX2NHSV0 U10191 ( .I0(n8053), .I1(n12090), .S(n12095), .ZN(n8054) );
  XOR2HSV0 U10192 ( .A1(n8054), .A2(n12096), .Z(n8055) );
  XOR2HSV0 U10193 ( .A1(n12097), .A2(n12091), .Z(n8056) );
  XOR2HSV0 U10194 ( .A1(n8055), .A2(n8056), .Z(n8057) );
  CLKNAND2HSV0 U10195 ( .A1(n8058), .A2(n8057), .ZN(n8059) );
  OAI21HSV0 U10196 ( .A1(n8057), .A2(n8058), .B(n8059), .ZN(n8060) );
  NAND2HSV0 U10197 ( .A1(\pe21/ti_7[3] ), .A2(\pe21/got [3]), .ZN(n8061) );
  CLKNAND2HSV0 U10198 ( .A1(n8061), .A2(n8060), .ZN(n8062) );
  OAI21HSV0 U10199 ( .A1(n8060), .A2(n8061), .B(n8062), .ZN(n8063) );
  NAND2HSV0 U10200 ( .A1(\pe21/got [4]), .A2(n12542), .ZN(n8064) );
  CLKNAND2HSV0 U10201 ( .A1(n8064), .A2(n8063), .ZN(n8065) );
  OAI21HSV2 U10202 ( .A1(n8063), .A2(n8064), .B(n8065), .ZN(n8066) );
  CLKNAND2HSV0 U10203 ( .A1(n8067), .A2(n8066), .ZN(n8068) );
  OAI21HSV2 U10204 ( .A1(n8066), .A2(n8067), .B(n8068), .ZN(n12098) );
  NAND2HSV0 U10205 ( .A1(\pe2/ti_7[1] ), .A2(\pe2/got [2]), .ZN(n8069) );
  CLKNHSV0 U10206 ( .I(n12667), .ZN(n8070) );
  XOR2HSV0 U10207 ( .A1(n11454), .A2(n11459), .Z(n8071) );
  XOR2HSV0 U10208 ( .A1(n11465), .A2(n11464), .Z(n8072) );
  NAND2HSV0 U10209 ( .A1(\pe12/got [3]), .A2(\pe12/ti_7[1] ), .ZN(n8073) );
  NAND2HSV0 U10210 ( .A1(\pe12/got [4]), .A2(n14255), .ZN(n8075) );
  NAND2HSV2 U10211 ( .A1(n8075), .A2(n8074), .ZN(n8076) );
  OAI21HSV2 U10212 ( .A1(n8074), .A2(n8075), .B(n8076), .ZN(n8077) );
  NAND2HSV2 U10213 ( .A1(n8078), .A2(n8077), .ZN(n8079) );
  OAI21HSV2 U10214 ( .A1(n8077), .A2(n8078), .B(n8079), .ZN(n8080) );
  CLKNHSV0 U10215 ( .I(n11512), .ZN(n8081) );
  INHSV2 U10216 ( .I(n11515), .ZN(n8082) );
  CLKNHSV0 U10217 ( .I(\pe7/got [3]), .ZN(n8086) );
  XOR2HSV0 U10218 ( .A1(n13616), .A2(n13615), .Z(n8087) );
  NAND2HSV0 U10219 ( .A1(\pe7/aot [3]), .A2(\pe7/bq[5] ), .ZN(n8089) );
  CLKNAND2HSV0 U10220 ( .A1(n8089), .A2(n13618), .ZN(n8090) );
  OAI21HSV0 U10221 ( .A1(n13618), .A2(n8089), .B(n8090), .ZN(n8091) );
  NAND2HSV0 U10222 ( .A1(\pe7/got [1]), .A2(\pe7/ti_7[1] ), .ZN(n8092) );
  CLKNAND2HSV0 U10223 ( .A1(n8092), .A2(n8091), .ZN(n8093) );
  OAI21HSV0 U10224 ( .A1(n8091), .A2(n8092), .B(n8093), .ZN(n8094) );
  NAND2HSV0 U10225 ( .A1(\pe7/got [2]), .A2(n14860), .ZN(n8095) );
  CLKNAND2HSV0 U10226 ( .A1(n8095), .A2(n8094), .ZN(n8096) );
  OAI21HSV0 U10227 ( .A1(n8094), .A2(n8095), .B(n8096), .ZN(n8097) );
  XOR2HSV0 U10228 ( .A1(n8088), .A2(n8097), .Z(n13619) );
  OAI21HSV4 U10229 ( .A1(n8098), .A2(n8099), .B(n8100), .ZN(n9512) );
  NAND2HSV0 U10230 ( .A1(n13844), .A2(n13316), .ZN(n8101) );
  NAND2HSV0 U10231 ( .A1(n8101), .A2(n13260), .ZN(n8102) );
  OAI21HSV0 U10232 ( .A1(n13260), .A2(n8101), .B(n8102), .ZN(\pov19[7] ) );
  CLKNHSV0 U10233 ( .I(\pe3/phq [7]), .ZN(n8103) );
  NAND2HSV2 U10234 ( .A1(\pe3/pvq [7]), .A2(n10979), .ZN(n8104) );
  MUX2NHSV1 U10235 ( .I0(\pe3/phq [7]), .I1(n8103), .S(n8104), .ZN(n10980) );
  NAND2HSV0 U10236 ( .A1(n12362), .A2(\pe20/pvq [7]), .ZN(n8105) );
  NAND2HSV0 U10237 ( .A1(n8105), .A2(\pe20/phq [7]), .ZN(n8106) );
  OAI21HSV0 U10238 ( .A1(\pe20/phq [7]), .A2(n8105), .B(n8106), .ZN(n11860) );
  INOR2HSV4 U10239 ( .A1(\pe4/ti_7t [1]), .B1(n14955), .ZN(n9613) );
  INOR2HSV0 U10240 ( .A1(\pe16/ti_7t [3]), .B1(n10796), .ZN(n11159) );
  INAND2HSV2 U10241 ( .A1(\pe6/ti_7t [4]), .B1(n15088), .ZN(n9312) );
  CLKNHSV0 U10242 ( .I(\pe3/phq [3]), .ZN(n8107) );
  INOR2HSV4 U10243 ( .A1(\pe11/ti_7t [1]), .B1(n10807), .ZN(n11914) );
  NAND2HSV0 U10244 ( .A1(n10943), .A2(n10994), .ZN(n8109) );
  NAND2HSV0 U10245 ( .A1(\pe21/aot [4]), .A2(\pe21/bq[1] ), .ZN(n8110) );
  NAND2HSV0 U10246 ( .A1(\pe21/bq[2] ), .A2(\pe21/aot [3]), .ZN(n8111) );
  CLKNAND2HSV0 U10247 ( .A1(n8111), .A2(n8110), .ZN(n8112) );
  OAI21HSV0 U10248 ( .A1(n8110), .A2(n8111), .B(n8112), .ZN(n8113) );
  NAND2HSV0 U10249 ( .A1(\pe21/aot [2]), .A2(\pe21/bq[3] ), .ZN(n8114) );
  CLKNAND2HSV0 U10250 ( .A1(n8114), .A2(n8113), .ZN(n8115) );
  OAI21HSV0 U10251 ( .A1(n8113), .A2(n8114), .B(n8115), .ZN(n8116) );
  NAND2HSV0 U10252 ( .A1(\pe21/aot [1]), .A2(\pe21/bq[4] ), .ZN(n8117) );
  CLKNAND2HSV0 U10253 ( .A1(n8117), .A2(n8116), .ZN(n8118) );
  OAI21HSV0 U10254 ( .A1(n8116), .A2(n8117), .B(n8118), .ZN(n8119) );
  NAND2HSV0 U10255 ( .A1(\pe21/got [1]), .A2(n12542), .ZN(n8120) );
  CLKNAND2HSV0 U10256 ( .A1(n8120), .A2(n8119), .ZN(n8121) );
  OAI21HSV0 U10257 ( .A1(n8119), .A2(n8120), .B(n8121), .ZN(n8122) );
  NAND2HSV0 U10258 ( .A1(\pe12/ti_7[1] ), .A2(\pe12/got [2]), .ZN(n8123) );
  NAND2HSV0 U10259 ( .A1(\pe12/got [3]), .A2(n14255), .ZN(n8124) );
  NAND2HSV0 U10260 ( .A1(n8124), .A2(n8123), .ZN(n8125) );
  OAI21HSV2 U10261 ( .A1(n8123), .A2(n8124), .B(n8125), .ZN(n12701) );
  INAND2HSV0 U10262 ( .A1(\pe2/ti_7t [3]), .B1(n9358), .ZN(n9359) );
  CLKNHSV0 U10263 ( .I(n12418), .ZN(n8126) );
  AOI22HSV0 U10264 ( .A1(\pe6/bq[7] ), .A2(\pe6/aot [1]), .B1(\pe6/bq[4] ), 
        .B2(\pe6/aot [4]), .ZN(n8127) );
  XOR2HSV0 U10265 ( .A1(n12414), .A2(n12415), .Z(n8128) );
  XOR2HSV0 U10266 ( .A1(n12413), .A2(n12412), .Z(n8129) );
  XOR2HSV0 U10267 ( .A1(n8128), .A2(n8129), .Z(n8130) );
  OAI21HSV0 U10268 ( .A1(n12417), .A2(n8127), .B(n8130), .ZN(n8131) );
  OAI31HSV0 U10269 ( .A1(n12417), .A2(n8130), .A3(n8127), .B(n8131), .ZN(n8132) );
  MUX2NHSV0 U10270 ( .I0(n8126), .I1(n12418), .S(n8132), .ZN(n8133) );
  NAND2HSV0 U10271 ( .A1(n14895), .A2(\pe6/got [1]), .ZN(n8134) );
  CLKNAND2HSV0 U10272 ( .A1(n8134), .A2(n8133), .ZN(n8135) );
  OAI21HSV0 U10273 ( .A1(n8133), .A2(n8134), .B(n8135), .ZN(n8136) );
  NAND2HSV0 U10274 ( .A1(n13034), .A2(\pe6/got [2]), .ZN(n8137) );
  NAND2HSV0 U10275 ( .A1(n8137), .A2(n8136), .ZN(n8138) );
  OAI21HSV2 U10276 ( .A1(n8136), .A2(n8137), .B(n8138), .ZN(n12420) );
  CLKNHSV0 U10277 ( .I(\pe1/got [6]), .ZN(n8139) );
  NAND2HSV0 U10278 ( .A1(\pe1/bq[5] ), .A2(\pe1/aot [6]), .ZN(n8140) );
  NAND2HSV0 U10279 ( .A1(n8140), .A2(n10618), .ZN(n8141) );
  OAI21HSV0 U10280 ( .A1(n10618), .A2(n8140), .B(n8141), .ZN(n8142) );
  XOR2HSV0 U10281 ( .A1(n10282), .A2(n8142), .Z(n8143) );
  XOR2HSV0 U10282 ( .A1(n10279), .A2(n10280), .Z(n8144) );
  XOR2HSV0 U10283 ( .A1(n8143), .A2(n8144), .Z(n8145) );
  NAND2HSV0 U10284 ( .A1(\pe1/got [4]), .A2(n10242), .ZN(n8146) );
  NAND2HSV2 U10285 ( .A1(n8146), .A2(n8145), .ZN(n8147) );
  NAND2HSV0 U10286 ( .A1(\pe1/got [5]), .A2(\pe1/ti_7[2] ), .ZN(n8148) );
  NAND2HSV0 U10287 ( .A1(n14703), .A2(n10283), .ZN(n8150) );
  OAI21HSV2 U10288 ( .A1(n8149), .A2(n8150), .B(n8151), .ZN(n13884) );
  NAND2HSV0 U10289 ( .A1(\pe4/bq[1] ), .A2(\pe4/aot [2]), .ZN(n8153) );
  NAND2HSV0 U10290 ( .A1(\pe4/aot [1]), .A2(\pe4/bq[2] ), .ZN(n8154) );
  CLKNAND2HSV0 U10291 ( .A1(n8154), .A2(n8153), .ZN(n8155) );
  OAI21HSV0 U10292 ( .A1(n8153), .A2(n8154), .B(n8155), .ZN(n8156) );
  XOR2HSV0 U10293 ( .A1(n8152), .A2(n8156), .Z(n8157) );
  NAND2HSV0 U10294 ( .A1(\pe4/got [2]), .A2(n6706), .ZN(n8158) );
  CLKNAND2HSV0 U10295 ( .A1(n8158), .A2(n8157), .ZN(n8159) );
  OAI21HSV0 U10296 ( .A1(n8157), .A2(n8158), .B(n8159), .ZN(\pe4/poht [6]) );
  NAND2HSV0 U10297 ( .A1(n10443), .A2(\pe9/got [4]), .ZN(n8160) );
  CLKNAND2HSV0 U10298 ( .A1(n8160), .A2(n11635), .ZN(n8161) );
  OAI21HSV0 U10299 ( .A1(n11635), .A2(n8160), .B(n8161), .ZN(n8162) );
  CLKNAND2HSV0 U10300 ( .A1(n8163), .A2(n8162), .ZN(n8164) );
  OAI21HSV0 U10301 ( .A1(n8162), .A2(n8163), .B(n8164), .ZN(n8165) );
  NAND2HSV0 U10302 ( .A1(n14963), .A2(\pe9/got [6]), .ZN(n8166) );
  XOR2HSV0 U10303 ( .A1(n13600), .A2(n13601), .Z(n8172) );
  NAND2HSV0 U10304 ( .A1(n15065), .A2(\pe13/got [4]), .ZN(n8173) );
  NAND2HSV0 U10305 ( .A1(\pe13/got [5]), .A2(n13587), .ZN(n8175) );
  OAI21HSV0 U10306 ( .A1(n8174), .A2(n8175), .B(n8176), .ZN(n8177) );
  NAND2HSV0 U10307 ( .A1(n13603), .A2(\pe13/got [6]), .ZN(n8178) );
  CLKNAND2HSV0 U10308 ( .A1(n8177), .A2(n8178), .ZN(n8179) );
  OAI21HSV0 U10309 ( .A1(n8177), .A2(n8178), .B(n8179), .ZN(n8180) );
  NAND2HSV0 U10310 ( .A1(n12997), .A2(\pe13/got [7]), .ZN(n8181) );
  CLKNAND2HSV0 U10311 ( .A1(n8181), .A2(n8180), .ZN(n8182) );
  OAI21HSV0 U10312 ( .A1(n8183), .A2(n8184), .B(n8185), .ZN(po13) );
  XOR2HSV0 U10313 ( .A1(n14028), .A2(n14027), .Z(n8186) );
  OAI21HSV0 U10314 ( .A1(n15167), .A2(n14309), .B(n8186), .ZN(n8187) );
  OAI31HSV0 U10315 ( .A1(n15167), .A2(n8186), .A3(n14309), .B(n8187), .ZN(
        n8188) );
  XOR2HSV0 U10316 ( .A1(n13748), .A2(n13747), .Z(n8189) );
  NAND2HSV0 U10317 ( .A1(n15184), .A2(\pe20/got [5]), .ZN(n8190) );
  CLKNAND2HSV0 U10318 ( .A1(n8190), .A2(n8189), .ZN(n8191) );
  OAI21HSV2 U10319 ( .A1(n8189), .A2(n8190), .B(n8191), .ZN(n8192) );
  OAI21HSV0 U10320 ( .A1(n8193), .A2(n8194), .B(n8195), .ZN(po20) );
  IOA21HSV2 U10321 ( .A1(n9500), .A2(n9541), .B(n9556), .ZN(\pe19/ti_7[1] ) );
  NAND2HSV2 U10322 ( .A1(n15160), .A2(\pe15/pvq [7]), .ZN(n8196) );
  NAND2HSV2 U10323 ( .A1(n8196), .A2(\pe15/phq [7]), .ZN(n8197) );
  OAI21HSV2 U10324 ( .A1(\pe15/phq [7]), .A2(n8196), .B(n8197), .ZN(n8198) );
  NAND2HSV0 U10325 ( .A1(n14587), .A2(\pe15/got [2]), .ZN(n8199) );
  NAND2HSV2 U10326 ( .A1(n8199), .A2(n8198), .ZN(n8200) );
  OAI21HSV2 U10327 ( .A1(n8198), .A2(n8199), .B(n8200), .ZN(n8201) );
  NAND2HSV0 U10328 ( .A1(\pe15/aot [2]), .A2(n14602), .ZN(n8202) );
  NAND2HSV2 U10329 ( .A1(n8202), .A2(n8201), .ZN(n8203) );
  OAI21HSV2 U10330 ( .A1(n8201), .A2(n8202), .B(n8203), .ZN(n12330) );
  NAND3HSV0 U10331 ( .A1(n11448), .A2(n11436), .A3(n11437), .ZN(n11435) );
  NAND2HSV4 U10332 ( .A1(\pe20/ti_1 ), .A2(\pe20/got [8]), .ZN(n8205) );
  OAI21HSV4 U10333 ( .A1(n8205), .A2(n8204), .B(n8206), .ZN(n9032) );
  INOR2HSV0 U10334 ( .A1(\pe10/ti_7t [4]), .B1(n10924), .ZN(n14119) );
  CLKNHSV0 U10335 ( .I(n14353), .ZN(n8208) );
  AOI22HSV0 U10336 ( .A1(\pe16/bq[3] ), .A2(\pe16/aot [3]), .B1(\pe16/aot [4]), 
        .B2(\pe16/bq[2] ), .ZN(n8209) );
  IAO21HSV2 U10337 ( .A1(n14352), .A2(n14351), .B(n8209), .ZN(n8210) );
  MUX2NHSV1 U10338 ( .I0(n14353), .I1(n8208), .S(n8210), .ZN(n14357) );
  OAI21HSV0 U10339 ( .A1(n11782), .A2(\pe7/ti_7t [5]), .B(n5967), .ZN(n8211)
         );
  AOI21HSV0 U10340 ( .A1(n12131), .A2(n12130), .B(n14008), .ZN(n8212) );
  OR2HSV1 U10341 ( .A1(n10787), .A2(n10786), .Z(n10110) );
  CLKNHSV0 U10342 ( .I(\pe11/got [2]), .ZN(n8215) );
  XOR2HSV0 U10343 ( .A1(n13758), .A2(n13757), .Z(n8216) );
  NAND2HSV0 U10344 ( .A1(\pe11/got [1]), .A2(n14365), .ZN(n8217) );
  CLKNAND2HSV0 U10345 ( .A1(n8217), .A2(n8216), .ZN(n8218) );
  OAI21HSV0 U10346 ( .A1(n8216), .A2(n8217), .B(n8218), .ZN(n8219) );
  OAI21HSV0 U10347 ( .A1(n14396), .A2(n8215), .B(n8219), .ZN(n8220) );
  OAI31HSV0 U10348 ( .A1(n14396), .A2(n8219), .A3(n8215), .B(n8220), .ZN(n8221) );
  NAND2HSV0 U10349 ( .A1(\pe11/got [3]), .A2(n14388), .ZN(n8222) );
  CLKNAND2HSV0 U10350 ( .A1(n8222), .A2(n8221), .ZN(n8223) );
  OAI21HSV0 U10351 ( .A1(n8224), .A2(n8225), .B(n8226), .ZN(\pe11/poht [4]) );
  CLKNHSV0 U10352 ( .I(n15077), .ZN(n8227) );
  NAND2HSV0 U10353 ( .A1(n8229), .A2(n8228), .ZN(n8230) );
  OAI21HSV0 U10354 ( .A1(n8228), .A2(n8229), .B(n8230), .ZN(\pe6/poht [3]) );
  CLKNHSV0 U10355 ( .I(\pe13/got [2]), .ZN(n8231) );
  XOR2HSV0 U10356 ( .A1(n12993), .A2(n12992), .Z(n8232) );
  XOR2HSV0 U10357 ( .A1(n12996), .A2(n8232), .Z(n8233) );
  NAND2HSV0 U10358 ( .A1(n13587), .A2(\pe13/got [1]), .ZN(n8234) );
  CLKNAND2HSV0 U10359 ( .A1(n8234), .A2(n8233), .ZN(n8235) );
  OAI21HSV0 U10360 ( .A1(n8233), .A2(n8234), .B(n8235), .ZN(n8236) );
  NAND2HSV0 U10361 ( .A1(n13826), .A2(n15093), .ZN(n8240) );
  OAI21HSV0 U10362 ( .A1(bo9[8]), .A2(n13826), .B(n8240), .ZN(n15133) );
  CLKNHSV0 U10363 ( .I(\pe8/ti_7t [7]), .ZN(n8241) );
  AOI21HSV0 U10364 ( .A1(n14189), .A2(n8241), .B(n15134), .ZN(n8242) );
  XOR2HSV0 U10365 ( .A1(n14210), .A2(n14211), .Z(n8243) );
  XOR2HSV0 U10366 ( .A1(n14195), .A2(n14194), .Z(n8244) );
  XOR2HSV0 U10367 ( .A1(n8243), .A2(n8244), .Z(n8245) );
  NAND2HSV0 U10368 ( .A1(n15066), .A2(\pe8/got [3]), .ZN(n8246) );
  CLKNAND2HSV0 U10369 ( .A1(n8246), .A2(n8245), .ZN(n8247) );
  OAI21HSV0 U10370 ( .A1(n8249), .A2(n8248), .B(n8250), .ZN(\pe8/poht [2]) );
  XOR2HSV0 U10371 ( .A1(n11287), .A2(n11288), .Z(n8251) );
  XOR2HSV0 U10372 ( .A1(n11286), .A2(n11285), .Z(n8252) );
  XOR2HSV0 U10373 ( .A1(n8251), .A2(n8252), .Z(n8253) );
  NAND2HSV0 U10374 ( .A1(n12631), .A2(\pe4/got [1]), .ZN(n8254) );
  CLKNAND2HSV0 U10375 ( .A1(n8254), .A2(n8253), .ZN(n8255) );
  OAI21HSV0 U10376 ( .A1(n8253), .A2(n8254), .B(n8255), .ZN(n8256) );
  NAND2HSV0 U10377 ( .A1(n14850), .A2(\pe4/got [2]), .ZN(n8257) );
  CLKNAND2HSV0 U10378 ( .A1(n8257), .A2(n8256), .ZN(n8258) );
  NAND2HSV0 U10379 ( .A1(n6181), .A2(\pe4/got [3]), .ZN(n8260) );
  CLKNAND2HSV0 U10380 ( .A1(n8260), .A2(n8259), .ZN(n8261) );
  NAND2HSV0 U10381 ( .A1(\pe4/got [4]), .A2(n6706), .ZN(n8263) );
  CLKNAND2HSV0 U10382 ( .A1(n8263), .A2(n8262), .ZN(n8264) );
  OAI21HSV0 U10383 ( .A1(n8262), .A2(n8263), .B(n8264), .ZN(\pe4/poht [4]) );
  NOR2HSV0 U10384 ( .A1(n10355), .A2(n12172), .ZN(n8265) );
  NOR2HSV0 U10385 ( .A1(n13693), .A2(n13692), .ZN(n8266) );
  AOI21HSV0 U10386 ( .A1(\pe20/got [2]), .A2(n13695), .B(n13694), .ZN(n8267)
         );
  AOI21HSV0 U10387 ( .A1(n13695), .A2(n8266), .B(n8267), .ZN(n8268) );
  NAND2HSV0 U10388 ( .A1(\pe20/got [4]), .A2(n6731), .ZN(n8269) );
  OAI21HSV0 U10389 ( .A1(n8270), .A2(n8271), .B(n8272), .ZN(\pe20/poht [3]) );
  CLKNHSV0 U10390 ( .I(n11565), .ZN(n8273) );
  NAND2HSV0 U10391 ( .A1(\pe8/aot [5]), .A2(\pe8/bq[6] ), .ZN(n8274) );
  AOI22HSV2 U10392 ( .A1(n11564), .A2(n8273), .B1(n11566), .B2(n8274), .ZN(
        n11569) );
  NAND2HSV0 U10393 ( .A1(n12476), .A2(\pe3/aot [4]), .ZN(n8275) );
  NAND2HSV0 U10394 ( .A1(\pe3/got [4]), .A2(n12475), .ZN(n8276) );
  NAND2HSV2 U10395 ( .A1(n8276), .A2(n8275), .ZN(n8277) );
  OAI21HSV2 U10396 ( .A1(n8275), .A2(n8276), .B(n8277), .ZN(n10205) );
  INAND2HSV0 U10397 ( .A1(\pe7/ti_7t [3]), .B1(n12311), .ZN(n12206) );
  NAND2HSV0 U10398 ( .A1(\pe4/aot [8]), .A2(\pe4/bq[5] ), .ZN(n8278) );
  NAND2HSV0 U10399 ( .A1(\pe4/aot [5]), .A2(\pe4/bq[8] ), .ZN(n8279) );
  NAND2HSV0 U10400 ( .A1(n8279), .A2(n8278), .ZN(n8280) );
  NAND2HSV0 U10401 ( .A1(\pe4/aot [6]), .A2(\pe4/bq[7] ), .ZN(n8281) );
  INAND2HSV0 U10402 ( .A1(\pe16/ti_7t [5]), .B1(n8957), .ZN(n11182) );
  NOR2HSV0 U10403 ( .A1(n14401), .A2(n14400), .ZN(n8282) );
  NAND2HSV0 U10404 ( .A1(\pe17/got [3]), .A2(n14399), .ZN(n8283) );
  NAND2HSV2 U10405 ( .A1(n8283), .A2(n8282), .ZN(n8284) );
  OAI21HSV2 U10406 ( .A1(n8282), .A2(n8283), .B(n8284), .ZN(n14424) );
  NAND2HSV0 U10407 ( .A1(\pe11/bq[3] ), .A2(\pe11/aot [4]), .ZN(n8285) );
  NAND2HSV0 U10408 ( .A1(\pe11/bq[4] ), .A2(\pe11/aot [3]), .ZN(n8286) );
  CLKNAND2HSV0 U10409 ( .A1(n8286), .A2(n8285), .ZN(n8287) );
  OAI21HSV0 U10410 ( .A1(n8285), .A2(n8286), .B(n8287), .ZN(n8288) );
  CLKNHSV0 U10411 ( .I(n14370), .ZN(n8289) );
  AOI22HSV0 U10412 ( .A1(n12562), .A2(\pe11/aot [1]), .B1(\pe11/aot [2]), .B2(
        \pe11/bq[5] ), .ZN(n8290) );
  AOI21HSV0 U10413 ( .A1(n12563), .A2(n8289), .B(n8290), .ZN(n8291) );
  CLKNAND2HSV0 U10414 ( .A1(n8291), .A2(n8288), .ZN(n8292) );
  OAI21HSV0 U10415 ( .A1(n8291), .A2(n8288), .B(n8292), .ZN(n8293) );
  NAND2HSV0 U10416 ( .A1(\pe11/bq[1] ), .A2(\pe11/aot [6]), .ZN(n8294) );
  CLKNAND2HSV0 U10417 ( .A1(n8294), .A2(n8293), .ZN(n8295) );
  OAI21HSV0 U10418 ( .A1(n8293), .A2(n8294), .B(n8295), .ZN(n8296) );
  NAND2HSV0 U10419 ( .A1(\pe11/bq[2] ), .A2(\pe11/aot [5]), .ZN(n8297) );
  CLKNAND2HSV0 U10420 ( .A1(n8297), .A2(n8296), .ZN(n8298) );
  OAI21HSV0 U10421 ( .A1(n8296), .A2(n8297), .B(n8298), .ZN(n8299) );
  NAND2HSV0 U10422 ( .A1(\pe11/got [1]), .A2(n12561), .ZN(n8300) );
  NAND2HSV0 U10423 ( .A1(n8300), .A2(n8299), .ZN(n8301) );
  OAI21HSV0 U10424 ( .A1(n8299), .A2(n8300), .B(n8301), .ZN(n12564) );
  CLKNHSV0 U10425 ( .I(\pe6/phq [1]), .ZN(n8302) );
  MUX2NHSV2 U10426 ( .I0(\pe6/phq [1]), .I1(n8302), .S(n8303), .ZN(n11949) );
  AOI21HSV0 U10427 ( .A1(n10939), .A2(n10943), .B(n10201), .ZN(n8304) );
  CLKNAND2HSV0 U10428 ( .A1(n8942), .A2(\pe20/ti_7t [1]), .ZN(n9062) );
  NAND2HSV0 U10429 ( .A1(\pe15/aot [3]), .A2(\pe15/bq[3] ), .ZN(n8305) );
  NAND2HSV0 U10430 ( .A1(\pe15/bq[1] ), .A2(\pe15/aot [5]), .ZN(n8306) );
  NAND2HSV0 U10431 ( .A1(n8306), .A2(n8305), .ZN(n8307) );
  OAI21HSV2 U10432 ( .A1(n8305), .A2(n8306), .B(n8307), .ZN(n12620) );
  CLKNHSV0 U10433 ( .I(n15087), .ZN(n8308) );
  CLKNHSV0 U10434 ( .I(n14818), .ZN(n8310) );
  NOR2HSV2 U10435 ( .A1(n14740), .A2(n14010), .ZN(n8311) );
  CLKNAND2HSV2 U10436 ( .A1(n8311), .A2(n12038), .ZN(n13874) );
  AOI21HSV0 U10437 ( .A1(n13931), .A2(n14866), .B(n13930), .ZN(n8312) );
  XOR2HSV0 U10438 ( .A1(n13929), .A2(n13928), .Z(n8313) );
  NAND2HSV0 U10439 ( .A1(n10443), .A2(\pe9/got [3]), .ZN(n8314) );
  CLKNAND2HSV0 U10440 ( .A1(n8314), .A2(n8313), .ZN(n8315) );
  OAI21HSV0 U10441 ( .A1(n8313), .A2(n8314), .B(n8315), .ZN(n8316) );
  NAND2HSV0 U10442 ( .A1(n13910), .A2(\pe9/got [4]), .ZN(n8317) );
  CLKNAND2HSV0 U10443 ( .A1(n8317), .A2(n8316), .ZN(n8318) );
  OAI21HSV0 U10444 ( .A1(n8316), .A2(n8317), .B(n8318), .ZN(n8319) );
  NAND2HSV0 U10445 ( .A1(n14963), .A2(\pe9/got [5]), .ZN(n8320) );
  CLKNAND2HSV0 U10446 ( .A1(n8320), .A2(n8319), .ZN(n8321) );
  OAI21HSV0 U10447 ( .A1(n8319), .A2(n8320), .B(n8321), .ZN(n8322) );
  OAI21HSV0 U10448 ( .A1(n14866), .A2(n6737), .B(n8312), .ZN(n8323) );
  CLKNAND2HSV0 U10449 ( .A1(n8323), .A2(n8322), .ZN(n8324) );
  NAND2HSV0 U10450 ( .A1(n9434), .A2(n7875), .ZN(n8326) );
  OAI21HSV0 U10451 ( .A1(n8325), .A2(n8326), .B(n8327), .ZN(\pe9/poht [1]) );
  NAND2HSV0 U10452 ( .A1(\pe6/ti_7[5] ), .A2(\pe6/got [6]), .ZN(n8329) );
  CLKNAND2HSV0 U10453 ( .A1(n8329), .A2(n8328), .ZN(n8330) );
  OAI21HSV0 U10454 ( .A1(n8331), .A2(n8332), .B(n8333), .ZN(po6) );
  AOI21HSV0 U10455 ( .A1(n15075), .A2(\pe10/got [8]), .B(n14828), .ZN(n8335)
         );
  CLKNHSV0 U10456 ( .I(n11523), .ZN(n8336) );
  CLKNHSV0 U10457 ( .I(\pe12/got [5]), .ZN(n8338) );
  NAND2HSV0 U10458 ( .A1(n14255), .A2(\pe12/got [2]), .ZN(n8339) );
  CLKNAND2HSV0 U10459 ( .A1(n8339), .A2(n14256), .ZN(n8340) );
  OAI21HSV0 U10460 ( .A1(n14256), .A2(n8339), .B(n8340), .ZN(n8341) );
  NAND2HSV0 U10461 ( .A1(n15190), .A2(\pe12/got [6]), .ZN(n8343) );
  NAND2HSV0 U10462 ( .A1(n14959), .A2(\pe12/got [7]), .ZN(n8346) );
  OAI21HSV0 U10463 ( .A1(n8345), .A2(n8346), .B(n8347), .ZN(\pe12/poht [1]) );
  OAI21HSV0 U10464 ( .A1(n12645), .A2(n10536), .B(n8348), .ZN(n8349) );
  AO31HSV2 U10465 ( .A1(\pe4/got [5]), .A2(n12631), .A3(n8350), .B(n8351), .Z(
        n8352) );
  NAND2HSV0 U10466 ( .A1(n12079), .A2(\pe4/got [6]), .ZN(n8353) );
  CLKNAND2HSV0 U10467 ( .A1(n8353), .A2(n8352), .ZN(n8354) );
  NAND2HSV0 U10468 ( .A1(n6181), .A2(\pe4/got [7]), .ZN(n8356) );
  CLKNAND2HSV0 U10469 ( .A1(n8356), .A2(n8355), .ZN(n8357) );
  NAND2HSV0 U10470 ( .A1(\pe4/got [8]), .A2(n6706), .ZN(n8359) );
  CLKNAND2HSV0 U10471 ( .A1(n8359), .A2(n8358), .ZN(n8360) );
  OAI21HSV0 U10472 ( .A1(n8358), .A2(n8359), .B(n8360), .ZN(po4) );
  XOR2HSV0 U10473 ( .A1(n13680), .A2(n13679), .Z(n8361) );
  NAND2HSV0 U10474 ( .A1(\pe20/aot [3]), .A2(\pe20/bq[1] ), .ZN(n8362) );
  CLKNAND2HSV0 U10475 ( .A1(n8362), .A2(n8361), .ZN(n8363) );
  OAI21HSV0 U10476 ( .A1(n8361), .A2(n8362), .B(n8363), .ZN(n8364) );
  CLKNAND2HSV0 U10477 ( .A1(n8365), .A2(n8364), .ZN(n8366) );
  OAI21HSV0 U10478 ( .A1(n8364), .A2(n8365), .B(n8366), .ZN(n8367) );
  NAND2HSV0 U10479 ( .A1(\pe20/ti_7[5] ), .A2(\pe20/got [1]), .ZN(n8368) );
  CLKNAND2HSV0 U10480 ( .A1(n8368), .A2(n8367), .ZN(n8369) );
  OAI21HSV0 U10481 ( .A1(n8370), .A2(n8371), .B(n8372), .ZN(\pe20/poht [5]) );
  AO22HSV2 U10482 ( .A1(\pe19/bq[5] ), .A2(n13317), .B1(\pe19/bq[2] ), .B2(
        n14915), .Z(n8373) );
  OAI21HSV2 U10483 ( .A1(n12152), .A2(n14224), .B(n8373), .ZN(n12153) );
  CLKNHSV0 U10484 ( .I(n14000), .ZN(n8374) );
  OAI21HSV0 U10485 ( .A1(n10616), .A2(n14539), .B(n8374), .ZN(n10617) );
  CLKNHSV0 U10486 ( .I(n9248), .ZN(n8375) );
  CLKNHSV0 U10487 ( .I(n9798), .ZN(n8376) );
  CLKNHSV0 U10488 ( .I(\pe8/bq[3] ), .ZN(n8377) );
  OAI21HSV0 U10489 ( .A1(n14207), .A2(n8377), .B(n14206), .ZN(n8378) );
  OAI21HSV0 U10490 ( .A1(n14209), .A2(n14208), .B(n8378), .ZN(n14210) );
  NAND2HSV0 U10491 ( .A1(\pe21/aot [4]), .A2(\pe21/bq[3] ), .ZN(n8379) );
  CLKNAND2HSV0 U10492 ( .A1(n8379), .A2(n10883), .ZN(n8380) );
  OAI21HSV0 U10493 ( .A1(n10883), .A2(n8379), .B(n8380), .ZN(n8381) );
  XOR2HSV0 U10494 ( .A1(n10882), .A2(n10881), .Z(n8382) );
  XOR2HSV0 U10495 ( .A1(n8381), .A2(n8382), .Z(n8383) );
  CLKNAND2HSV0 U10496 ( .A1(n8384), .A2(n8383), .ZN(n8385) );
  OAI21HSV0 U10497 ( .A1(n8383), .A2(n8384), .B(n8385), .ZN(n8386) );
  NAND2HSV0 U10498 ( .A1(\pe21/ti_7[3] ), .A2(\pe21/got [2]), .ZN(n8387) );
  CLKNAND2HSV0 U10499 ( .A1(n8387), .A2(n8386), .ZN(n8388) );
  OAI21HSV0 U10500 ( .A1(n8386), .A2(n8387), .B(n8388), .ZN(n8389) );
  NAND2HSV0 U10501 ( .A1(n15175), .A2(\pe21/got [3]), .ZN(n8390) );
  CLKNAND2HSV0 U10502 ( .A1(n8390), .A2(n8389), .ZN(n8391) );
  OAI21HSV0 U10503 ( .A1(n8389), .A2(n8390), .B(n8391), .ZN(n8392) );
  OAI21HSV2 U10504 ( .A1(n8392), .A2(n8393), .B(n8394), .ZN(n10884) );
  INAND3HSV2 U10505 ( .A1(n13884), .B1(n10601), .B2(n10602), .ZN(n8395) );
  NAND2HSV0 U10506 ( .A1(n10603), .A2(\pe1/got [8]), .ZN(n8396) );
  CLKNAND2HSV0 U10507 ( .A1(ctro3), .A2(\pe3/ti_7t [1]), .ZN(n10213) );
  NAND3HSV2 U10508 ( .A1(n10583), .A2(n10584), .A3(n11284), .ZN(n10588) );
  IOA21HSV2 U10509 ( .A1(\pe6/aot [4]), .A2(\pe6/bq[3] ), .B(n12936), .ZN(
        n8397) );
  OAI21HSV0 U10510 ( .A1(n13048), .A2(n12999), .B(n8397), .ZN(n8398) );
  AO22HSV2 U10511 ( .A1(\pe6/aot [1]), .A2(n13827), .B1(\pe6/bq[4] ), .B2(
        \pe6/aot [3]), .Z(n8399) );
  OAI21HSV2 U10512 ( .A1(n13000), .A2(n13049), .B(n8399), .ZN(n8400) );
  NAND2HSV2 U10513 ( .A1(n8400), .A2(n8398), .ZN(n8401) );
  OAI21HSV2 U10514 ( .A1(n8400), .A2(n8398), .B(n8401), .ZN(n8402) );
  NAND2HSV0 U10515 ( .A1(\pe6/bq[2] ), .A2(\pe6/aot [5]), .ZN(n8403) );
  NAND2HSV2 U10516 ( .A1(n8403), .A2(n8402), .ZN(n8404) );
  OAI21HSV2 U10517 ( .A1(n8402), .A2(n8403), .B(n8404), .ZN(n8405) );
  NAND2HSV0 U10518 ( .A1(\pe6/bq[1] ), .A2(\pe6/aot [6]), .ZN(n8406) );
  NAND2HSV2 U10519 ( .A1(n8406), .A2(n8405), .ZN(n8407) );
  OAI21HSV2 U10520 ( .A1(n8405), .A2(n8406), .B(n8407), .ZN(n12937) );
  CLKNAND2HSV4 U10521 ( .A1(n15168), .A2(n8408), .ZN(n14681) );
  NAND2HSV0 U10522 ( .A1(\pe14/got [3]), .A2(n15195), .ZN(n8411) );
  CLKNAND2HSV0 U10523 ( .A1(n8411), .A2(n8410), .ZN(n8412) );
  OAI21HSV0 U10524 ( .A1(n8410), .A2(n8411), .B(n8412), .ZN(n8413) );
  NAND2HSV0 U10525 ( .A1(\pe14/got [5]), .A2(n13086), .ZN(n8415) );
  CLKNAND2HSV0 U10526 ( .A1(n8415), .A2(n8414), .ZN(n8416) );
  OAI21HSV0 U10527 ( .A1(n8418), .A2(n8417), .B(n8419), .ZN(\pe14/poht [2]) );
  XOR2HSV0 U10528 ( .A1(n12510), .A2(n12509), .Z(n8420) );
  OAI21HSV0 U10529 ( .A1(n13100), .A2(n13761), .B(n8420), .ZN(n8421) );
  NAND2HSV0 U10530 ( .A1(\pe2/ti_7[5] ), .A2(\pe2/got [4]), .ZN(n8423) );
  NAND2HSV2 U10531 ( .A1(n8423), .A2(n8422), .ZN(n8424) );
  OAI21HSV2 U10532 ( .A1(n8422), .A2(n8423), .B(n8424), .ZN(n8425) );
  AND2HSV2 U10533 ( .A1(\pe9/ti_7t [7]), .A2(n9790), .Z(n8428) );
  AOI211HSV0 U10534 ( .A1(n9790), .A2(\pe9/ti_7t [7]), .B(n9792), .C(n9793), 
        .ZN(n8429) );
  XOR2HSV0 U10535 ( .A1(n13335), .A2(n13334), .Z(n8431) );
  NAND2HSV0 U10536 ( .A1(\pe19/got [4]), .A2(n14219), .ZN(n8432) );
  CLKNAND2HSV0 U10537 ( .A1(n8432), .A2(n8431), .ZN(n8433) );
  OAI21HSV0 U10538 ( .A1(n8431), .A2(n8432), .B(n8433), .ZN(n8434) );
  CLKNHSV0 U10539 ( .I(n13336), .ZN(n8435) );
  XOR2HSV0 U10540 ( .A1(n13033), .A2(n13032), .Z(n8436) );
  AOI21HSV0 U10541 ( .A1(\pe5/got [2]), .A2(n14952), .B(n8436), .ZN(n8437) );
  AO31HSV2 U10542 ( .A1(\pe5/got [2]), .A2(n14952), .A3(n8436), .B(n8437), .Z(
        n8438) );
  NAND2HSV0 U10543 ( .A1(\pe5/got [3]), .A2(n14916), .ZN(n8439) );
  CLKNAND2HSV0 U10544 ( .A1(n8439), .A2(n8438), .ZN(n8440) );
  OAI21HSV0 U10545 ( .A1(n8438), .A2(n8439), .B(n8440), .ZN(n8441) );
  NAND2HSV0 U10546 ( .A1(\pe5/got [4]), .A2(n6922), .ZN(n8442) );
  CLKNAND2HSV0 U10547 ( .A1(n8442), .A2(n8441), .ZN(n8443) );
  OAI21HSV0 U10548 ( .A1(n8441), .A2(n8442), .B(n8443), .ZN(n8444) );
  NAND2HSV0 U10549 ( .A1(\pe5/got [5]), .A2(n14846), .ZN(n8445) );
  NAND2HSV0 U10550 ( .A1(n8445), .A2(n8444), .ZN(n8446) );
  OAI21HSV0 U10551 ( .A1(n8444), .A2(n8445), .B(n8446), .ZN(n8447) );
  OAI21HSV0 U10552 ( .A1(n13809), .A2(n13280), .B(n8447), .ZN(n8448) );
  OAI31HSV0 U10553 ( .A1(n8447), .A2(n13809), .A3(n13280), .B(n8448), .ZN(
        n8449) );
  NAND2HSV0 U10554 ( .A1(\pe5/got [7]), .A2(\pe5/ti_7[7] ), .ZN(n8450) );
  CLKNAND2HSV0 U10555 ( .A1(n8450), .A2(n8449), .ZN(n8451) );
  OAI21HSV0 U10556 ( .A1(n8450), .A2(n8449), .B(n8451), .ZN(\pe5/poht [1]) );
  NAND2HSV0 U10557 ( .A1(\pe21/bq[8] ), .A2(\pe21/aot [3]), .ZN(n8452) );
  NAND2HSV0 U10558 ( .A1(\pe21/aot [7]), .A2(\pe21/bq[4] ), .ZN(n8453) );
  NAND2HSV0 U10559 ( .A1(n8453), .A2(n8452), .ZN(n8454) );
  OAI21HSV0 U10560 ( .A1(n8452), .A2(n8453), .B(n8454), .ZN(n10819) );
  AOI21HSV2 U10561 ( .A1(n14951), .A2(n8456), .B(n10051), .ZN(n10032) );
  CLKNAND2HSV0 U10562 ( .A1(\pe2/pvq [7]), .A2(n14558), .ZN(n8457) );
  NAND2HSV2 U10563 ( .A1(n8457), .A2(\pe2/phq [7]), .ZN(n8458) );
  OAI21HSV2 U10564 ( .A1(\pe2/phq [7]), .A2(n8457), .B(n8458), .ZN(n11247) );
  CLKNHSV0 U10565 ( .I(\pe19/bq[7] ), .ZN(n8459) );
  NAND2HSV0 U10566 ( .A1(\pe19/aot [7]), .A2(\pe19/bq[5] ), .ZN(n8460) );
  OAI21HSV0 U10567 ( .A1(n15099), .A2(n8459), .B(n8460), .ZN(n8461) );
  OAI31HSV2 U10568 ( .A1(n15099), .A2(n8460), .A3(n8459), .B(n8461), .ZN(n9552) );
  NAND2HSV0 U10569 ( .A1(n14949), .A2(\pe17/bq[5] ), .ZN(n8465) );
  NAND2HSV0 U10570 ( .A1(\pe14/bq[7] ), .A2(\pe14/aot [8]), .ZN(n8467) );
  OAI21HSV2 U10571 ( .A1(n8466), .A2(n8467), .B(n8468), .ZN(n9095) );
  NAND2HSV0 U10572 ( .A1(\pe13/pvq [6]), .A2(n14552), .ZN(n8469) );
  NAND2HSV2 U10573 ( .A1(n8469), .A2(\pe13/phq [6]), .ZN(n8470) );
  AOI22HSV0 U10574 ( .A1(\pe2/aot [1]), .A2(\pe2/bq[5] ), .B1(\pe2/aot [3]), 
        .B2(\pe2/bq[3] ), .ZN(n8471) );
  IAO21HSV2 U10575 ( .A1(n13093), .A2(n13092), .B(n8471), .ZN(n13097) );
  INOR2HSV0 U10576 ( .A1(\pe1/ti_7t [6]), .B1(n10228), .ZN(n10603) );
  NOR2HSV0 U10577 ( .A1(n8472), .A2(n13338), .ZN(n8473) );
  AOI211HSV1 U10578 ( .A1(n8472), .A2(n13338), .B(n13801), .C(n8473), .ZN(
        n8474) );
  XOR2HSV0 U10579 ( .A1(n13528), .A2(n13530), .Z(n8476) );
  NAND2HSV0 U10580 ( .A1(n14857), .A2(\pe8/got [4]), .ZN(n8478) );
  CLKNAND2HSV0 U10581 ( .A1(n8478), .A2(n8477), .ZN(n8479) );
  OAI21HSV0 U10582 ( .A1(n8477), .A2(n8478), .B(n8479), .ZN(n8480) );
  NAND2HSV0 U10583 ( .A1(n15066), .A2(\pe8/got [5]), .ZN(n8481) );
  CLKNAND2HSV0 U10584 ( .A1(n8481), .A2(n8480), .ZN(n8482) );
  OAI21HSV0 U10585 ( .A1(n8480), .A2(n8481), .B(n8482), .ZN(n8483) );
  NAND2HSV0 U10586 ( .A1(n14893), .A2(\pe8/got [6]), .ZN(n8484) );
  CLKNAND2HSV0 U10587 ( .A1(n8484), .A2(n8483), .ZN(n8485) );
  OAI21HSV0 U10588 ( .A1(n8483), .A2(n8484), .B(n8485), .ZN(n8486) );
  NAND2HSV0 U10589 ( .A1(n15182), .A2(\pe8/got [7]), .ZN(n8487) );
  CLKNAND2HSV0 U10590 ( .A1(n8487), .A2(n8486), .ZN(n8488) );
  OAI21HSV0 U10591 ( .A1(n8486), .A2(n8487), .B(n8488), .ZN(n8489) );
  NAND2HSV0 U10592 ( .A1(\pe8/got [8]), .A2(n15091), .ZN(n8490) );
  CLKNAND2HSV0 U10593 ( .A1(n8490), .A2(n8489), .ZN(n8491) );
  OAI21HSV0 U10594 ( .A1(n8489), .A2(n8490), .B(n8491), .ZN(po8) );
  XOR2HSV0 U10595 ( .A1(n13785), .A2(n13784), .Z(n8492) );
  OAI21HSV0 U10596 ( .A1(n13760), .A2(n13761), .B(n8492), .ZN(n8493) );
  OAI31HSV0 U10597 ( .A1(n13760), .A2(n8492), .A3(n13761), .B(n8493), .ZN(
        n8494) );
  AOI21HSV0 U10598 ( .A1(n6721), .A2(n14935), .B(n8494), .ZN(n8495) );
  AO31HSV2 U10599 ( .A1(n6721), .A2(n14935), .A3(n8494), .B(n8495), .Z(n8496)
         );
  NAND2HSV0 U10600 ( .A1(n14822), .A2(\pe2/ti_7[5] ), .ZN(n8498) );
  OAI21HSV2 U10601 ( .A1(n8497), .A2(n8498), .B(n8499), .ZN(n8500) );
  NAND2HSV0 U10602 ( .A1(n14061), .A2(n14818), .ZN(n8501) );
  OAI21HSV0 U10603 ( .A1(n8500), .A2(n8501), .B(n8502), .ZN(po2) );
  CLKNHSV0 U10604 ( .I(n11174), .ZN(n8503) );
  AOI21HSV0 U10605 ( .A1(n11897), .A2(n11948), .B(n11745), .ZN(n8504) );
  NOR2HSV0 U10606 ( .A1(n10260), .A2(n10255), .ZN(n8509) );
  NAND2HSV2 U10607 ( .A1(n8509), .A2(n10264), .ZN(n8510) );
  XOR2HSV0 U10608 ( .A1(n14226), .A2(n14225), .Z(n8511) );
  AOI21HSV0 U10609 ( .A1(\pe19/got [2]), .A2(n12148), .B(n8511), .ZN(n8512) );
  AO31HSV2 U10610 ( .A1(\pe19/got [2]), .A2(n12148), .A3(n8511), .B(n8512), 
        .Z(n8513) );
  NAND2HSV0 U10611 ( .A1(n14862), .A2(\pe19/got [6]), .ZN(n8515) );
  CLKNAND2HSV0 U10612 ( .A1(n8515), .A2(n8514), .ZN(n8516) );
  OAI21HSV0 U10613 ( .A1(n8514), .A2(n8515), .B(n8516), .ZN(\pe19/poht [2]) );
  NAND2HSV0 U10614 ( .A1(\pe7/bq[3] ), .A2(\pe7/aot [1]), .ZN(n8517) );
  AOI21HSV0 U10615 ( .A1(\pe7/bq[2] ), .A2(\pe7/aot [2]), .B(n8517), .ZN(n8518) );
  AO31HSV2 U10616 ( .A1(\pe7/bq[2] ), .A2(\pe7/aot [2]), .A3(n8517), .B(n8518), 
        .Z(n8519) );
  NAND2HSV0 U10617 ( .A1(\pe7/bq[1] ), .A2(\pe7/aot [3]), .ZN(n8520) );
  CLKNAND2HSV0 U10618 ( .A1(n8520), .A2(n8519), .ZN(n8521) );
  OAI21HSV0 U10619 ( .A1(n8519), .A2(n8520), .B(n8521), .ZN(n8522) );
  CLKNAND2HSV0 U10620 ( .A1(n8523), .A2(n8522), .ZN(n8524) );
  OAI21HSV0 U10621 ( .A1(n8522), .A2(n8523), .B(n8524), .ZN(n8525) );
  NAND2HSV0 U10622 ( .A1(\pe7/got [2]), .A2(n14487), .ZN(n8526) );
  CLKNAND2HSV0 U10623 ( .A1(n8525), .A2(n8526), .ZN(n8527) );
  OAI21HSV0 U10624 ( .A1(n8525), .A2(n8526), .B(n8527), .ZN(n8528) );
  NAND2HSV0 U10625 ( .A1(n13605), .A2(\pe7/got [3]), .ZN(n8529) );
  NAND2HSV0 U10626 ( .A1(n8529), .A2(n8528), .ZN(n8530) );
  OAI21HSV0 U10627 ( .A1(n8528), .A2(n8529), .B(n8530), .ZN(\pe7/poht [5]) );
  CLKNHSV0 U10628 ( .I(\pe5/got [4]), .ZN(n8531) );
  XOR2HSV0 U10629 ( .A1(n13392), .A2(n13393), .Z(n8532) );
  NAND2HSV0 U10630 ( .A1(\pe5/got [2]), .A2(n12780), .ZN(n8534) );
  OAI21HSV2 U10631 ( .A1(n8533), .A2(n8534), .B(n8535), .ZN(n8536) );
  NAND2HSV0 U10632 ( .A1(n8537), .A2(n8536), .ZN(n8538) );
  OAI21HSV0 U10633 ( .A1(n8536), .A2(n8537), .B(n8538), .ZN(n8539) );
  OAI21HSV0 U10634 ( .A1(n13401), .A2(n8531), .B(n8539), .ZN(n8540) );
  OAI31HSV0 U10635 ( .A1(n13401), .A2(n8539), .A3(n8531), .B(n8540), .ZN(n8541) );
  NAND2HSV0 U10636 ( .A1(\pe5/ti_7[7] ), .A2(\pe5/got [5]), .ZN(n8542) );
  CLKNAND2HSV0 U10637 ( .A1(n8542), .A2(n8541), .ZN(n8543) );
  OAI21HSV0 U10638 ( .A1(n8541), .A2(n8542), .B(n8543), .ZN(\pe5/poht [3]) );
  AOI22HSV0 U10639 ( .A1(\pe21/bq[4] ), .A2(\pe21/aot [6]), .B1(\pe21/aot [8]), 
        .B2(\pe21/bq[2] ), .ZN(n8545) );
  NAND2HSV0 U10640 ( .A1(\pe3/ctrq ), .A2(\pe3/pvq [6]), .ZN(n8546) );
  NAND2HSV2 U10641 ( .A1(n8546), .A2(\pe3/phq [6]), .ZN(n8547) );
  OAI21HSV2 U10642 ( .A1(\pe3/phq [6]), .A2(n8546), .B(n8547), .ZN(n10952) );
  NAND2HSV0 U10643 ( .A1(\pe16/bq[5] ), .A2(\pe16/aot [8]), .ZN(n8549) );
  CLKNHSV0 U10644 ( .I(\pe9/bq[5] ), .ZN(n8550) );
  IOA22HSV1 U10645 ( .B1(n9438), .B2(n8550), .A1(n14942), .A2(\pe9/bq[4] ), 
        .ZN(n9439) );
  CLKNHSV0 U10646 ( .I(n11316), .ZN(n8551) );
  AOI21HSV0 U10647 ( .A1(n11316), .A2(n12320), .B(n14584), .ZN(n8552) );
  OAI21HSV4 U10648 ( .A1(n15235), .A2(n8551), .B(n8552), .ZN(n11318) );
  NAND2HSV2 U10649 ( .A1(n8553), .A2(\pe2/phq [4]), .ZN(n8554) );
  NAND2HSV0 U10650 ( .A1(\pe2/aot [5]), .A2(\pe2/bq[8] ), .ZN(n8555) );
  AOI22HSV0 U10651 ( .A1(\pe8/aot [1]), .A2(\pe8/bq[5] ), .B1(\pe8/bq[4] ), 
        .B2(\pe8/aot [2]), .ZN(n8556) );
  IAO21HSV2 U10652 ( .A1(n14206), .A2(n14203), .B(n8556), .ZN(n13542) );
  CLKNHSV0 U10653 ( .I(\pe4/phq [1]), .ZN(n8557) );
  NAND2HSV2 U10654 ( .A1(\pe4/aot [8]), .A2(\pe4/bq[8] ), .ZN(n8558) );
  MUX2NHSV4 U10655 ( .I0(\pe4/phq [1]), .I1(n8557), .S(n8558), .ZN(n9611) );
  NAND2HSV0 U10656 ( .A1(\pe3/aot [3]), .A2(\pe3/bq[3] ), .ZN(n8559) );
  CLKNAND2HSV0 U10657 ( .A1(n8559), .A2(n12980), .ZN(n8560) );
  OAI21HSV0 U10658 ( .A1(n12980), .A2(n8559), .B(n8560), .ZN(n8561) );
  XOR2HSV0 U10659 ( .A1(n12979), .A2(n8561), .Z(n8562) );
  NAND2HSV0 U10660 ( .A1(n14820), .A2(\pe3/got [1]), .ZN(n8563) );
  CLKNAND2HSV0 U10661 ( .A1(n8563), .A2(n8562), .ZN(n8564) );
  OAI21HSV0 U10662 ( .A1(n8562), .A2(n8563), .B(n8564), .ZN(n8565) );
  NAND2HSV0 U10663 ( .A1(n14941), .A2(\pe3/got [4]), .ZN(n8570) );
  OAI21HSV0 U10664 ( .A1(n8569), .A2(n8570), .B(n8571), .ZN(n8572) );
  NAND2HSV0 U10665 ( .A1(\pe3/got [5]), .A2(n14819), .ZN(n8573) );
  OAI21HSV0 U10666 ( .A1(n8572), .A2(n8573), .B(n8574), .ZN(\pe3/poht [3]) );
  NAND2HSV0 U10667 ( .A1(\pe15/bq[3] ), .A2(\pe15/aot [1]), .ZN(n8575) );
  AOI21HSV0 U10668 ( .A1(\pe15/aot [3]), .A2(\pe15/bq[1] ), .B(n8575), .ZN(
        n8576) );
  AO31HSV2 U10669 ( .A1(\pe15/aot [3]), .A2(\pe15/bq[1] ), .A3(n8575), .B(
        n8576), .Z(n8577) );
  NAND2HSV0 U10670 ( .A1(\pe15/aot [2]), .A2(\pe15/bq[2] ), .ZN(n8578) );
  CLKNAND2HSV0 U10671 ( .A1(n8578), .A2(n8577), .ZN(n8579) );
  OAI21HSV0 U10672 ( .A1(n8577), .A2(n8578), .B(n8579), .ZN(n8580) );
  NAND2HSV0 U10673 ( .A1(\pe15/ti_7[5] ), .A2(\pe15/got [1]), .ZN(n8582) );
  NAND2HSV0 U10674 ( .A1(n8585), .A2(n8584), .ZN(n8586) );
  OAI21HSV0 U10675 ( .A1(n8584), .A2(n8585), .B(n8586), .ZN(\pe15/poht [5]) );
  XOR2HSV0 U10676 ( .A1(n14485), .A2(n14486), .Z(n8587) );
  XOR2HSV0 U10677 ( .A1(n14467), .A2(n14466), .Z(n8588) );
  XOR2HSV0 U10678 ( .A1(n8587), .A2(n8588), .Z(n8589) );
  OAI21HSV0 U10679 ( .A1(n14465), .A2(n14464), .B(n8589), .ZN(n8590) );
  AO31HSV2 U10680 ( .A1(n15081), .A2(n8591), .A3(\pe7/got [5]), .B(n8592), .Z(
        n8593) );
  NAND2HSV0 U10681 ( .A1(\pe7/ti_7[5] ), .A2(\pe7/got [6]), .ZN(n8594) );
  CLKNAND2HSV0 U10682 ( .A1(n8594), .A2(n8593), .ZN(n8595) );
  NAND2HSV0 U10683 ( .A1(n14829), .A2(n14487), .ZN(n8597) );
  CLKNAND2HSV0 U10684 ( .A1(n8597), .A2(n8596), .ZN(n8598) );
  OAI21HSV0 U10685 ( .A1(n8596), .A2(n8597), .B(n8598), .ZN(n8599) );
  NAND2HSV0 U10686 ( .A1(n8600), .A2(n8599), .ZN(n8601) );
  OAI21HSV0 U10687 ( .A1(n8599), .A2(n8600), .B(n8601), .ZN(po7) );
  NAND2HSV0 U10688 ( .A1(\pe10/got [3]), .A2(n6033), .ZN(n8602) );
  CLKNAND2HSV0 U10689 ( .A1(n8602), .A2(n10105), .ZN(n8603) );
  NAND2HSV0 U10690 ( .A1(n14940), .A2(\pe10/got [4]), .ZN(n8605) );
  CLKNAND2HSV0 U10691 ( .A1(n8605), .A2(n8604), .ZN(n8606) );
  NAND3HSV0 U10692 ( .A1(n10110), .A2(n10109), .A3(n10108), .ZN(n8608) );
  CLKNHSV0 U10693 ( .I(n13258), .ZN(n8611) );
  MUX2NHSV1 U10694 ( .I0(n8612), .I1(n13257), .S(n13256), .ZN(n8613) );
  MUX2NHSV0 U10695 ( .I0(n8611), .I1(n13258), .S(n8613), .ZN(pov1[7]) );
  IOA21HSV2 U10696 ( .A1(n15258), .A2(n12353), .B(n12354), .ZN(n14366) );
  INOR2HSV0 U10697 ( .A1(n10588), .B1(n10587), .ZN(n8615) );
  XOR2HSV0 U10698 ( .A1(n12382), .A2(n12384), .Z(n8617) );
  XOR2HSV0 U10699 ( .A1(n12383), .A2(n8617), .Z(n8618) );
  AOI21HSV0 U10700 ( .A1(\pe19/got [1]), .A2(n12148), .B(n8618), .ZN(n8619) );
  AO31HSV2 U10701 ( .A1(\pe19/got [1]), .A2(n12148), .A3(n8618), .B(n8619), 
        .Z(n8620) );
  NAND2HSV0 U10702 ( .A1(n14219), .A2(\pe19/got [2]), .ZN(n8621) );
  CLKNAND2HSV0 U10703 ( .A1(n8621), .A2(n8620), .ZN(n8622) );
  OAI21HSV0 U10704 ( .A1(n8620), .A2(n8621), .B(n8622), .ZN(n8623) );
  NAND2HSV0 U10705 ( .A1(n13315), .A2(\pe19/got [5]), .ZN(n8628) );
  CLKNAND2HSV0 U10706 ( .A1(n8628), .A2(n8627), .ZN(n8629) );
  OAI21HSV0 U10707 ( .A1(n8627), .A2(n8628), .B(n8629), .ZN(\pe19/poht [3]) );
  CLKNHSV0 U10708 ( .I(\pe5/got [3]), .ZN(n8630) );
  XOR2HSV0 U10709 ( .A1(n13382), .A2(n13381), .Z(n8631) );
  XOR2HSV0 U10710 ( .A1(n13384), .A2(n8631), .Z(n8632) );
  NAND2HSV0 U10711 ( .A1(n12780), .A2(\pe5/got [1]), .ZN(n8633) );
  CLKNAND2HSV0 U10712 ( .A1(n8633), .A2(n8632), .ZN(n8634) );
  OAI21HSV0 U10713 ( .A1(n8632), .A2(n8633), .B(n8634), .ZN(n8635) );
  OAI21HSV0 U10714 ( .A1(n8636), .A2(n8637), .B(n8638), .ZN(\pe5/poht [4]) );
  MUX2HSV0 U10715 ( .I0(\pe7/pq ), .I1(n14480), .S(n12067), .Z(\pe7/ti_1t ) );
  AOI22HSV0 U10716 ( .A1(\pe21/bq[1] ), .A2(\pe21/aot [7]), .B1(\pe21/bq[3] ), 
        .B2(\pe21/aot [5]), .ZN(n8639) );
  IAO21HSV2 U10717 ( .A1(n12089), .A2(n12552), .B(n8639), .ZN(n12091) );
  INAND2HSV0 U10718 ( .A1(\pe4/ti_7t [3]), .B1(n9714), .ZN(n9644) );
  NOR2HSV0 U10719 ( .A1(n13238), .A2(n13270), .ZN(n8640) );
  NAND2HSV0 U10720 ( .A1(\pe17/bq[1] ), .A2(\pe17/aot [5]), .ZN(n8641) );
  AOI21HSV2 U10721 ( .A1(n8641), .A2(n14017), .B(n8640), .ZN(n13242) );
  AOI21HSV0 U10722 ( .A1(n14831), .A2(n11415), .B(n11442), .ZN(n8642) );
  INOR2HSV0 U10723 ( .A1(\pe10/ti_7t [6]), .B1(n10070), .ZN(n10930) );
  NAND2HSV0 U10724 ( .A1(n10853), .A2(n6208), .ZN(n8645) );
  NAND2HSV0 U10725 ( .A1(n8645), .A2(poh21[4]), .ZN(n8646) );
  OAI21HSV2 U10726 ( .A1(poh21[4]), .A2(n8645), .B(n8646), .ZN(po[5]) );
  NAND2HSV0 U10727 ( .A1(n11296), .A2(n15233), .ZN(n8647) );
  OAI21HSV2 U10728 ( .A1(n11292), .A2(n11296), .B(n8647), .ZN(\pe15/ti_7[3] )
         );
  NAND2HSV0 U10729 ( .A1(n12362), .A2(n14839), .ZN(n8648) );
  OAI21HSV0 U10730 ( .A1(\pe20/pq ), .A2(n12362), .B(n8648), .ZN(\pe20/ti_1t )
         );
  CLKNHSV0 U10731 ( .I(\pe15/got [2]), .ZN(n8649) );
  XOR2HSV0 U10732 ( .A1(n13234), .A2(n13235), .Z(n8650) );
  XOR2HSV0 U10733 ( .A1(n13233), .A2(n13232), .Z(n8651) );
  XOR2HSV0 U10734 ( .A1(n8650), .A2(n8651), .Z(n8652) );
  NAND2HSV0 U10735 ( .A1(n14708), .A2(\pe15/got [1]), .ZN(n8653) );
  CLKNAND2HSV0 U10736 ( .A1(n8653), .A2(n8652), .ZN(n8654) );
  OAI21HSV2 U10737 ( .A1(n8652), .A2(n8653), .B(n8654), .ZN(n8655) );
  OAI21HSV0 U10738 ( .A1(n8656), .A2(n8657), .B(n8658), .ZN(\pe15/poht [4]) );
  CLKNHSV0 U10739 ( .I(\pe11/got [1]), .ZN(n8659) );
  XOR2HSV0 U10740 ( .A1(n14395), .A2(n14394), .Z(n8660) );
  NAND2HSV0 U10741 ( .A1(\pe11/aot [3]), .A2(\pe11/bq[1] ), .ZN(n8661) );
  CLKNAND2HSV0 U10742 ( .A1(n8661), .A2(n8660), .ZN(n8662) );
  OAI21HSV0 U10743 ( .A1(n8660), .A2(n8661), .B(n8662), .ZN(n8663) );
  OAI21HSV0 U10744 ( .A1(n14396), .A2(n8659), .B(n8663), .ZN(n8664) );
  OAI31HSV0 U10745 ( .A1(n14396), .A2(n8663), .A3(n8659), .B(n8664), .ZN(n8665) );
  NAND2HSV0 U10746 ( .A1(n14830), .A2(\pe11/got [2]), .ZN(n8666) );
  CLKNAND2HSV0 U10747 ( .A1(n8666), .A2(n8665), .ZN(n8667) );
  OAI21HSV0 U10748 ( .A1(n8668), .A2(n8669), .B(n8670), .ZN(\pe11/poht [5]) );
  NAND2HSV0 U10749 ( .A1(n14865), .A2(n6731), .ZN(n8671) );
  NAND2HSV0 U10750 ( .A1(n8671), .A2(n13794), .ZN(n8672) );
  OAI21HSV0 U10751 ( .A1(n13794), .A2(n8671), .B(n8672), .ZN(n15206) );
  MUX2HSV2 U10752 ( .I0(\pe1/ti_7t [1]), .I1(n14956), .S(n10606), .Z(n10242)
         );
  NAND2HSV0 U10753 ( .A1(\pe19/bq[3] ), .A2(\pe19/aot [1]), .ZN(n8673) );
  CLKNAND2HSV0 U10754 ( .A1(n8673), .A2(n13314), .ZN(n8674) );
  OAI21HSV0 U10755 ( .A1(n13314), .A2(n8673), .B(n8674), .ZN(n8675) );
  XOR2HSV0 U10756 ( .A1(n14343), .A2(n14345), .Z(n8676) );
  NAND2HSV0 U10757 ( .A1(\pe17/ti_7[3] ), .A2(\pe17/got [3]), .ZN(n8677) );
  OAI21HSV0 U10758 ( .A1(n15167), .A2(n14347), .B(n8678), .ZN(n8679) );
  CLKNHSV0 U10759 ( .I(n13610), .ZN(n8681) );
  XOR2HSV0 U10760 ( .A1(n12946), .A2(n12948), .Z(n8682) );
  XOR2HSV0 U10761 ( .A1(n12947), .A2(n8682), .Z(n8683) );
  MUX2NHSV0 U10762 ( .I0(n13610), .I1(n8681), .S(n8683), .ZN(n8684) );
  OAI21HSV0 U10763 ( .A1(n14465), .A2(n12943), .B(n8684), .ZN(n8685) );
  OAI31HSV0 U10764 ( .A1(n14465), .A2(n8684), .A3(n12943), .B(n8685), .ZN(
        n8686) );
  CLKNAND2HSV0 U10765 ( .A1(n8687), .A2(n8686), .ZN(n8688) );
  OAI21HSV0 U10766 ( .A1(n8686), .A2(n8687), .B(n8688), .ZN(n8689) );
  NAND2HSV0 U10767 ( .A1(\pe7/ti_7[5] ), .A2(\pe7/got [3]), .ZN(n8690) );
  CLKNAND2HSV0 U10768 ( .A1(n8690), .A2(n8689), .ZN(n8691) );
  OAI21HSV0 U10769 ( .A1(n8689), .A2(n8690), .B(n8691), .ZN(n8692) );
  NAND2HSV0 U10770 ( .A1(n6038), .A2(n14487), .ZN(n8693) );
  CLKNAND2HSV0 U10771 ( .A1(n8693), .A2(n8692), .ZN(n8694) );
  OAI21HSV0 U10772 ( .A1(n8692), .A2(n8693), .B(n8694), .ZN(n8695) );
  CLKNAND2HSV0 U10773 ( .A1(n8695), .A2(n8696), .ZN(n8697) );
  OAI21HSV0 U10774 ( .A1(n8695), .A2(n8696), .B(n8697), .ZN(\pe7/poht [3]) );
  CLKNHSV0 U10775 ( .I(\pe5/got [1]), .ZN(n8698) );
  NAND2HSV0 U10776 ( .A1(\pe5/bq[1] ), .A2(\pe5/aot [2]), .ZN(n8699) );
  AOI21HSV0 U10777 ( .A1(\pe5/bq[2] ), .A2(\pe5/aot [1]), .B(n8699), .ZN(n8700) );
  AO31HSV2 U10778 ( .A1(\pe5/bq[2] ), .A2(\pe5/aot [1]), .A3(n8699), .B(n8700), 
        .Z(n8701) );
  NAND2HSV0 U10779 ( .A1(\pe5/ti_7[7] ), .A2(\pe5/got [2]), .ZN(n8704) );
  NAND2HSV0 U10780 ( .A1(n8704), .A2(n8703), .ZN(n8705) );
  OAI21HSV0 U10781 ( .A1(n8703), .A2(n8704), .B(n8705), .ZN(\pe5/poht [6]) );
  CLKNHSV0 U10782 ( .I(n13098), .ZN(n8706) );
  MUX2NHSV0 U10783 ( .I0(n8706), .I1(n13098), .S(n13097), .ZN(n8707) );
  CLKNHSV0 U10784 ( .I(n13100), .ZN(n8708) );
  OAI21HSV2 U10785 ( .A1(n8709), .A2(n8710), .B(n8711), .ZN(\pe2/poht [3]) );
  NAND2HSV0 U10786 ( .A1(n5997), .A2(\pe18/ti_7[1] ), .ZN(n8712) );
  CLKNHSV0 U10787 ( .I(bo18[5]), .ZN(n8713) );
  MUX2NHSV0 U10788 ( .I0(n8713), .I1(n14563), .S(n14564), .ZN(n15050) );
  MUX2HSV0 U10789 ( .I0(\pe12/pq ), .I1(n13830), .S(n14938), .Z(\pe12/ti_1t )
         );
  NAND2HSV0 U10790 ( .A1(\pe10/got [8]), .A2(n6033), .ZN(n8714) );
  NAND2HSV0 U10791 ( .A1(n8714), .A2(n13840), .ZN(n8715) );
  OAI21HSV2 U10792 ( .A1(n13840), .A2(n8714), .B(n8715), .ZN(n15263) );
  NAND2HSV0 U10793 ( .A1(\pe9/got [8]), .A2(n6209), .ZN(n8716) );
  NAND2HSV0 U10794 ( .A1(n8716), .A2(n9745), .ZN(n8717) );
  OAI21HSV0 U10795 ( .A1(n9745), .A2(n8716), .B(n8717), .ZN(pov9[5]) );
  CLKNHSV0 U10796 ( .I(bo7[8]), .ZN(n8718) );
  MUX2NHSV0 U10797 ( .I0(n8718), .I1(n11801), .S(n12067), .ZN(n15121) );
  NAND2HSV0 U10798 ( .A1(\pe4/got [8]), .A2(\pe4/ti_7[1] ), .ZN(n8719) );
  NAND2HSV0 U10799 ( .A1(n8719), .A2(n13851), .ZN(n8720) );
  OAI21HSV2 U10800 ( .A1(n13851), .A2(n8719), .B(n8720), .ZN(n15284) );
  NAND2HSV0 U10801 ( .A1(\pe21/aot [2]), .A2(\pe21/bq[8] ), .ZN(n8721) );
  NAND2HSV2 U10802 ( .A1(n8721), .A2(\pe21/phq [7]), .ZN(n8722) );
  OAI21HSV2 U10803 ( .A1(\pe21/phq [7]), .A2(n8721), .B(n8722), .ZN(n10844) );
  CLKNAND2HSV0 U10804 ( .A1(\pe8/pvq [7]), .A2(n14758), .ZN(n8723) );
  NAND2HSV2 U10805 ( .A1(n8723), .A2(\pe8/phq [7]), .ZN(n8724) );
  OAI21HSV2 U10806 ( .A1(\pe8/phq [7]), .A2(n8723), .B(n8724), .ZN(n11546) );
  CLKNHSV0 U10807 ( .I(\pe15/phq [6]), .ZN(n8725) );
  INAND2HSV0 U10808 ( .A1(\pe11/ti_7t [3]), .B1(n15090), .ZN(n11721) );
  NAND2HSV0 U10809 ( .A1(\pe16/got [5]), .A2(n11200), .ZN(n8726) );
  AO31HSV2 U10810 ( .A1(n13041), .A2(\pe6/pvq [5]), .A3(\pe6/phq [5]), .B(
        n8727), .Z(n9278) );
  OA21HSV4 U10811 ( .A1(n8976), .A2(n8977), .B(n8975), .Z(n8980) );
  INAND2HSV0 U10812 ( .A1(\pe18/ti_7t [3]), .B1(n13146), .ZN(n9200) );
  NAND2HSV0 U10813 ( .A1(\pe6/aot [4]), .A2(\pe6/bq[1] ), .ZN(n8728) );
  NAND2HSV0 U10814 ( .A1(\pe6/bq[2] ), .A2(\pe6/aot [3]), .ZN(n8729) );
  NAND2HSV0 U10815 ( .A1(n8729), .A2(n8728), .ZN(n8730) );
  OAI21HSV0 U10816 ( .A1(n8728), .A2(n8729), .B(n8730), .ZN(n13001) );
  CLKNHSV0 U10817 ( .I(n14336), .ZN(n8731) );
  AOI22HSV0 U10818 ( .A1(\pe17/aot [1]), .A2(n14412), .B1(\pe17/bq[3] ), .B2(
        \pe17/aot [5]), .ZN(n8732) );
  IAO21HSV2 U10819 ( .A1(n14335), .A2(n14334), .B(n8732), .ZN(n8733) );
  MUX2NHSV0 U10820 ( .I0(n14336), .I1(n8731), .S(n8733), .ZN(n14345) );
  NAND2HSV0 U10821 ( .A1(\pe1/bq[3] ), .A2(\pe1/aot [4]), .ZN(n8734) );
  OAI21HSV0 U10822 ( .A1(n14500), .A2(n13969), .B(n8734), .ZN(n8735) );
  OAI31HSV0 U10823 ( .A1(n14500), .A2(n8734), .A3(n13969), .B(n8735), .ZN(
        n13941) );
  CLKNHSV0 U10824 ( .I(n8905), .ZN(n8736) );
  OAI21HSV0 U10825 ( .A1(n13853), .A2(n13852), .B(n13854), .ZN(n8739) );
  OAI31HSV0 U10826 ( .A1(n13853), .A2(n13854), .A3(n13852), .B(n8739), .ZN(
        n15239) );
  NAND2HSV2 U10827 ( .A1(n12474), .A2(n14834), .ZN(n8740) );
  OAI21HSV2 U10828 ( .A1(bo3[8]), .A2(n12474), .B(n8740), .ZN(n15054) );
  NAND2HSV0 U10829 ( .A1(n12362), .A2(n14954), .ZN(n8741) );
  OAI21HSV0 U10830 ( .A1(bo20[8]), .A2(n12362), .B(n8741), .ZN(n8916) );
  NAND2HSV0 U10831 ( .A1(n5997), .A2(n14669), .ZN(n8742) );
  NAND2HSV0 U10832 ( .A1(n13255), .A2(n8742), .ZN(n8743) );
  OAI21HSV0 U10833 ( .A1(n8742), .A2(n13255), .B(n8743), .ZN(n15214) );
  CLKNHSV0 U10834 ( .I(n15178), .ZN(n8744) );
  NAND2HSV0 U10835 ( .A1(n14750), .A2(n15188), .ZN(n8745) );
  NAND2HSV0 U10836 ( .A1(n8745), .A2(n13259), .ZN(n8746) );
  OAI21HSV0 U10837 ( .A1(n13259), .A2(n8745), .B(n8746), .ZN(n15240) );
  XOR2HSV0 U10838 ( .A1(n13666), .A2(n13665), .Z(n8747) );
  XOR2HSV0 U10839 ( .A1(n13664), .A2(n8747), .Z(n8748) );
  NAND2HSV0 U10840 ( .A1(\pe20/got [5]), .A2(n6731), .ZN(n8752) );
  CLKNAND2HSV0 U10841 ( .A1(n8752), .A2(n8751), .ZN(n8753) );
  OAI21HSV0 U10842 ( .A1(n8751), .A2(n8752), .B(n8753), .ZN(n8754) );
  OAI21HSV0 U10843 ( .A1(n8754), .A2(n8755), .B(n8756), .ZN(\pe20/poht [2]) );
  NAND2HSV0 U10844 ( .A1(\pe19/bq[2] ), .A2(\pe19/aot [1]), .ZN(n8757) );
  NAND2HSV0 U10845 ( .A1(\pe19/aot [2]), .A2(\pe19/bq[1] ), .ZN(n8758) );
  CLKNAND2HSV0 U10846 ( .A1(n8758), .A2(n8757), .ZN(n8759) );
  OAI21HSV0 U10847 ( .A1(n8757), .A2(n8758), .B(n8759), .ZN(n8760) );
  XOR2HSV0 U10848 ( .A1(n14496), .A2(n14495), .Z(n8761) );
  XOR2HSV0 U10849 ( .A1(n14494), .A2(n8761), .Z(n8762) );
  CLKNAND2HSV0 U10850 ( .A1(n8763), .A2(n8762), .ZN(n8764) );
  OAI21HSV0 U10851 ( .A1(n8762), .A2(n8763), .B(n8764), .ZN(n8765) );
  NAND2HSV0 U10852 ( .A1(\pe14/got [2]), .A2(n15195), .ZN(n8766) );
  CLKNAND2HSV0 U10853 ( .A1(n8766), .A2(n8765), .ZN(n8767) );
  OAI21HSV0 U10854 ( .A1(n8765), .A2(n8766), .B(n8767), .ZN(n8768) );
  OAI21HSV0 U10855 ( .A1(n14489), .A2(n14488), .B(n8768), .ZN(n8769) );
  OAI31HSV0 U10856 ( .A1(n14489), .A2(n8768), .A3(n14488), .B(n8769), .ZN(
        n8770) );
  CLKNAND2HSV0 U10857 ( .A1(n8771), .A2(n8770), .ZN(n8772) );
  OAI21HSV0 U10858 ( .A1(n8770), .A2(n8771), .B(n8772), .ZN(n8773) );
  OAI21HSV0 U10859 ( .A1(n8774), .A2(n8773), .B(n8775), .ZN(\pe14/poht [3]) );
  CLKNHSV0 U10860 ( .I(\pe10/got [2]), .ZN(n8776) );
  XOR2HSV0 U10861 ( .A1(n13474), .A2(n13475), .Z(n8777) );
  NAND2HSV0 U10862 ( .A1(\pe10/ti_7[5] ), .A2(\pe10/got [3]), .ZN(n8778) );
  NAND2HSV0 U10863 ( .A1(\pe10/ti_7[6] ), .A2(\pe10/got [4]), .ZN(n8779) );
  CLKNHSV0 U10864 ( .I(n14208), .ZN(n8780) );
  MUX2NHSV0 U10865 ( .I0(n14208), .I1(n8780), .S(n13486), .ZN(n8781) );
  CLKNHSV0 U10866 ( .I(n14203), .ZN(n8782) );
  MUX2NHSV0 U10867 ( .I0(n8782), .I1(n14203), .S(n13487), .ZN(n8783) );
  XOR2HSV0 U10868 ( .A1(n8783), .A2(n8781), .Z(n8784) );
  AOI21HSV0 U10869 ( .A1(n15066), .A2(\pe8/got [1]), .B(n8784), .ZN(n8785) );
  AO31HSV2 U10870 ( .A1(n8784), .A2(n15066), .A3(\pe8/got [1]), .B(n8785), .Z(
        n8786) );
  NAND2HSV0 U10871 ( .A1(n14196), .A2(\pe8/got [2]), .ZN(n8787) );
  CLKNAND2HSV0 U10872 ( .A1(n8787), .A2(n8786), .ZN(n8788) );
  OAI21HSV0 U10873 ( .A1(n8786), .A2(n8787), .B(n8788), .ZN(n8789) );
  NAND2HSV0 U10874 ( .A1(n15182), .A2(\pe8/got [3]), .ZN(n8790) );
  CLKNAND2HSV0 U10875 ( .A1(n8790), .A2(n8789), .ZN(n8791) );
  OAI21HSV0 U10876 ( .A1(n8789), .A2(n8790), .B(n8791), .ZN(n8792) );
  NAND2HSV0 U10877 ( .A1(n15091), .A2(\pe8/got [4]), .ZN(n8793) );
  CLKNAND2HSV0 U10878 ( .A1(n8793), .A2(n8792), .ZN(n8794) );
  OAI21HSV0 U10879 ( .A1(n8792), .A2(n8793), .B(n8794), .ZN(\pe8/poht [4]) );
  XOR2HSV0 U10880 ( .A1(n12938), .A2(n12937), .Z(n8795) );
  XOR2HSV0 U10881 ( .A1(n12939), .A2(n8795), .Z(n8796) );
  NAND2HSV0 U10882 ( .A1(n15077), .A2(\pe6/got [3]), .ZN(n8797) );
  CLKNAND2HSV0 U10883 ( .A1(n8797), .A2(n8796), .ZN(n8798) );
  OAI21HSV0 U10884 ( .A1(n8796), .A2(n8797), .B(n8798), .ZN(n8799) );
  NAND2HSV0 U10885 ( .A1(\pe6/ti_7[5] ), .A2(\pe6/got [4]), .ZN(n8800) );
  CLKNAND2HSV0 U10886 ( .A1(n8800), .A2(n8799), .ZN(n8801) );
  OAI21HSV0 U10887 ( .A1(n8799), .A2(n8800), .B(n8801), .ZN(n8802) );
  CLKNAND2HSV0 U10888 ( .A1(n8803), .A2(n8802), .ZN(n8804) );
  NAND2HSV0 U10889 ( .A1(n14179), .A2(\pe6/got [6]), .ZN(n8806) );
  NAND2HSV0 U10890 ( .A1(n8806), .A2(n8805), .ZN(n8807) );
  OAI21HSV0 U10891 ( .A1(n8805), .A2(n8806), .B(n8807), .ZN(\pe6/poht [2]) );
  CLKNHSV0 U10892 ( .I(\pe1/got [3]), .ZN(n8808) );
  NAND2HSV0 U10893 ( .A1(n10242), .A2(\pe1/got [1]), .ZN(n8809) );
  CLKNAND2HSV0 U10894 ( .A1(n8809), .A2(n14004), .ZN(n8810) );
  OAI21HSV0 U10895 ( .A1(n14004), .A2(n8809), .B(n8810), .ZN(n8811) );
  XOR2HSV0 U10896 ( .A1(n13997), .A2(n13996), .Z(n8812) );
  XOR2HSV0 U10897 ( .A1(n8811), .A2(n8812), .Z(n8813) );
  OAI21HSV0 U10898 ( .A1(n14005), .A2(n8808), .B(n8813), .ZN(n8814) );
  OAI31HSV0 U10899 ( .A1(n14005), .A2(n8813), .A3(n8808), .B(n8814), .ZN(n8815) );
  NAND2HSV0 U10900 ( .A1(n14847), .A2(\pe1/got [4]), .ZN(n8816) );
  CLKNAND2HSV0 U10901 ( .A1(n8816), .A2(n8815), .ZN(n8817) );
  OAI21HSV0 U10902 ( .A1(n8815), .A2(n8816), .B(n8817), .ZN(n8818) );
  CLKNAND2HSV0 U10903 ( .A1(\pe1/ti_7[5] ), .A2(\pe1/got [5]), .ZN(n8819) );
  OAI21HSV2 U10904 ( .A1(n8818), .A2(n8819), .B(n8820), .ZN(n8821) );
  NAND2HSV0 U10905 ( .A1(\pe1/ti_7[6] ), .A2(\pe1/got [6]), .ZN(n8822) );
  CLKNAND2HSV0 U10906 ( .A1(n8825), .A2(n8824), .ZN(n8826) );
  OAI21HSV0 U10907 ( .A1(n8824), .A2(n8825), .B(n8826), .ZN(\pe1/poht [1]) );
  CLKNHSV0 U10908 ( .I(\pe21/pq ), .ZN(n8827) );
  MUX2NHSV0 U10909 ( .I0(n8827), .I1(n10847), .S(n14574), .ZN(\pe21/ti_1t ) );
  MUX2HSV0 U10910 ( .I0(\pe18/pq ), .I1(n13818), .S(n14790), .Z(\pe18/ti_1t )
         );
  CLKNHSV0 U10911 ( .I(n13875), .ZN(n8828) );
  INOR3HSV2 U10912 ( .A1(n13874), .B1(n13873), .B2(n13872), .ZN(n8829) );
  MUX2NHSV0 U10913 ( .I0(n8828), .I1(n13875), .S(n8829), .ZN(n15221) );
  NAND2HSV0 U10914 ( .A1(n13832), .A2(\pe16/pq ), .ZN(n8830) );
  OAI21HSV0 U10915 ( .A1(n13833), .A2(n13832), .B(n8830), .ZN(\pe16/ti_1t ) );
  MUX2HSV0 U10916 ( .I0(bo16[4]), .I1(\pe16/bq[4] ), .S(n14743), .Z(n15162) );
  MUX2HSV0 U10917 ( .I0(\pe13/pq ), .I1(n13819), .S(n13820), .Z(\pe13/ti_1t )
         );
  NAND2HSV0 U10918 ( .A1(n15179), .A2(\pe11/ti_7[1] ), .ZN(n8831) );
  NAND2HSV0 U10919 ( .A1(n8831), .A2(n13856), .ZN(n8832) );
  OAI21HSV0 U10920 ( .A1(n13856), .A2(n8831), .B(n8832), .ZN(n15259) );
  MUX2HSV0 U10921 ( .I0(bo10[8]), .I1(n12272), .S(n14554), .Z(n15028) );
  NAND2HSV0 U10922 ( .A1(\pe8/got [8]), .A2(\pe8/ti_7[1] ), .ZN(n8833) );
  NAND2HSV0 U10923 ( .A1(n8833), .A2(n6700), .ZN(n8834) );
  MUX2HSV0 U10924 ( .I0(bo7[5]), .I1(\pe7/bq[5] ), .S(n12067), .Z(n15122) );
  NAND2HSV0 U10925 ( .A1(n13861), .A2(n10346), .ZN(n8835) );
  NAND2HSV0 U10926 ( .A1(n8835), .A2(n13855), .ZN(n8836) );
  OAI21HSV2 U10927 ( .A1(n13855), .A2(n8835), .B(n8836), .ZN(n15279) );
  MUX2HSV0 U10928 ( .I0(bo5[7]), .I1(\pe5/bq[7] ), .S(n11818), .Z(n15110) );
  CLKNHSV0 U10929 ( .I(\pe4/pq ), .ZN(n8837) );
  MUX2NHSV0 U10930 ( .I0(n8837), .I1(n13813), .S(n13822), .ZN(\pe4/ti_1t ) );
  NAND2HSV0 U10931 ( .A1(n11708), .A2(n11707), .ZN(n8838) );
  NAND2HSV0 U10932 ( .A1(n8838), .A2(n10964), .ZN(n8839) );
  OAI21HSV0 U10933 ( .A1(n11709), .A2(n8838), .B(n8839), .ZN(n15286) );
  CLKNHSV0 U10934 ( .I(n13795), .ZN(n8840) );
  MUX2NHSV0 U10935 ( .I0(n8840), .I1(n13795), .S(n13796), .ZN(n15291) );
  AND2HSV0 U10936 ( .A1(\pe14/bq[6] ), .A2(\pe14/aot [5]), .Z(n11097) );
  CLKNAND2HSV0 U10937 ( .A1(n14953), .A2(\pe3/bq[4] ), .ZN(n8841) );
  AND2HSV0 U10938 ( .A1(n5973), .A2(\pe17/bq[1] ), .Z(n14409) );
  INAND2HSV0 U10939 ( .A1(n12139), .B1(n12138), .ZN(n12143) );
  INAND2HSV0 U10940 ( .A1(\pe9/ti_7t [3]), .B1(n9734), .ZN(n9735) );
  CLKNHSV0 U10941 ( .I(n12234), .ZN(n8842) );
  CLKNAND2HSV0 U10942 ( .A1(\pe7/pvq [6]), .A2(\pe7/ctrq ), .ZN(n8843) );
  CLKNAND2HSV0 U10943 ( .A1(n8843), .A2(\pe7/phq [6]), .ZN(n8844) );
  INOR2HSV0 U10944 ( .A1(\pe7/ti_7t [7]), .B1(n12308), .ZN(n14054) );
  AND2HSV0 U10945 ( .A1(\pe14/bq[5] ), .A2(n14891), .Z(n9108) );
  CLKNAND2HSV0 U10946 ( .A1(n10875), .A2(n10874), .ZN(n8846) );
  CLKNAND2HSV0 U10947 ( .A1(n8846), .A2(poh21[5]), .ZN(n8847) );
  OAI21HSV0 U10948 ( .A1(poh21[5]), .A2(n8846), .B(n8847), .ZN(po[6]) );
  CLKNAND2HSV0 U10949 ( .A1(n11780), .A2(n11781), .ZN(n8848) );
  CLKNAND2HSV0 U10950 ( .A1(n8848), .A2(poh21[1]), .ZN(n8849) );
  OAI21HSV0 U10951 ( .A1(poh21[1]), .A2(n8848), .B(n8849), .ZN(po[2]) );
  CLKNAND2HSV0 U10952 ( .A1(n8955), .A2(n14855), .ZN(n8850) );
  CLKNAND2HSV0 U10953 ( .A1(n15179), .A2(n14830), .ZN(n8851) );
  CLKNAND2HSV0 U10954 ( .A1(n8851), .A2(n13889), .ZN(n8852) );
  OAI21HSV0 U10955 ( .A1(n13889), .A2(n8851), .B(n8852), .ZN(n15254) );
  AOI21HSV0 U10956 ( .A1(n15089), .A2(n13897), .B(n13898), .ZN(n8853) );
  AO31HSV0 U10957 ( .A1(n15089), .A2(n13897), .A3(n13898), .B(n8853), .Z(
        n15274) );
  CLKNAND2HSV0 U10958 ( .A1(n15180), .A2(n14941), .ZN(n8854) );
  CLKNAND2HSV0 U10959 ( .A1(n8854), .A2(n13888), .ZN(n8855) );
  OAI21HSV0 U10960 ( .A1(n12500), .A2(n8854), .B(n8855), .ZN(n15285) );
  OAI21HSV0 U10961 ( .A1(n8856), .A2(n8857), .B(n8858), .ZN(po21) );
  CLKNAND2HSV0 U10962 ( .A1(n8859), .A2(n13337), .ZN(n8860) );
  OAI21HSV0 U10963 ( .A1(n13337), .A2(n8859), .B(n8860), .ZN(\pe13/poht [7])
         );
  XOR2HSV0 U10964 ( .A1(n12056), .A2(n12055), .Z(n8861) );
  OAI21HSV0 U10965 ( .A1(n12645), .A2(n12049), .B(n8861), .ZN(n8862) );
  OAI31HSV0 U10966 ( .A1(n12645), .A2(n8861), .A3(n12049), .B(n8862), .ZN(
        n8863) );
  CLKNAND2HSV0 U10967 ( .A1(n12631), .A2(\pe4/got [2]), .ZN(n8864) );
  CLKNAND2HSV0 U10968 ( .A1(n8864), .A2(n8863), .ZN(n8865) );
  OAI21HSV0 U10969 ( .A1(n8863), .A2(n8864), .B(n8865), .ZN(n8866) );
  CLKNAND2HSV0 U10970 ( .A1(n14850), .A2(\pe4/got [3]), .ZN(n8867) );
  CLKNAND2HSV0 U10971 ( .A1(n8867), .A2(n8866), .ZN(n8868) );
  CLKNAND2HSV0 U10972 ( .A1(\pe4/got [4]), .A2(n6181), .ZN(n8870) );
  CLKNAND2HSV0 U10973 ( .A1(n8873), .A2(n8872), .ZN(n8874) );
  OAI21HSV0 U10974 ( .A1(n8873), .A2(n8872), .B(n8874), .ZN(\pe4/poht [3]) );
  CLKNHSV0 U10975 ( .I(bo21[3]), .ZN(n8875) );
  MUX2NHSV0 U10976 ( .I0(n8875), .I1(n14560), .S(n14574), .ZN(n15048) );
  CLKNAND2HSV0 U10977 ( .A1(n8876), .A2(n13848), .ZN(n8877) );
  OAI21HSV0 U10978 ( .A1(n13848), .A2(n8876), .B(n8877), .ZN(n15209) );
  CLKNHSV0 U10979 ( .I(n10596), .ZN(n8878) );
  OAI21HSV0 U10980 ( .A1(n10595), .A2(n8878), .B(n10598), .ZN(n8879) );
  OAI31HSV0 U10981 ( .A1(n10595), .A2(n10598), .A3(n8878), .B(n8879), .ZN(
        n15207) );
  MUX2HSV0 U10982 ( .I0(bo20[1]), .I1(\pe20/bq[1] ), .S(n12362), .Z(n15013) );
  CLKNHSV0 U10983 ( .I(\pe19/pq ), .ZN(n8880) );
  MUX2NHSV0 U10984 ( .I0(n8880), .I1(n12155), .S(n14501), .ZN(\pe19/ti_1t ) );
  INAND3HSV0 U10985 ( .A1(n13868), .B1(n13869), .B2(n13870), .ZN(n8881) );
  OAI21HSV0 U10986 ( .A1(n13871), .A2(n8881), .B(n8882), .ZN(n15227) );
  CLKNHSV0 U10987 ( .I(bo16[7]), .ZN(n8883) );
  MUX2NHSV0 U10988 ( .I0(n8883), .I1(n14565), .S(n6599), .ZN(n15051) );
  NAND3HSV0 U10989 ( .A1(n11699), .A2(n11698), .A3(n11700), .ZN(n8884) );
  CLKNAND2HSV0 U10990 ( .A1(n8884), .A2(n11701), .ZN(n8885) );
  OAI21HSV0 U10991 ( .A1(n11701), .A2(n8884), .B(n8885), .ZN(n15202) );
  MUX2HSV0 U10992 ( .I0(\pe15/pq ), .I1(n14587), .S(n13815), .Z(\pe15/ti_1t )
         );
  MUX2HSV0 U10993 ( .I0(bo15[4]), .I1(\pe15/bq[4] ), .S(n12343), .Z(n15022) );
  CLKNAND2HSV0 U10994 ( .A1(n14750), .A2(\pe13/ti_7[1] ), .ZN(n8886) );
  CLKNAND2HSV0 U10995 ( .A1(n8886), .A2(n13847), .ZN(n8887) );
  OAI21HSV0 U10996 ( .A1(n13847), .A2(n8886), .B(n8887), .ZN(n15245) );
  CLKNHSV0 U10997 ( .I(bo13[5]), .ZN(n8888) );
  MUX2NHSV0 U10998 ( .I0(n8888), .I1(n11832), .S(n14795), .ZN(n15151) );
  CLKNHSV0 U10999 ( .I(bo12[7]), .ZN(n8889) );
  MUX2NHSV0 U11000 ( .I0(n8889), .I1(n14577), .S(n14578), .ZN(n15062) );
  MUX2HSV0 U11001 ( .I0(\pe11/pq ), .I1(n13811), .S(n13812), .Z(\pe11/ti_1t )
         );
  CLKNHSV0 U11002 ( .I(bo10[5]), .ZN(n8890) );
  MUX2NHSV0 U11003 ( .I0(n8890), .I1(n10029), .S(n14554), .ZN(n14989) );
  CLKNAND2HSV0 U11004 ( .A1(\pe9/got [8]), .A2(\pe9/ti_7[1] ), .ZN(n8891) );
  CLKNAND2HSV0 U11005 ( .A1(n8891), .A2(n7880), .ZN(n8892) );
  OAI21HSV0 U11006 ( .A1(n7880), .A2(n8891), .B(n8892), .ZN(n15265) );
  CLKNHSV0 U11007 ( .I(\pe9/pq ), .ZN(n8893) );
  MUX2NHSV0 U11008 ( .I0(n8893), .I1(n8943), .S(n13826), .ZN(\pe9/ti_1t ) );
  CLKNHSV0 U11009 ( .I(n13876), .ZN(n8894) );
  OAI21HSV0 U11010 ( .A1(n8894), .A2(n13877), .B(\pe8/got [8]), .ZN(n8895) );
  CLKNAND2HSV0 U11011 ( .A1(n8895), .A2(n13878), .ZN(n8896) );
  OAI21HSV0 U11012 ( .A1(n8895), .A2(n13878), .B(n8896), .ZN(n15204) );
  CLKNAND2HSV0 U11013 ( .A1(n10459), .A2(\pe7/ti_7[1] ), .ZN(n8897) );
  MUX2HSV0 U11014 ( .I0(bo7[1]), .I1(\pe7/bq[1] ), .S(n12067), .Z(n15037) );
  MUX2HSV0 U11015 ( .I0(\pe6/pq ), .I1(n13824), .S(n13828), .Z(\pe6/ti_1t ) );
  AOI21HSV0 U11016 ( .A1(n14916), .A2(n13861), .B(n6704), .ZN(n8898) );
  AO31HSV0 U11017 ( .A1(n14916), .A2(n13861), .A3(n6704), .B(n8898), .Z(n15277) );
  MUX2HSV0 U11018 ( .I0(bo4[7]), .I1(\pe4/bq[7] ), .S(n13822), .Z(\pe4/bqt[7] ) );
  MUX2HSV0 U11019 ( .I0(bo3[5]), .I1(\pe3/bq[5] ), .S(n12474), .Z(n15043) );
  CLKNHSV0 U11020 ( .I(\pe2/pq ), .ZN(n8899) );
  MUX2NHSV0 U11021 ( .I0(n8899), .I1(n13775), .S(n14523), .ZN(\pe2/ti_1t ) );
  CLKNHSV0 U11022 ( .I(bo1[7]), .ZN(n8900) );
  MUX2NHSV0 U11023 ( .I0(n8900), .I1(n14503), .S(\pe1/ctrq ), .ZN(n14975) );
  BUFHSV4 U11024 ( .I(ctro14), .Z(n11093) );
  INHSV4 U11025 ( .I(ctro7), .ZN(n11782) );
  INHSV4 U11026 ( .I(ctro7), .ZN(n12308) );
  INHSV4 U11027 ( .I(n12311), .ZN(n12252) );
  INHSV12 U11028 ( .I(ctro19), .ZN(n9541) );
  INHSV4 U11029 ( .I(ctro8), .ZN(n11591) );
  INHSV4 U11030 ( .I(ctro8), .ZN(n10508) );
  CLKNHSV0 U11031 ( .I(n11956), .ZN(n14788) );
  INHSV2 U11032 ( .I(\pe8/got [8]), .ZN(n11603) );
  INHSV6 U11033 ( .I(ctro3), .ZN(n10405) );
  INHSV4 U11034 ( .I(n10405), .ZN(n10939) );
  INHSV6 U11035 ( .I(n10405), .ZN(n10994) );
  CLKNHSV6 U11036 ( .I(n10863), .ZN(n10873) );
  INHSV4 U11037 ( .I(n11780), .ZN(n9398) );
  INHSV8 U11038 ( .I(n11795), .ZN(n12362) );
  INHSV8 U11039 ( .I(ctro15), .ZN(n10521) );
  INHSV4 U11040 ( .I(n12266), .ZN(n10459) );
  INHSV6 U11041 ( .I(n14904), .ZN(n10562) );
  INHSV6 U11042 ( .I(n14904), .ZN(n13822) );
  INHSV6 U11043 ( .I(n11943), .ZN(n11948) );
  INHSV12 U11044 ( .I(n14926), .ZN(n13826) );
  CLKNHSV0 U11045 ( .I(n11954), .ZN(n14832) );
  CLKNHSV6 U11046 ( .I(ctro5), .ZN(n10307) );
  INHSV2 U11047 ( .I(n10307), .ZN(n13015) );
  INHSV6 U11048 ( .I(n11156), .ZN(n14702) );
  INHSV4 U11049 ( .I(n9629), .ZN(n9714) );
  INHSV4 U11050 ( .I(n10073), .ZN(n10040) );
  CLKNHSV0 U11051 ( .I(\pe21/got [6]), .ZN(n10852) );
  INHSV6 U11052 ( .I(n13146), .ZN(n13145) );
  INHSV6 U11053 ( .I(n13145), .ZN(n13143) );
  INHSV4 U11054 ( .I(n9921), .ZN(n9881) );
  INHSV6 U11055 ( .I(ctro13), .ZN(n9977) );
  INHSV2 U11056 ( .I(n15090), .ZN(n11765) );
  BUFHSV4 U11057 ( .I(ctro11), .Z(n9609) );
  INHSV4 U11058 ( .I(n9203), .ZN(n11988) );
  INHSV4 U11059 ( .I(n10508), .ZN(n11521) );
  INHSV4 U11060 ( .I(n10796), .ZN(n10689) );
  INHSV4 U11061 ( .I(n11782), .ZN(n12267) );
  CLKNAND2HSV4 U11062 ( .A1(n9880), .A2(n9879), .ZN(n9920) );
  INHSV2 U11063 ( .I(n5977), .ZN(n9797) );
  CLKNHSV0 U11064 ( .I(\pe5/ti_1 ), .ZN(n10316) );
  INHSV2 U11065 ( .I(n10522), .ZN(n11296) );
  INHSV4 U11066 ( .I(n14404), .ZN(n14571) );
  CLKNHSV6 U11067 ( .I(n12187), .ZN(n14554) );
  INHSV4 U11068 ( .I(n11848), .ZN(n14572) );
  INHSV4 U11069 ( .I(n11848), .ZN(n14758) );
  INHSV6 U11070 ( .I(n11812), .ZN(n11818) );
  INHSV4 U11071 ( .I(n14540), .ZN(n11786) );
  INHSV4 U11072 ( .I(n14540), .ZN(n14574) );
  INHSV6 U11073 ( .I(n14543), .ZN(n14501) );
  INHSV12 U11074 ( .I(n10803), .ZN(n12067) );
  BUFHSV4 U11075 ( .I(n11790), .Z(n12357) );
  INHSV4 U11076 ( .I(n9977), .ZN(n9921) );
  INHSV4 U11077 ( .I(n9977), .ZN(n9988) );
  INHSV2 U11078 ( .I(\pe1/aot [7]), .ZN(n10616) );
  INHSV2 U11079 ( .I(n10307), .ZN(n13018) );
  NOR2HSV4 U11080 ( .A1(n11603), .A2(n11521), .ZN(n11602) );
  INHSV2 U11081 ( .I(ctro20), .ZN(n13676) );
  INHSV4 U11082 ( .I(n13676), .ZN(n8942) );
  BUFHSV8 U11083 ( .I(ctro20), .Z(n15177) );
  CLKNHSV0 U11084 ( .I(\pe16/got [4]), .ZN(n13189) );
  CLKNHSV0 U11085 ( .I(\pe4/bq[1] ), .ZN(n12771) );
  NOR2HSV2 U11086 ( .A1(n13141), .A2(n13146), .ZN(n9149) );
  INHSV4 U11087 ( .I(n12830), .ZN(n14735) );
  INHSV2 U11088 ( .I(n10525), .ZN(n11447) );
  CLKNAND2HSV2 U11089 ( .A1(ctro14), .A2(\pe14/ti_7t [4]), .ZN(n11113) );
  INHSV2 U11090 ( .I(n11113), .ZN(n11091) );
  CLKAND2HSV2 U11091 ( .A1(n12206), .A2(n10459), .Z(n8905) );
  CLKNHSV0 U11092 ( .I(\pe10/bq[1] ), .ZN(n12338) );
  INHSV6 U11093 ( .I(ctro4), .ZN(n9629) );
  INHSV4 U11094 ( .I(n14861), .ZN(n10510) );
  INHSV4 U11095 ( .I(\pe11/ctrq ), .ZN(n11838) );
  CLKNHSV0 U11096 ( .I(\pe16/got [6]), .ZN(n14070) );
  INHSV4 U11097 ( .I(n14701), .ZN(n12713) );
  CLKNAND2HSV2 U11098 ( .A1(n9517), .A2(n9516), .ZN(n11777) );
  AND2HSV2 U11099 ( .A1(n11211), .A2(n14064), .Z(n8906) );
  BUFHSV2 U11100 ( .I(ctro14), .Z(n11090) );
  CLKNHSV0 U11101 ( .I(\pe10/bq[3] ), .ZN(n12188) );
  INHSV4 U11102 ( .I(n10435), .ZN(n14429) );
  INHSV4 U11103 ( .I(n15134), .ZN(n13488) );
  INHSV4 U11104 ( .I(\pe7/ctrq ), .ZN(n10803) );
  CLKNHSV0 U11105 ( .I(\pe13/bq[2] ), .ZN(n9960) );
  CLKNHSV0 U11106 ( .I(\pe14/bq[3] ), .ZN(n13560) );
  INHSV4 U11107 ( .I(n9884), .ZN(n9882) );
  INHSV2 U11108 ( .I(n9399), .ZN(n9734) );
  NAND2HSV4 U11109 ( .A1(n14828), .A2(\pe10/ti_7t [3]), .ZN(n10127) );
  INHSV4 U11110 ( .I(n14836), .ZN(n14837) );
  XOR2HSV0 U11111 ( .A1(n9512), .A2(n9511), .Z(n9555) );
  AND2HSV2 U11112 ( .A1(n10800), .A2(n9307), .Z(n8910) );
  CLKNHSV0 U11113 ( .I(\pe4/bq[2] ), .ZN(n12190) );
  CLKNHSV0 U11114 ( .I(\pe3/bq[3] ), .ZN(n12355) );
  CLKNHSV0 U11115 ( .I(\pe15/bq[2] ), .ZN(n12344) );
  CLKNHSV0 U11116 ( .I(n9533), .ZN(n13104) );
  NAND2HSV2 U11117 ( .A1(n9842), .A2(\pe6/ti_7t [3]), .ZN(n9533) );
  AND2HSV2 U11118 ( .A1(n12017), .A2(n12016), .Z(n8911) );
  INHSV4 U11119 ( .I(\pe10/phq [2]), .ZN(n10041) );
  XOR2HSV4 U11120 ( .A1(n9234), .A2(n9233), .Z(n8912) );
  INHSV4 U11121 ( .I(n10853), .ZN(n10402) );
  INHSV4 U11122 ( .I(n11834), .ZN(n14552) );
  INHSV4 U11123 ( .I(n9720), .ZN(n9420) );
  INHSV4 U11124 ( .I(\pe16/ctrq ), .ZN(n13832) );
  INHSV6 U11125 ( .I(ctro17), .ZN(n13268) );
  INHSV2 U11126 ( .I(n13268), .ZN(n13269) );
  INHSV2 U11127 ( .I(n13268), .ZN(n14013) );
  OR2HSV1 U11128 ( .A1(n13346), .A2(n13345), .Z(n8913) );
  NAND2HSV2 U11129 ( .A1(ctro2), .A2(\pe2/ti_7t [6]), .ZN(n8914) );
  INHSV2 U11130 ( .I(n11691), .ZN(n9794) );
  INHSV2 U11131 ( .I(n12308), .ZN(n12309) );
  INHSV6 U11132 ( .I(n10796), .ZN(n8957) );
  INHSV4 U11133 ( .I(n8957), .ZN(n11220) );
  INHSV2 U11134 ( .I(n9358), .ZN(n11266) );
  INHSV4 U11135 ( .I(ctro1), .ZN(n10228) );
  INHSV2 U11136 ( .I(n13143), .ZN(n11976) );
  INHSV4 U11137 ( .I(n9461), .ZN(n13718) );
  CLKNHSV0 U11138 ( .I(n11590), .ZN(n11597) );
  AND2HSV2 U11139 ( .A1(n15177), .A2(\pe20/ti_7t [6]), .Z(n8915) );
  INHSV2 U11140 ( .I(n9541), .ZN(n14700) );
  INHSV4 U11141 ( .I(n9736), .ZN(n9434) );
  MUX2HSV2 U11142 ( .I0(bo21[8]), .I1(n13810), .S(n6014), .Z(n8917) );
  MUX2HSV2 U11143 ( .I0(bo9[7]), .I1(n5976), .S(n13826), .Z(n8918) );
  MUX2HSV2 U11144 ( .I0(bo6[7]), .I1(n8933), .S(n14870), .Z(n8919) );
  INHSV2 U11145 ( .I(\pe2/got [1]), .ZN(n13776) );
  CLKNHSV0 U11146 ( .I(n9286), .ZN(n9288) );
  INHSV4 U11147 ( .I(n15074), .ZN(n9790) );
  INHSV6 U11148 ( .I(n15074), .ZN(n14866) );
  NOR2HSV2 U11149 ( .A1(n11668), .A2(n11667), .ZN(n8920) );
  OR2HSV1 U11150 ( .A1(n12311), .A2(n10459), .Z(n8921) );
  NAND2HSV0 U11151 ( .A1(n11691), .A2(n9434), .ZN(n8922) );
  NAND2HSV2 U11152 ( .A1(n9734), .A2(\pe9/ti_7t [5]), .ZN(n8923) );
  BUFHSV4 U11153 ( .I(\pe3/ti_1 ), .Z(n12475) );
  CLKNHSV0 U11154 ( .I(n12155), .ZN(n13821) );
  CLKNAND2HSV2 U11155 ( .A1(\pe7/aot [5]), .A2(\pe7/bq[6] ), .ZN(n12234) );
  INHSV2 U11156 ( .I(n8934), .ZN(n8925) );
  NAND2HSV0 U11157 ( .A1(\pe7/aot [8]), .A2(\pe7/bq[5] ), .ZN(n12063) );
  NAND2HSV2 U11158 ( .A1(\pe4/bq[7] ), .A2(\pe4/aot [8]), .ZN(n9125) );
  INHSV4 U11159 ( .I(n8931), .ZN(n14502) );
  INHSV2 U11160 ( .I(\pe4/ti_1 ), .ZN(n8926) );
  INHSV2 U11161 ( .I(n8926), .ZN(n8927) );
  INHSV4 U11162 ( .I(n14013), .ZN(n8928) );
  CLKNHSV0 U11163 ( .I(\pe7/bq[6] ), .ZN(n8929) );
  INHSV2 U11164 ( .I(n8929), .ZN(n8930) );
  INHSV4 U11165 ( .I(\pe1/bq[8] ), .ZN(n8931) );
  NAND2HSV2 U11166 ( .A1(\pe21/bq[8] ), .A2(\pe21/aot [5]), .ZN(n10395) );
  NAND2HSV2 U11167 ( .A1(\pe16/aot [2]), .A2(\pe16/bq[6] ), .ZN(n14083) );
  INAND2HSV2 U11168 ( .A1(n11692), .B1(n8920), .ZN(n11672) );
  NOR2HSV0 U11169 ( .A1(n14582), .A2(n14866), .ZN(n11690) );
  CLKNHSV0 U11170 ( .I(\pe6/bq[7] ), .ZN(n8932) );
  CLKNHSV0 U11171 ( .I(n8932), .ZN(n8933) );
  NAND2HSV0 U11172 ( .A1(\pe21/got [6]), .A2(\pe21/ti_7[5] ), .ZN(n13135) );
  CLKNAND2HSV2 U11173 ( .A1(\pe6/aot [1]), .A2(\pe6/bq[4] ), .ZN(n13000) );
  INHSV4 U11174 ( .I(\pe6/ctrq ), .ZN(n8934) );
  CLKNHSV6 U11175 ( .I(n8934), .ZN(n8935) );
  NAND2HSV0 U11176 ( .A1(\pe6/bq[7] ), .A2(\pe6/aot [8]), .ZN(n9251) );
  CLKNHSV0 U11177 ( .I(\pe20/aot [7]), .ZN(n8936) );
  INHSV2 U11178 ( .I(n8936), .ZN(n8937) );
  NAND2HSV0 U11179 ( .A1(\pe3/got [5]), .A2(\pe3/ti_1 ), .ZN(n10199) );
  INHSV6 U11180 ( .I(n14512), .ZN(n14790) );
  CLKNHSV0 U11181 ( .I(n11952), .ZN(n8938) );
  INHSV2 U11182 ( .I(n10405), .ZN(n10168) );
  NAND2HSV0 U11183 ( .A1(\pe10/ti_7[5] ), .A2(\pe10/got [1]), .ZN(n14114) );
  CLKNHSV0 U11184 ( .I(\pe10/got [1]), .ZN(n13899) );
  NAND2HSV0 U11185 ( .A1(n14940), .A2(\pe10/got [1]), .ZN(n13461) );
  INHSV2 U11186 ( .I(n10521), .ZN(n10522) );
  BUFHSV2 U11187 ( .I(\pe6/ti_1 ), .Z(n13824) );
  NAND2HSV2 U11188 ( .A1(n12022), .A2(n12021), .ZN(n12109) );
  INHSV4 U11189 ( .I(n13268), .ZN(n12021) );
  OAI21HSV0 U11190 ( .A1(n15201), .A2(n13902), .B(n13901), .ZN(n13904) );
  INHSV2 U11191 ( .I(n13677), .ZN(n8939) );
  NAND2HSV0 U11192 ( .A1(n14523), .A2(\pe2/pq ), .ZN(n13768) );
  CLKNHSV0 U11193 ( .I(n10451), .ZN(n8940) );
  INHSV4 U11194 ( .I(n14199), .ZN(n8941) );
  INHSV4 U11195 ( .I(\pe8/bq[6] ), .ZN(n14199) );
  CLKNAND2HSV2 U11196 ( .A1(n11094), .A2(n8948), .ZN(n11115) );
  NAND3HSV2 U11197 ( .A1(n11064), .A2(n11062), .A3(n8948), .ZN(n11061) );
  NAND2HSV0 U11198 ( .A1(\pe13/aot [8]), .A2(\pe13/bq[5] ), .ZN(n9891) );
  BUFHSV2 U11199 ( .I(\pe13/aot [8]), .Z(n14939) );
  NAND2HSV0 U11200 ( .A1(\pe9/bq[2] ), .A2(\pe9/aot [6]), .ZN(n13915) );
  NAND2HSV0 U11201 ( .A1(\pe9/aot [6]), .A2(\pe9/bq[6] ), .ZN(n9445) );
  NAND2HSV0 U11202 ( .A1(\pe18/bq[5] ), .A2(\pe18/aot [8]), .ZN(n9158) );
  CLKNAND2HSV2 U11203 ( .A1(n9823), .A2(n13897), .ZN(n9306) );
  NAND2HSV0 U11204 ( .A1(n9823), .A2(\pe6/got [4]), .ZN(n9299) );
  CLKNHSV0 U11205 ( .I(\pe9/ti_1 ), .ZN(n8943) );
  INHSV2 U11206 ( .I(n8943), .ZN(n8944) );
  NAND2HSV0 U11207 ( .A1(\pe16/aot [8]), .A2(\pe16/bq[4] ), .ZN(n10698) );
  CLKNHSV0 U11208 ( .I(n14503), .ZN(n8945) );
  INHSV4 U11209 ( .I(\pe1/bq[7] ), .ZN(n14503) );
  AOI21HSV2 U11210 ( .A1(n12260), .A2(n9420), .B(n9734), .ZN(n9005) );
  CLKNHSV0 U11211 ( .I(n13766), .ZN(n8946) );
  NAND2HSV0 U11212 ( .A1(\pe13/aot [6]), .A2(\pe13/bq[7] ), .ZN(n9890) );
  NAND2HSV0 U11213 ( .A1(\pe3/aot [3]), .A2(\pe3/bq[5] ), .ZN(n12748) );
  NAND2HSV0 U11214 ( .A1(\pe3/bq[5] ), .A2(\pe3/aot [8]), .ZN(n10194) );
  NAND2HSV0 U11215 ( .A1(\pe3/aot [6]), .A2(\pe3/bq[6] ), .ZN(n10207) );
  NAND2HSV2 U11216 ( .A1(\pe3/bq[6] ), .A2(\pe3/aot [2]), .ZN(n12750) );
  NAND2HSV0 U11217 ( .A1(\pe3/aot [6]), .A2(\pe3/bq[7] ), .ZN(n10195) );
  NAND2HSV0 U11218 ( .A1(n14820), .A2(\pe3/got [4]), .ZN(n12493) );
  NAND2HSV2 U11219 ( .A1(n13733), .A2(\pe20/bq[6] ), .ZN(n9019) );
  NAND2HSV0 U11220 ( .A1(n10784), .A2(\pe10/got [8]), .ZN(n10785) );
  NAND2HSV0 U11221 ( .A1(\pe20/bq[6] ), .A2(\pe20/aot [5]), .ZN(n9476) );
  NAND2HSV2 U11222 ( .A1(\pe20/bq[7] ), .A2(\pe20/aot [8]), .ZN(n9027) );
  NAND2HSV2 U11223 ( .A1(\pe13/aot [1]), .A2(\pe13/bq[5] ), .ZN(n12924) );
  AND2HSV2 U11224 ( .A1(\pe13/aot [1]), .A2(\pe13/bq[1] ), .Z(n13337) );
  NAND2HSV0 U11225 ( .A1(n12609), .A2(\pe4/got [4]), .ZN(n12605) );
  NAND2HSV0 U11226 ( .A1(n12631), .A2(\pe4/got [4]), .ZN(n12655) );
  CLKNHSV0 U11227 ( .I(\pe4/got [4]), .ZN(n10536) );
  CLKNHSV0 U11228 ( .I(\pe9/aot [5]), .ZN(n8949) );
  INHSV2 U11229 ( .I(n8949), .ZN(n8950) );
  NAND2HSV0 U11230 ( .A1(n7875), .A2(\pe9/got [4]), .ZN(n9795) );
  NAND2HSV0 U11231 ( .A1(n7875), .A2(\pe9/got [3]), .ZN(n11644) );
  NAND2HSV0 U11232 ( .A1(n7875), .A2(\pe9/got [6]), .ZN(n11666) );
  NAND2HSV0 U11233 ( .A1(n6731), .A2(\pe20/got [1]), .ZN(n14176) );
  NAND2HSV0 U11234 ( .A1(n11854), .A2(\pe20/got [1]), .ZN(n13691) );
  INHSV4 U11235 ( .I(n14546), .ZN(n14512) );
  INHSV4 U11236 ( .I(n14512), .ZN(n14564) );
  NAND2HSV0 U11237 ( .A1(\pe21/bq[6] ), .A2(\pe21/aot [2]), .ZN(n12090) );
  NAND2HSV0 U11238 ( .A1(\pe21/bq[6] ), .A2(\pe21/aot [5]), .ZN(n10813) );
  NAND2HSV0 U11239 ( .A1(n9763), .A2(\pe9/got [5]), .ZN(n9788) );
  NAND2HSV0 U11240 ( .A1(n14896), .A2(\pe9/got [5]), .ZN(n9414) );
  CLKNHSV0 U11241 ( .I(n14822), .ZN(n8953) );
  INHSV2 U11242 ( .I(n8953), .ZN(n8954) );
  NAND2HSV0 U11243 ( .A1(\pe18/got [5]), .A2(\pe18/ti_1 ), .ZN(n9157) );
  NAND2HSV2 U11244 ( .A1(n14851), .A2(\pe18/got [5]), .ZN(n13173) );
  INHSV2 U11245 ( .I(\pe18/got [5]), .ZN(n14621) );
  INHSV4 U11246 ( .I(n14955), .ZN(n14861) );
  INHSV4 U11247 ( .I(n11089), .ZN(n8955) );
  INHSV4 U11248 ( .I(n11220), .ZN(n8956) );
  NAND2HSV4 U11249 ( .A1(n11387), .A2(\pe15/got [7]), .ZN(n11290) );
  MUX2NHSV4 U11250 ( .I0(n8960), .I1(n8958), .S(n9324), .ZN(n8965) );
  NAND3HSV2 U11251 ( .A1(n9395), .A2(\pe21/aot [8]), .A3(\pe21/bq[8] ), .ZN(
        n9397) );
  CLKXOR2HSV4 U11252 ( .A1(n9100), .A2(n11081), .Z(n9102) );
  NAND2HSV2 U11253 ( .A1(\pe4/aot [6]), .A2(\pe4/bq[5] ), .ZN(n9693) );
  CLKNAND2HSV8 U11254 ( .A1(n10373), .A2(n10372), .ZN(n10400) );
  INHSV4 U11255 ( .I(n9733), .ZN(n10355) );
  CLKNAND2HSV2 U11256 ( .A1(n13089), .A2(n8955), .ZN(n13090) );
  NOR2HSV4 U11257 ( .A1(n12981), .A2(n10168), .ZN(n11000) );
  INHSV4 U11259 ( .I(n13766), .ZN(n9324) );
  INHSV2 U11260 ( .I(\pe2/pvq [1]), .ZN(n8959) );
  NAND2HSV2 U11261 ( .A1(n8960), .A2(n8959), .ZN(n8963) );
  INHSV2 U11262 ( .I(ctro2), .ZN(n9378) );
  INHSV2 U11263 ( .I(\pe2/ti_7t [1]), .ZN(n8966) );
  NOR2HSV4 U11264 ( .A1(n9378), .A2(n8966), .ZN(n8967) );
  INHSV2 U11265 ( .I(n8967), .ZN(n9338) );
  INHSV4 U11266 ( .I(ctro2), .ZN(n9381) );
  NAND2HSV2 U11267 ( .A1(n9338), .A2(n9358), .ZN(n8987) );
  CLKNAND2HSV1 U11268 ( .A1(n8987), .A2(\pe2/got [7]), .ZN(n8968) );
  INHSV2 U11269 ( .I(n10708), .ZN(n14818) );
  INHSV2 U11270 ( .I(\pe2/phq [2]), .ZN(n8969) );
  AOI21HSV2 U11271 ( .A1(n8974), .A2(n8973), .B(n8972), .ZN(n8976) );
  INHSV2 U11272 ( .I(n8980), .ZN(n8978) );
  NOR2HSV1 U11273 ( .A1(n10708), .A2(ctro2), .ZN(n11242) );
  CLKNHSV0 U11274 ( .I(n11242), .ZN(n8979) );
  CLKAND2HSV2 U11275 ( .A1(n9358), .A2(\pe2/ti_7t [2]), .Z(n8981) );
  XNOR2HSV4 U11276 ( .A1(n8983), .A2(n9345), .ZN(n8985) );
  AOI21HSV4 U11277 ( .A1(n8985), .A2(n11266), .B(n8984), .ZN(n8994) );
  CLKNAND2HSV1 U11278 ( .A1(\pe2/aot [7]), .A2(\pe2/bq[6] ), .ZN(n8989) );
  NAND2HSV0 U11279 ( .A1(n14858), .A2(\pe2/bq[5] ), .ZN(n8988) );
  XNOR2HSV4 U11280 ( .A1(n8992), .A2(n8991), .ZN(n8993) );
  XNOR2HSV4 U11281 ( .A1(n8994), .A2(n8993), .ZN(n15070) );
  CLKNAND2HSV2 U11282 ( .A1(\pe9/ti_1 ), .A2(\pe9/got [8]), .ZN(n8996) );
  NAND2HSV4 U11283 ( .A1(\pe9/aot [8]), .A2(\pe9/bq[8] ), .ZN(n8995) );
  CLKNAND2HSV4 U11284 ( .A1(\pe9/ctrq ), .A2(\pe9/pvq [1]), .ZN(n8997) );
  INHSV2 U11285 ( .I(\pe9/got [8]), .ZN(n9451) );
  NOR2HSV2 U11286 ( .A1(ctro9), .A2(n9451), .ZN(n11691) );
  NAND2HSV2 U11287 ( .A1(\pe9/ti_1 ), .A2(\pe9/got [7]), .ZN(n8999) );
  INHSV2 U11288 ( .I(\pe9/phq [2]), .ZN(n8998) );
  CLKNHSV2 U11289 ( .I(\pe9/ti_7t [2]), .ZN(n9003) );
  NOR2HSV4 U11290 ( .A1(n9450), .A2(n9003), .ZN(n9004) );
  INHSV2 U11291 ( .I(\pe9/got [8]), .ZN(n9720) );
  CLKNAND2HSV2 U11292 ( .A1(n7880), .A2(n9005), .ZN(n9006) );
  NAND2HSV2 U11293 ( .A1(ctro9), .A2(\pe9/ti_7t [1]), .ZN(n9400) );
  INHSV1 U11294 ( .I(n9400), .ZN(n9008) );
  INHSV2 U11295 ( .I(ctro9), .ZN(n9399) );
  CLKNAND2HSV0 U11296 ( .A1(n9400), .A2(n9734), .ZN(n9429) );
  INHSV2 U11297 ( .I(\pe9/got [7]), .ZN(n9736) );
  INHSV2 U11298 ( .I(n9736), .ZN(n9449) );
  CLKNAND2HSV1 U11299 ( .A1(n9429), .A2(n9449), .ZN(n9009) );
  CLKNHSV2 U11300 ( .I(\pe20/phq [1]), .ZN(n9010) );
  XNOR2HSV4 U11301 ( .A1(n9032), .A2(n9031), .ZN(n12352) );
  INHSV2 U11302 ( .I(n9062), .ZN(n9011) );
  NOR2HSV4 U11303 ( .A1(n12352), .A2(n9011), .ZN(n9038) );
  NAND2HSV0 U11304 ( .A1(n9062), .A2(ctro20), .ZN(n9040) );
  BUFHSV2 U11305 ( .I(\pe20/got [7]), .Z(n14890) );
  INHSV2 U11306 ( .I(n14890), .ZN(n9461) );
  CLKNAND2HSV1 U11307 ( .A1(n9040), .A2(n13718), .ZN(n9012) );
  INHSV2 U11308 ( .I(\pe20/phq [3]), .ZN(n9013) );
  NAND3HSV2 U11309 ( .A1(\pe20/phq [3]), .A2(\pe20/aot [7]), .A3(\pe20/bq[7] ), 
        .ZN(n9014) );
  BUFHSV8 U11310 ( .I(\pe20/aot [8]), .Z(n13733) );
  XNOR2HSV4 U11311 ( .A1(n9017), .A2(n9016), .ZN(n9018) );
  INHSV4 U11312 ( .I(\pe20/phq [2]), .ZN(n9024) );
  OAI21HSV4 U11313 ( .A1(n9024), .A2(n9023), .B(n9022), .ZN(n9026) );
  INHSV4 U11314 ( .I(n14954), .ZN(n13734) );
  NAND2HSV2 U11315 ( .A1(n13734), .A2(\pe20/aot [7]), .ZN(n9025) );
  XNOR2HSV4 U11316 ( .A1(n9026), .A2(n9025), .ZN(n9030) );
  CLKNAND2HSV0 U11317 ( .A1(\pe20/pvq [2]), .A2(\pe20/ctrq ), .ZN(n9028) );
  XOR2HSV0 U11318 ( .A1(n9028), .A2(n9027), .Z(n9029) );
  XNOR2HSV4 U11319 ( .A1(n9030), .A2(n9029), .ZN(n13848) );
  XNOR2HSV4 U11320 ( .A1(n9032), .A2(n9031), .ZN(n9061) );
  INHSV2 U11321 ( .I(\pe20/got [8]), .ZN(n9034) );
  NOR2HSV2 U11322 ( .A1(n9034), .A2(ctro20), .ZN(n11888) );
  CLKNHSV0 U11323 ( .I(ctro20), .ZN(n13645) );
  INHSV2 U11324 ( .I(n9034), .ZN(n14865) );
  AOI21HSV2 U11325 ( .A1(n9061), .A2(n14865), .B(n15177), .ZN(n9035) );
  XOR2HSV4 U11326 ( .A1(n9058), .A2(n9057), .Z(n9037) );
  CLKNHSV2 U11327 ( .I(n8942), .ZN(n10412) );
  INHSV2 U11328 ( .I(n9034), .ZN(n11880) );
  INHSV2 U11329 ( .I(\pe20/ti_7t [3]), .ZN(n10410) );
  NAND2HSV2 U11330 ( .A1(n10410), .A2(n15177), .ZN(n9465) );
  AOI21HSV4 U11331 ( .A1(n9037), .A2(n10412), .B(n9036), .ZN(n9056) );
  INHSV2 U11332 ( .I(n9038), .ZN(n9039) );
  CLKNHSV2 U11333 ( .I(n9039), .ZN(n9042) );
  CLKNAND2HSV0 U11334 ( .A1(n9040), .A2(\pe20/got [6]), .ZN(n9041) );
  NOR2HSV4 U11335 ( .A1(n9042), .A2(n9041), .ZN(n9052) );
  CLKNHSV2 U11336 ( .I(n9043), .ZN(n9047) );
  NAND2HSV2 U11337 ( .A1(\pe20/bq[5] ), .A2(\pe20/aot [8]), .ZN(n9044) );
  NAND2HSV2 U11338 ( .A1(n13734), .A2(\pe20/aot [5]), .ZN(n9049) );
  NAND2HSV2 U11339 ( .A1(n12362), .A2(\pe20/pvq [4]), .ZN(n9050) );
  INHSV4 U11340 ( .I(n9055), .ZN(n9053) );
  NAND2HSV2 U11341 ( .A1(n8942), .A2(\pe20/ti_7t [4]), .ZN(n9462) );
  CLKNAND2HSV1 U11342 ( .A1(n9465), .A2(n13718), .ZN(n9059) );
  NAND2HSV2 U11343 ( .A1(n13734), .A2(\pe20/aot [4]), .ZN(n9064) );
  NAND2HSV0 U11344 ( .A1(\pe20/aot [5]), .A2(\pe20/bq[7] ), .ZN(n9063) );
  XOR2HSV0 U11345 ( .A1(n9064), .A2(n9063), .Z(n9067) );
  NAND2HSV0 U11346 ( .A1(\pe20/aot [7]), .A2(\pe20/bq[5] ), .ZN(n9066) );
  NAND2HSV0 U11347 ( .A1(\pe20/got [4]), .A2(n13738), .ZN(n9065) );
  BUFHSV8 U11348 ( .I(\pe20/aot [6]), .Z(n14946) );
  NAND2HSV2 U11349 ( .A1(n14946), .A2(\pe20/bq[6] ), .ZN(n9069) );
  CLKNAND2HSV1 U11350 ( .A1(n13733), .A2(\pe20/bq[4] ), .ZN(n9068) );
  INHSV2 U11351 ( .I(n10521), .ZN(n14704) );
  XNOR2HSV4 U11352 ( .A1(n9074), .A2(n9073), .ZN(n9078) );
  BUFHSV4 U11353 ( .I(\pe14/ctrq ), .Z(n14516) );
  CLKNAND2HSV2 U11354 ( .A1(n14516), .A2(\pe14/pvq [3]), .ZN(n9076) );
  NAND2HSV0 U11355 ( .A1(\pe14/bq[7] ), .A2(\pe14/aot [7]), .ZN(n9075) );
  XNOR2HSV4 U11356 ( .A1(n9076), .A2(n9075), .ZN(n9077) );
  XNOR2HSV4 U11357 ( .A1(n9078), .A2(n9077), .ZN(n11037) );
  CLKNAND2HSV1 U11358 ( .A1(\pe14/pvq [1]), .A2(\pe14/ctrq ), .ZN(n9079) );
  INHSV2 U11359 ( .I(\pe14/got [7]), .ZN(n13580) );
  INHSV2 U11360 ( .I(n13580), .ZN(n13085) );
  CLKAND2HSV1 U11361 ( .A1(n11156), .A2(n13085), .Z(n9080) );
  INHSV2 U11362 ( .I(\pe14/ti_7t [1]), .ZN(n9081) );
  NOR2HSV2 U11363 ( .A1(n11156), .A2(n9081), .ZN(n11784) );
  CLKNAND2HSV0 U11364 ( .A1(n11784), .A2(\pe14/got [7]), .ZN(n9082) );
  CLKNAND2HSV4 U11365 ( .A1(n9083), .A2(n9082), .ZN(n11038) );
  XNOR2HSV4 U11366 ( .A1(n11037), .A2(n11038), .ZN(n9100) );
  INHSV2 U11367 ( .I(\pe14/got [8]), .ZN(n13852) );
  NOR2HSV2 U11368 ( .A1(n11093), .A2(n13852), .ZN(n11120) );
  INHSV2 U11369 ( .I(n9084), .ZN(n9092) );
  INHSV4 U11370 ( .I(\pe14/phq [2]), .ZN(n9087) );
  CLKNAND2HSV3 U11371 ( .A1(n9086), .A2(n9087), .ZN(n9085) );
  OAI21HSV4 U11372 ( .A1(n9087), .A2(n9086), .B(n9085), .ZN(n9090) );
  BUFHSV2 U11373 ( .I(\pe14/ctrq ), .Z(n9088) );
  NAND2HSV2 U11374 ( .A1(n9088), .A2(\pe14/pvq [2]), .ZN(n9089) );
  XNOR2HSV4 U11375 ( .A1(n9090), .A2(n9089), .ZN(n9096) );
  XNOR2HSV4 U11376 ( .A1(n9096), .A2(n9095), .ZN(n9091) );
  AOI22HSV4 U11377 ( .A1(n14702), .A2(\pe14/ti_7t [2]), .B1(n9092), .B2(n9091), 
        .ZN(n9099) );
  XNOR2HSV4 U11378 ( .A1(n9094), .A2(n9093), .ZN(n9103) );
  AOI21HSV2 U11379 ( .A1(n15176), .A2(\pe14/got [8]), .B(n11090), .ZN(n9097)
         );
  CLKXOR2HSV4 U11380 ( .A1(n9096), .A2(n9095), .Z(n13854) );
  CLKNAND2HSV2 U11381 ( .A1(n9097), .A2(n13854), .ZN(n9098) );
  CLKNAND2HSV4 U11382 ( .A1(n9099), .A2(n9098), .ZN(n11081) );
  INHSV2 U11383 ( .I(\pe14/ti_7t [3]), .ZN(n11039) );
  NAND2HSV2 U11384 ( .A1(n11090), .A2(n11039), .ZN(n11059) );
  CLKNAND2HSV1 U11385 ( .A1(n11059), .A2(\pe14/got [8]), .ZN(n9101) );
  AOI21HSV4 U11386 ( .A1(n9103), .A2(n8948), .B(n11784), .ZN(n11110) );
  INHSV2 U11387 ( .I(\pe14/got [6]), .ZN(n13059) );
  NOR2HSV4 U11388 ( .A1(n11110), .A2(n13059), .ZN(n9113) );
  NAND2HSV2 U11389 ( .A1(\pe14/got [5]), .A2(\pe14/ti_1 ), .ZN(n9105) );
  NAND2HSV0 U11390 ( .A1(\pe14/bq[8] ), .A2(\pe14/aot [5]), .ZN(n9104) );
  XOR2HSV2 U11391 ( .A1(n9105), .A2(n9104), .Z(n9107) );
  XNOR2HSV4 U11392 ( .A1(n9107), .A2(n9106), .ZN(n9111) );
  NAND2HSV2 U11393 ( .A1(\pe14/aot [6]), .A2(\pe14/bq[7] ), .ZN(n9109) );
  BUFHSV8 U11394 ( .I(\pe14/aot [8]), .Z(n14891) );
  XOR3HSV2 U11395 ( .A1(\pe14/phq [4]), .A2(n9109), .A3(n9108), .Z(n9110) );
  XNOR2HSV4 U11396 ( .A1(n9111), .A2(n9110), .ZN(n9112) );
  XNOR2HSV4 U11397 ( .A1(n9113), .A2(n9112), .ZN(n9115) );
  BUFHSV4 U11398 ( .I(n11081), .Z(n14944) );
  INHSV2 U11399 ( .I(n9629), .ZN(n9680) );
  CLKNAND2HSV2 U11400 ( .A1(\pe4/ti_1 ), .A2(\pe4/got [8]), .ZN(n9117) );
  CLKNAND2HSV2 U11401 ( .A1(\pe4/ctrq ), .A2(\pe4/pvq [1]), .ZN(n9116) );
  XNOR2HSV4 U11402 ( .A1(n9117), .A2(n9116), .ZN(n9612) );
  XNOR2HSV4 U11403 ( .A1(n9612), .A2(n9611), .ZN(n9129) );
  INHSV2 U11404 ( .I(n9629), .ZN(n12597) );
  NOR2HSV2 U11405 ( .A1(n15083), .A2(n12597), .ZN(n10586) );
  INHSV2 U11406 ( .I(n9118), .ZN(n9128) );
  NAND2HSV2 U11407 ( .A1(\pe4/bq[8] ), .A2(\pe4/aot [7]), .ZN(n9121) );
  CLKNAND2HSV2 U11408 ( .A1(\pe4/aot [7]), .A2(\pe4/bq[8] ), .ZN(n9119) );
  CLKNAND2HSV2 U11409 ( .A1(n9119), .A2(\pe4/phq [2]), .ZN(n9120) );
  OAI21HSV4 U11410 ( .A1(n9121), .A2(\pe4/phq [2]), .B(n9120), .ZN(n9123) );
  NAND2HSV0 U11411 ( .A1(\pe4/got [7]), .A2(\pe4/ti_1 ), .ZN(n9122) );
  XNOR2HSV4 U11412 ( .A1(n9123), .A2(n9122), .ZN(n9127) );
  CLKNAND2HSV2 U11413 ( .A1(\pe4/pvq [2]), .A2(\pe4/ctrq ), .ZN(n9124) );
  XOR2HSV2 U11414 ( .A1(n9125), .A2(n9124), .Z(n9126) );
  INHSV2 U11415 ( .I(n9629), .ZN(n10535) );
  AOI21HSV2 U11416 ( .A1(n9129), .A2(\pe4/got [8]), .B(n10535), .ZN(n9130) );
  XNOR2HSV4 U11417 ( .A1(n9132), .A2(n9131), .ZN(n9138) );
  CLKBUFHSV4 U11418 ( .I(ctro18), .Z(n9133) );
  INHSV2 U11419 ( .I(n9133), .ZN(n9217) );
  INHSV2 U11420 ( .I(\pe17/phq [1]), .ZN(n9134) );
  CLKNHSV0 U11421 ( .I(\pe18/ctrq ), .ZN(n10802) );
  BUFHSV2 U11422 ( .I(ctro18), .Z(n13342) );
  CLKNAND2HSV1 U11423 ( .A1(n9139), .A2(n13342), .ZN(n9166) );
  NAND2HSV2 U11424 ( .A1(n9166), .A2(\pe18/got [7]), .ZN(n9140) );
  CLKNAND2HSV3 U11425 ( .A1(n9142), .A2(\pe18/phq [2]), .ZN(n9141) );
  OAI21HSV4 U11426 ( .A1(n9142), .A2(\pe18/phq [2]), .B(n9141), .ZN(n9144) );
  CLKBUFHSV4 U11427 ( .I(\pe18/bq[8] ), .Z(n14511) );
  XNOR2HSV4 U11428 ( .A1(n9144), .A2(n9143), .ZN(n9148) );
  CLKNAND2HSV2 U11429 ( .A1(\pe18/pvq [2]), .A2(\pe18/ctrq ), .ZN(n9146) );
  XOR2HSV2 U11430 ( .A1(n9146), .A2(n9145), .Z(n9147) );
  XNOR2HSV4 U11431 ( .A1(n9148), .A2(n9147), .ZN(n9152) );
  INHSV2 U11432 ( .I(\pe18/got [8]), .ZN(n13141) );
  CLKBUFHSV4 U11433 ( .I(ctro18), .Z(n13146) );
  INHSV2 U11434 ( .I(n9149), .ZN(n12010) );
  CLKAND2HSV2 U11435 ( .A1(n13342), .A2(\pe18/ti_7t [2]), .Z(n9151) );
  CLKNAND2HSV1 U11436 ( .A1(n9200), .A2(\pe18/got [8]), .ZN(n9153) );
  NAND2HSV2 U11437 ( .A1(\pe18/aot [5]), .A2(\pe18/bq[8] ), .ZN(n9156) );
  NAND2HSV0 U11438 ( .A1(\pe18/aot [7]), .A2(\pe18/bq[6] ), .ZN(n9155) );
  XOR2HSV0 U11439 ( .A1(n9156), .A2(n9155), .Z(n9160) );
  XOR2HSV2 U11440 ( .A1(n9160), .A2(n9159), .Z(n9164) );
  BUFHSV8 U11441 ( .I(\pe18/bq[7] ), .Z(n14513) );
  NAND2HSV0 U11442 ( .A1(\pe18/aot [6]), .A2(n14513), .ZN(n9161) );
  XNOR2HSV1 U11443 ( .A1(n9162), .A2(n9161), .ZN(n9163) );
  XNOR2HSV4 U11444 ( .A1(n9169), .A2(n9168), .ZN(n9173) );
  NAND2HSV2 U11445 ( .A1(ctro18), .A2(\pe18/ti_7t [4]), .ZN(n13142) );
  INHSV2 U11446 ( .I(n13142), .ZN(n13140) );
  INHSV2 U11447 ( .I(\pe18/got [7]), .ZN(n9201) );
  AOI21HSV1 U11448 ( .A1(n13142), .A2(n13143), .B(n9201), .ZN(n9174) );
  CLKNAND2HSV0 U11449 ( .A1(\pe18/ti_7[1] ), .A2(\pe18/got [4]), .ZN(n9192) );
  NAND2HSV0 U11450 ( .A1(\pe18/aot [5]), .A2(\pe18/bq[6] ), .ZN(n9176) );
  NAND2HSV0 U11451 ( .A1(\pe18/aot [3]), .A2(\pe18/bq[8] ), .ZN(n9175) );
  XOR2HSV0 U11452 ( .A1(n9176), .A2(n9175), .Z(n9180) );
  NAND2HSV2 U11453 ( .A1(\pe18/aot [7]), .A2(\pe18/bq[4] ), .ZN(n9178) );
  NAND2HSV0 U11454 ( .A1(\pe18/aot [8]), .A2(\pe18/bq[3] ), .ZN(n9177) );
  XOR2HSV0 U11455 ( .A1(n9178), .A2(n9177), .Z(n9179) );
  XOR2HSV2 U11456 ( .A1(n9180), .A2(n9179), .Z(n9184) );
  NAND2HSV2 U11457 ( .A1(\pe18/bq[5] ), .A2(\pe18/aot [6]), .ZN(n9182) );
  BUFHSV8 U11458 ( .I(\pe18/ti_1 ), .Z(n13818) );
  CLKNAND2HSV0 U11459 ( .A1(n13818), .A2(\pe18/got [3]), .ZN(n9181) );
  XOR2HSV0 U11460 ( .A1(n9182), .A2(n9181), .Z(n9183) );
  XNOR2HSV1 U11461 ( .A1(n9184), .A2(n9183), .ZN(n9189) );
  XNOR2HSV1 U11462 ( .A1(n9185), .A2(\pe18/phq [6]), .ZN(n9187) );
  CLKNAND2HSV0 U11463 ( .A1(\pe18/aot [4]), .A2(n14513), .ZN(n9186) );
  XNOR2HSV1 U11464 ( .A1(n9187), .A2(n9186), .ZN(n9188) );
  NAND2HSV2 U11465 ( .A1(n11996), .A2(\pe18/got [5]), .ZN(n9190) );
  XOR3HSV2 U11466 ( .A1(n9192), .A2(n9191), .A3(n9190), .Z(n9197) );
  NAND2HSV2 U11467 ( .A1(n9133), .A2(\pe18/ti_7t [3]), .ZN(n9455) );
  CLKNHSV0 U11468 ( .I(n9455), .ZN(n9195) );
  INHSV2 U11469 ( .I(n6039), .ZN(n13147) );
  AOI21HSV1 U11470 ( .A1(ctro18), .A2(n9455), .B(n13147), .ZN(n9194) );
  OAI21HSV2 U11471 ( .A1(n15218), .A2(n9195), .B(n9194), .ZN(n9196) );
  XNOR2HSV1 U11472 ( .A1(n9197), .A2(n9196), .ZN(n9198) );
  XNOR2HSV4 U11473 ( .A1(n9199), .A2(n9198), .ZN(n9220) );
  XNOR2HSV1 U11474 ( .A1(n9202), .A2(\pe18/phq [5]), .ZN(n9213) );
  INHSV2 U11475 ( .I(\pe18/aot [8]), .ZN(n9203) );
  NAND2HSV0 U11476 ( .A1(n11988), .A2(\pe18/bq[4] ), .ZN(n9205) );
  CLKNHSV1 U11477 ( .I(\pe18/aot [7]), .ZN(n14625) );
  INHSV2 U11478 ( .I(\pe18/bq[5] ), .ZN(n14563) );
  NOR2HSV2 U11479 ( .A1(n14625), .A2(n14563), .ZN(n9204) );
  XOR2HSV2 U11480 ( .A1(n9205), .A2(n9204), .Z(n9212) );
  NAND2HSV0 U11481 ( .A1(\pe18/got [4]), .A2(\pe18/ti_1 ), .ZN(n9207) );
  NAND2HSV0 U11482 ( .A1(\pe18/aot [6]), .A2(\pe18/bq[6] ), .ZN(n9206) );
  XOR2HSV2 U11483 ( .A1(n9207), .A2(n9206), .Z(n9211) );
  NAND2HSV0 U11484 ( .A1(\pe18/aot [4]), .A2(n14511), .ZN(n9209) );
  NAND2HSV0 U11485 ( .A1(n14513), .A2(\pe18/aot [5]), .ZN(n9208) );
  XOR2HSV2 U11486 ( .A1(n9209), .A2(n9208), .Z(n9210) );
  XOR4HSV2 U11487 ( .A1(n9213), .A2(n9212), .A3(n9211), .A4(n9210), .Z(n9214)
         );
  NAND2HSV2 U11488 ( .A1(n6039), .A2(n11996), .ZN(n9215) );
  NOR2HSV2 U11489 ( .A1(n9217), .A2(\pe18/ti_7t [5]), .ZN(n13346) );
  NOR2HSV2 U11490 ( .A1(n13346), .A2(n13141), .ZN(n9218) );
  XNOR2HSV4 U11491 ( .A1(n9220), .A2(n9219), .ZN(n15215) );
  NAND2HSV2 U11492 ( .A1(\pe6/aot [7]), .A2(\pe6/bq[7] ), .ZN(n9222) );
  XOR2HSV4 U11493 ( .A1(n9222), .A2(n9221), .Z(n9226) );
  NAND2HSV2 U11494 ( .A1(\pe6/aot [8]), .A2(\pe6/bq[6] ), .ZN(n9224) );
  CLKNAND2HSV2 U11495 ( .A1(\pe6/aot [6]), .A2(\pe6/bq[8] ), .ZN(n9223) );
  XOR2HSV4 U11496 ( .A1(n9224), .A2(n9223), .Z(n9225) );
  XNOR2HSV4 U11497 ( .A1(n9226), .A2(n9225), .ZN(n9229) );
  BUFHSV8 U11498 ( .I(n8935), .Z(n13041) );
  NAND2HSV2 U11499 ( .A1(n13041), .A2(\pe6/pvq [3]), .ZN(n9227) );
  XOR2HSV0 U11500 ( .A1(n9227), .A2(\pe6/phq [3]), .Z(n9228) );
  CLKNAND2HSV2 U11501 ( .A1(\pe6/ctrq ), .A2(\pe6/pvq [1]), .ZN(n9230) );
  XNOR2HSV4 U11502 ( .A1(n9231), .A2(n9230), .ZN(n11950) );
  XNOR2HSV4 U11503 ( .A1(n11950), .A2(n11949), .ZN(n9242) );
  INHSV4 U11504 ( .I(ctro6), .ZN(n10799) );
  INHSV2 U11505 ( .I(n10799), .ZN(n9802) );
  NOR2HSV4 U11506 ( .A1(n9242), .A2(n9802), .ZN(n9244) );
  OAI21HSV0 U11507 ( .A1(n10799), .A2(\pe6/ti_7t [1]), .B(\pe6/got [7]), .ZN(
        n9232) );
  INHSV2 U11508 ( .I(n14863), .ZN(n13829) );
  NAND2HSV2 U11509 ( .A1(n13829), .A2(\pe6/aot [7]), .ZN(n9234) );
  CLKNAND2HSV2 U11510 ( .A1(n8925), .A2(\pe6/pvq [2]), .ZN(n9233) );
  INHSV2 U11511 ( .I(n8912), .ZN(n9241) );
  INHSV4 U11512 ( .I(\pe6/phq [2]), .ZN(n9237) );
  CLKNAND2HSV3 U11513 ( .A1(n9236), .A2(n9237), .ZN(n9235) );
  OAI21HSV4 U11514 ( .A1(n9237), .A2(n9236), .B(n9235), .ZN(n9239) );
  CLKNHSV2 U11515 ( .I(n9251), .ZN(n9238) );
  XNOR2HSV4 U11516 ( .A1(n9239), .A2(n9238), .ZN(n9240) );
  INHSV4 U11517 ( .I(ctro6), .ZN(n9285) );
  NOR2HSV2 U11518 ( .A1(n10799), .A2(\pe6/ti_7t [2]), .ZN(n9291) );
  NOR2HSV2 U11519 ( .A1(n9291), .A2(n15095), .ZN(n9243) );
  CLKNAND2HSV1 U11520 ( .A1(n6725), .A2(n9244), .ZN(n9245) );
  INHSV2 U11521 ( .I(n9245), .ZN(n9246) );
  CLKNHSV3 U11522 ( .I(n9285), .ZN(n9842) );
  NAND2HSV2 U11523 ( .A1(\pe6/pvq [4]), .A2(n8925), .ZN(n9250) );
  NAND2HSV0 U11524 ( .A1(\pe6/got [5]), .A2(\pe6/ti_1 ), .ZN(n9249) );
  XOR2HSV2 U11525 ( .A1(n9250), .A2(n9249), .Z(n9256) );
  NOR2HSV2 U11526 ( .A1(n9251), .A2(n9298), .ZN(n9254) );
  INHSV4 U11527 ( .I(n14885), .ZN(n9252) );
  AOI22HSV0 U11528 ( .A1(n9252), .A2(\pe6/bq[5] ), .B1(\pe6/bq[7] ), .B2(
        \pe6/aot [6]), .ZN(n9253) );
  NOR2HSV2 U11529 ( .A1(n9254), .A2(n9253), .ZN(n9255) );
  XNOR2HSV4 U11530 ( .A1(n9257), .A2(\pe6/phq [4]), .ZN(n9259) );
  NAND2HSV0 U11531 ( .A1(\pe6/aot [7]), .A2(\pe6/bq[6] ), .ZN(n9258) );
  XNOR2HSV4 U11532 ( .A1(n9259), .A2(n9258), .ZN(n9260) );
  INHSV1 U11533 ( .I(n9291), .ZN(n9266) );
  NAND2HSV0 U11534 ( .A1(n9266), .A2(n5977), .ZN(n9261) );
  CLKNHSV0 U11535 ( .I(n9285), .ZN(n15088) );
  CLKAND2HSV1 U11536 ( .A1(n9312), .A2(\pe6/got [8]), .Z(n9264) );
  BUFHSV2 U11537 ( .I(\pe6/got [8]), .Z(n13897) );
  NAND2HSV0 U11538 ( .A1(n9266), .A2(\pe6/got [6]), .ZN(n9267) );
  NAND2HSV2 U11539 ( .A1(\pe6/aot [6]), .A2(\pe6/bq[6] ), .ZN(n9271) );
  NAND2HSV0 U11540 ( .A1(\pe6/bq[4] ), .A2(\pe6/aot [8]), .ZN(n9270) );
  XOR2HSV0 U11541 ( .A1(n9271), .A2(n9270), .Z(n9275) );
  NAND2HSV0 U11542 ( .A1(\pe6/aot [7]), .A2(\pe6/bq[5] ), .ZN(n9273) );
  NAND2HSV0 U11543 ( .A1(\pe6/got [4]), .A2(\pe6/ti_1 ), .ZN(n9272) );
  XOR2HSV0 U11544 ( .A1(n9273), .A2(n9272), .Z(n9274) );
  XOR2HSV0 U11545 ( .A1(n9275), .A2(n9274), .Z(n9281) );
  NAND2HSV0 U11546 ( .A1(\pe6/aot [5]), .A2(\pe6/bq[7] ), .ZN(n9277) );
  NAND2HSV0 U11547 ( .A1(\pe6/aot [4]), .A2(\pe6/bq[8] ), .ZN(n9276) );
  XOR2HSV0 U11548 ( .A1(n9277), .A2(n9276), .Z(n9279) );
  CLKXOR2HSV4 U11549 ( .A1(n9279), .A2(n9278), .Z(n9280) );
  XOR2HSV4 U11550 ( .A1(n9281), .A2(n9280), .Z(n9283) );
  NAND2HSV2 U11551 ( .A1(n9823), .A2(\pe6/got [5]), .ZN(n9282) );
  INHSV2 U11552 ( .I(n9285), .ZN(n9798) );
  INHSV2 U11553 ( .I(n9798), .ZN(n9536) );
  OAI21HSV0 U11554 ( .A1(n9832), .A2(\pe6/ti_7t [5]), .B(n13897), .ZN(n9286)
         );
  AOI21HSV2 U11555 ( .A1(n9287), .A2(n9536), .B(n9286), .ZN(n9320) );
  NAND2HSV2 U11556 ( .A1(n9287), .A2(n9832), .ZN(n9289) );
  CLKNAND2HSV2 U11557 ( .A1(n9289), .A2(n9288), .ZN(n9319) );
  INHSV2 U11558 ( .I(\pe6/got [6]), .ZN(n12410) );
  CLKNHSV0 U11559 ( .I(\pe6/got [5]), .ZN(n9290) );
  NOR2HSV1 U11560 ( .A1(n9291), .A2(n9290), .ZN(n9307) );
  AND2HSV2 U11561 ( .A1(n9307), .A2(ctro6), .Z(n9303) );
  CLKNHSV0 U11562 ( .I(n9307), .ZN(n9302) );
  NAND2HSV0 U11563 ( .A1(\pe6/aot [7]), .A2(\pe6/bq[4] ), .ZN(n9293) );
  CLKNAND2HSV1 U11564 ( .A1(\pe6/aot [3]), .A2(\pe6/bq[8] ), .ZN(n9292) );
  XOR2HSV0 U11565 ( .A1(n9293), .A2(n9292), .Z(n9297) );
  NAND2HSV0 U11566 ( .A1(\pe6/aot [8]), .A2(\pe6/bq[3] ), .ZN(n9295) );
  NAND2HSV0 U11567 ( .A1(\pe6/aot [5]), .A2(\pe6/bq[6] ), .ZN(n9294) );
  XOR2HSV0 U11568 ( .A1(n9295), .A2(n9294), .Z(n9296) );
  XOR2HSV0 U11569 ( .A1(n9297), .A2(n9296), .Z(n9301) );
  NAND2HSV2 U11570 ( .A1(\pe6/aot [4]), .A2(\pe6/bq[7] ), .ZN(n12416) );
  INHSV2 U11571 ( .I(n6724), .ZN(n9305) );
  XNOR2HSV4 U11572 ( .A1(n9306), .A2(n9305), .ZN(n10800) );
  INHSV2 U11573 ( .I(n10800), .ZN(n15071) );
  NAND2HSV0 U11574 ( .A1(n13105), .A2(n9832), .ZN(n9309) );
  CLKNHSV0 U11575 ( .I(n9309), .ZN(n9311) );
  CLKNAND2HSV1 U11576 ( .A1(n9832), .A2(n13897), .ZN(n9840) );
  NOR2HSV0 U11577 ( .A1(n13105), .A2(n9840), .ZN(n9310) );
  MUX2NHSV2 U11578 ( .I0(n9311), .I1(n9310), .S(n13057), .ZN(n9315) );
  NOR2HSV0 U11579 ( .A1(ctro6), .A2(\pe6/got [8]), .ZN(n9843) );
  CLKNAND2HSV0 U11580 ( .A1(n9312), .A2(n5977), .ZN(n9313) );
  AOI21HSV2 U11581 ( .A1(n7521), .A2(n9843), .B(n9313), .ZN(n9314) );
  CLKNAND2HSV2 U11582 ( .A1(n9315), .A2(n9314), .ZN(n9316) );
  XNOR2HSV4 U11583 ( .A1(n9317), .A2(n9316), .ZN(n9318) );
  NAND2HSV2 U11584 ( .A1(n9358), .A2(\pe2/ti_7t [4]), .ZN(n10709) );
  INHSV2 U11585 ( .I(n10709), .ZN(n10711) );
  AOI21HSV2 U11586 ( .A1(n10709), .A2(n9358), .B(n9360), .ZN(n9321) );
  OAI21HSV4 U11587 ( .A1(n15070), .A2(n10711), .B(n9321), .ZN(n9357) );
  NAND2HSV0 U11588 ( .A1(\pe2/aot [6]), .A2(\pe2/bq[5] ), .ZN(n9323) );
  NAND2HSV0 U11589 ( .A1(\pe2/aot [7]), .A2(\pe2/bq[4] ), .ZN(n9322) );
  XOR2HSV0 U11590 ( .A1(n9323), .A2(n9322), .Z(n9337) );
  XNOR2HSV4 U11591 ( .A1(n9325), .A2(\pe2/phq [6]), .ZN(n9327) );
  CLKNAND2HSV0 U11592 ( .A1(\pe2/aot [5]), .A2(\pe2/bq[6] ), .ZN(n9326) );
  XNOR2HSV4 U11593 ( .A1(n9327), .A2(n9326), .ZN(n9336) );
  NAND2HSV0 U11594 ( .A1(\pe2/aot [3]), .A2(\pe2/bq[8] ), .ZN(n9330) );
  NAND2HSV0 U11595 ( .A1(\pe2/ti_1 ), .A2(\pe2/got [3]), .ZN(n9332) );
  NAND2HSV0 U11596 ( .A1(\pe2/aot [4]), .A2(\pe2/bq[7] ), .ZN(n9331) );
  XOR2HSV0 U11597 ( .A1(n9332), .A2(n9331), .Z(n9333) );
  XOR3HSV2 U11598 ( .A1(n9337), .A2(n9336), .A3(n9335), .Z(n9340) );
  CLKNAND2HSV0 U11599 ( .A1(\pe2/ti_7[1] ), .A2(\pe2/got [4]), .ZN(n9339) );
  XNOR2HSV4 U11600 ( .A1(n9340), .A2(n9339), .ZN(n9344) );
  BUFHSV8 U11601 ( .I(n9345), .Z(n13762) );
  XNOR2HSV4 U11602 ( .A1(n9344), .A2(n9343), .ZN(n9355) );
  XNOR2HSV4 U11603 ( .A1(n9347), .A2(n9346), .ZN(n10797) );
  NAND2HSV0 U11604 ( .A1(n9359), .A2(n14822), .ZN(n9349) );
  NOR2HSV2 U11605 ( .A1(n9348), .A2(n9349), .ZN(n9354) );
  CLKNHSV2 U11606 ( .I(n9363), .ZN(n9350) );
  INHSV1 U11607 ( .I(n9350), .ZN(n9353) );
  NOR2HSV2 U11608 ( .A1(n9350), .A2(n9349), .ZN(n9351) );
  AOI31HSV2 U11609 ( .A1(n9355), .A2(n9354), .A3(n9353), .B(n9352), .ZN(n9356)
         );
  XNOR2HSV4 U11610 ( .A1(n9357), .A2(n9356), .ZN(n9383) );
  NOR2HSV4 U11611 ( .A1(n13795), .A2(n9358), .ZN(n9382) );
  CLKNHSV0 U11612 ( .I(n9359), .ZN(n9361) );
  NOR2HSV1 U11613 ( .A1(n9361), .A2(n9360), .ZN(n9362) );
  CLKNAND2HSV0 U11614 ( .A1(\pe2/aot [7]), .A2(\pe2/bq[5] ), .ZN(n9366) );
  NAND2HSV0 U11615 ( .A1(\pe2/aot [4]), .A2(\pe2/bq[8] ), .ZN(n9365) );
  XOR2HSV0 U11616 ( .A1(n9366), .A2(n9365), .Z(n9370) );
  CLKNAND2HSV1 U11617 ( .A1(\pe2/aot [6]), .A2(\pe2/bq[6] ), .ZN(n9368) );
  XOR2HSV0 U11618 ( .A1(n9370), .A2(n9369), .Z(n9376) );
  CLKNAND2HSV0 U11619 ( .A1(\pe2/ctrq ), .A2(\pe2/pvq [5]), .ZN(n9372) );
  XOR2HSV0 U11620 ( .A1(n9372), .A2(\pe2/phq [5]), .Z(n9373) );
  XOR2HSV0 U11621 ( .A1(n9374), .A2(n9373), .Z(n9375) );
  NOR2HSV1 U11622 ( .A1(n9378), .A2(\pe2/ti_7t [5]), .ZN(n11261) );
  NOR2HSV1 U11623 ( .A1(n11261), .A2(n10708), .ZN(n9384) );
  INHSV2 U11624 ( .I(n9384), .ZN(n9379) );
  NAND2HSV2 U11625 ( .A1(n9383), .A2(n8914), .ZN(n9392) );
  AND2HSV2 U11626 ( .A1(n9384), .A2(n9378), .Z(n9385) );
  INAND2HSV2 U11627 ( .A1(n11267), .B1(n11266), .ZN(n9387) );
  INHSV2 U11628 ( .I(n9387), .ZN(n9389) );
  AOI22HSV4 U11629 ( .A1(n9390), .A2(n8914), .B1(n9389), .B2(n9388), .ZN(n9391) );
  XNOR2HSV4 U11630 ( .A1(n9394), .A2(n9393), .ZN(n10371) );
  INHSV2 U11631 ( .I(\pe21/phq [1]), .ZN(n9395) );
  CLKNAND2HSV3 U11632 ( .A1(n9397), .A2(n9396), .ZN(n10370) );
  BUFHSV2 U11633 ( .I(ctro21), .Z(n11780) );
  NAND2HSV2 U11634 ( .A1(n10874), .A2(\pe21/ti_7t [1]), .ZN(n10385) );
  NAND2HSV2 U11635 ( .A1(n9734), .A2(\pe9/ti_7t [3]), .ZN(n10441) );
  CLKNAND2HSV1 U11636 ( .A1(\pe9/ti_7[1] ), .A2(\pe9/got [4]), .ZN(n9416) );
  BUFHSV8 U11637 ( .I(\pe9/bq[7] ), .Z(n13911) );
  NAND2HSV0 U11638 ( .A1(\pe9/aot [4]), .A2(n5976), .ZN(n9402) );
  NAND2HSV0 U11639 ( .A1(\pe9/aot [6]), .A2(\pe9/bq[5] ), .ZN(n9401) );
  XOR2HSV0 U11640 ( .A1(n9402), .A2(n9401), .Z(n9413) );
  NAND2HSV2 U11641 ( .A1(n13826), .A2(\pe9/pvq [6]), .ZN(n9403) );
  XNOR2HSV1 U11642 ( .A1(n9403), .A2(\pe9/phq [6]), .ZN(n9404) );
  INHSV2 U11643 ( .I(n6303), .ZN(n9438) );
  INHSV2 U11644 ( .I(\pe9/bq[4] ), .ZN(n9772) );
  NOR2HSV4 U11645 ( .A1(n9438), .A2(n9772), .ZN(n13920) );
  XNOR2HSV1 U11646 ( .A1(n9404), .A2(n13920), .ZN(n9412) );
  NAND2HSV0 U11647 ( .A1(\pe9/aot [3]), .A2(\pe9/bq[8] ), .ZN(n9406) );
  BUFHSV2 U11648 ( .I(\pe9/bq[6] ), .Z(n11647) );
  NAND2HSV0 U11649 ( .A1(n11647), .A2(\pe9/aot [5]), .ZN(n9405) );
  XOR2HSV0 U11650 ( .A1(n9406), .A2(n9405), .Z(n9410) );
  BUFHSV2 U11651 ( .I(\pe9/aot [8]), .Z(n14942) );
  NAND2HSV2 U11652 ( .A1(n14942), .A2(\pe9/bq[3] ), .ZN(n9408) );
  NAND2HSV2 U11653 ( .A1(n8944), .A2(\pe9/got [3]), .ZN(n9407) );
  XOR2HSV0 U11654 ( .A1(n9408), .A2(n9407), .Z(n9409) );
  XOR2HSV0 U11655 ( .A1(n9410), .A2(n9409), .Z(n9411) );
  XOR3HSV2 U11656 ( .A1(n9413), .A2(n9412), .A3(n9411), .Z(n9415) );
  XOR3HSV2 U11657 ( .A1(n9416), .A2(n9415), .A3(n9414), .Z(n9417) );
  XNOR2HSV4 U11658 ( .A1(n9418), .A2(n9417), .ZN(n9436) );
  INHSV2 U11659 ( .I(n14866), .ZN(n9739) );
  NAND2HSV0 U11660 ( .A1(\pe9/aot [6]), .A2(\pe9/bq[7] ), .ZN(n9423) );
  NAND2HSV0 U11661 ( .A1(\pe9/aot [5]), .A2(\pe9/bq[8] ), .ZN(n9422) );
  XOR2HSV0 U11662 ( .A1(n9423), .A2(n9422), .Z(n9427) );
  NAND2HSV0 U11663 ( .A1(\pe9/aot [7]), .A2(\pe9/bq[6] ), .ZN(n9425) );
  XOR2HSV0 U11664 ( .A1(n9425), .A2(n9424), .Z(n9426) );
  CLKNAND2HSV2 U11665 ( .A1(n14942), .A2(\pe9/bq[5] ), .ZN(n9440) );
  CLKNAND2HSV0 U11666 ( .A1(n9429), .A2(\pe9/got [6]), .ZN(n9431) );
  NOR2HSV0 U11667 ( .A1(n9736), .A2(ctro9), .ZN(n9435) );
  BUFHSV2 U11668 ( .I(n9744), .Z(n15069) );
  CLKNAND2HSV2 U11669 ( .A1(n13826), .A2(\pe9/pvq [5]), .ZN(n9437) );
  XNOR2HSV1 U11670 ( .A1(n9437), .A2(\pe9/phq [5]), .ZN(n9442) );
  INHSV1 U11671 ( .I(n13920), .ZN(n9441) );
  NAND2HSV0 U11672 ( .A1(\pe9/aot [4]), .A2(\pe9/bq[8] ), .ZN(n9767) );
  NAND2HSV2 U11673 ( .A1(n13911), .A2(\pe9/aot [5]), .ZN(n9443) );
  NAND2HSV0 U11674 ( .A1(\pe9/got [4]), .A2(\pe9/ti_1 ), .ZN(n9444) );
  XOR2HSV0 U11675 ( .A1(n9445), .A2(n9444), .Z(n9446) );
  NAND2HSV0 U11676 ( .A1(n9783), .A2(\pe9/got [6]), .ZN(n9447) );
  CLKNHSV1 U11677 ( .I(ctro9), .ZN(n9450) );
  INHSV1 U11678 ( .I(\pe9/ti_7t [5]), .ZN(n9452) );
  AOI21HSV2 U11679 ( .A1(n9452), .A2(n9790), .B(n9451), .ZN(n9453) );
  INHSV2 U11680 ( .I(\pe9/ti_7t [6]), .ZN(n13931) );
  NAND2HSV2 U11681 ( .A1(n13931), .A2(n14866), .ZN(n9791) );
  INHSV2 U11682 ( .I(n9791), .ZN(n11668) );
  CLKNHSV0 U11683 ( .I(\pe20/ti_7t [5]), .ZN(n9458) );
  CLKNAND2HSV1 U11684 ( .A1(n9458), .A2(n15177), .ZN(n13641) );
  CLKNAND2HSV0 U11685 ( .A1(n13641), .A2(n11880), .ZN(n10592) );
  CLKNAND2HSV2 U11686 ( .A1(n12048), .A2(n8939), .ZN(n9460) );
  NOR2HSV4 U11687 ( .A1(n9460), .A2(n9459), .ZN(n10594) );
  CLKNHSV1 U11688 ( .I(n9462), .ZN(n9464) );
  AOI21HSV2 U11689 ( .A1(n9462), .A2(n15177), .B(n9461), .ZN(n9463) );
  OAI21HSV4 U11690 ( .A1(n14821), .A2(n9464), .B(n9463), .ZN(n9487) );
  CLKNAND2HSV0 U11691 ( .A1(n9465), .A2(\pe20/got [6]), .ZN(n9466) );
  CLKNHSV2 U11692 ( .I(n9466), .ZN(n9467) );
  CLKNAND2HSV0 U11693 ( .A1(\pe20/pvq [6]), .A2(n12362), .ZN(n9468) );
  CLKNAND2HSV1 U11694 ( .A1(n13733), .A2(\pe20/bq[3] ), .ZN(n9469) );
  XNOR2HSV4 U11695 ( .A1(n9470), .A2(n9469), .ZN(n9474) );
  NAND2HSV0 U11696 ( .A1(n14946), .A2(\pe20/bq[5] ), .ZN(n9472) );
  NAND2HSV0 U11697 ( .A1(\pe20/aot [7]), .A2(\pe20/bq[4] ), .ZN(n9471) );
  XOR2HSV0 U11698 ( .A1(n9472), .A2(n9471), .Z(n9473) );
  XNOR2HSV4 U11699 ( .A1(n9474), .A2(n9473), .ZN(n9484) );
  NAND2HSV0 U11700 ( .A1(\pe20/aot [3]), .A2(\pe20/bq[8] ), .ZN(n9475) );
  XOR2HSV0 U11701 ( .A1(n9476), .A2(n9475), .Z(n9478) );
  NAND2HSV0 U11702 ( .A1(\pe20/aot [4]), .A2(\pe20/bq[7] ), .ZN(n9477) );
  XOR3HSV2 U11703 ( .A1(n9484), .A2(n9483), .A3(n9482), .Z(n9485) );
  XNOR2HSV4 U11704 ( .A1(n9487), .A2(n9486), .ZN(n10598) );
  XNOR2HSV4 U11705 ( .A1(n9512), .A2(n9511), .ZN(n9500) );
  INHSV2 U11706 ( .I(\pe19/ti_7t [1]), .ZN(n9488) );
  NOR2HSV2 U11707 ( .A1(n9541), .A2(n9488), .ZN(n9489) );
  NOR2HSV4 U11708 ( .A1(n9500), .A2(n9489), .ZN(n9527) );
  INHSV2 U11709 ( .I(n9489), .ZN(n9556) );
  INHSV2 U11710 ( .I(n9541), .ZN(n12172) );
  NAND2HSV2 U11711 ( .A1(n9556), .A2(n14700), .ZN(n9525) );
  CLKNAND2HSV1 U11712 ( .A1(n9525), .A2(\pe19/got [7]), .ZN(n9490) );
  NOR2HSV4 U11713 ( .A1(n9527), .A2(n9490), .ZN(n9499) );
  CLKBUFHSV4 U11714 ( .I(\pe19/aot [8]), .Z(n14915) );
  NAND2HSV2 U11715 ( .A1(n14915), .A2(\pe19/bq[6] ), .ZN(n9497) );
  XNOR2HSV4 U11716 ( .A1(n9491), .A2(\pe19/phq [3]), .ZN(n9496) );
  BUFHSV6 U11717 ( .I(\pe19/bq[8] ), .Z(n14506) );
  NAND2HSV2 U11718 ( .A1(n14506), .A2(\pe19/aot [6]), .ZN(n9495) );
  NAND2HSV2 U11719 ( .A1(\pe19/bq[7] ), .A2(\pe19/aot [7]), .ZN(n9492) );
  XNOR2HSV4 U11720 ( .A1(n9493), .A2(n9492), .ZN(n9494) );
  XOR4HSV2 U11721 ( .A1(n9497), .A2(n9496), .A3(n9495), .A4(n9494), .Z(n9498)
         );
  INHSV4 U11722 ( .I(\pe19/got [8]), .ZN(n12135) );
  INHSV2 U11723 ( .I(n12135), .ZN(n13844) );
  INHSV2 U11724 ( .I(n9541), .ZN(n9721) );
  CLKNAND2HSV4 U11725 ( .A1(\pe19/aot [7]), .A2(\pe19/bq[8] ), .ZN(n9503) );
  INHSV4 U11726 ( .I(\pe19/phq [2]), .ZN(n9502) );
  CLKNAND2HSV3 U11727 ( .A1(n9503), .A2(n9502), .ZN(n9501) );
  OAI21HSV4 U11728 ( .A1(n9502), .A2(n9503), .B(n9501), .ZN(n9506) );
  NAND2HSV0 U11729 ( .A1(\pe19/aot [8]), .A2(\pe19/bq[7] ), .ZN(n9504) );
  INHSV2 U11730 ( .I(n9504), .ZN(n9505) );
  XNOR2HSV4 U11731 ( .A1(n9506), .A2(n9505), .ZN(n9510) );
  NAND2HSV2 U11732 ( .A1(\pe19/ti_1 ), .A2(\pe19/got [7]), .ZN(n9508) );
  NAND2HSV0 U11733 ( .A1(\pe19/ctrq ), .A2(\pe19/pvq [2]), .ZN(n9507) );
  XOR2HSV0 U11734 ( .A1(n9508), .A2(n9507), .Z(n9509) );
  XNOR2HSV4 U11735 ( .A1(n9510), .A2(n9509), .ZN(n9514) );
  OR2HSV1 U11736 ( .A1(n12135), .A2(n14700), .Z(n9513) );
  NOR2HSV0 U11737 ( .A1(n9541), .A2(\pe19/ti_7t [3]), .ZN(n9542) );
  NOR2HSV2 U11738 ( .A1(n9542), .A2(n12135), .ZN(n9722) );
  NAND2HSV2 U11739 ( .A1(n9581), .A2(\pe19/got [7]), .ZN(n9532) );
  NAND2HSV2 U11740 ( .A1(\pe19/bq[8] ), .A2(\pe19/aot [5]), .ZN(n9519) );
  NAND2HSV0 U11741 ( .A1(\pe19/got [5]), .A2(\pe19/ti_1 ), .ZN(n9518) );
  XOR3HSV2 U11742 ( .A1(\pe19/phq [4]), .A2(n9519), .A3(n9518), .Z(n9530) );
  NAND2HSV0 U11743 ( .A1(\pe19/ctrq ), .A2(\pe19/pvq [4]), .ZN(n9520) );
  XNOR2HSV2 U11744 ( .A1(n12152), .A2(n9520), .ZN(n9524) );
  NAND2HSV0 U11745 ( .A1(\pe19/aot [6]), .A2(\pe19/bq[7] ), .ZN(n9522) );
  NAND2HSV0 U11746 ( .A1(\pe19/aot [7]), .A2(\pe19/bq[6] ), .ZN(n9521) );
  XOR2HSV2 U11747 ( .A1(n9522), .A2(n9521), .Z(n9523) );
  XNOR2HSV4 U11748 ( .A1(n9524), .A2(n9523), .ZN(n9529) );
  NAND2HSV0 U11749 ( .A1(n9525), .A2(\pe19/got [6]), .ZN(n9526) );
  NOR2HSV4 U11750 ( .A1(n9527), .A2(n9526), .ZN(n9528) );
  XNOR3HSV2 U11751 ( .A1(n9530), .A2(n9529), .A3(n9528), .ZN(n9531) );
  CLKNAND2HSV1 U11752 ( .A1(ctro6), .A2(\pe6/ti_7t [5]), .ZN(n9799) );
  CLKNHSV0 U11753 ( .I(n9722), .ZN(n9538) );
  NOR2HSV2 U11754 ( .A1(n9538), .A2(n9721), .ZN(n9539) );
  NAND3HSV3 U11755 ( .A1(n9727), .A2(n9725), .A3(n9539), .ZN(n9730) );
  INHSV2 U11756 ( .I(n9541), .ZN(n10357) );
  INHSV2 U11757 ( .I(\pe19/got [7]), .ZN(n12139) );
  NOR2HSV2 U11758 ( .A1(n9542), .A2(n12139), .ZN(n9543) );
  NAND2HSV2 U11759 ( .A1(\pe19/bq[6] ), .A2(\pe19/aot [6]), .ZN(n9545) );
  NAND2HSV0 U11760 ( .A1(\pe19/aot [8]), .A2(\pe19/bq[4] ), .ZN(n9544) );
  XOR2HSV0 U11761 ( .A1(n9545), .A2(n9544), .Z(n9549) );
  NAND2HSV0 U11762 ( .A1(\pe19/got [4]), .A2(\pe19/ti_1 ), .ZN(n9547) );
  NAND2HSV0 U11763 ( .A1(\pe19/aot [4]), .A2(\pe19/bq[8] ), .ZN(n9546) );
  XOR2HSV0 U11764 ( .A1(n9547), .A2(n9546), .Z(n9548) );
  XOR2HSV0 U11765 ( .A1(n9549), .A2(n9548), .Z(n9554) );
  CLKNHSV0 U11766 ( .I(\pe19/aot [5]), .ZN(n15099) );
  NAND2HSV0 U11767 ( .A1(\pe19/ctrq ), .A2(\pe19/pvq [5]), .ZN(n9550) );
  XOR2HSV0 U11768 ( .A1(n9550), .A2(\pe19/phq [5]), .Z(n9551) );
  NAND2HSV0 U11769 ( .A1(\pe19/ti_7[1] ), .A2(\pe19/got [5]), .ZN(n9557) );
  INHSV2 U11770 ( .I(n9558), .ZN(n9559) );
  CLKAND2HSV1 U11771 ( .A1(n12138), .A2(n13844), .Z(n9561) );
  OAI21HSV2 U11772 ( .A1(n10356), .A2(n9562), .B(n9561), .ZN(n9563) );
  INHSV2 U11773 ( .I(\pe19/ti_7t [4]), .ZN(n9564) );
  NOR2HSV2 U11774 ( .A1(n9541), .A2(n9564), .ZN(n9565) );
  INHSV2 U11775 ( .I(n9565), .ZN(n9723) );
  NAND2HSV2 U11776 ( .A1(n14700), .A2(\pe19/ti_7t [3]), .ZN(n10468) );
  INAND2HSV2 U11777 ( .A1(n15212), .B1(n10468), .ZN(n9585) );
  NAND3HSV0 U11778 ( .A1(n15212), .A2(\pe19/got [6]), .A3(n9541), .ZN(n9584)
         );
  CLKBUFHSV4 U11779 ( .I(\pe19/bq[7] ), .Z(n14576) );
  CLKNAND2HSV1 U11780 ( .A1(\pe19/aot [4]), .A2(n14576), .ZN(n9567) );
  CLKBUFHSV4 U11781 ( .I(\pe19/aot [5]), .Z(n13317) );
  NAND2HSV0 U11782 ( .A1(n13317), .A2(\pe19/bq[6] ), .ZN(n9566) );
  XOR2HSV0 U11783 ( .A1(n9567), .A2(n9566), .Z(n9578) );
  NAND2HSV0 U11784 ( .A1(n14506), .A2(\pe19/aot [3]), .ZN(n9568) );
  XNOR2HSV1 U11785 ( .A1(n9569), .A2(n9568), .ZN(n9577) );
  NAND2HSV0 U11786 ( .A1(\pe19/got [3]), .A2(\pe19/ti_1 ), .ZN(n9571) );
  NAND2HSV0 U11787 ( .A1(\pe19/aot [7]), .A2(\pe19/bq[4] ), .ZN(n9570) );
  XOR2HSV0 U11788 ( .A1(n9571), .A2(n9570), .Z(n9575) );
  NAND2HSV0 U11789 ( .A1(\pe19/aot [8]), .A2(\pe19/bq[3] ), .ZN(n9573) );
  NAND2HSV0 U11790 ( .A1(\pe19/aot [6]), .A2(\pe19/bq[5] ), .ZN(n9572) );
  XOR2HSV0 U11791 ( .A1(n9573), .A2(n9572), .Z(n9574) );
  XOR2HSV0 U11792 ( .A1(n9575), .A2(n9574), .Z(n9576) );
  XOR3HSV2 U11793 ( .A1(n9578), .A2(n9577), .A3(n9576), .Z(n9580) );
  NAND2HSV0 U11794 ( .A1(\pe19/ti_7[1] ), .A2(\pe19/got [4]), .ZN(n9579) );
  XNOR2HSV4 U11795 ( .A1(n9580), .A2(n9579), .ZN(n9583) );
  NAND2HSV0 U11796 ( .A1(n9581), .A2(\pe19/got [5]), .ZN(n9582) );
  XNOR2HSV4 U11797 ( .A1(n9583), .A2(n9582), .ZN(n9587) );
  CLKNHSV0 U11798 ( .I(\pe19/got [6]), .ZN(n13336) );
  AOI21HSV0 U11799 ( .A1(n10468), .A2(n10357), .B(n13336), .ZN(n9589) );
  CLKNHSV0 U11800 ( .I(n10468), .ZN(n9586) );
  NAND2HSV0 U11801 ( .A1(n9586), .A2(\pe19/got [6]), .ZN(n9588) );
  CLKNAND2HSV2 U11802 ( .A1(\pe11/aot [7]), .A2(\pe11/bq[8] ), .ZN(n9590) );
  NAND2HSV4 U11803 ( .A1(n9590), .A2(\pe11/phq [2]), .ZN(n9593) );
  INHSV3 U11804 ( .I(\pe11/phq [2]), .ZN(n9591) );
  NAND3HSV4 U11805 ( .A1(n9591), .A2(\pe11/aot [7]), .A3(\pe11/bq[8] ), .ZN(
        n9592) );
  CLKNAND2HSV3 U11806 ( .A1(n9593), .A2(n9592), .ZN(n9595) );
  NAND2HSV1 U11807 ( .A1(\pe11/aot [8]), .A2(\pe11/bq[7] ), .ZN(n9594) );
  XNOR2HSV4 U11808 ( .A1(n9595), .A2(n9594), .ZN(n9599) );
  NAND2HSV2 U11809 ( .A1(\pe11/got [7]), .A2(\pe11/ti_1 ), .ZN(n9597) );
  CLKNAND2HSV2 U11810 ( .A1(\pe11/ctrq ), .A2(\pe11/pvq [2]), .ZN(n9596) );
  XOR2HSV2 U11811 ( .A1(n9597), .A2(n9596), .Z(n9598) );
  XNOR2HSV4 U11812 ( .A1(n9599), .A2(n9598), .ZN(n9605) );
  INHSV2 U11813 ( .I(\pe11/got [8]), .ZN(n11896) );
  NOR2HSV2 U11814 ( .A1(n11896), .A2(n9609), .ZN(n11942) );
  NAND2HSV4 U11815 ( .A1(\pe11/got [8]), .A2(\pe11/ti_1 ), .ZN(n9601) );
  CLKNAND2HSV2 U11816 ( .A1(\pe11/bq[8] ), .A2(\pe11/aot [8]), .ZN(n9600) );
  AND2HSV4 U11817 ( .A1(\pe11/pvq [1]), .A2(\pe11/phq [1]), .Z(n9603) );
  AOI21HSV2 U11818 ( .A1(\pe11/ctrq ), .A2(\pe11/pvq [1]), .B(\pe11/phq [1]), 
        .ZN(n9602) );
  CLKAND2HSV2 U11819 ( .A1(ctro11), .A2(\pe11/ti_7t [2]), .Z(n9604) );
  AOI31HSV2 U11820 ( .A1(n9605), .A2(n11942), .A3(n15260), .B(n9604), .ZN(
        n9608) );
  AOI21HSV2 U11821 ( .A1(n15260), .A2(\pe11/got [8]), .B(n15090), .ZN(n9606)
         );
  INHSV2 U11822 ( .I(n9605), .ZN(n13856) );
  CLKNAND2HSV2 U11823 ( .A1(n9606), .A2(n13856), .ZN(n9607) );
  INHSV2 U11824 ( .I(ctro11), .ZN(n10807) );
  INHSV2 U11825 ( .I(n11914), .ZN(n11916) );
  NAND2HSV2 U11826 ( .A1(n11916), .A2(n9609), .ZN(n11732) );
  CLKNAND2HSV1 U11827 ( .A1(n11732), .A2(\pe11/got [7]), .ZN(n9610) );
  XNOR2HSV4 U11828 ( .A1(n9612), .A2(n9611), .ZN(n10528) );
  NOR2HSV4 U11829 ( .A1(n10528), .A2(n9613), .ZN(n9635) );
  INHSV2 U11830 ( .I(n9613), .ZN(n9659) );
  CLKNAND2HSV1 U11831 ( .A1(n9659), .A2(n10535), .ZN(n9636) );
  NAND2HSV2 U11832 ( .A1(\pe4/aot [6]), .A2(\pe4/bq[8] ), .ZN(n9615) );
  XNOR2HSV4 U11833 ( .A1(n9615), .A2(n9614), .ZN(n9623) );
  CLKNHSV2 U11834 ( .I(n9616), .ZN(n9618) );
  CLKNHSV2 U11835 ( .I(\pe4/phq [3]), .ZN(n9617) );
  CLKNAND2HSV2 U11836 ( .A1(n9618), .A2(n9617), .ZN(n9621) );
  NAND2HSV2 U11837 ( .A1(n9619), .A2(\pe4/phq [3]), .ZN(n9620) );
  XNOR2HSV4 U11838 ( .A1(n9623), .A2(n9622), .ZN(n9627) );
  CLKNAND2HSV1 U11839 ( .A1(\pe4/pvq [3]), .A2(\pe4/ctrq ), .ZN(n9625) );
  NAND2HSV0 U11840 ( .A1(\pe4/aot [7]), .A2(\pe4/bq[7] ), .ZN(n9624) );
  XNOR2HSV4 U11841 ( .A1(n9627), .A2(n9626), .ZN(n9642) );
  XNOR2HSV4 U11842 ( .A1(n9643), .A2(n9642), .ZN(n9628) );
  XNOR2HSV4 U11843 ( .A1(n9628), .A2(n14733), .ZN(n9631) );
  NAND2HSV2 U11844 ( .A1(n9644), .A2(\pe4/got [8]), .ZN(n9630) );
  AOI21HSV4 U11845 ( .A1(n9631), .A2(n10510), .B(n9630), .ZN(n9638) );
  CLKNAND2HSV2 U11846 ( .A1(n13822), .A2(\pe4/pvq [4]), .ZN(n9632) );
  NAND2HSV0 U11847 ( .A1(\pe4/got [5]), .A2(\pe4/ti_1 ), .ZN(n9634) );
  NAND2HSV0 U11848 ( .A1(\pe4/aot [7]), .A2(\pe4/bq[6] ), .ZN(n9633) );
  CLKAND2HSV1 U11849 ( .A1(n9636), .A2(\pe4/got [6]), .Z(n9637) );
  INHSV3 U11850 ( .I(n9639), .ZN(n9640) );
  INHSV2 U11851 ( .I(n9714), .ZN(n9712) );
  NAND2HSV2 U11852 ( .A1(n9680), .A2(\pe4/ti_7t [4]), .ZN(n9674) );
  CLKNAND2HSV2 U11853 ( .A1(n14733), .A2(\pe4/got [8]), .ZN(n9679) );
  XNOR2HSV4 U11854 ( .A1(n9643), .A2(n9642), .ZN(n9678) );
  XNOR2HSV4 U11855 ( .A1(n9679), .A2(n9678), .ZN(n15283) );
  INHSV2 U11856 ( .I(n9644), .ZN(n9684) );
  INHSV2 U11857 ( .I(\pe4/got [7]), .ZN(n9673) );
  NOR2HSV2 U11858 ( .A1(n9684), .A2(n9673), .ZN(n9645) );
  OAI21HSV4 U11859 ( .A1(n15283), .A2(n12597), .B(n9645), .ZN(n9667) );
  CLKNHSV0 U11860 ( .I(\pe4/ti_1 ), .ZN(n13813) );
  NOR2HSV2 U11861 ( .A1(n10536), .A2(n13813), .ZN(n9647) );
  CLKBUFHSV2 U11862 ( .I(\pe4/aot [7]), .Z(n12636) );
  NAND2HSV0 U11863 ( .A1(n12636), .A2(\pe4/bq[5] ), .ZN(n9646) );
  XOR2HSV0 U11864 ( .A1(n9647), .A2(n9646), .Z(n9650) );
  NAND2HSV2 U11865 ( .A1(\pe4/pvq [5]), .A2(n10562), .ZN(n9648) );
  XOR2HSV0 U11866 ( .A1(n9648), .A2(\pe4/phq [5]), .Z(n9649) );
  CLKXOR2HSV4 U11867 ( .A1(n9650), .A2(n9649), .Z(n9658) );
  NAND2HSV0 U11868 ( .A1(\pe4/aot [6]), .A2(\pe4/bq[6] ), .ZN(n9652) );
  INHSV4 U11869 ( .I(n14842), .ZN(n14843) );
  NAND2HSV0 U11870 ( .A1(n14843), .A2(\pe4/bq[4] ), .ZN(n9651) );
  XOR2HSV0 U11871 ( .A1(n9652), .A2(n9651), .Z(n9656) );
  NAND2HSV0 U11872 ( .A1(\pe4/aot [5]), .A2(\pe4/bq[7] ), .ZN(n9654) );
  INHSV4 U11873 ( .I(n14875), .ZN(n13823) );
  CLKNAND2HSV1 U11874 ( .A1(n13823), .A2(\pe4/aot [4]), .ZN(n9653) );
  XOR2HSV0 U11875 ( .A1(n9654), .A2(n9653), .Z(n9655) );
  XOR2HSV0 U11876 ( .A1(n9656), .A2(n9655), .Z(n9657) );
  XNOR2HSV4 U11877 ( .A1(n9658), .A2(n9657), .ZN(n9662) );
  NAND2HSV2 U11878 ( .A1(n9712), .A2(n10528), .ZN(n9660) );
  NAND2HSV4 U11879 ( .A1(n9660), .A2(n9659), .ZN(\pe4/ti_7[1] ) );
  CLKNAND2HSV1 U11880 ( .A1(\pe4/ti_7[1] ), .A2(\pe4/got [5]), .ZN(n9661) );
  CLKXOR2HSV4 U11881 ( .A1(n9662), .A2(n9661), .Z(n9665) );
  NAND2HSV0 U11882 ( .A1(n14733), .A2(\pe4/got [6]), .ZN(n9663) );
  INHSV2 U11883 ( .I(n9663), .ZN(n9664) );
  XNOR2HSV4 U11884 ( .A1(n9665), .A2(n9664), .ZN(n9666) );
  CLKNHSV0 U11885 ( .I(n14933), .ZN(n9668) );
  CLKNHSV2 U11886 ( .I(n10583), .ZN(n9669) );
  NAND2HSV2 U11887 ( .A1(n9668), .A2(n9669), .ZN(n9671) );
  NAND2HSV2 U11888 ( .A1(n9669), .A2(n15083), .ZN(n9670) );
  CLKNHSV1 U11889 ( .I(n9674), .ZN(n9676) );
  AOI21HSV2 U11890 ( .A1(n9674), .A2(n14861), .B(n9673), .ZN(n9675) );
  NOR2HSV0 U11891 ( .A1(n9679), .A2(n14861), .ZN(n9677) );
  NAND2HSV2 U11892 ( .A1(n9677), .A2(n9678), .ZN(n9703) );
  INHSV2 U11893 ( .I(n9678), .ZN(n9683) );
  CLKNHSV0 U11894 ( .I(n9679), .ZN(n9681) );
  NOR2HSV1 U11895 ( .A1(n9681), .A2(n9680), .ZN(n9682) );
  NAND2HSV2 U11896 ( .A1(n9683), .A2(n9682), .ZN(n9704) );
  INHSV2 U11897 ( .I(\pe4/got [6]), .ZN(n12596) );
  NOR2HSV1 U11898 ( .A1(n9684), .A2(n12596), .ZN(n9705) );
  CLKNAND2HSV1 U11899 ( .A1(n14843), .A2(\pe4/bq[3] ), .ZN(n9686) );
  BUFHSV4 U11900 ( .I(\pe4/bq[6] ), .Z(n12581) );
  NAND2HSV2 U11901 ( .A1(\pe4/aot [5]), .A2(n12581), .ZN(n9685) );
  XOR2HSV0 U11902 ( .A1(n9686), .A2(n9685), .Z(n9698) );
  CLKNAND2HSV1 U11903 ( .A1(\pe4/ctrq ), .A2(\pe4/pvq [6]), .ZN(n9687) );
  XNOR2HSV1 U11904 ( .A1(n9687), .A2(\pe4/phq [6]), .ZN(n9689) );
  NAND2HSV0 U11905 ( .A1(\pe4/aot [4]), .A2(\pe4/bq[7] ), .ZN(n9688) );
  XNOR2HSV1 U11906 ( .A1(n9689), .A2(n9688), .ZN(n9697) );
  NAND2HSV2 U11907 ( .A1(\pe4/got [3]), .A2(n8927), .ZN(n9691) );
  NAND2HSV0 U11908 ( .A1(\pe4/bq[4] ), .A2(\pe4/aot [7]), .ZN(n9690) );
  XOR2HSV0 U11909 ( .A1(n9693), .A2(n9692), .Z(n9694) );
  XOR2HSV0 U11910 ( .A1(n9695), .A2(n9694), .Z(n9696) );
  XOR3HSV2 U11911 ( .A1(n9698), .A2(n9697), .A3(n9696), .Z(n9700) );
  NAND2HSV0 U11912 ( .A1(\pe4/ti_7[1] ), .A2(\pe4/got [4]), .ZN(n9699) );
  XNOR2HSV1 U11913 ( .A1(n9700), .A2(n9699), .ZN(n9702) );
  CLKBUFHSV2 U11914 ( .I(n14733), .Z(n10537) );
  NAND2HSV2 U11915 ( .A1(n10537), .A2(\pe4/got [5]), .ZN(n9701) );
  XNOR2HSV4 U11916 ( .A1(n9702), .A2(n9701), .ZN(n9709) );
  INHSV2 U11917 ( .I(n9703), .ZN(n9708) );
  INHSV2 U11918 ( .I(n9704), .ZN(n9707) );
  INHSV1 U11919 ( .I(n9705), .ZN(n9706) );
  CLKNHSV0 U11920 ( .I(\pe4/ti_7t [5]), .ZN(n9710) );
  AO21HSV1 U11921 ( .A1(n9710), .A2(n12597), .B(n15083), .Z(n9711) );
  CLKNHSV2 U11922 ( .I(n13879), .ZN(n9716) );
  CLKNAND2HSV3 U11923 ( .A1(n9716), .A2(n6722), .ZN(n9717) );
  NAND2HSV2 U11924 ( .A1(n10535), .A2(\pe4/ti_7t [6]), .ZN(n9719) );
  OR2HSV1 U11925 ( .A1(n9722), .A2(n9721), .Z(n9724) );
  INHSV2 U11926 ( .I(n9726), .ZN(n9732) );
  INHSV2 U11927 ( .I(n9727), .ZN(n9729) );
  NAND3HSV4 U11928 ( .A1(n9732), .A2(n9731), .A3(n9730), .ZN(n9733) );
  CLKNHSV2 U11929 ( .I(n7881), .ZN(n9740) );
  CLKNHSV0 U11930 ( .I(n9735), .ZN(n9737) );
  OR2HSV1 U11931 ( .A1(n9737), .A2(n9736), .Z(n9738) );
  AOI21HSV4 U11932 ( .A1(n9740), .A2(n9739), .B(n9738), .ZN(n9742) );
  NOR2HSV1 U11933 ( .A1(n9420), .A2(ctro9), .ZN(n9793) );
  CLKNHSV2 U11934 ( .I(n9793), .ZN(n9743) );
  INHSV2 U11935 ( .I(n9746), .ZN(n9747) );
  NAND2HSV0 U11936 ( .A1(\pe9/aot [4]), .A2(\pe9/bq[1] ), .ZN(n13918) );
  NAND2HSV0 U11937 ( .A1(\pe9/aot [2]), .A2(\pe9/bq[3] ), .ZN(n9749) );
  XNOR2HSV1 U11938 ( .A1(n13918), .A2(n9749), .ZN(n9751) );
  CLKNHSV0 U11939 ( .I(\pe9/got [2]), .ZN(n9750) );
  NOR2HSV2 U11940 ( .A1(n9751), .A2(n9750), .ZN(n9753) );
  CLKNAND2HSV2 U11941 ( .A1(n9754), .A2(\pe9/got [2]), .ZN(n9752) );
  CLKNAND2HSV0 U11942 ( .A1(\pe9/aot [3]), .A2(\pe9/bq[2] ), .ZN(n9756) );
  NAND2HSV0 U11943 ( .A1(\pe9/bq[4] ), .A2(\pe9/aot [1]), .ZN(n9755) );
  XOR2HSV0 U11944 ( .A1(n9756), .A2(n9755), .Z(n9757) );
  XNOR2HSV1 U11945 ( .A1(n9758), .A2(n9757), .ZN(n9759) );
  CLKNAND2HSV0 U11946 ( .A1(\pe9/ti_7[1] ), .A2(\pe9/got [3]), .ZN(n9786) );
  NAND2HSV0 U11947 ( .A1(n14942), .A2(\pe9/bq[2] ), .ZN(n9765) );
  NAND2HSV0 U11948 ( .A1(n5976), .A2(\pe9/aot [3]), .ZN(n9764) );
  XOR2HSV0 U11949 ( .A1(n9765), .A2(n9764), .Z(n9782) );
  NAND2HSV2 U11950 ( .A1(n13826), .A2(\pe9/pvq [7]), .ZN(n9766) );
  XNOR2HSV1 U11951 ( .A1(n9766), .A2(\pe9/phq [7]), .ZN(n9771) );
  NAND2HSV0 U11952 ( .A1(\pe9/aot [2]), .A2(\pe9/bq[6] ), .ZN(n13922) );
  NOR2HSV2 U11953 ( .A1(n9767), .A2(n13922), .ZN(n9769) );
  AOI22HSV0 U11954 ( .A1(\pe9/aot [4]), .A2(n11647), .B1(\pe9/bq[8] ), .B2(
        \pe9/aot [2]), .ZN(n9768) );
  NOR2HSV1 U11955 ( .A1(n9769), .A2(n9768), .ZN(n9770) );
  NOR2HSV1 U11956 ( .A1(n9773), .A2(n9772), .ZN(n9775) );
  NAND2HSV2 U11957 ( .A1(\pe9/got [2]), .A2(n8944), .ZN(n9774) );
  XOR2HSV0 U11958 ( .A1(n9775), .A2(n9774), .Z(n9779) );
  NAND2HSV2 U11959 ( .A1(\pe9/bq[5] ), .A2(\pe9/aot [5]), .ZN(n9777) );
  NAND2HSV0 U11960 ( .A1(\pe9/bq[3] ), .A2(\pe9/aot [7]), .ZN(n9776) );
  XOR2HSV0 U11961 ( .A1(n9777), .A2(n9776), .Z(n9778) );
  XOR2HSV0 U11962 ( .A1(n9779), .A2(n9778), .Z(n9780) );
  XOR3HSV2 U11963 ( .A1(n9782), .A2(n9781), .A3(n9780), .Z(n9785) );
  NAND2HSV0 U11964 ( .A1(n14896), .A2(\pe9/got [4]), .ZN(n9784) );
  XNOR3HSV2 U11965 ( .A1(n9786), .A2(n9785), .A3(n9784), .ZN(n9787) );
  INOR2HSV0 U11966 ( .A1(n15074), .B1(n9791), .ZN(n9792) );
  INHSV1 U11967 ( .I(n9799), .ZN(n9801) );
  AOI21HSV2 U11968 ( .A1(n9799), .A2(n9798), .B(n9797), .ZN(n9800) );
  NAND2HSV2 U11969 ( .A1(n9802), .A2(\pe6/ti_7t [2]), .ZN(n10801) );
  CLKNHSV0 U11970 ( .I(n10801), .ZN(n9805) );
  CLKNHSV0 U11971 ( .I(\pe6/got [4]), .ZN(n9803) );
  AOI21HSV1 U11972 ( .A1(n10801), .A2(n9842), .B(n9803), .ZN(n9804) );
  OA21HSV4 U11973 ( .A1(n10800), .A2(n9805), .B(n9804), .Z(n9827) );
  NAND2HSV0 U11974 ( .A1(\pe6/aot [5]), .A2(\pe6/bq[5] ), .ZN(n9807) );
  NAND2HSV0 U11975 ( .A1(\pe6/aot [4]), .A2(\pe6/bq[6] ), .ZN(n9806) );
  XOR2HSV0 U11976 ( .A1(n9807), .A2(n9806), .Z(n9811) );
  NAND2HSV0 U11977 ( .A1(\pe6/aot [3]), .A2(\pe6/bq[7] ), .ZN(n9809) );
  NAND2HSV0 U11978 ( .A1(\pe6/aot [6]), .A2(\pe6/bq[4] ), .ZN(n9808) );
  XOR2HSV0 U11979 ( .A1(n9809), .A2(n9808), .Z(n9810) );
  XOR2HSV0 U11980 ( .A1(n9811), .A2(n9810), .Z(n9815) );
  CLKNAND2HSV0 U11981 ( .A1(n13829), .A2(\pe6/aot [2]), .ZN(n9813) );
  NAND2HSV0 U11982 ( .A1(\pe6/bq[2] ), .A2(\pe6/aot [8]), .ZN(n9812) );
  XOR2HSV0 U11983 ( .A1(n9813), .A2(n9812), .Z(n9814) );
  XNOR2HSV4 U11984 ( .A1(n9815), .A2(n9814), .ZN(n9822) );
  NAND2HSV0 U11985 ( .A1(\pe6/aot [7]), .A2(\pe6/bq[3] ), .ZN(n9817) );
  NAND2HSV0 U11986 ( .A1(\pe6/got [2]), .A2(n13824), .ZN(n9816) );
  XOR2HSV0 U11987 ( .A1(n9817), .A2(n9816), .Z(n9820) );
  CLKNAND2HSV1 U11988 ( .A1(n13041), .A2(\pe6/pvq [7]), .ZN(n9818) );
  XOR2HSV0 U11989 ( .A1(n9818), .A2(\pe6/phq [7]), .Z(n9819) );
  XNOR2HSV1 U11990 ( .A1(n9820), .A2(n9819), .ZN(n9821) );
  XNOR2HSV4 U11991 ( .A1(n9822), .A2(n9821), .ZN(n9825) );
  BUFHSV4 U11992 ( .I(n6445), .Z(n14895) );
  NAND2HSV2 U11993 ( .A1(n14895), .A2(\pe6/got [3]), .ZN(n9824) );
  XNOR2HSV4 U11994 ( .A1(n9825), .A2(n9824), .ZN(n9826) );
  XNOR2HSV4 U11995 ( .A1(n9827), .A2(n9826), .ZN(n9831) );
  NAND2HSV2 U11996 ( .A1(n9829), .A2(\pe6/got [5]), .ZN(n9830) );
  XNOR2HSV4 U11997 ( .A1(n9831), .A2(n9830), .ZN(n9837) );
  NOR2HSV2 U11998 ( .A1(n7813), .A2(n15095), .ZN(n13103) );
  NAND2HSV2 U11999 ( .A1(n9834), .A2(n9832), .ZN(n9833) );
  XNOR2HSV4 U12000 ( .A1(n9837), .A2(n9836), .ZN(n9838) );
  INHSV2 U12001 ( .I(n9840), .ZN(n9841) );
  INHSV1 U12002 ( .I(n9843), .ZN(n9845) );
  CLKNAND2HSV1 U12003 ( .A1(n15088), .A2(\pe6/ti_7t [7]), .ZN(n9844) );
  NAND2HSV0 U12004 ( .A1(n13057), .A2(\pe6/got [1]), .ZN(n9857) );
  NAND2HSV0 U12005 ( .A1(\pe6/aot [4]), .A2(\pe6/bq[2] ), .ZN(n9855) );
  NAND2HSV2 U12006 ( .A1(\pe6/aot [2]), .A2(\pe6/bq[5] ), .ZN(n12936) );
  INHSV2 U12007 ( .I(n12936), .ZN(n9850) );
  CLKNHSV0 U12008 ( .I(n13000), .ZN(n9849) );
  AOI22HSV0 U12009 ( .A1(\pe6/aot [2]), .A2(\pe6/bq[4] ), .B1(\pe6/bq[5] ), 
        .B2(\pe6/aot [1]), .ZN(n9848) );
  AOI21HSV2 U12010 ( .A1(n9850), .A2(n9849), .B(n9848), .ZN(n9854) );
  NAND2HSV2 U12011 ( .A1(\pe6/aot [5]), .A2(\pe6/bq[3] ), .ZN(n12418) );
  CLKNAND2HSV1 U12012 ( .A1(\pe6/aot [3]), .A2(\pe6/bq[1] ), .ZN(n12984) );
  NOR2HSV0 U12013 ( .A1(n12418), .A2(n12984), .ZN(n9852) );
  AOI22HSV0 U12014 ( .A1(\pe6/aot [5]), .A2(\pe6/bq[1] ), .B1(\pe6/aot [3]), 
        .B2(\pe6/bq[3] ), .ZN(n9851) );
  NOR2HSV2 U12015 ( .A1(n9852), .A2(n9851), .ZN(n9853) );
  XOR3HSV2 U12016 ( .A1(n9855), .A2(n9854), .A3(n9853), .Z(n9856) );
  XNOR2HSV1 U12017 ( .A1(n9857), .A2(n9856), .ZN(n9860) );
  BUFHSV6 U12018 ( .I(n9858), .Z(n15077) );
  NAND2HSV0 U12019 ( .A1(n15077), .A2(\pe6/got [2]), .ZN(n9859) );
  CLKNHSV2 U12020 ( .I(n9859), .ZN(n9861) );
  INHSV1 U12021 ( .I(\pe6/got [2]), .ZN(n12998) );
  CLKNAND2HSV0 U12022 ( .A1(\pe13/pvq [3]), .A2(\pe13/ctrq ), .ZN(n9862) );
  CLKBUFHSV4 U12023 ( .I(\pe13/bq[7] ), .Z(n13591) );
  NAND2HSV2 U12024 ( .A1(n13591), .A2(\pe13/aot [7]), .ZN(n13590) );
  NAND2HSV0 U12025 ( .A1(\pe13/ti_1 ), .A2(\pe13/got [6]), .ZN(n9863) );
  XOR2HSV0 U12026 ( .A1(n13590), .A2(n9863), .Z(n9864) );
  XNOR2HSV4 U12027 ( .A1(n9865), .A2(n9864), .ZN(n9905) );
  INHSV2 U12028 ( .I(\pe13/ti_7t [1]), .ZN(n9866) );
  NOR2HSV2 U12029 ( .A1(n9977), .A2(n9866), .ZN(n9867) );
  NOR2HSV4 U12030 ( .A1(n15246), .A2(n9867), .ZN(n9900) );
  INHSV2 U12031 ( .I(n9867), .ZN(n9916) );
  CLKNAND2HSV1 U12032 ( .A1(n9916), .A2(n9988), .ZN(n9898) );
  XNOR2HSV4 U12033 ( .A1(n9905), .A2(n9904), .ZN(n9885) );
  INHSV2 U12034 ( .I(\pe13/got [8]), .ZN(n9956) );
  NOR2HSV2 U12035 ( .A1(n9956), .A2(n9921), .ZN(n9978) );
  INHSV2 U12036 ( .I(\pe13/aot [7]), .ZN(n9869) );
  INHSV2 U12037 ( .I(\pe13/bq[8] ), .ZN(n9868) );
  NOR2HSV2 U12038 ( .A1(n9869), .A2(n9868), .ZN(n9870) );
  XNOR2HSV4 U12039 ( .A1(n9871), .A2(n9870), .ZN(n9875) );
  CLKNAND2HSV1 U12040 ( .A1(\pe13/got [7]), .A2(\pe13/ti_1 ), .ZN(n9873) );
  NAND2HSV0 U12041 ( .A1(\pe13/ctrq ), .A2(\pe13/pvq [2]), .ZN(n9872) );
  XOR2HSV0 U12042 ( .A1(n9873), .A2(n9872), .Z(n9874) );
  XNOR2HSV4 U12043 ( .A1(n9875), .A2(n9874), .ZN(n9877) );
  CLKAND2HSV2 U12044 ( .A1(n9921), .A2(\pe13/ti_7t [2]), .Z(n9876) );
  AOI21HSV4 U12045 ( .A1(n8907), .A2(n9877), .B(n9876), .ZN(n9880) );
  AOI21HSV2 U12046 ( .A1(n15246), .A2(\pe13/got [8]), .B(n15087), .ZN(n9878)
         );
  INHSV4 U12047 ( .I(n9877), .ZN(n13847) );
  CLKNAND2HSV3 U12048 ( .A1(n13847), .A2(n9878), .ZN(n9879) );
  INHSV3 U12049 ( .I(n9920), .ZN(n9884) );
  NOR2HSV2 U12050 ( .A1(n9977), .A2(\pe13/ti_7t [3]), .ZN(n9908) );
  NOR2HSV2 U12051 ( .A1(n9908), .A2(n9956), .ZN(n9883) );
  CLKNAND2HSV0 U12052 ( .A1(n9884), .A2(n9977), .ZN(n9887) );
  INHSV2 U12053 ( .I(n9885), .ZN(n9886) );
  NAND2HSV2 U12054 ( .A1(\pe13/aot [7]), .A2(\pe13/bq[6] ), .ZN(n9889) );
  NAND2HSV0 U12055 ( .A1(\pe13/got [5]), .A2(\pe13/ti_1 ), .ZN(n9888) );
  XOR2HSV2 U12056 ( .A1(n9889), .A2(n9888), .Z(n9892) );
  NAND2HSV2 U12057 ( .A1(\pe13/ctrq ), .A2(\pe13/pvq [4]), .ZN(n9893) );
  XNOR2HSV4 U12058 ( .A1(n9893), .A2(\pe13/phq [4]), .ZN(n9895) );
  XNOR2HSV1 U12059 ( .A1(n9895), .A2(n9894), .ZN(n9896) );
  XNOR2HSV4 U12060 ( .A1(n9897), .A2(n9896), .ZN(n9902) );
  CLKNAND2HSV0 U12061 ( .A1(n9898), .A2(\pe13/got [6]), .ZN(n9899) );
  NOR2HSV4 U12062 ( .A1(n9900), .A2(n9899), .ZN(n9901) );
  NAND2HSV2 U12063 ( .A1(n9988), .A2(\pe13/ti_7t [4]), .ZN(n9949) );
  INHSV2 U12064 ( .I(n9949), .ZN(n9951) );
  INHSV3 U12065 ( .I(n9956), .ZN(n14750) );
  XNOR2HSV4 U12066 ( .A1(n9905), .A2(n9904), .ZN(n9907) );
  INHSV2 U12067 ( .I(\pe13/got [7]), .ZN(n9948) );
  NOR2HSV2 U12068 ( .A1(n9908), .A2(n9948), .ZN(n9909) );
  NAND2HSV0 U12069 ( .A1(\pe13/ti_1 ), .A2(\pe13/got [4]), .ZN(n9911) );
  NAND2HSV0 U12070 ( .A1(\pe13/aot [7]), .A2(\pe13/bq[5] ), .ZN(n9910) );
  XOR2HSV0 U12071 ( .A1(n9911), .A2(n9910), .Z(n9914) );
  NAND2HSV0 U12072 ( .A1(\pe13/bq[6] ), .A2(\pe13/aot [6]), .ZN(n10009) );
  NAND2HSV0 U12073 ( .A1(\pe13/bq[7] ), .A2(\pe13/aot [5]), .ZN(n9912) );
  XOR2HSV0 U12074 ( .A1(n10009), .A2(n9912), .Z(n9913) );
  XOR2HSV0 U12075 ( .A1(n9914), .A2(n9913), .Z(n9915) );
  INHSV3 U12076 ( .I(\pe13/ctrq ), .ZN(n11834) );
  CLKNAND2HSV0 U12077 ( .A1(n9977), .A2(n15246), .ZN(n9917) );
  NAND2HSV2 U12078 ( .A1(n9917), .A2(n9916), .ZN(\pe13/ti_7[1] ) );
  XNOR2HSV4 U12079 ( .A1(n9999), .A2(n9979), .ZN(n15242) );
  CLKNAND2HSV1 U12080 ( .A1(n9921), .A2(\pe13/ti_7t [5]), .ZN(n9922) );
  NAND2HSV2 U12081 ( .A1(n15244), .A2(n9881), .ZN(n9925) );
  NAND2HSV0 U12082 ( .A1(n15087), .A2(\pe13/ti_7t [3]), .ZN(n9924) );
  BUFHSV2 U12083 ( .I(n9957), .Z(n15065) );
  CLKNAND2HSV0 U12084 ( .A1(n15065), .A2(\pe13/got [2]), .ZN(n9930) );
  CLKNAND2HSV0 U12085 ( .A1(n9882), .A2(\pe13/got [1]), .ZN(n9929) );
  CLKNHSV0 U12086 ( .I(\pe13/aot [2]), .ZN(n9926) );
  NOR2HSV2 U12087 ( .A1(n9926), .A2(n9960), .ZN(n13592) );
  CLKNHSV0 U12088 ( .I(\pe13/aot [5]), .ZN(n9927) );
  INHSV2 U12089 ( .I(\pe13/bq[5] ), .ZN(n11832) );
  NOR2HSV2 U12090 ( .A1(n9927), .A2(n11832), .ZN(n12922) );
  NAND2HSV0 U12091 ( .A1(\pe13/ti_7[1] ), .A2(\pe13/got [4]), .ZN(n9945) );
  BUFHSV2 U12092 ( .I(\pe13/ti_1 ), .Z(n13819) );
  NAND2HSV0 U12093 ( .A1(n13819), .A2(\pe13/got [3]), .ZN(n9934) );
  NAND2HSV0 U12094 ( .A1(\pe13/bq[5] ), .A2(\pe13/aot [6]), .ZN(n9933) );
  XOR2HSV0 U12095 ( .A1(n9934), .A2(n9933), .Z(n9943) );
  CLKNAND2HSV0 U12096 ( .A1(n13591), .A2(\pe13/aot [4]), .ZN(n9935) );
  CLKNAND2HSV0 U12097 ( .A1(\pe13/aot [7]), .A2(\pe13/bq[4] ), .ZN(n9937) );
  NAND2HSV0 U12098 ( .A1(n14939), .A2(\pe13/bq[3] ), .ZN(n9936) );
  XOR2HSV0 U12099 ( .A1(n9937), .A2(n9936), .Z(n9941) );
  NAND2HSV0 U12100 ( .A1(\pe13/aot [5]), .A2(\pe13/bq[6] ), .ZN(n9939) );
  NAND2HSV0 U12101 ( .A1(\pe13/aot [3]), .A2(\pe13/bq[8] ), .ZN(n9938) );
  XOR2HSV0 U12102 ( .A1(n9939), .A2(n9938), .Z(n9940) );
  XOR2HSV0 U12103 ( .A1(n9941), .A2(n9940), .Z(n9942) );
  CLKNAND2HSV1 U12104 ( .A1(n9920), .A2(\pe13/got [5]), .ZN(n9944) );
  AOI21HSV1 U12105 ( .A1(n9949), .A2(n9921), .B(n9948), .ZN(n9950) );
  NOR2HSV1 U12106 ( .A1(n15243), .A2(n15087), .ZN(n9955) );
  NOR2HSV1 U12107 ( .A1(n9977), .A2(\pe13/ti_7t [5]), .ZN(n9996) );
  NAND2HSV2 U12108 ( .A1(n15087), .A2(\pe13/ti_7t [6]), .ZN(n9990) );
  CLKNAND2HSV1 U12109 ( .A1(n9957), .A2(\pe13/got [5]), .ZN(n9976) );
  CLKNAND2HSV1 U12110 ( .A1(n9882), .A2(\pe13/got [4]), .ZN(n9959) );
  NAND2HSV0 U12111 ( .A1(\pe13/ti_7[1] ), .A2(\pe13/got [3]), .ZN(n9958) );
  CLKNAND2HSV1 U12112 ( .A1(n13591), .A2(\pe13/aot [3]), .ZN(n10016) );
  XOR2HSV0 U12113 ( .A1(n12922), .A2(n10016), .Z(n9974) );
  CLKNAND2HSV0 U12114 ( .A1(n14939), .A2(\pe13/bq[2] ), .ZN(n9962) );
  NAND2HSV0 U12115 ( .A1(\pe13/got [2]), .A2(n13819), .ZN(n9961) );
  XOR2HSV0 U12116 ( .A1(n9962), .A2(n9961), .Z(n9965) );
  CLKNAND2HSV1 U12117 ( .A1(n14552), .A2(\pe13/pvq [7]), .ZN(n9963) );
  XNOR2HSV1 U12118 ( .A1(n9963), .A2(\pe13/phq [7]), .ZN(n9964) );
  XNOR2HSV1 U12119 ( .A1(n9965), .A2(n9964), .ZN(n9973) );
  NAND2HSV0 U12120 ( .A1(\pe13/aot [7]), .A2(\pe13/bq[3] ), .ZN(n9967) );
  NAND2HSV0 U12121 ( .A1(\pe13/bq[4] ), .A2(\pe13/aot [6]), .ZN(n9966) );
  XOR2HSV0 U12122 ( .A1(n9967), .A2(n9966), .Z(n9971) );
  NAND2HSV0 U12123 ( .A1(\pe13/aot [4]), .A2(\pe13/bq[6] ), .ZN(n9969) );
  XOR2HSV0 U12124 ( .A1(n9969), .A2(n9968), .Z(n9970) );
  XOR2HSV0 U12125 ( .A1(n9971), .A2(n9970), .Z(n9972) );
  XOR3HSV2 U12126 ( .A1(n9974), .A2(n9973), .A3(n9972), .Z(n9975) );
  NAND3HSV2 U12127 ( .A1(n9979), .A2(\pe13/ti_7[4] ), .A3(n9978), .ZN(n9984)
         );
  NOR2HSV2 U12128 ( .A1(ctro13), .A2(\pe13/got [8]), .ZN(n9987) );
  CLKNHSV0 U12129 ( .I(n9996), .ZN(n9980) );
  CLKNAND2HSV0 U12130 ( .A1(n9980), .A2(\pe13/got [7]), .ZN(n9981) );
  AOI21HSV2 U12131 ( .A1(n9982), .A2(n9987), .B(n9981), .ZN(n9983) );
  OAI211HSV2 U12132 ( .A1(\pe13/ti_7[4] ), .A2(n10000), .B(n9984), .C(n9983), 
        .ZN(n9985) );
  CLKNHSV0 U12133 ( .I(n9999), .ZN(n9994) );
  NOR2HSV0 U12134 ( .A1(n9992), .A2(n15087), .ZN(n9993) );
  NAND2HSV2 U12135 ( .A1(n9994), .A2(n9993), .ZN(n10003) );
  INHSV2 U12136 ( .I(n10003), .ZN(n9998) );
  CLKNAND2HSV1 U12137 ( .A1(n13587), .A2(\pe13/got [4]), .ZN(n10001) );
  CLKNHSV0 U12138 ( .I(\pe13/got [5]), .ZN(n9995) );
  NOR2HSV0 U12139 ( .A1(n9996), .A2(n9995), .ZN(n10002) );
  CLKNAND2HSV0 U12140 ( .A1(n10001), .A2(n10002), .ZN(n9997) );
  NOR2HSV2 U12141 ( .A1(n9998), .A2(n9997), .ZN(n10006) );
  INAND2HSV2 U12142 ( .A1(n10000), .B1(n9999), .ZN(n10005) );
  AOI31HSV2 U12143 ( .A1(n10003), .A2(n10002), .A3(n10005), .B(n10001), .ZN(
        n10004) );
  NAND2HSV0 U12144 ( .A1(n15065), .A2(\pe13/got [3]), .ZN(n10026) );
  NAND2HSV0 U12145 ( .A1(\pe13/ti_7[1] ), .A2(\pe13/got [1]), .ZN(n10022) );
  NAND2HSV0 U12146 ( .A1(\pe13/aot [4]), .A2(\pe13/bq[4] ), .ZN(n10008) );
  NAND2HSV0 U12147 ( .A1(\pe13/aot [7]), .A2(\pe13/bq[1] ), .ZN(n10007) );
  XOR2HSV0 U12148 ( .A1(n10008), .A2(n10007), .Z(n10013) );
  CLKNHSV0 U12149 ( .I(n10009), .ZN(n10011) );
  AOI22HSV0 U12150 ( .A1(\pe13/aot [6]), .A2(\pe13/bq[2] ), .B1(\pe13/bq[6] ), 
        .B2(\pe13/aot [2]), .ZN(n10010) );
  AOI21HSV0 U12151 ( .A1(n13592), .A2(n10011), .B(n10010), .ZN(n10012) );
  XNOR2HSV1 U12152 ( .A1(n10013), .A2(n10012), .ZN(n10020) );
  CLKNHSV0 U12153 ( .I(\pe13/aot [3]), .ZN(n10014) );
  OAI21HSV0 U12154 ( .A1(n12924), .A2(n10016), .B(n10015), .ZN(n10018) );
  NAND2HSV0 U12155 ( .A1(\pe13/aot [5]), .A2(\pe13/bq[3] ), .ZN(n10017) );
  XNOR2HSV1 U12156 ( .A1(n10018), .A2(n10017), .ZN(n10019) );
  XNOR2HSV1 U12157 ( .A1(n10020), .A2(n10019), .ZN(n10021) );
  XNOR2HSV1 U12158 ( .A1(n10022), .A2(n10021), .ZN(n10024) );
  NAND2HSV0 U12159 ( .A1(n9882), .A2(\pe13/got [2]), .ZN(n10023) );
  XNOR2HSV1 U12160 ( .A1(n10024), .A2(n10023), .ZN(n10025) );
  XOR2HSV0 U12161 ( .A1(n10026), .A2(n10025), .Z(n10027) );
  INHSV2 U12162 ( .I(ctro10), .ZN(n10070) );
  INHSV2 U12163 ( .I(n10070), .ZN(n10058) );
  INHSV2 U12164 ( .I(n10070), .ZN(n10073) );
  INHSV2 U12165 ( .I(n10073), .ZN(n10924) );
  NAND2HSV2 U12166 ( .A1(n10058), .A2(\pe10/ti_7t [1]), .ZN(n10088) );
  BUFHSV8 U12167 ( .I(\pe10/aot [8]), .Z(n14951) );
  NAND2HSV2 U12168 ( .A1(\pe10/bq[6] ), .A2(\pe10/aot [7]), .ZN(n10030) );
  INHSV2 U12169 ( .I(n10030), .ZN(n10051) );
  NAND2HSV2 U12170 ( .A1(\pe10/bq[5] ), .A2(\pe10/aot [7]), .ZN(n10077) );
  NOR2HSV1 U12171 ( .A1(n10077), .A2(n10053), .ZN(n10031) );
  NOR2HSV2 U12172 ( .A1(n10032), .A2(n10031), .ZN(n10034) );
  XNOR2HSV4 U12173 ( .A1(n10034), .A2(n10033), .ZN(n10039) );
  INHSV4 U12174 ( .I(\pe10/ctrq ), .ZN(n10035) );
  XOR3HSV2 U12175 ( .A1(\pe10/phq [4]), .A2(n10037), .A3(n10036), .Z(n10038)
         );
  INHSV2 U12176 ( .I(ctro10), .ZN(n10925) );
  CLKNAND2HSV1 U12177 ( .A1(\pe10/got [7]), .A2(\pe10/ti_1 ), .ZN(n10044) );
  NAND2HSV2 U12178 ( .A1(\pe10/ti_1 ), .A2(\pe10/got [7]), .ZN(n10042) );
  NOR2HSV4 U12179 ( .A1(n10042), .A2(n10041), .ZN(n10043) );
  INHSV2 U12180 ( .I(n10047), .ZN(n10046) );
  INHSV2 U12181 ( .I(n10052), .ZN(n10045) );
  NAND2HSV0 U12182 ( .A1(n10073), .A2(\pe10/ti_7t [2]), .ZN(n10060) );
  INHSV2 U12183 ( .I(n10060), .ZN(n10048) );
  NOR2HSV4 U12184 ( .A1(n10049), .A2(n10048), .ZN(n10050) );
  NOR2HSV2 U12185 ( .A1(n15098), .A2(ctro10), .ZN(n10148) );
  INHSV2 U12186 ( .I(\pe10/aot [7]), .ZN(n10804) );
  OAI21HSV4 U12187 ( .A1(n6312), .A2(n10804), .B(n10053), .ZN(n10054) );
  AOI21HSV1 U12188 ( .A1(n15096), .A2(n10058), .B(n15140), .ZN(n10059) );
  OR2HSV1 U12189 ( .A1(n10060), .A2(n15098), .Z(n10061) );
  NAND2HSV4 U12190 ( .A1(n10062), .A2(n10061), .ZN(n10063) );
  INHSV2 U12191 ( .I(n10925), .ZN(n10119) );
  INHSV2 U12192 ( .I(n10070), .ZN(n14828) );
  NOR2HSV2 U12193 ( .A1(n10599), .A2(\pe10/ti_7t [4]), .ZN(n10125) );
  NOR2HSV2 U12194 ( .A1(n10125), .A2(n15098), .ZN(n10072) );
  INHSV2 U12195 ( .I(n10127), .ZN(n10784) );
  AOI21HSV1 U12196 ( .A1(n10073), .A2(n10127), .B(n15140), .ZN(n10074) );
  CLKNAND2HSV0 U12197 ( .A1(\pe10/aot [6]), .A2(\pe10/bq[6] ), .ZN(n10076) );
  XOR2HSV0 U12198 ( .A1(n10077), .A2(n10076), .Z(n10081) );
  NAND2HSV0 U12199 ( .A1(\pe10/aot [5]), .A2(\pe10/bq[7] ), .ZN(n10078) );
  XOR2HSV0 U12200 ( .A1(n10079), .A2(n10078), .Z(n10080) );
  XNOR2HSV4 U12201 ( .A1(n10085), .A2(n10084), .ZN(n10087) );
  INHSV2 U12202 ( .I(\pe10/ti_7t [5]), .ZN(n10112) );
  INHSV2 U12203 ( .I(n14122), .ZN(n10926) );
  NAND2HSV0 U12204 ( .A1(n10926), .A2(ctro10), .ZN(n14125) );
  BUFHSV2 U12205 ( .I(\pe10/aot [6]), .Z(n14133) );
  CLKNAND2HSV1 U12206 ( .A1(n14133), .A2(\pe10/bq[4] ), .ZN(n10090) );
  NAND2HSV0 U12207 ( .A1(\pe10/aot [2]), .A2(n12272), .ZN(n10089) );
  XOR2HSV0 U12208 ( .A1(n10090), .A2(n10089), .Z(n10104) );
  NAND2HSV0 U12209 ( .A1(\pe10/got [2]), .A2(\pe10/ti_1 ), .ZN(n10091) );
  XOR2HSV0 U12210 ( .A1(n10092), .A2(n10091), .Z(n10095) );
  XNOR2HSV1 U12211 ( .A1(n10093), .A2(\pe10/phq [7]), .ZN(n10094) );
  NAND2HSV0 U12212 ( .A1(\pe10/aot [7]), .A2(\pe10/bq[3] ), .ZN(n10097) );
  NAND2HSV0 U12213 ( .A1(\pe10/aot [5]), .A2(\pe10/bq[5] ), .ZN(n10096) );
  XOR2HSV0 U12214 ( .A1(n10097), .A2(n10096), .Z(n10101) );
  CLKNAND2HSV0 U12215 ( .A1(\pe10/aot [4]), .A2(\pe10/bq[6] ), .ZN(n10099) );
  NAND2HSV0 U12216 ( .A1(\pe10/aot [3]), .A2(\pe10/bq[7] ), .ZN(n10098) );
  XOR2HSV0 U12217 ( .A1(n10099), .A2(n10098), .Z(n10100) );
  XOR2HSV0 U12218 ( .A1(n10101), .A2(n10100), .Z(n10102) );
  CLKBUFHSV4 U12219 ( .I(n10145), .Z(n14940) );
  NAND2HSV0 U12220 ( .A1(n10599), .A2(\pe10/got [8]), .ZN(n10106) );
  INAND2HSV2 U12221 ( .A1(n10106), .B1(n15075), .ZN(n10786) );
  INHSV2 U12222 ( .I(n6701), .ZN(n10787) );
  NAND2HSV0 U12223 ( .A1(n10786), .A2(n10107), .ZN(n10109) );
  CLKNAND2HSV0 U12224 ( .A1(n10111), .A2(\pe10/got [7]), .ZN(n10117) );
  NOR2HSV0 U12225 ( .A1(\pe10/got [7]), .A2(n14828), .ZN(n10113) );
  AO21HSV1 U12226 ( .A1(n10112), .A2(n14828), .B(n15098), .Z(n10120) );
  NOR2HSV1 U12227 ( .A1(n10125), .A2(n15140), .ZN(n10126) );
  AOI21HSV0 U12228 ( .A1(n10127), .A2(ctro10), .B(n15097), .ZN(n10128) );
  NAND2HSV2 U12229 ( .A1(n14951), .A2(\pe10/bq[3] ), .ZN(n10130) );
  NAND2HSV0 U12230 ( .A1(\pe10/aot [4]), .A2(\pe10/bq[7] ), .ZN(n10129) );
  XOR2HSV0 U12231 ( .A1(n10130), .A2(n10129), .Z(n10134) );
  CLKNAND2HSV1 U12232 ( .A1(\pe10/bq[4] ), .A2(\pe10/aot [7]), .ZN(n10132) );
  NAND2HSV0 U12233 ( .A1(\pe10/got [3]), .A2(\pe10/ti_1 ), .ZN(n10131) );
  XOR2HSV0 U12234 ( .A1(n10132), .A2(n10131), .Z(n10133) );
  XOR2HSV0 U12235 ( .A1(n10134), .A2(n10133), .Z(n10142) );
  NAND2HSV0 U12236 ( .A1(\pe10/ctrq ), .A2(\pe10/pvq [6]), .ZN(n10140) );
  XNOR2HSV4 U12237 ( .A1(n10135), .A2(\pe10/phq [6]), .ZN(n10139) );
  CLKNAND2HSV1 U12238 ( .A1(\pe10/aot [5]), .A2(\pe10/bq[6] ), .ZN(n10137) );
  NAND2HSV0 U12239 ( .A1(\pe10/aot [3]), .A2(\pe10/bq[8] ), .ZN(n10136) );
  XOR2HSV0 U12240 ( .A1(n10137), .A2(n10136), .Z(n10138) );
  XOR3HSV2 U12241 ( .A1(n10140), .A2(n10139), .A3(n10138), .Z(n10141) );
  XNOR2HSV4 U12242 ( .A1(n10142), .A2(n10141), .ZN(n10144) );
  NAND2HSV2 U12243 ( .A1(n14874), .A2(\pe10/got [4]), .ZN(n10143) );
  XNOR2HSV4 U12244 ( .A1(n10144), .A2(n10143), .ZN(n10147) );
  NAND2HSV2 U12245 ( .A1(n10145), .A2(\pe10/got [5]), .ZN(n10146) );
  NAND2HSV0 U12246 ( .A1(n15177), .A2(\pe20/ti_7t [5]), .ZN(n10149) );
  NAND2HSV2 U12247 ( .A1(\pe3/pvq [3]), .A2(\pe3/ctrq ), .ZN(n10152) );
  XNOR2HSV4 U12248 ( .A1(n10152), .A2(n10151), .ZN(n10153) );
  CLKNAND2HSV1 U12249 ( .A1(n10153), .A2(n10154), .ZN(n10158) );
  INHSV2 U12250 ( .I(n10153), .ZN(n10156) );
  INHSV2 U12251 ( .I(n10154), .ZN(n10155) );
  CLKNAND2HSV3 U12252 ( .A1(n10156), .A2(n10155), .ZN(n10157) );
  CLKNAND2HSV3 U12253 ( .A1(n10157), .A2(n10158), .ZN(n10162) );
  CLKNAND2HSV1 U12254 ( .A1(n12475), .A2(\pe3/got [6]), .ZN(n10160) );
  NAND2HSV0 U12255 ( .A1(\pe3/aot [7]), .A2(\pe3/bq[7] ), .ZN(n10159) );
  XNOR2HSV1 U12256 ( .A1(n10160), .A2(n10159), .ZN(n10161) );
  XNOR2HSV4 U12257 ( .A1(n10164), .A2(n10163), .ZN(n10166) );
  XNOR2HSV4 U12258 ( .A1(n10166), .A2(n10165), .ZN(n12351) );
  INHSV2 U12259 ( .I(n10213), .ZN(n10167) );
  NOR2HSV4 U12260 ( .A1(n12351), .A2(n10167), .ZN(n10191) );
  CLKNAND2HSV1 U12261 ( .A1(n10213), .A2(n10168), .ZN(n10189) );
  CLKNAND2HSV1 U12262 ( .A1(n10189), .A2(\pe3/got [7]), .ZN(n10169) );
  INHSV2 U12263 ( .I(ctro3), .ZN(n10188) );
  INHSV2 U12264 ( .I(n10188), .ZN(n10942) );
  INHSV2 U12265 ( .I(n15180), .ZN(n10201) );
  NOR2HSV2 U12266 ( .A1(n10939), .A2(n10201), .ZN(n10995) );
  NAND2HSV2 U12267 ( .A1(n12351), .A2(n10995), .ZN(n10170) );
  CLKNAND2HSV3 U12268 ( .A1(\pe3/got [7]), .A2(\pe3/ti_1 ), .ZN(n10172) );
  INHSV4 U12269 ( .I(\pe3/phq [2]), .ZN(n10171) );
  CLKNAND2HSV3 U12270 ( .A1(n10172), .A2(n10171), .ZN(n10178) );
  NOR2HSV4 U12271 ( .A1(n10172), .A2(n10171), .ZN(n10174) );
  CLKNAND2HSV2 U12272 ( .A1(\pe3/aot [7]), .A2(\pe3/bq[8] ), .ZN(n10175) );
  OAI21HSV4 U12273 ( .A1(n10173), .A2(n10174), .B(n10175), .ZN(n10180) );
  INHSV2 U12274 ( .I(n10175), .ZN(n10176) );
  NAND3HSV3 U12275 ( .A1(n10177), .A2(n10178), .A3(n10176), .ZN(n10179) );
  CLKNAND2HSV3 U12276 ( .A1(n10180), .A2(n10179), .ZN(n10184) );
  XNOR2HSV4 U12277 ( .A1(n10182), .A2(n10181), .ZN(n10183) );
  XNOR2HSV4 U12278 ( .A1(n10184), .A2(n10183), .ZN(n13842) );
  BUFHSV8 U12279 ( .I(\pe3/got [8]), .Z(n15180) );
  AOI21HSV2 U12280 ( .A1(n12351), .A2(n15180), .B(n10939), .ZN(n10187) );
  INHSV3 U12281 ( .I(n13842), .ZN(n10186) );
  CLKAND2HSV2 U12282 ( .A1(n10946), .A2(n15180), .Z(n10406) );
  CLKNAND2HSV0 U12283 ( .A1(n10189), .A2(\pe3/got [6]), .ZN(n10190) );
  NOR2HSV2 U12284 ( .A1(n10191), .A2(n10190), .ZN(n10200) );
  NAND2HSV2 U12285 ( .A1(\pe3/aot [7]), .A2(\pe3/bq[6] ), .ZN(n10193) );
  XNOR2HSV4 U12286 ( .A1(n10193), .A2(n10192), .ZN(n10197) );
  XNOR2HSV4 U12287 ( .A1(n10195), .A2(n10194), .ZN(n10196) );
  BUFHSV4 U12288 ( .I(\pe3/bq[8] ), .Z(n12476) );
  NAND2HSV2 U12289 ( .A1(n12476), .A2(\pe3/aot [5]), .ZN(n10198) );
  BUFHSV6 U12290 ( .I(\pe3/got [7]), .Z(n14931) );
  NAND2HSV2 U12291 ( .A1(n10994), .A2(\pe3/ti_7t [4]), .ZN(n10943) );
  INHSV2 U12292 ( .I(n10943), .ZN(n10944) );
  CLKNHSV0 U12293 ( .I(\pe3/ctrq ), .ZN(n10978) );
  CLKBUFHSV4 U12294 ( .I(\pe3/aot [8]), .Z(n14953) );
  NAND2HSV0 U12295 ( .A1(\pe3/aot [7]), .A2(\pe3/bq[5] ), .ZN(n10206) );
  XOR2HSV0 U12296 ( .A1(n10207), .A2(n10206), .Z(n10210) );
  NAND2HSV0 U12297 ( .A1(\pe3/aot [5]), .A2(\pe3/bq[7] ), .ZN(n10208) );
  XNOR2HSV1 U12298 ( .A1(n10208), .A2(\pe3/phq [5]), .ZN(n10209) );
  XNOR2HSV1 U12299 ( .A1(n10210), .A2(n10209), .ZN(n10211) );
  XNOR2HSV4 U12300 ( .A1(n10212), .A2(n10211), .ZN(n10215) );
  NAND2HSV0 U12301 ( .A1(n10405), .A2(n12351), .ZN(n10214) );
  CLKNAND2HSV1 U12302 ( .A1(n10939), .A2(\pe3/ti_7t [5]), .ZN(n10217) );
  INHSV2 U12303 ( .I(\pe1/got [8]), .ZN(n10260) );
  INHSV4 U12304 ( .I(ctro1), .ZN(n10606) );
  NOR2HSV4 U12305 ( .A1(n10222), .A2(n8931), .ZN(n14956) );
  CLKNAND2HSV1 U12306 ( .A1(n10242), .A2(\pe1/got [7]), .ZN(n10221) );
  NOR2HSV2 U12307 ( .A1(n10616), .A2(n14503), .ZN(n10223) );
  INHSV4 U12308 ( .I(\pe1/bq[6] ), .ZN(n13968) );
  NOR2HSV2 U12309 ( .A1(n10222), .A2(n13968), .ZN(n10238) );
  NAND2HSV2 U12310 ( .A1(\pe1/aot [7]), .A2(\pe1/bq[6] ), .ZN(n10253) );
  OAI22HSV2 U12311 ( .A1(n10223), .A2(n10238), .B1(n10253), .B2(n10225), .ZN(
        n10219) );
  XNOR2HSV4 U12312 ( .A1(n10221), .A2(n10220), .ZN(n10264) );
  NAND2HSV0 U12313 ( .A1(\pe1/aot [7]), .A2(\pe1/bq[8] ), .ZN(n10224) );
  INHSV2 U12314 ( .I(n10226), .ZN(n13838) );
  NOR2HSV2 U12315 ( .A1(n10260), .A2(ctro1), .ZN(n10601) );
  AOI21HSV0 U12316 ( .A1(n14956), .A2(\pe1/got [8]), .B(ctro1), .ZN(n10227) );
  INHSV2 U12317 ( .I(n10228), .ZN(n14868) );
  CLKNAND2HSV1 U12318 ( .A1(n14868), .A2(\pe1/ti_7t [2]), .ZN(n10229) );
  AOI21HSV4 U12319 ( .A1(n13838), .A2(n10232), .B(n10231), .ZN(n10255) );
  INHSV2 U12320 ( .I(\pe1/got [7]), .ZN(n10633) );
  INOR2HSV1 U12321 ( .A1(n10606), .B1(n10633), .ZN(n10233) );
  CLKNAND2HSV1 U12322 ( .A1(pov1[3]), .A2(n10233), .ZN(n10235) );
  AND2HSV2 U12323 ( .A1(ctro1), .A2(\pe1/ti_7t [3]), .Z(n10624) );
  INHSV2 U12324 ( .I(n10633), .ZN(n14703) );
  CLKNAND2HSV0 U12325 ( .A1(n10624), .A2(n14703), .ZN(n10234) );
  NAND2HSV2 U12326 ( .A1(n10235), .A2(n10234), .ZN(n10249) );
  INHSV4 U12327 ( .I(n10255), .ZN(\pe1/ti_7[2] ) );
  NAND2HSV0 U12328 ( .A1(\pe1/ti_7[2] ), .A2(\pe1/got [6]), .ZN(n10241) );
  CLKNHSV0 U12329 ( .I(\pe1/aot [6]), .ZN(n10236) );
  INHSV2 U12330 ( .I(\pe1/bq[4] ), .ZN(n14500) );
  NOR2HSV2 U12331 ( .A1(n10236), .A2(n14500), .ZN(n14000) );
  AOI22HSV0 U12332 ( .A1(\pe1/aot [6]), .A2(\pe1/bq[6] ), .B1(\pe1/aot [8]), 
        .B2(\pe1/bq[4] ), .ZN(n10237) );
  XOR2HSV0 U12333 ( .A1(n10239), .A2(n13971), .Z(n10240) );
  CLKNAND2HSV0 U12334 ( .A1(n10242), .A2(\pe1/got [5]), .ZN(n10245) );
  NAND2HSV2 U12335 ( .A1(\pe1/aot [5]), .A2(n8945), .ZN(n13993) );
  NAND2HSV0 U12336 ( .A1(\pe1/aot [7]), .A2(\pe1/bq[5] ), .ZN(n10243) );
  XOR2HSV0 U12337 ( .A1(n13993), .A2(n10243), .Z(n10244) );
  XOR2HSV0 U12338 ( .A1(n10245), .A2(n10244), .Z(n10246) );
  XNOR2HSV4 U12339 ( .A1(n10249), .A2(n10248), .ZN(n10278) );
  NAND2HSV0 U12340 ( .A1(\pe1/aot [8]), .A2(\pe1/bq[5] ), .ZN(n10251) );
  NAND2HSV0 U12341 ( .A1(\pe1/bq[8] ), .A2(\pe1/aot [5]), .ZN(n10250) );
  NAND2HSV2 U12342 ( .A1(n10242), .A2(\pe1/got [6]), .ZN(n10257) );
  XOR3HSV2 U12343 ( .A1(n10257), .A2(n10258), .A3(n10256), .Z(n10273) );
  NOR2HSV0 U12344 ( .A1(\pe1/ti_7[2] ), .A2(ctro1), .ZN(n10259) );
  NAND2HSV2 U12345 ( .A1(n10259), .A2(n10264), .ZN(n10276) );
  CLKNHSV0 U12346 ( .I(\pe1/ti_7t [3]), .ZN(n10261) );
  AOI21HSV0 U12347 ( .A1(n10261), .A2(ctro1), .B(n10260), .ZN(n10274) );
  CLKNHSV0 U12348 ( .I(n10274), .ZN(n10262) );
  NOR2HSV0 U12349 ( .A1(n10262), .A2(ctro1), .ZN(n10263) );
  NAND2HSV0 U12350 ( .A1(\pe1/ti_7[2] ), .A2(n10606), .ZN(n10266) );
  NAND2HSV0 U12351 ( .A1(ctro1), .A2(\pe1/ti_7t [4]), .ZN(n10270) );
  INHSV2 U12352 ( .I(n10273), .ZN(n13859) );
  NAND3HSV2 U12353 ( .A1(n10276), .A2(n10275), .A3(n10274), .ZN(n13860) );
  NAND2HSV2 U12354 ( .A1(n10627), .A2(n10626), .ZN(n10283) );
  NAND2HSV2 U12355 ( .A1(n10283), .A2(\pe1/got [8]), .ZN(n10277) );
  XNOR2HSV4 U12356 ( .A1(n10278), .A2(n10277), .ZN(pov1[5]) );
  CLKNAND2HSV1 U12357 ( .A1(\pe1/got [8]), .A2(pov1[5]), .ZN(n10602) );
  INHSV2 U12358 ( .I(n10606), .ZN(n10605) );
  INHSV2 U12359 ( .I(n10605), .ZN(n10631) );
  NAND2HSV0 U12360 ( .A1(\pe1/aot [5]), .A2(\pe1/bq[6] ), .ZN(n10280) );
  NAND2HSV0 U12361 ( .A1(\pe1/aot [4]), .A2(\pe1/bq[7] ), .ZN(n10279) );
  CLKNHSV0 U12362 ( .I(\pe1/aot [3]), .ZN(n13969) );
  INHSV2 U12363 ( .I(\pe1/bq[3] ), .ZN(n14539) );
  NOR2HSV2 U12364 ( .A1(n13969), .A2(n14539), .ZN(n12866) );
  CLKNAND2HSV1 U12365 ( .A1(\pe1/aot [7]), .A2(\pe1/bq[4] ), .ZN(n10618) );
  INHSV2 U12366 ( .I(n13884), .ZN(n10284) );
  NAND3HSV2 U12367 ( .A1(n10602), .A2(n10284), .A3(n10631), .ZN(n10286) );
  CLKBUFHSV4 U12368 ( .I(pov1[5]), .Z(n10608) );
  INHSV2 U12369 ( .I(n10603), .ZN(n10285) );
  NAND3HSV4 U12370 ( .A1(n10286), .A2(n10604), .A3(n10285), .ZN(\pe1/ti_7[6] )
         );
  INHSV2 U12371 ( .I(\pe5/ti_7t [1]), .ZN(n10320) );
  CLKNAND2HSV2 U12372 ( .A1(\pe5/ctrq ), .A2(\pe5/pvq [1]), .ZN(n10288) );
  XNOR2HSV4 U12373 ( .A1(n10288), .A2(n10287), .ZN(n10293) );
  CLKNAND2HSV1 U12374 ( .A1(\pe5/got [8]), .A2(\pe5/ti_1 ), .ZN(n10291) );
  CLKNAND2HSV1 U12375 ( .A1(n10289), .A2(\pe5/phq [1]), .ZN(n10290) );
  OAI21HSV2 U12376 ( .A1(\pe5/phq [1]), .A2(n10291), .B(n10290), .ZN(n10292)
         );
  XNOR2HSV4 U12377 ( .A1(n10293), .A2(n10292), .ZN(n10527) );
  NAND2HSV2 U12378 ( .A1(n10346), .A2(\pe5/got [6]), .ZN(n10306) );
  CLKNAND2HSV0 U12379 ( .A1(\pe5/aot [8]), .A2(\pe5/bq[5] ), .ZN(n10295) );
  NAND2HSV0 U12380 ( .A1(\pe5/aot [5]), .A2(\pe5/bq[8] ), .ZN(n10294) );
  XOR2HSV0 U12381 ( .A1(n10295), .A2(n10294), .Z(n10299) );
  NAND2HSV2 U12382 ( .A1(\pe5/got [5]), .A2(\pe5/ti_1 ), .ZN(n10297) );
  NAND2HSV0 U12383 ( .A1(\pe5/bq[7] ), .A2(\pe5/aot [6]), .ZN(n10296) );
  XOR2HSV0 U12384 ( .A1(n10297), .A2(n10296), .Z(n10298) );
  NAND2HSV2 U12385 ( .A1(\pe5/pvq [4]), .A2(\pe5/ctrq ), .ZN(n10300) );
  XNOR2HSV1 U12386 ( .A1(n10300), .A2(\pe5/phq [4]), .ZN(n10302) );
  NAND2HSV0 U12387 ( .A1(\pe5/aot [7]), .A2(\pe5/bq[6] ), .ZN(n10301) );
  XNOR2HSV1 U12388 ( .A1(n10302), .A2(n10301), .ZN(n10303) );
  INHSV2 U12389 ( .I(n10307), .ZN(n10322) );
  NAND2HSV2 U12390 ( .A1(\pe5/aot [7]), .A2(\pe5/bq[8] ), .ZN(n10309) );
  CLKNAND2HSV1 U12391 ( .A1(\pe5/ti_1 ), .A2(\pe5/got [7]), .ZN(n10308) );
  XNOR2HSV1 U12392 ( .A1(n10309), .A2(n10308), .ZN(n10310) );
  XNOR2HSV4 U12393 ( .A1(n10311), .A2(n10310), .ZN(n10312) );
  INHSV2 U12394 ( .I(\pe5/got [8]), .ZN(n10326) );
  NOR2HSV2 U12395 ( .A1(n10326), .A2(ctro5), .ZN(n11473) );
  INHSV4 U12396 ( .I(n10312), .ZN(n13855) );
  INHSV2 U12397 ( .I(n10326), .ZN(n15067) );
  AOI21HSV2 U12398 ( .A1(n10527), .A2(n15067), .B(n10322), .ZN(n10313) );
  NAND2HSV2 U12399 ( .A1(n11492), .A2(\pe5/got [7]), .ZN(n10314) );
  XNOR2HSV4 U12400 ( .A1(n10315), .A2(n10314), .ZN(n11475) );
  INHSV4 U12401 ( .I(n6704), .ZN(n11476) );
  BUFHSV2 U12402 ( .I(\pe5/got [8]), .Z(n13861) );
  NAND2HSV0 U12403 ( .A1(\pe5/ti_1 ), .A2(\pe5/got [6]), .ZN(n10318) );
  NAND2HSV0 U12404 ( .A1(\pe5/aot [6]), .A2(\pe5/bq[8] ), .ZN(n10317) );
  XOR2HSV0 U12405 ( .A1(n10318), .A2(n10317), .Z(n10319) );
  INHSV2 U12406 ( .I(\pe5/got [7]), .ZN(n13429) );
  AOI21HSV2 U12407 ( .A1(n10320), .A2(n10322), .B(n13429), .ZN(n10321) );
  OAI21HSV2 U12408 ( .A1(n10527), .A2(n10322), .B(n10321), .ZN(n10323) );
  NAND2HSV0 U12409 ( .A1(n15067), .A2(n10307), .ZN(n10324) );
  NOR2HSV0 U12410 ( .A1(n15278), .A2(n10324), .ZN(n10325) );
  CLKNAND2HSV0 U12411 ( .A1(n11476), .A2(n10325), .ZN(n10330) );
  CLKAND2HSV1 U12412 ( .A1(n15278), .A2(n11473), .Z(n10328) );
  NAND2HSV2 U12413 ( .A1(n13015), .A2(\pe5/ti_7t [4]), .ZN(n11474) );
  NOR2HSV0 U12414 ( .A1(n11474), .A2(n10326), .ZN(n10327) );
  OR2HSV1 U12415 ( .A1(n13018), .A2(n13861), .Z(n11472) );
  CLKNHSV1 U12416 ( .I(n10332), .ZN(n10352) );
  NAND2HSV0 U12417 ( .A1(\pe5/bq[5] ), .A2(\pe5/aot [7]), .ZN(n10334) );
  NAND2HSV0 U12418 ( .A1(\pe5/aot [4]), .A2(\pe5/bq[8] ), .ZN(n10333) );
  XOR2HSV0 U12419 ( .A1(n10334), .A2(n10333), .Z(n10338) );
  NAND2HSV0 U12420 ( .A1(\pe5/ti_1 ), .A2(\pe5/got [4]), .ZN(n10336) );
  NAND2HSV0 U12421 ( .A1(\pe5/aot [5]), .A2(\pe5/bq[7] ), .ZN(n10335) );
  XOR2HSV0 U12422 ( .A1(n10336), .A2(n10335), .Z(n10337) );
  XOR2HSV0 U12423 ( .A1(n10338), .A2(n10337), .Z(n10345) );
  NAND2HSV0 U12424 ( .A1(\pe5/aot [6]), .A2(\pe5/bq[6] ), .ZN(n10340) );
  NAND2HSV0 U12425 ( .A1(\pe5/aot [8]), .A2(\pe5/bq[4] ), .ZN(n10339) );
  XOR2HSV0 U12426 ( .A1(n10340), .A2(n10339), .Z(n10343) );
  NAND2HSV0 U12427 ( .A1(\pe5/pvq [5]), .A2(\pe5/ctrq ), .ZN(n10341) );
  XOR2HSV0 U12428 ( .A1(n10341), .A2(\pe5/phq [5]), .Z(n10342) );
  XOR2HSV0 U12429 ( .A1(n10343), .A2(n10342), .Z(n10344) );
  XOR2HSV0 U12430 ( .A1(n10345), .A2(n10344), .Z(n10348) );
  NAND2HSV2 U12431 ( .A1(n10346), .A2(\pe5/got [5]), .ZN(n10347) );
  XNOR2HSV4 U12432 ( .A1(n10348), .A2(n10347), .ZN(n10350) );
  NAND2HSV0 U12433 ( .A1(n11492), .A2(\pe5/got [6]), .ZN(n10349) );
  NAND2HSV2 U12434 ( .A1(n13018), .A2(\pe5/ti_7t [5]), .ZN(n13284) );
  NOR2HSV2 U12435 ( .A1(n10355), .A2(n12135), .ZN(n10354) );
  INHSV2 U12436 ( .I(n10354), .ZN(n12141) );
  INHSV2 U12437 ( .I(n10356), .ZN(n12140) );
  INHSV2 U12438 ( .I(n12140), .ZN(n11712) );
  OAI21HSV4 U12439 ( .A1(n10359), .A2(n10360), .B(n10358), .ZN(n10363) );
  INHSV4 U12440 ( .I(n10361), .ZN(n13810) );
  NAND2HSV2 U12441 ( .A1(n13810), .A2(\pe21/aot [7]), .ZN(n10362) );
  XNOR2HSV4 U12442 ( .A1(n10363), .A2(n10362), .ZN(n10369) );
  INHSV4 U12443 ( .I(n10369), .ZN(n10367) );
  NAND2HSV0 U12444 ( .A1(\pe21/ti_1 ), .A2(\pe21/got [7]), .ZN(n10365) );
  CLKNAND2HSV3 U12445 ( .A1(n10369), .A2(n10368), .ZN(n10376) );
  INHSV2 U12446 ( .I(\pe21/got [8]), .ZN(n10862) );
  NOR2HSV2 U12447 ( .A1(n10862), .A2(n10863), .ZN(n10869) );
  INHSV2 U12448 ( .I(n10400), .ZN(n10389) );
  CLKBUFHSV4 U12449 ( .I(ctro21), .Z(n10863) );
  INHSV2 U12450 ( .I(\pe21/got [8]), .ZN(n10837) );
  CLKNAND2HSV4 U12451 ( .A1(n10379), .A2(n10378), .ZN(n10401) );
  CLKNHSV0 U12452 ( .I(n10401), .ZN(n10380) );
  INHSV4 U12453 ( .I(\pe21/ctrq ), .ZN(n14540) );
  NAND2HSV2 U12454 ( .A1(n11786), .A2(\pe21/pvq [3]), .ZN(n10382) );
  NAND2HSV0 U12455 ( .A1(\pe21/bq[8] ), .A2(\pe21/aot [6]), .ZN(n10381) );
  XOR2HSV0 U12456 ( .A1(n10382), .A2(n10381), .Z(n10383) );
  XNOR2HSV4 U12457 ( .A1(n10384), .A2(n10383), .ZN(n10414) );
  XNOR2HSV4 U12458 ( .A1(n10414), .A2(n10413), .ZN(n10392) );
  NOR2HSV2 U12459 ( .A1(n10389), .A2(n10388), .ZN(n10391) );
  INHSV2 U12460 ( .I(n10837), .ZN(n10415) );
  CLKNAND2HSV1 U12461 ( .A1(n10644), .A2(n10415), .ZN(n10390) );
  INHSV2 U12462 ( .I(n10873), .ZN(n10853) );
  NAND2HSV2 U12463 ( .A1(\pe21/ti_7t [4]), .A2(n10403), .ZN(n10854) );
  NAND2HSV2 U12464 ( .A1(n6207), .A2(n10854), .ZN(n15175) );
  AND2HSV2 U12465 ( .A1(n10789), .A2(n10406), .Z(n10407) );
  AND2HSV2 U12466 ( .A1(n8942), .A2(n10410), .Z(n10411) );
  BUFHSV8 U12467 ( .I(n6710), .Z(n14916) );
  XNOR2HSV4 U12468 ( .A1(n10414), .A2(n10413), .ZN(n10809) );
  NAND2HSV2 U12469 ( .A1(n11780), .A2(\pe21/ti_7t [3]), .ZN(n10841) );
  OAI21HSV4 U12470 ( .A1(n10865), .A2(n6435), .B(n10841), .ZN(\pe21/ti_7[3] )
         );
  INHSV4 U12471 ( .I(ctro17), .ZN(n12014) );
  INHSV2 U12472 ( .I(n10418), .ZN(n10526) );
  INHSV2 U12473 ( .I(n12014), .ZN(n12130) );
  CLKNAND2HSV1 U12474 ( .A1(n10526), .A2(n12130), .ZN(n10431) );
  INHSV2 U12475 ( .I(\pe17/got [7]), .ZN(n10435) );
  NAND2HSV2 U12476 ( .A1(n10431), .A2(n14429), .ZN(n10419) );
  NAND2HSV0 U12477 ( .A1(\pe17/got [6]), .A2(\pe17/ti_1 ), .ZN(n10420) );
  XNOR2HSV4 U12478 ( .A1(n10473), .A2(n10472), .ZN(n10423) );
  INHSV2 U12479 ( .I(n12130), .ZN(n13252) );
  INHSV2 U12480 ( .I(\pe17/got [8]), .ZN(n14397) );
  NOR2HSV2 U12481 ( .A1(n12021), .A2(n14397), .ZN(n14007) );
  NAND2HSV2 U12482 ( .A1(n12021), .A2(\pe17/ti_7t [2]), .ZN(n10469) );
  NOR2HSV1 U12483 ( .A1(n8928), .A2(\pe17/ti_7t [3]), .ZN(n10716) );
  CLKBUFHSV4 U12484 ( .I(\pe17/aot [8]), .Z(n14949) );
  NAND2HSV2 U12485 ( .A1(\pe17/ctrq ), .A2(\pe17/pvq [4]), .ZN(n10424) );
  XNOR2HSV4 U12486 ( .A1(n10424), .A2(\pe17/phq [4]), .ZN(n10428) );
  CLKNHSV1 U12487 ( .I(\pe17/aot [5]), .ZN(n10426) );
  CLKNHSV0 U12488 ( .I(\pe17/bq[8] ), .ZN(n10425) );
  NOR2HSV2 U12489 ( .A1(n10426), .A2(n10425), .ZN(n10427) );
  XNOR2HSV1 U12490 ( .A1(n10428), .A2(n10427), .ZN(n10429) );
  CLKNAND2HSV0 U12491 ( .A1(n10431), .A2(\pe17/got [6]), .ZN(n10432) );
  NOR2HSV2 U12492 ( .A1(n10433), .A2(n10432), .ZN(n10434) );
  INHSV2 U12493 ( .I(n13268), .ZN(n14010) );
  INHSV2 U12494 ( .I(n14010), .ZN(n12043) );
  AND2HSV2 U12495 ( .A1(n12043), .A2(n14429), .Z(n10437) );
  INHSV2 U12496 ( .I(\pe17/got [7]), .ZN(n14333) );
  NOR2HSV1 U12497 ( .A1(n10469), .A2(n14333), .ZN(n10436) );
  INHSV2 U12498 ( .I(n10471), .ZN(n10439) );
  NOR2HSV2 U12499 ( .A1(n12014), .A2(n15080), .ZN(n12132) );
  INHSV2 U12500 ( .I(n12132), .ZN(n12131) );
  INHSV2 U12501 ( .I(n12131), .ZN(n10440) );
  NAND2HSV2 U12502 ( .A1(n10442), .A2(n10441), .ZN(n10443) );
  INHSV2 U12503 ( .I(n15273), .ZN(n10445) );
  BUFHSV4 U12504 ( .I(ctro7), .Z(n12311) );
  INHSV2 U12505 ( .I(n5967), .ZN(n12266) );
  NOR2HSV2 U12506 ( .A1(n12311), .A2(n12266), .ZN(n12273) );
  INHSV1 U12507 ( .I(n12273), .ZN(n10444) );
  NOR2HSV4 U12508 ( .A1(n10445), .A2(n10444), .ZN(n10457) );
  INHSV4 U12509 ( .I(\pe7/phq [2]), .ZN(n10448) );
  CLKNAND2HSV3 U12510 ( .A1(n10447), .A2(n10448), .ZN(n10446) );
  OAI21HSV4 U12511 ( .A1(n10448), .A2(n10447), .B(n10446), .ZN(n10450) );
  NAND2HSV0 U12512 ( .A1(\pe7/ctrq ), .A2(\pe7/pvq [2]), .ZN(n10449) );
  XNOR2HSV4 U12513 ( .A1(n10450), .A2(n10449), .ZN(n10455) );
  INHSV2 U12514 ( .I(\pe7/bq[8] ), .ZN(n11801) );
  INHSV2 U12515 ( .I(\pe7/aot [7]), .ZN(n10451) );
  NOR2HSV2 U12516 ( .A1(n11801), .A2(n10451), .ZN(n10453) );
  NAND2HSV0 U12517 ( .A1(\pe7/bq[7] ), .A2(\pe7/aot [8]), .ZN(n10452) );
  XNOR2HSV4 U12518 ( .A1(n10455), .A2(n10454), .ZN(n10458) );
  CLKAND2HSV2 U12519 ( .A1(n12267), .A2(\pe7/ti_7t [2]), .Z(n10456) );
  AOI21HSV4 U12520 ( .A1(n10457), .A2(n10458), .B(n10456), .ZN(n12060) );
  INHSV4 U12521 ( .I(n12201), .ZN(n12204) );
  INHSV2 U12522 ( .I(\pe7/ti_7t [1]), .ZN(n10460) );
  NOR2HSV2 U12523 ( .A1(n11782), .A2(n10460), .ZN(n10461) );
  NOR2HSV4 U12524 ( .A1(n15273), .A2(n10461), .ZN(n12074) );
  INHSV2 U12525 ( .I(n10461), .ZN(n11783) );
  CLKNAND2HSV1 U12526 ( .A1(n11783), .A2(n12267), .ZN(n12072) );
  CLKNAND2HSV1 U12527 ( .A1(n12072), .A2(\pe7/got [7]), .ZN(n10462) );
  NOR2HSV4 U12528 ( .A1(n12074), .A2(n10462), .ZN(n12058) );
  NAND2HSV0 U12529 ( .A1(\pe7/aot [6]), .A2(\pe7/bq[8] ), .ZN(n10467) );
  NAND2HSV2 U12530 ( .A1(\pe7/ctrq ), .A2(\pe7/pvq [3]), .ZN(n10463) );
  XOR2HSV2 U12531 ( .A1(n10463), .A2(\pe7/phq [3]), .Z(n10466) );
  BUFHSV4 U12532 ( .I(\pe7/ti_1 ), .Z(n14480) );
  CLKNAND2HSV1 U12533 ( .A1(n14480), .A2(\pe7/got [6]), .ZN(n10465) );
  XOR4HSV4 U12534 ( .A1(n10467), .A2(n10466), .A3(n10465), .A4(n10464), .Z(
        n12057) );
  XNOR2HSV4 U12535 ( .A1(n12058), .A2(n12057), .ZN(n12203) );
  XNOR2HSV4 U12536 ( .A1(n12204), .A2(n12203), .ZN(n15271) );
  CLKNAND2HSV1 U12537 ( .A1(n12311), .A2(\pe7/ti_7t [3]), .ZN(n12280) );
  INHSV2 U12538 ( .I(n12020), .ZN(n12022) );
  INHSV2 U12539 ( .I(\pe17/got [2]), .ZN(n14400) );
  INHSV4 U12540 ( .I(\pe8/phq [2]), .ZN(n10476) );
  CLKNAND2HSV2 U12541 ( .A1(n10475), .A2(n10476), .ZN(n10474) );
  OAI21HSV4 U12542 ( .A1(n10476), .A2(n10475), .B(n10474), .ZN(n10478) );
  BUFHSV8 U12543 ( .I(\pe8/ctrq ), .Z(n11574) );
  NAND2HSV2 U12544 ( .A1(n11574), .A2(\pe8/pvq [2]), .ZN(n10477) );
  XNOR2HSV4 U12545 ( .A1(n10478), .A2(n10477), .ZN(n10482) );
  INHSV2 U12546 ( .I(\pe8/aot [7]), .ZN(n10496) );
  INHSV2 U12547 ( .I(\pe8/bq[8] ), .ZN(n13516) );
  CLKNAND2HSV0 U12548 ( .A1(\pe8/got [7]), .A2(\pe8/ti_1 ), .ZN(n10479) );
  XNOR2HSV4 U12549 ( .A1(n10482), .A2(n10481), .ZN(n10489) );
  NAND2HSV2 U12550 ( .A1(\pe8/bq[8] ), .A2(\pe8/aot [8]), .ZN(n10483) );
  AOI21HSV2 U12551 ( .A1(\pe8/ctrq ), .A2(\pe8/pvq [1]), .B(\pe8/phq [1]), 
        .ZN(n10485) );
  AOI21HSV2 U12552 ( .A1(n11796), .A2(\pe8/got [8]), .B(n12372), .ZN(n10487)
         );
  CLKNAND2HSV2 U12553 ( .A1(n6700), .A2(n10487), .ZN(n10506) );
  INHSV2 U12554 ( .I(ctro8), .ZN(n15082) );
  INHSV2 U12555 ( .I(n15082), .ZN(n12372) );
  NAND2HSV2 U12556 ( .A1(n11602), .A2(n11796), .ZN(n10488) );
  INHSV2 U12557 ( .I(n10488), .ZN(n10490) );
  AOI22HSV4 U12558 ( .A1(n12372), .A2(\pe8/ti_7t [2]), .B1(n10490), .B2(n10489), .ZN(n10507) );
  NAND3HSV2 U12559 ( .A1(n10506), .A2(n10507), .A3(n11591), .ZN(n11515) );
  INHSV2 U12560 ( .I(n10508), .ZN(n14189) );
  NOR2HSV2 U12561 ( .A1(\pe8/got [8]), .A2(n14189), .ZN(n11538) );
  INHSV2 U12562 ( .I(n14838), .ZN(n10491) );
  NAND2HSV2 U12563 ( .A1(n10491), .A2(\pe8/bq[6] ), .ZN(n10493) );
  CLKNAND2HSV1 U12564 ( .A1(\pe8/ti_1 ), .A2(\pe8/got [6]), .ZN(n10492) );
  XNOR2HSV4 U12565 ( .A1(n10493), .A2(n10492), .ZN(n10495) );
  CLKNAND2HSV1 U12566 ( .A1(\pe8/aot [6]), .A2(\pe8/bq[8] ), .ZN(n13518) );
  XNOR2HSV4 U12567 ( .A1(n13518), .A2(\pe8/phq [3]), .ZN(n10494) );
  XNOR2HSV4 U12568 ( .A1(n10495), .A2(n10494), .ZN(n10501) );
  INHSV1 U12569 ( .I(n10496), .ZN(n10497) );
  INHSV2 U12570 ( .I(n15132), .ZN(n13825) );
  NAND2HSV2 U12571 ( .A1(n10497), .A2(n13825), .ZN(n10499) );
  INHSV2 U12572 ( .I(\pe8/ctrq ), .ZN(n11848) );
  XNOR2HSV4 U12573 ( .A1(n10499), .A2(n10498), .ZN(n10500) );
  XNOR2HSV4 U12574 ( .A1(n10501), .A2(n10500), .ZN(n10505) );
  CLKNHSV0 U12575 ( .I(\pe8/ti_7t [1]), .ZN(n10502) );
  INHSV2 U12576 ( .I(\pe8/got [7]), .ZN(n11513) );
  AOI21HSV2 U12577 ( .A1(n10502), .A2(n11521), .B(n11513), .ZN(n10503) );
  OAI21HSV2 U12578 ( .A1(n11796), .A2(n14189), .B(n10503), .ZN(n10504) );
  XNOR2HSV4 U12579 ( .A1(n10505), .A2(n10504), .ZN(n11523) );
  NAND2HSV2 U12580 ( .A1(n12372), .A2(\pe8/ti_7t [3]), .ZN(n11512) );
  INHSV2 U12581 ( .I(n11523), .ZN(n11511) );
  NAND2HSV4 U12582 ( .A1(n10507), .A2(n10506), .ZN(n11580) );
  INHSV2 U12583 ( .I(n11580), .ZN(n15079) );
  INHSV2 U12584 ( .I(n10508), .ZN(n14190) );
  OR2HSV1 U12585 ( .A1(n11603), .A2(n14190), .Z(n10509) );
  NAND2HSV2 U12586 ( .A1(n11511), .A2(n11516), .ZN(n11563) );
  CLKNAND2HSV1 U12587 ( .A1(n9680), .A2(\pe4/ti_7t [3]), .ZN(n10511) );
  CLKNAND2HSV1 U12588 ( .A1(\pe15/pvq [2]), .A2(\pe15/ctrq ), .ZN(n10513) );
  XNOR2HSV4 U12589 ( .A1(n10514), .A2(n10513), .ZN(n10518) );
  NAND2HSV0 U12590 ( .A1(\pe15/got [7]), .A2(\pe15/ti_1 ), .ZN(n10516) );
  NAND2HSV0 U12591 ( .A1(\pe15/bq[7] ), .A2(\pe15/aot [8]), .ZN(n10515) );
  XOR2HSV2 U12592 ( .A1(n10516), .A2(n10515), .Z(n10517) );
  XNOR2HSV4 U12593 ( .A1(n10518), .A2(n10517), .ZN(n13857) );
  INHSV2 U12594 ( .I(\pe15/ti_7t [2]), .ZN(n10520) );
  INHSV2 U12595 ( .I(\pe15/got [8]), .ZN(n11405) );
  NOR2HSV0 U12596 ( .A1(n14704), .A2(n11405), .ZN(n10519) );
  NOR2HSV2 U12597 ( .A1(n10522), .A2(n11405), .ZN(n12336) );
  CLKNHSV0 U12598 ( .I(n11390), .ZN(n12830) );
  INHSV2 U12599 ( .I(\pe16/got [8]), .ZN(n14297) );
  NOR2HSV2 U12600 ( .A1(n14297), .A2(n8957), .ZN(n14064) );
  NAND2HSV2 U12601 ( .A1(n10689), .A2(\pe16/ti_7t [2]), .ZN(n10678) );
  INHSV2 U12602 ( .I(\pe16/got [8]), .ZN(n11181) );
  INHSV2 U12603 ( .I(n11181), .ZN(n12194) );
  INHSV1 U12604 ( .I(ctro12), .ZN(n10525) );
  NAND2HSV2 U12605 ( .A1(n11447), .A2(\pe12/ti_7t [1]), .ZN(n10729) );
  INHSV2 U12606 ( .I(n15090), .ZN(n12353) );
  CLKNHSV1 U12607 ( .I(n10527), .ZN(n14881) );
  INHSV1 U12608 ( .I(n10528), .ZN(n14901) );
  INHSV2 U12609 ( .I(\pe16/got [7]), .ZN(n10676) );
  INHSV2 U12610 ( .I(n10676), .ZN(n14873) );
  BUFHSV2 U12611 ( .I(\pe15/ctrq ), .Z(n15160) );
  CLKNHSV0 U12612 ( .I(\pe15/bq[8] ), .ZN(n10529) );
  INHSV2 U12613 ( .I(n10529), .ZN(n14602) );
  MUX2HSV2 U12614 ( .I0(bo15[8]), .I1(n14602), .S(n15160), .Z(n15155) );
  BUFHSV2 U12615 ( .I(\pe15/aot [8]), .Z(n14937) );
  BUFHSV2 U12616 ( .I(\pe15/aot [7]), .Z(n14936) );
  INHSV2 U12617 ( .I(\pe12/aot [8]), .ZN(n10735) );
  CLKNHSV0 U12618 ( .I(n10735), .ZN(n14876) );
  INHSV2 U12619 ( .I(n14869), .ZN(n14870) );
  CLKBUFHSV2 U12620 ( .I(\pe7/aot [6]), .Z(n14705) );
  CLKBUFHSV2 U12621 ( .I(\pe8/aot [6]), .Z(n14947) );
  NAND2HSV2 U12622 ( .A1(n15188), .A2(\pe13/got [1]), .ZN(n10533) );
  CLKNAND2HSV1 U12623 ( .A1(\pe13/aot [1]), .A2(\pe13/bq[2] ), .ZN(n10531) );
  CLKNAND2HSV0 U12624 ( .A1(\pe13/bq[1] ), .A2(\pe13/aot [2]), .ZN(n10530) );
  XOR2HSV0 U12625 ( .A1(n10531), .A2(n10530), .Z(n10532) );
  XOR2HSV0 U12626 ( .A1(n10533), .A2(n10532), .Z(n10534) );
  NAND2HSV2 U12627 ( .A1(n10535), .A2(\pe4/ti_7t [5]), .ZN(n12604) );
  INHSV2 U12628 ( .I(n12604), .ZN(n10582) );
  INHSV2 U12629 ( .I(n10582), .ZN(n11284) );
  BUFHSV4 U12630 ( .I(n14933), .Z(n12631) );
  NAND2HSV0 U12631 ( .A1(n10537), .A2(\pe4/got [3]), .ZN(n10539) );
  NAND2HSV0 U12632 ( .A1(\pe4/ti_7[1] ), .A2(\pe4/got [2]), .ZN(n10538) );
  CLKNAND2HSV0 U12633 ( .A1(n10562), .A2(\pe4/pq ), .ZN(n10541) );
  NAND2HSV0 U12634 ( .A1(\pe4/aot [7]), .A2(\pe4/bq[2] ), .ZN(n10540) );
  XOR2HSV0 U12635 ( .A1(n10541), .A2(n10540), .Z(n10545) );
  CLKNAND2HSV0 U12636 ( .A1(n12581), .A2(\pe4/aot [3]), .ZN(n10543) );
  NAND2HSV0 U12637 ( .A1(\pe4/aot [2]), .A2(\pe4/bq[7] ), .ZN(n10542) );
  XOR2HSV0 U12638 ( .A1(n10543), .A2(n10542), .Z(n10544) );
  XOR2HSV0 U12639 ( .A1(n10545), .A2(n10544), .Z(n10549) );
  NAND2HSV0 U12640 ( .A1(\pe4/bq[4] ), .A2(\pe4/aot [5]), .ZN(n10547) );
  NAND2HSV0 U12641 ( .A1(\pe4/bq[5] ), .A2(\pe4/aot [4]), .ZN(n10546) );
  XOR2HSV0 U12642 ( .A1(n10547), .A2(n10546), .Z(n10548) );
  XNOR2HSV1 U12643 ( .A1(n10549), .A2(n10548), .ZN(n10557) );
  NAND2HSV0 U12644 ( .A1(\pe4/aot [6]), .A2(\pe4/bq[3] ), .ZN(n10551) );
  NAND2HSV0 U12645 ( .A1(n8927), .A2(\pe4/got [1]), .ZN(n10550) );
  XOR2HSV0 U12646 ( .A1(n10551), .A2(n10550), .Z(n10555) );
  NAND2HSV0 U12647 ( .A1(n14843), .A2(\pe4/bq[1] ), .ZN(n10553) );
  NAND2HSV0 U12648 ( .A1(n13823), .A2(\pe4/aot [1]), .ZN(n10552) );
  XOR2HSV0 U12649 ( .A1(n10553), .A2(n10552), .Z(n10554) );
  XOR2HSV0 U12650 ( .A1(n10555), .A2(n10554), .Z(n10556) );
  XNOR2HSV1 U12651 ( .A1(n10557), .A2(n10556), .ZN(n10558) );
  NAND2HSV2 U12652 ( .A1(n14933), .A2(\pe4/got [6]), .ZN(n10580) );
  NAND2HSV0 U12653 ( .A1(\pe4/ti_7[1] ), .A2(\pe4/got [3]), .ZN(n10577) );
  NAND2HSV0 U12654 ( .A1(n14733), .A2(\pe4/got [4]), .ZN(n10576) );
  CLKNAND2HSV1 U12655 ( .A1(\pe4/aot [5]), .A2(\pe4/bq[5] ), .ZN(n12633) );
  NAND2HSV0 U12656 ( .A1(\pe4/aot [3]), .A2(\pe4/bq[7] ), .ZN(n10559) );
  XOR2HSV0 U12657 ( .A1(n12633), .A2(n10559), .Z(n10574) );
  NAND2HSV0 U12658 ( .A1(\pe4/aot [6]), .A2(\pe4/bq[4] ), .ZN(n10561) );
  NAND2HSV0 U12659 ( .A1(n12636), .A2(\pe4/bq[3] ), .ZN(n10560) );
  XOR2HSV0 U12660 ( .A1(n10561), .A2(n10560), .Z(n10565) );
  NAND2HSV2 U12661 ( .A1(\pe4/pvq [7]), .A2(n10562), .ZN(n10563) );
  XNOR2HSV1 U12662 ( .A1(n10563), .A2(\pe4/phq [7]), .ZN(n10564) );
  XNOR2HSV1 U12663 ( .A1(n10565), .A2(n10564), .ZN(n10573) );
  NAND2HSV0 U12664 ( .A1(\pe4/aot [4]), .A2(\pe4/bq[6] ), .ZN(n10567) );
  NAND2HSV0 U12665 ( .A1(n8927), .A2(\pe4/got [2]), .ZN(n10566) );
  XOR2HSV0 U12666 ( .A1(n10567), .A2(n10566), .Z(n10571) );
  CLKNAND2HSV0 U12667 ( .A1(n14843), .A2(\pe4/bq[2] ), .ZN(n10569) );
  NAND2HSV0 U12668 ( .A1(n13823), .A2(\pe4/aot [2]), .ZN(n10568) );
  XOR2HSV0 U12669 ( .A1(n10569), .A2(n10568), .Z(n10570) );
  XOR2HSV0 U12670 ( .A1(n10571), .A2(n10570), .Z(n10572) );
  XOR3HSV2 U12671 ( .A1(n10574), .A2(n10573), .A3(n10572), .Z(n10575) );
  XOR3HSV2 U12672 ( .A1(n10577), .A2(n10575), .A3(n10576), .Z(n10578) );
  XNOR2HSV4 U12673 ( .A1(n10579), .A2(n10578), .ZN(n10581) );
  CLKNAND2HSV0 U12674 ( .A1(\pe4/got [8]), .A2(n12271), .ZN(n10584) );
  CLKNAND2HSV0 U12675 ( .A1(n12604), .A2(n9680), .ZN(n12656) );
  NAND2HSV2 U12676 ( .A1(n12656), .A2(\pe4/got [7]), .ZN(n10587) );
  NAND2HSV2 U12677 ( .A1(n14861), .A2(\pe4/ti_7t [7]), .ZN(n12598) );
  INHSV2 U12678 ( .I(n12598), .ZN(n12591) );
  NAND2HSV0 U12679 ( .A1(n10058), .A2(\pe10/ti_7t [7]), .ZN(n13900) );
  INHSV2 U12680 ( .I(n13900), .ZN(n13902) );
  INHSV2 U12681 ( .I(n13902), .ZN(n10590) );
  NAND2HSV0 U12682 ( .A1(n12602), .A2(\pe4/got [8]), .ZN(n10600) );
  XNOR2HSV0 U12683 ( .A1(n10600), .A2(n12595), .ZN(n15280) );
  CLKAND2HSV2 U12684 ( .A1(n10605), .A2(\pe1/ti_7t [5]), .Z(n10628) );
  OA21HSV2 U12685 ( .A1(n10628), .A2(n10606), .B(n14703), .Z(n10607) );
  OAI21HSV4 U12686 ( .A1(n10608), .A2(n10628), .B(n10607), .ZN(n13258) );
  NAND2HSV0 U12687 ( .A1(\pe1/aot [8]), .A2(\pe1/bq[2] ), .ZN(n10610) );
  NAND2HSV0 U12688 ( .A1(\pe1/aot [5]), .A2(\pe1/bq[5] ), .ZN(n10609) );
  XOR2HSV0 U12689 ( .A1(n10610), .A2(n10609), .Z(n10614) );
  CLKNAND2HSV0 U12690 ( .A1(\pe1/aot [4]), .A2(\pe1/bq[6] ), .ZN(n10612) );
  NAND2HSV0 U12691 ( .A1(\pe1/aot [3]), .A2(\pe1/bq[7] ), .ZN(n10611) );
  XOR2HSV0 U12692 ( .A1(n10612), .A2(n10611), .Z(n10613) );
  XOR2HSV0 U12693 ( .A1(n10614), .A2(n10613), .Z(n10615) );
  OAI21HSV2 U12694 ( .A1(n13965), .A2(n10618), .B(n10617), .ZN(n10620) );
  NAND2HSV0 U12695 ( .A1(\pe1/aot [2]), .A2(\pe1/bq[8] ), .ZN(n10619) );
  XNOR2HSV1 U12696 ( .A1(n10620), .A2(n10619), .ZN(n10622) );
  NAND2HSV0 U12697 ( .A1(n10242), .A2(\pe1/got [3]), .ZN(n10621) );
  XOR2HSV0 U12698 ( .A1(n10622), .A2(n10621), .Z(n10623) );
  INHSV2 U12699 ( .I(\pe1/got [5]), .ZN(n10625) );
  INHSV2 U12700 ( .I(n10634), .ZN(n13256) );
  NAND2HSV2 U12701 ( .A1(pov1[5]), .A2(n10631), .ZN(n10630) );
  INHSV2 U12702 ( .I(n10628), .ZN(n10629) );
  NAND2HSV4 U12703 ( .A1(n10630), .A2(n10629), .ZN(\pe1/ti_7[5] ) );
  OAI21HSV1 U12704 ( .A1(n10634), .A2(n14703), .B(n10631), .ZN(n10632) );
  NOR2HSV1 U12705 ( .A1(n13256), .A2(n10633), .ZN(n10636) );
  NOR2HSV1 U12706 ( .A1(\pe1/ti_7[5] ), .A2(n10634), .ZN(n10635) );
  AOI21HSV1 U12707 ( .A1(n10636), .A2(\pe1/ti_7[5] ), .B(n10635), .ZN(n10637)
         );
  NAND2HSV2 U12708 ( .A1(n14868), .A2(\pe1/ti_7t [7]), .ZN(n10638) );
  NOR2HSV0 U12709 ( .A1(n10853), .A2(n10862), .ZN(n10641) );
  INHSV2 U12710 ( .I(\pe21/ti_7t [4]), .ZN(n10835) );
  OR2HSV1 U12711 ( .A1(n10873), .A2(n10835), .Z(n10808) );
  OR2HSV1 U12712 ( .A1(n10808), .A2(n10862), .Z(n10642) );
  INHSV2 U12713 ( .I(\pe21/got [7]), .ZN(n10860) );
  INHSV2 U12714 ( .I(n10860), .ZN(n13107) );
  NAND2HSV0 U12715 ( .A1(\pe21/bq[6] ), .A2(\pe21/aot [6]), .ZN(n10647) );
  NAND2HSV0 U12716 ( .A1(\pe21/ti_1 ), .A2(\pe21/got [4]), .ZN(n10646) );
  XOR2HSV2 U12717 ( .A1(n10647), .A2(n10646), .Z(n10656) );
  NAND2HSV0 U12718 ( .A1(\pe21/bq[4] ), .A2(\pe21/aot [8]), .ZN(n10842) );
  XOR2HSV2 U12719 ( .A1(n10648), .A2(n10842), .Z(n10655) );
  NAND2HSV0 U12720 ( .A1(\pe21/bq[5] ), .A2(\pe21/aot [7]), .ZN(n10650) );
  NAND2HSV2 U12721 ( .A1(\pe21/aot [4]), .A2(n13810), .ZN(n10649) );
  XNOR2HSV4 U12722 ( .A1(n10650), .A2(n10649), .ZN(n10653) );
  XNOR2HSV4 U12723 ( .A1(n10651), .A2(\pe21/phq [5]), .ZN(n10652) );
  XNOR2HSV4 U12724 ( .A1(n10653), .A2(n10652), .ZN(n10654) );
  XNOR2HSV4 U12725 ( .A1(n10659), .A2(n10658), .ZN(n10660) );
  CLKNAND2HSV3 U12726 ( .A1(n14570), .A2(\pe16/pvq [3]), .ZN(n10663) );
  XNOR2HSV4 U12727 ( .A1(n10663), .A2(n10662), .ZN(n10666) );
  XNOR2HSV1 U12728 ( .A1(n10664), .A2(\pe16/phq [3]), .ZN(n10665) );
  XNOR2HSV4 U12729 ( .A1(n10666), .A2(n10665), .ZN(n10670) );
  CLKNAND2HSV1 U12730 ( .A1(\pe16/aot [8]), .A2(\pe16/bq[6] ), .ZN(n10668) );
  CLKBUFHSV2 U12731 ( .I(\pe16/ti_1 ), .Z(n14266) );
  CLKNAND2HSV1 U12732 ( .A1(\pe16/got [6]), .A2(n14266), .ZN(n10667) );
  XOR2HSV0 U12733 ( .A1(n10668), .A2(n10667), .Z(n10669) );
  INHSV2 U12734 ( .I(n8957), .ZN(n11207) );
  NOR2HSV2 U12735 ( .A1(n10796), .A2(\pe16/ti_7t [3]), .ZN(n10706) );
  NOR2HSV2 U12736 ( .A1(n10706), .A2(n14297), .ZN(n11205) );
  INHSV2 U12737 ( .I(n10676), .ZN(n14292) );
  INHSV2 U12738 ( .I(n14292), .ZN(n13229) );
  INHSV1 U12739 ( .I(n10680), .ZN(n10681) );
  INHSV2 U12740 ( .I(\pe16/phq [4]), .ZN(n10685) );
  INHSV2 U12741 ( .I(\pe16/ctrq ), .ZN(n11827) );
  INHSV2 U12742 ( .I(\pe16/pvq [4]), .ZN(n10683) );
  INHSV2 U12743 ( .I(\pe16/got [5]), .ZN(n14363) );
  INHSV2 U12744 ( .I(\pe16/ti_1 ), .ZN(n13833) );
  NOR2HSV2 U12745 ( .A1(n14363), .A2(n13833), .ZN(n10684) );
  CLKNAND2HSV1 U12746 ( .A1(n10686), .A2(\pe16/got [6]), .ZN(n10687) );
  INHSV4 U12747 ( .I(n10689), .ZN(n14066) );
  NAND2HSV2 U12748 ( .A1(n10689), .A2(\pe16/ti_7t [4]), .ZN(n11157) );
  INHSV2 U12749 ( .I(n14297), .ZN(n11179) );
  CLKNAND2HSV1 U12750 ( .A1(\pe16/bq[6] ), .A2(\pe16/aot [6]), .ZN(n10692) );
  NAND2HSV0 U12751 ( .A1(\pe16/aot [5]), .A2(\pe16/bq[7] ), .ZN(n10691) );
  XOR2HSV0 U12752 ( .A1(n10692), .A2(n10691), .Z(n10696) );
  NAND2HSV0 U12753 ( .A1(\pe16/aot [4]), .A2(\pe16/bq[8] ), .ZN(n10694) );
  NAND2HSV0 U12754 ( .A1(\pe16/got [4]), .A2(\pe16/ti_1 ), .ZN(n10693) );
  XOR2HSV0 U12755 ( .A1(n10693), .A2(n10694), .Z(n10695) );
  NAND2HSV0 U12756 ( .A1(\pe16/aot [7]), .A2(\pe16/bq[5] ), .ZN(n10697) );
  CLKNAND2HSV1 U12757 ( .A1(\pe16/pvq [5]), .A2(\pe16/ctrq ), .ZN(n10699) );
  XOR2HSV0 U12758 ( .A1(n10699), .A2(\pe16/phq [5]), .Z(n10700) );
  XOR2HSV0 U12759 ( .A1(n10701), .A2(n10700), .Z(n10702) );
  NOR2HSV1 U12760 ( .A1(n10706), .A2(n13229), .ZN(n10707) );
  MUX2HSV2 U12761 ( .I0(\pe16/ti_7t [5]), .I1(n15228), .S(n11220), .Z(n14835)
         );
  AOI21HSV2 U12762 ( .A1(n10709), .A2(n9358), .B(n10708), .ZN(n10710) );
  OAI21HSV2 U12763 ( .A1(n15070), .A2(n10711), .B(n10710), .ZN(n11265) );
  XNOR2HSV1 U12764 ( .A1(n11265), .A2(n11267), .ZN(n15292) );
  INHSV2 U12765 ( .I(n13102), .ZN(\pe2/ti_7[5] ) );
  CLKNAND2HSV1 U12766 ( .A1(n10713), .A2(n10712), .ZN(n14399) );
  NOR2HSV2 U12767 ( .A1(n10716), .A2(n14333), .ZN(n10717) );
  NAND2HSV2 U12768 ( .A1(n14949), .A2(\pe17/bq[4] ), .ZN(n10719) );
  NAND2HSV0 U12769 ( .A1(\pe17/got [4]), .A2(\pe17/ti_1 ), .ZN(n10718) );
  NAND2HSV2 U12770 ( .A1(\pe12/aot [8]), .A2(\pe12/bq[6] ), .ZN(n10723) );
  CLKNAND2HSV1 U12771 ( .A1(\pe12/got [6]), .A2(\pe12/ti_1 ), .ZN(n10726) );
  NAND2HSV0 U12772 ( .A1(\pe12/aot [6]), .A2(\pe12/bq[8] ), .ZN(n10725) );
  XOR2HSV0 U12773 ( .A1(n10726), .A2(n10725), .Z(n10727) );
  INHSV2 U12774 ( .I(ctro12), .ZN(n10728) );
  INHSV4 U12775 ( .I(n10728), .ZN(n14831) );
  CLKNAND2HSV0 U12776 ( .A1(n10729), .A2(n11447), .ZN(n10760) );
  CLKNAND2HSV1 U12777 ( .A1(n10760), .A2(\pe12/got [7]), .ZN(n10730) );
  INHSV2 U12778 ( .I(ctro12), .ZN(n11446) );
  INHSV1 U12779 ( .I(n11446), .ZN(n14246) );
  INHSV2 U12780 ( .I(\pe12/got [8]), .ZN(n11442) );
  NOR2HSV2 U12781 ( .A1(n11442), .A2(n14831), .ZN(n11469) );
  INHSV2 U12782 ( .I(n10731), .ZN(n10742) );
  INHSV2 U12783 ( .I(\pe12/phq [2]), .ZN(n10734) );
  OAI21HSV4 U12784 ( .A1(n10734), .A2(n10733), .B(n10732), .ZN(n10737) );
  INHSV2 U12785 ( .I(\pe12/bq[7] ), .ZN(n14577) );
  NOR2HSV2 U12786 ( .A1(n10735), .A2(n14577), .ZN(n10736) );
  XNOR2HSV4 U12787 ( .A1(n10737), .A2(n10736), .ZN(n10741) );
  CLKNAND2HSV1 U12788 ( .A1(\pe12/ti_1 ), .A2(\pe12/got [7]), .ZN(n10739) );
  XOR2HSV0 U12789 ( .A1(n10739), .A2(n10738), .Z(n10740) );
  XNOR2HSV4 U12790 ( .A1(n10741), .A2(n10740), .ZN(n10743) );
  AOI22HSV4 U12791 ( .A1(\pe12/ti_7t [2]), .A2(n14246), .B1(n10742), .B2(
        n10743), .ZN(n10764) );
  INHSV2 U12792 ( .I(n11448), .ZN(n11471) );
  INHSV4 U12793 ( .I(n10743), .ZN(n13849) );
  CLKNAND2HSV3 U12794 ( .A1(n10744), .A2(n13849), .ZN(n10765) );
  CLKNAND2HSV3 U12795 ( .A1(n10764), .A2(n10765), .ZN(n15192) );
  CLKNHSV0 U12796 ( .I(\pe12/ti_7t [3]), .ZN(n10745) );
  NAND2HSV0 U12797 ( .A1(n10745), .A2(n14831), .ZN(n10768) );
  CLKNAND2HSV1 U12798 ( .A1(n10768), .A2(\pe12/got [8]), .ZN(n10746) );
  CLKBUFHSV4 U12799 ( .I(\pe12/bq[8] ), .Z(n14507) );
  NAND2HSV2 U12800 ( .A1(n14507), .A2(\pe12/aot [5]), .ZN(n10749) );
  NAND2HSV0 U12801 ( .A1(\pe12/got [5]), .A2(\pe12/ti_1 ), .ZN(n10748) );
  NAND2HSV0 U12802 ( .A1(\pe12/aot [6]), .A2(\pe12/bq[7] ), .ZN(n10751) );
  XNOR2HSV1 U12803 ( .A1(n10751), .A2(n10750), .ZN(n10752) );
  XNOR2HSV1 U12804 ( .A1(n10753), .A2(n10752), .ZN(n10758) );
  NAND2HSV0 U12805 ( .A1(\pe12/bq[6] ), .A2(\pe12/aot [7]), .ZN(n10754) );
  XOR2HSV0 U12806 ( .A1(n10754), .A2(\pe12/phq [4]), .Z(n10756) );
  BUFHSV8 U12807 ( .I(\pe12/ctrq ), .Z(n14578) );
  CLKNAND2HSV1 U12808 ( .A1(n14578), .A2(\pe12/pvq [4]), .ZN(n10755) );
  XNOR2HSV1 U12809 ( .A1(n10756), .A2(n10755), .ZN(n10757) );
  XNOR2HSV1 U12810 ( .A1(n10758), .A2(n10757), .ZN(n10763) );
  INHSV2 U12811 ( .I(n10759), .ZN(n10761) );
  NAND3HSV2 U12812 ( .A1(n10761), .A2(\pe12/got [6]), .A3(n10760), .ZN(n10762)
         );
  NAND2HSV2 U12813 ( .A1(n14831), .A2(\pe12/ti_7t [4]), .ZN(n11415) );
  INHSV2 U12814 ( .I(n11415), .ZN(n11417) );
  CLKNAND2HSV3 U12815 ( .A1(n15192), .A2(\pe12/got [8]), .ZN(n11436) );
  CLKNHSV0 U12816 ( .I(n10768), .ZN(n11438) );
  INHSV2 U12817 ( .I(\pe12/got [7]), .ZN(n11414) );
  NOR2HSV2 U12818 ( .A1(n11438), .A2(n11414), .ZN(n10769) );
  NAND2HSV0 U12819 ( .A1(\pe12/got [4]), .A2(\pe12/ti_1 ), .ZN(n10771) );
  NAND2HSV0 U12820 ( .A1(\pe12/bq[5] ), .A2(\pe12/aot [7]), .ZN(n10770) );
  XOR2HSV0 U12821 ( .A1(n10771), .A2(n10770), .Z(n10773) );
  NAND2HSV0 U12822 ( .A1(\pe12/ctrq ), .A2(\pe12/pvq [5]), .ZN(n10772) );
  NAND2HSV0 U12823 ( .A1(\pe12/aot [8]), .A2(\pe12/bq[4] ), .ZN(n10775) );
  NAND2HSV0 U12824 ( .A1(\pe12/aot [6]), .A2(\pe12/bq[6] ), .ZN(n10774) );
  XOR2HSV0 U12825 ( .A1(n10775), .A2(n10774), .Z(n10779) );
  CLKNAND2HSV0 U12826 ( .A1(\pe12/aot [5]), .A2(\pe12/bq[7] ), .ZN(n10777) );
  NAND2HSV0 U12827 ( .A1(\pe12/aot [4]), .A2(\pe12/bq[8] ), .ZN(n10776) );
  XOR2HSV0 U12828 ( .A1(n10777), .A2(n10776), .Z(n10778) );
  XOR2HSV0 U12829 ( .A1(n10779), .A2(n10778), .Z(n10780) );
  CLKNHSV0 U12830 ( .I(\pe12/ti_7t [5]), .ZN(n10782) );
  NAND2HSV0 U12831 ( .A1(n11471), .A2(n10782), .ZN(n10783) );
  OAI21HSV4 U12832 ( .A1(n15249), .A2(n11471), .B(n10783), .ZN(n14237) );
  INHSV4 U12833 ( .I(n14237), .ZN(n14701) );
  NAND2HSV2 U12834 ( .A1(n10786), .A2(n10785), .ZN(n10788) );
  XNOR2HSV4 U12835 ( .A1(n10788), .A2(n10787), .ZN(n15200) );
  INHSV1 U12836 ( .I(n13057), .ZN(n14877) );
  CLKBUFHSV4 U12837 ( .I(n12907), .Z(n14935) );
  INHSV1 U12838 ( .I(ctro3), .ZN(n10789) );
  CLKNAND2HSV1 U12839 ( .A1(n10994), .A2(\pe3/ti_7t [3]), .ZN(n10971) );
  NAND2HSV2 U12840 ( .A1(n10972), .A2(n10971), .ZN(n14820) );
  INHSV2 U12841 ( .I(\pe15/ti_7t [3]), .ZN(n11292) );
  CLKBUFHSV4 U12842 ( .I(\pe15/got [8]), .Z(n15178) );
  INHSV2 U12843 ( .I(n10521), .ZN(n12320) );
  CLKNAND2HSV1 U12844 ( .A1(n12320), .A2(\pe15/ti_7t [1]), .ZN(n11316) );
  CLKNAND2HSV3 U12845 ( .A1(n10790), .A2(n11316), .ZN(n11387) );
  INHSV2 U12846 ( .I(\pe15/ctrq ), .ZN(n11844) );
  INHSV4 U12847 ( .I(n11844), .ZN(n13815) );
  NAND2HSV2 U12848 ( .A1(\pe15/pvq [3]), .A2(n13815), .ZN(n10791) );
  XNOR2HSV1 U12849 ( .A1(n10791), .A2(\pe15/phq [3]), .ZN(n10792) );
  XNOR2HSV4 U12850 ( .A1(n10793), .A2(n10792), .ZN(n11289) );
  XNOR2HSV4 U12851 ( .A1(n11290), .A2(n11289), .ZN(n11295) );
  CLKNAND2HSV3 U12852 ( .A1(n11977), .A2(n13142), .ZN(n14851) );
  INHSV2 U12853 ( .I(n11159), .ZN(n11160) );
  CLKNAND2HSV0 U12854 ( .A1(n11447), .A2(\pe12/ti_7t [3]), .ZN(n14247) );
  INHSV2 U12855 ( .I(n13034), .ZN(n14880) );
  BUFHSV2 U12856 ( .I(n11387), .Z(n15072) );
  INHSV2 U12857 ( .I(ctro8), .ZN(n12316) );
  CLKNHSV0 U12858 ( .I(n14755), .ZN(n12346) );
  CLKNHSV0 U12859 ( .I(n12346), .ZN(n14761) );
  CLKNHSV0 U12860 ( .I(n10978), .ZN(n11790) );
  MUX2HSV2 U12861 ( .I0(bo7[4]), .I1(\pe7/bq[4] ), .S(n12067), .Z(n15126) );
  INHSV2 U12862 ( .I(n10804), .ZN(n14844) );
  MUX2HSV2 U12863 ( .I0(bo3[1]), .I1(\pe3/bq[1] ), .S(n10805), .Z(n15101) );
  CLKBUFHSV2 U12864 ( .I(\pe16/aot [6]), .Z(n14932) );
  CLKBUFHSV4 U12865 ( .I(\pe8/aot [8]), .Z(n14950) );
  MUX2HSV1 U12866 ( .I0(bo9[3]), .I1(\pe9/bq[3] ), .S(n13826), .Z(n15137) );
  MUX2HSV1 U12867 ( .I0(bo9[5]), .I1(\pe9/bq[5] ), .S(n13826), .Z(n15136) );
  CLKNHSV0 U12868 ( .I(\pe2/aot [6]), .ZN(n10806) );
  INHSV2 U12869 ( .I(n10806), .ZN(n14741) );
  INHSV4 U12870 ( .I(n10807), .ZN(n15090) );
  INHSV2 U12871 ( .I(n14540), .ZN(n15092) );
  MUX2HSV1 U12872 ( .I0(bo9[6]), .I1(n11647), .S(n13826), .Z(n15135) );
  CLKBUFHSV4 U12873 ( .I(\pe12/aot [7]), .Z(n14948) );
  CLKBUFHSV2 U12874 ( .I(\pe14/aot [6]), .Z(n14889) );
  BUFHSV2 U12875 ( .I(\pe15/got [7]), .Z(n14864) );
  BUFHSV2 U12876 ( .I(\pe19/got [7]), .Z(n14841) );
  CLKNHSV0 U12877 ( .I(n11958), .ZN(n14721) );
  NAND3HSV0 U12878 ( .A1(n10809), .A2(n10810), .A3(n10841), .ZN(n10832) );
  CLKNHSV0 U12879 ( .I(n10832), .ZN(n10829) );
  CLKNAND2HSV0 U12880 ( .A1(n10841), .A2(n11780), .ZN(n10840) );
  CLKNAND2HSV0 U12881 ( .A1(n10840), .A2(\pe21/got [6]), .ZN(n10830) );
  NAND2HSV0 U12882 ( .A1(\pe21/ti_7[1] ), .A2(\pe21/got [4]), .ZN(n10824) );
  CLKNAND2HSV0 U12883 ( .A1(n15092), .A2(\pe21/pvq [6]), .ZN(n10816) );
  XNOR2HSV4 U12884 ( .A1(n10811), .A2(\pe21/phq [6]), .ZN(n10815) );
  NAND2HSV0 U12885 ( .A1(\pe21/bq[5] ), .A2(\pe21/aot [6]), .ZN(n10812) );
  XOR2HSV0 U12886 ( .A1(n10813), .A2(n10812), .Z(n10814) );
  XOR3HSV2 U12887 ( .A1(n10816), .A2(n10815), .A3(n10814), .Z(n10822) );
  NAND2HSV2 U12888 ( .A1(\pe21/bq[7] ), .A2(\pe21/aot [4]), .ZN(n10818) );
  XOR2HSV0 U12889 ( .A1(n10818), .A2(n10817), .Z(n10820) );
  XOR2HSV0 U12890 ( .A1(n10820), .A2(n10819), .Z(n10821) );
  XOR2HSV2 U12891 ( .A1(n10824), .A2(n10823), .Z(n10828) );
  CLKNHSV0 U12892 ( .I(n10830), .ZN(n10831) );
  CLKNAND2HSV0 U12893 ( .A1(n10832), .A2(n10831), .ZN(n10833) );
  NOR2HSV2 U12894 ( .A1(n10833), .A2(n8901), .ZN(n10834) );
  NOR2HSV1 U12895 ( .A1(n9398), .A2(\pe21/ti_7t [5]), .ZN(n10861) );
  NOR2HSV1 U12896 ( .A1(n10861), .A2(n10837), .ZN(n10838) );
  AND2HSV2 U12897 ( .A1(\pe21/bq[2] ), .A2(\pe21/aot [6]), .Z(n12092) );
  CLKNAND2HSV1 U12898 ( .A1(\pe21/bq[3] ), .A2(\pe21/aot [7]), .ZN(n12089) );
  NAND2HSV0 U12899 ( .A1(\pe21/bq[7] ), .A2(\pe21/aot [3]), .ZN(n10846) );
  NAND2HSV0 U12900 ( .A1(\pe21/bq[5] ), .A2(\pe21/aot [5]), .ZN(n10845) );
  XOR2HSV0 U12901 ( .A1(n10846), .A2(n10845), .Z(n10851) );
  NAND2HSV0 U12902 ( .A1(\pe21/bq[6] ), .A2(\pe21/aot [4]), .ZN(n10849) );
  CLKNHSV0 U12903 ( .I(\pe21/ti_1 ), .ZN(n10847) );
  INHSV2 U12904 ( .I(n10847), .ZN(n13834) );
  CLKNAND2HSV0 U12905 ( .A1(n13834), .A2(\pe21/got [2]), .ZN(n10848) );
  XOR2HSV0 U12906 ( .A1(n10849), .A2(n10848), .Z(n10850) );
  INHSV1 U12907 ( .I(n10854), .ZN(n10856) );
  AOI21HSV2 U12908 ( .A1(n10854), .A2(n10853), .B(n10852), .ZN(n10855) );
  OAI21HSV4 U12909 ( .A1(n6208), .A2(n10856), .B(n10855), .ZN(n10857) );
  INHSV2 U12910 ( .I(n10874), .ZN(n13801) );
  INHSV2 U12911 ( .I(n10862), .ZN(n13797) );
  NOR2HSV0 U12912 ( .A1(n13797), .A2(n10863), .ZN(n10864) );
  NAND2HSV0 U12913 ( .A1(\pe21/ti_7t [7]), .A2(n10865), .ZN(n10866) );
  INHSV3 U12914 ( .I(n10868), .ZN(n13338) );
  NAND2HSV2 U12915 ( .A1(\pe21/bq[1] ), .A2(\pe21/aot [2]), .ZN(n10871) );
  NAND2HSV0 U12916 ( .A1(\pe21/bq[2] ), .A2(\pe21/aot [1]), .ZN(n10870) );
  XOR2HSV0 U12917 ( .A1(n10871), .A2(n10870), .Z(n10872) );
  NAND2HSV2 U12918 ( .A1(n15085), .A2(\pe21/got [6]), .ZN(n10887) );
  NAND2HSV0 U12919 ( .A1(\pe21/bq[2] ), .A2(\pe21/aot [5]), .ZN(n10878) );
  NAND2HSV0 U12920 ( .A1(\pe21/bq[1] ), .A2(\pe21/aot [6]), .ZN(n10877) );
  XOR2HSV0 U12921 ( .A1(n10878), .A2(n10877), .Z(n10882) );
  NAND2HSV0 U12922 ( .A1(\pe21/bq[5] ), .A2(\pe21/aot [1]), .ZN(n12543) );
  NOR2HSV0 U12923 ( .A1(n12543), .A2(n12090), .ZN(n10880) );
  AOI22HSV0 U12924 ( .A1(\pe21/bq[6] ), .A2(\pe21/aot [1]), .B1(\pe21/bq[5] ), 
        .B2(\pe21/aot [2]), .ZN(n10879) );
  NOR2HSV1 U12925 ( .A1(n10880), .A2(n10879), .ZN(n10881) );
  NAND2HSV0 U12926 ( .A1(\pe21/bq[4] ), .A2(\pe21/aot [3]), .ZN(n10883) );
  XNOR2HSV4 U12927 ( .A1(n10885), .A2(n10884), .ZN(n10886) );
  XOR2HSV0 U12928 ( .A1(n10887), .A2(n10886), .Z(\pe21/poht [2]) );
  CLKNAND2HSV2 U12929 ( .A1(n7519), .A2(\pe21/got [3]), .ZN(n10889) );
  NAND2HSV2 U12930 ( .A1(n15085), .A2(\pe21/got [3]), .ZN(n10899) );
  CLKNAND2HSV2 U12931 ( .A1(n7519), .A2(\pe21/got [2]), .ZN(n10897) );
  NAND2HSV2 U12932 ( .A1(\pe21/got [1]), .A2(\pe21/ti_7[5] ), .ZN(n10895) );
  CLKNAND2HSV0 U12933 ( .A1(\pe21/bq[1] ), .A2(\pe21/aot [3]), .ZN(n10892) );
  NAND2HSV0 U12934 ( .A1(\pe21/bq[2] ), .A2(\pe21/aot [2]), .ZN(n10891) );
  XOR2HSV0 U12935 ( .A1(n10892), .A2(n10891), .Z(n10893) );
  CLKNAND2HSV1 U12936 ( .A1(\pe21/bq[3] ), .A2(\pe21/aot [1]), .ZN(n12547) );
  XNOR2HSV1 U12937 ( .A1(n10893), .A2(n12547), .ZN(n10894) );
  XOR2HSV0 U12938 ( .A1(n10899), .A2(n10898), .Z(\pe21/poht [5]) );
  NAND2HSV2 U12939 ( .A1(n8952), .A2(\pe10/got [8]), .ZN(n10933) );
  CLKNAND2HSV0 U12940 ( .A1(n14940), .A2(\pe10/got [3]), .ZN(n10901) );
  NAND2HSV0 U12941 ( .A1(n6033), .A2(\pe10/got [2]), .ZN(n10900) );
  XNOR2HSV1 U12942 ( .A1(n10901), .A2(n10900), .ZN(n10921) );
  CLKNHSV2 U12943 ( .I(\pe10/ctrq ), .ZN(n12187) );
  CLKNAND2HSV0 U12944 ( .A1(\pe10/pq ), .A2(n14554), .ZN(n10903) );
  NAND2HSV0 U12945 ( .A1(n14951), .A2(\pe10/bq[1] ), .ZN(n10902) );
  XOR2HSV0 U12946 ( .A1(n10903), .A2(n10902), .Z(n10907) );
  NAND2HSV0 U12947 ( .A1(\pe10/bq[5] ), .A2(\pe10/aot [4]), .ZN(n10905) );
  NAND2HSV0 U12948 ( .A1(\pe10/got [1]), .A2(\pe10/ti_1 ), .ZN(n10904) );
  XOR2HSV0 U12949 ( .A1(n10905), .A2(n10904), .Z(n10906) );
  XOR2HSV0 U12950 ( .A1(n10907), .A2(n10906), .Z(n10911) );
  BUFHSV2 U12951 ( .I(\pe10/bq[7] ), .Z(n14567) );
  NAND2HSV0 U12952 ( .A1(\pe10/aot [2]), .A2(n14567), .ZN(n10909) );
  NAND2HSV0 U12953 ( .A1(\pe10/aot [1]), .A2(n12272), .ZN(n10908) );
  XOR2HSV0 U12954 ( .A1(n10909), .A2(n10908), .Z(n10910) );
  XNOR2HSV1 U12955 ( .A1(n10911), .A2(n10910), .ZN(n10919) );
  NAND2HSV0 U12956 ( .A1(n14844), .A2(\pe10/bq[2] ), .ZN(n10913) );
  NAND2HSV0 U12957 ( .A1(n14133), .A2(\pe10/bq[3] ), .ZN(n10912) );
  XOR2HSV0 U12958 ( .A1(n10913), .A2(n10912), .Z(n10917) );
  NAND2HSV0 U12959 ( .A1(\pe10/aot [5]), .A2(\pe10/bq[4] ), .ZN(n10915) );
  NAND2HSV0 U12960 ( .A1(\pe10/aot [3]), .A2(\pe10/bq[6] ), .ZN(n10914) );
  XOR2HSV0 U12961 ( .A1(n10915), .A2(n10914), .Z(n10916) );
  XOR2HSV0 U12962 ( .A1(n10917), .A2(n10916), .Z(n10918) );
  XNOR2HSV1 U12963 ( .A1(n10919), .A2(n10918), .ZN(n10920) );
  XNOR2HSV1 U12964 ( .A1(n10921), .A2(n10920), .ZN(n10923) );
  NAND2HSV0 U12965 ( .A1(n14856), .A2(\pe10/got [4]), .ZN(n10922) );
  XOR2HSV0 U12966 ( .A1(n10923), .A2(n10922), .Z(n10929) );
  AOI21HSV4 U12967 ( .A1(n15200), .A2(n10925), .B(n14119), .ZN(n13476) );
  INHSV1 U12968 ( .I(\pe10/got [5]), .ZN(n13466) );
  NOR2HSV2 U12969 ( .A1(n13476), .A2(n13466), .ZN(n10928) );
  XOR3HSV2 U12970 ( .A1(n10929), .A2(n10928), .A3(n10927), .Z(n10932) );
  NOR2HSV0 U12971 ( .A1(n10930), .A2(n10040), .ZN(n13467) );
  NOR3HSV2 U12972 ( .A1(n13468), .A2(n13467), .A3(n15140), .ZN(n10931) );
  XOR2HSV0 U12973 ( .A1(n10932), .A2(n10931), .Z(n10934) );
  CLKNAND2HSV1 U12974 ( .A1(n10933), .A2(n10934), .ZN(n10938) );
  CLKNHSV0 U12975 ( .I(n10934), .ZN(n10935) );
  CLKNAND2HSV1 U12976 ( .A1(n10938), .A2(n10937), .ZN(po10) );
  INHSV2 U12977 ( .I(n10945), .ZN(n11773) );
  CLKNAND2HSV0 U12978 ( .A1(n10946), .A2(\pe3/got [6]), .ZN(n10947) );
  NOR2HSV2 U12979 ( .A1(n10948), .A2(n10947), .ZN(n10963) );
  NAND2HSV0 U12980 ( .A1(\pe3/ti_7[1] ), .A2(\pe3/got [4]), .ZN(n10962) );
  NAND2HSV0 U12981 ( .A1(\pe3/aot [7]), .A2(\pe3/bq[4] ), .ZN(n10950) );
  NAND2HSV0 U12982 ( .A1(\pe3/bq[5] ), .A2(\pe3/aot [6]), .ZN(n10949) );
  XOR2HSV0 U12983 ( .A1(n10950), .A2(n10949), .Z(n10961) );
  NAND2HSV0 U12984 ( .A1(\pe3/aot [5]), .A2(\pe3/bq[6] ), .ZN(n10951) );
  CLKNAND2HSV1 U12985 ( .A1(n12476), .A2(\pe3/aot [3]), .ZN(n10954) );
  NAND2HSV0 U12986 ( .A1(\pe3/aot [4]), .A2(\pe3/bq[7] ), .ZN(n10953) );
  XOR2HSV0 U12987 ( .A1(n10954), .A2(n10953), .Z(n10958) );
  CLKNAND2HSV0 U12988 ( .A1(n14953), .A2(\pe3/bq[3] ), .ZN(n10956) );
  CLKNAND2HSV1 U12989 ( .A1(n12475), .A2(\pe3/got [3]), .ZN(n10955) );
  XOR2HSV0 U12990 ( .A1(n10956), .A2(n10955), .Z(n10957) );
  XOR2HSV0 U12991 ( .A1(n10958), .A2(n10957), .Z(n10959) );
  XNOR2HSV4 U12992 ( .A1(n10968), .A2(n10967), .ZN(n10964) );
  MUX2NHSV4 U12993 ( .I0(n10966), .I1(n10965), .S(n10964), .ZN(n10999) );
  CLKNHSV1 U12994 ( .I(n11707), .ZN(n10970) );
  CLKAND2HSV2 U12995 ( .A1(n10994), .A2(\pe3/ti_7t [6]), .Z(n10969) );
  AOI21HSV4 U12996 ( .A1(n11709), .A2(n10970), .B(n10969), .ZN(n10998) );
  NOR2HSV2 U12997 ( .A1(n10994), .A2(n15180), .ZN(n12501) );
  NAND2HSV0 U12998 ( .A1(n5949), .A2(\pe3/got [3]), .ZN(n10973) );
  NAND2HSV0 U12999 ( .A1(\pe3/aot [4]), .A2(\pe3/bq[6] ), .ZN(n10975) );
  CLKNAND2HSV0 U13000 ( .A1(n14953), .A2(\pe3/bq[2] ), .ZN(n10974) );
  XOR2HSV0 U13001 ( .A1(n10975), .A2(n10974), .Z(n10990) );
  NAND2HSV0 U13002 ( .A1(\pe3/bq[4] ), .A2(\pe3/aot [6]), .ZN(n10977) );
  NAND2HSV0 U13003 ( .A1(\pe3/got [2]), .A2(n12475), .ZN(n10976) );
  XOR2HSV0 U13004 ( .A1(n10977), .A2(n10976), .Z(n10981) );
  CLKNHSV0 U13005 ( .I(n10978), .ZN(n10979) );
  XNOR2HSV1 U13006 ( .A1(n10981), .A2(n10980), .ZN(n10989) );
  NAND2HSV0 U13007 ( .A1(\pe3/aot [5]), .A2(\pe3/bq[5] ), .ZN(n10983) );
  NAND2HSV0 U13008 ( .A1(\pe3/aot [2]), .A2(n12476), .ZN(n10982) );
  XOR2HSV0 U13009 ( .A1(n10983), .A2(n10982), .Z(n10987) );
  NAND2HSV0 U13010 ( .A1(\pe3/aot [7]), .A2(\pe3/bq[3] ), .ZN(n10985) );
  NAND2HSV0 U13011 ( .A1(\pe3/aot [3]), .A2(\pe3/bq[7] ), .ZN(n10984) );
  XOR2HSV0 U13012 ( .A1(n10985), .A2(n10984), .Z(n10986) );
  XOR2HSV0 U13013 ( .A1(n10987), .A2(n10986), .Z(n10988) );
  XOR3HSV2 U13014 ( .A1(n10990), .A2(n10989), .A3(n10988), .Z(n10991) );
  CLKNAND2HSV0 U13015 ( .A1(n11006), .A2(n14931), .ZN(n10996) );
  CLKNAND2HSV3 U13016 ( .A1(n10999), .A2(n10998), .ZN(n12981) );
  AOI22HSV4 U13017 ( .A1(n10994), .A2(\pe3/ti_7t [7]), .B1(n13888), .B2(n11000), .ZN(n12502) );
  NAND2HSV4 U13018 ( .A1(n12503), .A2(n12502), .ZN(n14819) );
  NAND2HSV2 U13019 ( .A1(\pe3/got [6]), .A2(n14819), .ZN(n11035) );
  CLKNAND2HSV1 U13020 ( .A1(n11005), .A2(n11001), .ZN(n11016) );
  NAND2HSV0 U13021 ( .A1(n11003), .A2(n10789), .ZN(n11004) );
  NOR2HSV2 U13022 ( .A1(n11005), .A2(n11004), .ZN(n11014) );
  CLKNHSV0 U13023 ( .I(n11006), .ZN(n11008) );
  CLKNHSV0 U13024 ( .I(\pe3/got [4]), .ZN(n11007) );
  NOR2HSV2 U13025 ( .A1(n11008), .A2(n11007), .ZN(n11011) );
  CLKNAND2HSV0 U13026 ( .A1(n11017), .A2(n11011), .ZN(n11009) );
  NOR2HSV1 U13027 ( .A1(n11014), .A2(n11009), .ZN(n11010) );
  INHSV1 U13028 ( .I(n11011), .ZN(n11013) );
  INHSV2 U13029 ( .I(n11017), .ZN(n11012) );
  OAI21HSV2 U13030 ( .A1(n11014), .A2(n11013), .B(n11012), .ZN(n11015) );
  NAND2HSV0 U13031 ( .A1(n14820), .A2(\pe3/got [2]), .ZN(n11031) );
  NAND2HSV0 U13032 ( .A1(\pe3/got [1]), .A2(n14872), .ZN(n11029) );
  NAND2HSV0 U13033 ( .A1(\pe3/aot [3]), .A2(\pe3/bq[4] ), .ZN(n11019) );
  NAND2HSV0 U13034 ( .A1(\pe3/aot [1]), .A2(n6723), .ZN(n11018) );
  XOR2HSV0 U13035 ( .A1(n11019), .A2(n11018), .Z(n11023) );
  NAND2HSV0 U13036 ( .A1(\pe3/aot [4]), .A2(\pe3/bq[3] ), .ZN(n11021) );
  NAND2HSV0 U13037 ( .A1(\pe3/aot [2]), .A2(\pe3/bq[5] ), .ZN(n11020) );
  XOR2HSV0 U13038 ( .A1(n11021), .A2(n11020), .Z(n11022) );
  XOR2HSV0 U13039 ( .A1(n11023), .A2(n11022), .Z(n11027) );
  NAND2HSV0 U13040 ( .A1(\pe3/bq[1] ), .A2(\pe3/aot [6]), .ZN(n11025) );
  NAND2HSV0 U13041 ( .A1(\pe3/aot [5]), .A2(\pe3/bq[2] ), .ZN(n11024) );
  XOR2HSV0 U13042 ( .A1(n11025), .A2(n11024), .Z(n11026) );
  XNOR2HSV1 U13043 ( .A1(n11027), .A2(n11026), .ZN(n11028) );
  XOR2HSV0 U13044 ( .A1(n11029), .A2(n11028), .Z(n11030) );
  XOR2HSV0 U13045 ( .A1(n11031), .A2(n11030), .Z(n11032) );
  NAND2HSV0 U13046 ( .A1(\pe3/got [5]), .A2(n12957), .ZN(n11033) );
  XOR2HSV0 U13047 ( .A1(n11034), .A2(n11035), .Z(\pe3/poht [2]) );
  INHSV2 U13048 ( .I(\pe14/got [4]), .ZN(n11144) );
  CLKNAND2HSV2 U13049 ( .A1(n11081), .A2(\pe14/got [8]), .ZN(n11062) );
  XNOR2HSV4 U13050 ( .A1(n6729), .A2(n11037), .ZN(n11064) );
  INHSV2 U13051 ( .I(\pe14/got [3]), .ZN(n14488) );
  NOR2HSV0 U13052 ( .A1(n11110), .A2(n14488), .ZN(n11058) );
  CLKNAND2HSV0 U13053 ( .A1(\pe14/aot [4]), .A2(\pe14/bq[6] ), .ZN(n11149) );
  NAND2HSV0 U13054 ( .A1(\pe14/aot [3]), .A2(\pe14/bq[7] ), .ZN(n11040) );
  XOR2HSV0 U13055 ( .A1(n11149), .A2(n11040), .Z(n11055) );
  CLKNHSV0 U13056 ( .I(\pe14/ctrq ), .ZN(n13067) );
  INHSV2 U13057 ( .I(n13067), .ZN(n14742) );
  NAND2HSV2 U13058 ( .A1(n14742), .A2(\pe14/pvq [7]), .ZN(n11041) );
  XNOR2HSV1 U13059 ( .A1(n11041), .A2(\pe14/phq [7]), .ZN(n11046) );
  CLKNAND2HSV0 U13060 ( .A1(\pe14/aot [2]), .A2(\pe14/bq[4] ), .ZN(n14492) );
  BUFHSV4 U13061 ( .I(\pe14/bq[8] ), .Z(n14505) );
  AOI22HSV0 U13062 ( .A1(n14505), .A2(\pe14/aot [2]), .B1(\pe14/aot [6]), .B2(
        \pe14/bq[4] ), .ZN(n11043) );
  NOR2HSV1 U13063 ( .A1(n11044), .A2(n11043), .ZN(n11045) );
  XNOR2HSV1 U13064 ( .A1(n11046), .A2(n11045), .ZN(n11054) );
  NAND2HSV0 U13065 ( .A1(n5968), .A2(\pe14/got [2]), .ZN(n11048) );
  NAND2HSV0 U13066 ( .A1(\pe14/bq[3] ), .A2(\pe14/aot [7]), .ZN(n11047) );
  XOR2HSV0 U13067 ( .A1(n11048), .A2(n11047), .Z(n11052) );
  CLKNAND2HSV0 U13068 ( .A1(n14891), .A2(\pe14/bq[2] ), .ZN(n11050) );
  NAND2HSV0 U13069 ( .A1(\pe14/bq[5] ), .A2(\pe14/aot [5]), .ZN(n11049) );
  XOR2HSV0 U13070 ( .A1(n11050), .A2(n11049), .Z(n11051) );
  XOR2HSV0 U13071 ( .A1(n11052), .A2(n11051), .Z(n11053) );
  XOR3HSV2 U13072 ( .A1(n11055), .A2(n11054), .A3(n11053), .Z(n11057) );
  CLKNAND2HSV1 U13073 ( .A1(n14944), .A2(\pe14/got [4]), .ZN(n11056) );
  INHSV2 U13074 ( .I(n11059), .ZN(n11095) );
  NOR2HSV2 U13075 ( .A1(n11095), .A2(n13580), .ZN(n11060) );
  NAND2HSV2 U13076 ( .A1(n11061), .A2(n11060), .ZN(n11087) );
  CLKNHSV0 U13077 ( .I(n11062), .ZN(n11063) );
  NOR2HSV3 U13078 ( .A1(n11065), .A2(n11064), .ZN(n11088) );
  NOR2HSV2 U13079 ( .A1(n11087), .A2(n11088), .ZN(n11084) );
  CLKNAND2HSV0 U13080 ( .A1(\pe14/aot [6]), .A2(\pe14/bq[6] ), .ZN(n11067) );
  NAND2HSV0 U13081 ( .A1(\pe14/aot [5]), .A2(\pe14/bq[7] ), .ZN(n11066) );
  XOR2HSV0 U13082 ( .A1(n11067), .A2(n11066), .Z(n11071) );
  NAND2HSV0 U13083 ( .A1(\pe14/aot [8]), .A2(\pe14/bq[4] ), .ZN(n11069) );
  NAND2HSV0 U13084 ( .A1(\pe14/got [4]), .A2(\pe14/ti_1 ), .ZN(n11068) );
  XOR2HSV0 U13085 ( .A1(n11069), .A2(n11068), .Z(n11070) );
  XNOR2HSV1 U13086 ( .A1(n11071), .A2(n11070), .ZN(n11078) );
  NAND2HSV2 U13087 ( .A1(n14516), .A2(\pe14/pvq [5]), .ZN(n11072) );
  XNOR2HSV4 U13088 ( .A1(n11072), .A2(\pe14/phq [5]), .ZN(n11076) );
  NAND2HSV0 U13089 ( .A1(\pe14/bq[5] ), .A2(\pe14/aot [7]), .ZN(n11074) );
  NAND2HSV0 U13090 ( .A1(\pe14/aot [4]), .A2(\pe14/bq[8] ), .ZN(n11073) );
  XOR2HSV0 U13091 ( .A1(n11074), .A2(n11073), .Z(n11075) );
  XNOR2HSV4 U13092 ( .A1(n11076), .A2(n11075), .ZN(n11077) );
  INHSV2 U13093 ( .I(\pe14/got [5]), .ZN(n13552) );
  NOR2HSV2 U13094 ( .A1(n11110), .A2(n13552), .ZN(n11079) );
  XNOR2HSV1 U13095 ( .A1(n11080), .A2(n11079), .ZN(n11083) );
  AND2HSV2 U13096 ( .A1(n11081), .A2(\pe14/got [6]), .Z(n11082) );
  XNOR2HSV4 U13097 ( .A1(n11083), .A2(n11082), .ZN(n11085) );
  INHSV2 U13098 ( .I(\pe14/got [8]), .ZN(n11089) );
  NOR2HSV1 U13099 ( .A1(n8948), .A2(\pe14/ti_7t [5]), .ZN(n11114) );
  CLKNHSV0 U13100 ( .I(n11114), .ZN(n11092) );
  NOR2HSV4 U13101 ( .A1(n11094), .A2(n11093), .ZN(n11117) );
  CLKNAND2HSV2 U13102 ( .A1(n14516), .A2(\pe14/pvq [6]), .ZN(n11096) );
  XOR3HSV2 U13103 ( .A1(\pe14/phq [6]), .A2(n11097), .A3(n11096), .Z(n11101)
         );
  CLKNAND2HSV1 U13104 ( .A1(n14891), .A2(\pe14/bq[3] ), .ZN(n11099) );
  NAND2HSV0 U13105 ( .A1(\pe14/bq[4] ), .A2(\pe14/aot [7]), .ZN(n11098) );
  XOR2HSV0 U13106 ( .A1(n11099), .A2(n11098), .Z(n11100) );
  XOR2HSV2 U13107 ( .A1(n11101), .A2(n11100), .Z(n11109) );
  CLKNAND2HSV0 U13108 ( .A1(\pe14/aot [6]), .A2(\pe14/bq[5] ), .ZN(n11103) );
  NAND2HSV0 U13109 ( .A1(\pe14/got [3]), .A2(n5968), .ZN(n11102) );
  XOR2HSV0 U13110 ( .A1(n11103), .A2(n11102), .Z(n11107) );
  NAND2HSV0 U13111 ( .A1(\pe14/aot [4]), .A2(\pe14/bq[7] ), .ZN(n11104) );
  XNOR2HSV4 U13112 ( .A1(n11105), .A2(n11104), .ZN(n11106) );
  XNOR2HSV4 U13113 ( .A1(n11107), .A2(n11106), .ZN(n11108) );
  XNOR2HSV4 U13114 ( .A1(n11109), .A2(n11108), .ZN(n11112) );
  BUFHSV4 U13115 ( .I(n11110), .Z(n13853) );
  NOR2HSV4 U13116 ( .A1(n13853), .A2(n11144), .ZN(n11111) );
  NAND2HSV2 U13117 ( .A1(n14702), .A2(\pe14/ti_7t [7]), .ZN(n13582) );
  XNOR2HSV4 U13118 ( .A1(n11122), .A2(n11121), .ZN(n15236) );
  CLKAND2HSV2 U13119 ( .A1(n14702), .A2(\pe14/ti_7t [5]), .Z(n11123) );
  AOI21HSV4 U13120 ( .A1(n15236), .A2(n8948), .B(n11123), .ZN(n14489) );
  CLKNHSV0 U13121 ( .I(\pe14/got [2]), .ZN(n11124) );
  NOR2HSV2 U13122 ( .A1(n14489), .A2(n11124), .ZN(n11134) );
  NAND2HSV0 U13123 ( .A1(\pe14/got [1]), .A2(n15195), .ZN(n11132) );
  NAND2HSV0 U13124 ( .A1(\pe14/aot [4]), .A2(\pe14/bq[1] ), .ZN(n11126) );
  NAND2HSV0 U13125 ( .A1(\pe14/aot [3]), .A2(\pe14/bq[2] ), .ZN(n11125) );
  XOR2HSV0 U13126 ( .A1(n11126), .A2(n11125), .Z(n11130) );
  NAND2HSV0 U13127 ( .A1(\pe14/aot [1]), .A2(\pe14/bq[4] ), .ZN(n11128) );
  NAND2HSV0 U13128 ( .A1(\pe14/aot [2]), .A2(\pe14/bq[3] ), .ZN(n11127) );
  XOR2HSV0 U13129 ( .A1(n11128), .A2(n11127), .Z(n11129) );
  XOR2HSV0 U13130 ( .A1(n11130), .A2(n11129), .Z(n11131) );
  XOR2HSV0 U13131 ( .A1(n11132), .A2(n11131), .Z(n11133) );
  XOR2HSV2 U13132 ( .A1(n11134), .A2(n11133), .Z(n11138) );
  CLKNHSV0 U13133 ( .I(n11226), .ZN(n11136) );
  AOI21HSV0 U13134 ( .A1(n11226), .A2(n14702), .B(n14488), .ZN(n11135) );
  NAND2HSV2 U13135 ( .A1(n11138), .A2(n11137), .ZN(n11142) );
  INHSV1 U13136 ( .I(n11138), .ZN(n11140) );
  NAND2HSV2 U13137 ( .A1(n11140), .A2(n11139), .ZN(n11141) );
  CLKNAND2HSV2 U13138 ( .A1(n11142), .A2(n11141), .ZN(n11143) );
  NAND2HSV0 U13139 ( .A1(\pe14/aot [2]), .A2(\pe14/bq[5] ), .ZN(n11146) );
  NAND2HSV0 U13140 ( .A1(\pe14/aot [3]), .A2(\pe14/bq[4] ), .ZN(n11145) );
  XOR2HSV0 U13141 ( .A1(n11146), .A2(n11145), .Z(n11151) );
  CLKNAND2HSV1 U13142 ( .A1(\pe14/bq[3] ), .A2(\pe14/aot [1]), .ZN(n11276) );
  CLKNHSV0 U13143 ( .I(\pe14/aot [4]), .ZN(n11147) );
  BUFHSV2 U13144 ( .I(\pe14/bq[6] ), .Z(n14518) );
  NAND2HSV0 U13145 ( .A1(\pe14/aot [1]), .A2(n14518), .ZN(n13554) );
  OAI21HSV0 U13146 ( .A1(n13560), .A2(n11147), .B(n13554), .ZN(n11148) );
  OAI21HSV0 U13147 ( .A1(n11276), .A2(n11149), .B(n11148), .ZN(n11150) );
  XNOR2HSV1 U13148 ( .A1(n11151), .A2(n11150), .ZN(n11155) );
  NAND2HSV0 U13149 ( .A1(n14889), .A2(\pe14/bq[1] ), .ZN(n11153) );
  NAND2HSV0 U13150 ( .A1(\pe14/bq[2] ), .A2(\pe14/aot [5]), .ZN(n11152) );
  XOR2HSV0 U13151 ( .A1(n11153), .A2(n11152), .Z(n11154) );
  CLKNAND2HSV0 U13152 ( .A1(n11160), .A2(n8957), .ZN(n11200) );
  CLKNHSV0 U13153 ( .I(\pe16/ti_7[1] ), .ZN(n11161) );
  INHSV4 U13154 ( .I(\pe16/got [3]), .ZN(n14096) );
  CLKNAND2HSV0 U13155 ( .A1(\pe16/aot [3]), .A2(n6004), .ZN(n13211) );
  CLKNHSV0 U13156 ( .I(\pe16/aot [2]), .ZN(n14271) );
  NAND2HSV2 U13157 ( .A1(\pe16/aot [2]), .A2(n5947), .ZN(n14273) );
  NAND2HSV0 U13158 ( .A1(\pe16/bq[6] ), .A2(\pe16/aot [4]), .ZN(n11163) );
  NAND2HSV0 U13159 ( .A1(\pe16/aot [7]), .A2(\pe16/bq[3] ), .ZN(n11162) );
  CLKNAND2HSV0 U13160 ( .A1(\pe16/aot [8]), .A2(\pe16/bq[2] ), .ZN(n11166) );
  NAND2HSV0 U13161 ( .A1(\pe16/aot [6]), .A2(\pe16/bq[4] ), .ZN(n11165) );
  NAND2HSV0 U13162 ( .A1(\pe16/aot [5]), .A2(\pe16/bq[5] ), .ZN(n11168) );
  NAND2HSV0 U13163 ( .A1(\pe16/got [2]), .A2(n14266), .ZN(n11167) );
  XOR2HSV2 U13164 ( .A1(n11170), .A2(n11169), .Z(n11171) );
  NOR2HSV0 U13165 ( .A1(n12194), .A2(n8957), .ZN(n11173) );
  CLKNAND2HSV0 U13166 ( .A1(n11182), .A2(n14873), .ZN(n11172) );
  INHSV2 U13167 ( .I(n11180), .ZN(n11176) );
  NAND2HSV2 U13168 ( .A1(n11182), .A2(n11179), .ZN(n13868) );
  NOR2HSV1 U13169 ( .A1(n13868), .A2(n8957), .ZN(n11183) );
  NOR2HSV2 U13170 ( .A1(n14096), .A2(n13833), .ZN(n11184) );
  XOR3HSV2 U13171 ( .A1(\pe16/phq [6]), .A2(n11185), .A3(n11184), .Z(n11189)
         );
  NAND2HSV0 U13172 ( .A1(\pe16/aot [5]), .A2(\pe16/bq[6] ), .ZN(n11186) );
  XNOR2HSV4 U13173 ( .A1(n11189), .A2(n11188), .ZN(n11197) );
  CLKNAND2HSV1 U13174 ( .A1(\pe16/aot [6]), .A2(\pe16/bq[5] ), .ZN(n11191) );
  NAND2HSV0 U13175 ( .A1(\pe16/aot [4]), .A2(\pe16/bq[7] ), .ZN(n11190) );
  XOR2HSV0 U13176 ( .A1(n11191), .A2(n11190), .Z(n11195) );
  NAND2HSV0 U13177 ( .A1(\pe16/aot [3]), .A2(\pe16/bq[8] ), .ZN(n11193) );
  NAND2HSV0 U13178 ( .A1(\pe16/aot [8]), .A2(\pe16/bq[3] ), .ZN(n11192) );
  XOR2HSV0 U13179 ( .A1(n11193), .A2(n11192), .Z(n11194) );
  XOR2HSV2 U13180 ( .A1(n11195), .A2(n11194), .Z(n11196) );
  XNOR2HSV4 U13181 ( .A1(n11197), .A2(n11196), .ZN(n11199) );
  NAND2HSV2 U13182 ( .A1(\pe16/ti_7[1] ), .A2(\pe16/got [4]), .ZN(n11198) );
  CLKNAND2HSV1 U13183 ( .A1(n11200), .A2(\pe16/got [6]), .ZN(n11202) );
  INHSV1 U13184 ( .I(n11202), .ZN(n11201) );
  NAND2HSV0 U13185 ( .A1(n11205), .A2(n11207), .ZN(n11206) );
  OAI21HSV1 U13186 ( .A1(n11207), .A2(\pe16/ti_7t [4]), .B(n14292), .ZN(n11208) );
  AOI21HSV0 U13187 ( .A1(n11211), .A2(n15185), .B(n13868), .ZN(n11212) );
  NAND2HSV2 U13188 ( .A1(n11212), .A2(n13870), .ZN(n11213) );
  INHSV2 U13189 ( .I(\pe16/ti_7t [7]), .ZN(n14071) );
  NAND2HSV2 U13190 ( .A1(n8956), .A2(n14071), .ZN(n13188) );
  NOR2HSV2 U13191 ( .A1(n14364), .A2(n14096), .ZN(n11225) );
  CLKNAND2HSV0 U13192 ( .A1(\pe16/aot [2]), .A2(\pe16/bq[2] ), .ZN(n11217) );
  NAND2HSV0 U13193 ( .A1(\pe16/aot [1]), .A2(\pe16/bq[3] ), .ZN(n11216) );
  XOR2HSV0 U13194 ( .A1(n11217), .A2(n11216), .Z(n11219) );
  NAND2HSV0 U13195 ( .A1(\pe16/aot [3]), .A2(\pe16/bq[1] ), .ZN(n11218) );
  XNOR2HSV1 U13196 ( .A1(n11219), .A2(n11218), .ZN(n11223) );
  INHSV4 U13197 ( .I(n15186), .ZN(n13190) );
  CLKNAND2HSV1 U13198 ( .A1(n14293), .A2(\pe16/got [1]), .ZN(n11221) );
  XOR3HSV2 U13199 ( .A1(n11223), .A2(n11221), .A3(n11222), .Z(n11224) );
  XOR2HSV0 U13200 ( .A1(n11225), .A2(n11224), .Z(\pe16/poht [5]) );
  NAND2HSV4 U13201 ( .A1(n11227), .A2(n11226), .ZN(n14855) );
  NAND2HSV2 U13202 ( .A1(n14855), .A2(\pe14/got [1]), .ZN(n11231) );
  CLKNAND2HSV1 U13203 ( .A1(\pe14/aot [1]), .A2(\pe14/bq[2] ), .ZN(n11229) );
  NAND2HSV0 U13204 ( .A1(\pe14/aot [2]), .A2(\pe14/bq[1] ), .ZN(n11228) );
  XOR2HSV0 U13205 ( .A1(n11229), .A2(n11228), .Z(n11230) );
  CLKXOR2HSV2 U13206 ( .A1(n11231), .A2(n11230), .Z(n11233) );
  XOR2HSV0 U13207 ( .A1(n11233), .A2(n11232), .Z(\pe14/poht [6]) );
  NAND2HSV0 U13208 ( .A1(\pe2/aot [3]), .A2(\pe2/bq[1] ), .ZN(n11235) );
  NAND2HSV0 U13209 ( .A1(\pe2/aot [2]), .A2(\pe2/bq[2] ), .ZN(n11234) );
  XOR2HSV0 U13210 ( .A1(n11235), .A2(n11234), .Z(n11236) );
  CLKNAND2HSV1 U13211 ( .A1(\pe2/aot [1]), .A2(\pe2/bq[3] ), .ZN(n13092) );
  XNOR2HSV1 U13212 ( .A1(n11236), .A2(n13092), .ZN(n11241) );
  CLKNAND2HSV0 U13213 ( .A1(\pe2/ti_7[5] ), .A2(\pe2/got [1]), .ZN(n11239) );
  XOR3HSV2 U13214 ( .A1(n11241), .A2(n11240), .A3(n11239), .Z(n11273) );
  NAND2HSV2 U13215 ( .A1(n12907), .A2(n14822), .ZN(n11260) );
  INHSV2 U13216 ( .I(\pe2/got [5]), .ZN(n12878) );
  NAND2HSV0 U13217 ( .A1(\pe2/ti_7[1] ), .A2(\pe2/got [3]), .ZN(n11243) );
  BUFHSV2 U13218 ( .I(\pe2/bq[6] ), .Z(n14510) );
  CLKNAND2HSV1 U13219 ( .A1(n14510), .A2(\pe2/aot [4]), .ZN(n12508) );
  BUFHSV4 U13220 ( .I(\pe2/bq[7] ), .Z(n14504) );
  CLKNAND2HSV0 U13221 ( .A1(\pe2/aot [3]), .A2(n14504), .ZN(n11244) );
  XOR2HSV0 U13222 ( .A1(n12508), .A2(n11244), .Z(n11257) );
  NAND2HSV0 U13223 ( .A1(\pe2/got [2]), .A2(n13831), .ZN(n11246) );
  NAND2HSV0 U13224 ( .A1(n14858), .A2(\pe2/bq[2] ), .ZN(n11245) );
  XOR2HSV0 U13225 ( .A1(n11246), .A2(n11245), .Z(n11248) );
  INHSV1 U13226 ( .I(n13766), .ZN(n14558) );
  XNOR2HSV1 U13227 ( .A1(n11248), .A2(n11247), .ZN(n11256) );
  NAND2HSV0 U13228 ( .A1(\pe2/aot [7]), .A2(\pe2/bq[3] ), .ZN(n11250) );
  NAND2HSV0 U13229 ( .A1(\pe2/bq[4] ), .A2(\pe2/aot [6]), .ZN(n11249) );
  XOR2HSV0 U13230 ( .A1(n11250), .A2(n11249), .Z(n11254) );
  NAND2HSV0 U13231 ( .A1(\pe2/aot [5]), .A2(\pe2/bq[5] ), .ZN(n11252) );
  NAND2HSV0 U13232 ( .A1(\pe2/aot [2]), .A2(n14559), .ZN(n11251) );
  XOR2HSV0 U13233 ( .A1(n11252), .A2(n11251), .Z(n11253) );
  XOR2HSV0 U13234 ( .A1(n11254), .A2(n11253), .Z(n11255) );
  XOR3HSV2 U13235 ( .A1(n11257), .A2(n11256), .A3(n11255), .Z(n11258) );
  CLKNHSV0 U13236 ( .I(n11261), .ZN(n11262) );
  CLKNAND2HSV0 U13237 ( .A1(n11262), .A2(\pe2/got [7]), .ZN(n11263) );
  AOI21HSV2 U13238 ( .A1(n11265), .A2(n11264), .B(n11263), .ZN(n11271) );
  INHSV2 U13239 ( .I(n11265), .ZN(n11269) );
  CLKNAND2HSV1 U13240 ( .A1(n11269), .A2(n11268), .ZN(n11270) );
  NAND2HSV2 U13241 ( .A1(n14957), .A2(\pe2/got [3]), .ZN(n11272) );
  CLKNHSV1 U13242 ( .I(\pe14/got [1]), .ZN(n13567) );
  NOR2HSV2 U13243 ( .A1(n14489), .A2(n13567), .ZN(n11279) );
  CLKNAND2HSV0 U13244 ( .A1(\pe14/aot [3]), .A2(\pe14/bq[1] ), .ZN(n11275) );
  NAND2HSV0 U13245 ( .A1(\pe14/aot [2]), .A2(\pe14/bq[2] ), .ZN(n11274) );
  XOR2HSV0 U13246 ( .A1(n11275), .A2(n11274), .Z(n11277) );
  XNOR2HSV1 U13247 ( .A1(n11277), .A2(n11276), .ZN(n11278) );
  NAND2HSV2 U13248 ( .A1(n13086), .A2(\pe14/got [2]), .ZN(n11280) );
  XOR2HSV2 U13249 ( .A1(n11281), .A2(n11280), .Z(n11283) );
  XOR2HSV0 U13250 ( .A1(n11283), .A2(n11282), .Z(\pe14/poht [5]) );
  NAND2HSV0 U13251 ( .A1(\pe4/aot [4]), .A2(\pe4/bq[1] ), .ZN(n11286) );
  NAND2HSV0 U13252 ( .A1(\pe4/aot [3]), .A2(\pe4/bq[2] ), .ZN(n11285) );
  NAND2HSV0 U13253 ( .A1(\pe4/aot [1]), .A2(\pe4/bq[4] ), .ZN(n11288) );
  NAND2HSV0 U13254 ( .A1(\pe4/aot [2]), .A2(\pe4/bq[3] ), .ZN(n11287) );
  INHSV2 U13255 ( .I(n11291), .ZN(n11294) );
  NAND2HSV2 U13256 ( .A1(n11292), .A2(n14704), .ZN(n11369) );
  NAND2HSV2 U13257 ( .A1(n11369), .A2(n15178), .ZN(n11293) );
  AOI21HSV4 U13258 ( .A1(n11340), .A2(n11294), .B(n11293), .ZN(n11334) );
  INHSV2 U13259 ( .I(n11295), .ZN(n11299) );
  CLKNHSV0 U13260 ( .I(n11323), .ZN(n11297) );
  INHSV2 U13261 ( .I(n11342), .ZN(n11298) );
  NAND2HSV4 U13262 ( .A1(n11299), .A2(n11298), .ZN(n11333) );
  INAND2HSV2 U13263 ( .A1(n12317), .B1(n11390), .ZN(n13864) );
  NAND2HSV2 U13264 ( .A1(\pe15/bq[6] ), .A2(\pe15/aot [7]), .ZN(n11301) );
  INHSV2 U13265 ( .I(n11301), .ZN(n11303) );
  NAND2HSV2 U13266 ( .A1(\pe15/bq[5] ), .A2(\pe15/aot [8]), .ZN(n11302) );
  INHSV2 U13267 ( .I(n11302), .ZN(n11300) );
  AOI22HSV2 U13268 ( .A1(\pe15/bq[7] ), .A2(\pe15/aot [6]), .B1(n14602), .B2(
        \pe15/aot [5]), .ZN(n11308) );
  NOR2HSV2 U13269 ( .A1(n11307), .A2(n11308), .ZN(n11306) );
  NAND2HSV2 U13270 ( .A1(\pe15/aot [5]), .A2(\pe15/bq[7] ), .ZN(n11347) );
  NOR2HSV2 U13271 ( .A1(n11304), .A2(n11347), .ZN(n11309) );
  INHSV2 U13272 ( .I(n11309), .ZN(n11305) );
  OAI21HSV2 U13273 ( .A1(n11309), .A2(n11308), .B(n11307), .ZN(n11310) );
  CLKNAND2HSV3 U13274 ( .A1(n11311), .A2(n11310), .ZN(n11315) );
  NAND2HSV2 U13275 ( .A1(\pe15/got [5]), .A2(\pe15/ti_1 ), .ZN(n11313) );
  NAND2HSV2 U13276 ( .A1(\pe15/pvq [4]), .A2(n13815), .ZN(n11312) );
  XOR3HSV2 U13277 ( .A1(\pe15/phq [4]), .A2(n11313), .A3(n11312), .Z(n11314)
         );
  XNOR2HSV4 U13278 ( .A1(n11315), .A2(n11314), .ZN(n11319) );
  INHSV2 U13279 ( .I(\pe15/got [6]), .ZN(n14584) );
  XNOR2HSV4 U13280 ( .A1(n11319), .A2(n11318), .ZN(n11330) );
  CLKNHSV0 U13281 ( .I(n11330), .ZN(n11317) );
  XNOR2HSV4 U13282 ( .A1(n11319), .A2(n11318), .ZN(n11327) );
  OAI21HSV2 U13283 ( .A1(n11330), .A2(n11390), .B(n10521), .ZN(n11362) );
  NOR2HSV0 U13284 ( .A1(n11327), .A2(\pe15/got [7]), .ZN(n11320) );
  NOR3HSV2 U13285 ( .A1(n11361), .A2(n11362), .A3(n11320), .ZN(n11321) );
  NAND2HSV2 U13286 ( .A1(n13865), .A2(n11321), .ZN(n11322) );
  INHSV4 U13287 ( .I(n11322), .ZN(n11337) );
  INHSV2 U13288 ( .I(\pe15/got [7]), .ZN(n12317) );
  CLKNHSV0 U13289 ( .I(n11323), .ZN(n11326) );
  CLKNHSV2 U13290 ( .I(n11324), .ZN(n11325) );
  NOR2HSV4 U13291 ( .A1(n11326), .A2(n11325), .ZN(n11394) );
  NAND2HSV2 U13292 ( .A1(n11394), .A2(n11327), .ZN(n11328) );
  CLKNAND2HSV2 U13293 ( .A1(n11329), .A2(n11328), .ZN(n11332) );
  NOR2HSV4 U13294 ( .A1(n11332), .A2(n11331), .ZN(n11335) );
  NAND3HSV4 U13295 ( .A1(n11335), .A2(n11334), .A3(n11333), .ZN(n11367) );
  NAND2HSV2 U13296 ( .A1(n14704), .A2(\pe15/ti_7t [4]), .ZN(n11366) );
  NAND2HSV0 U13297 ( .A1(n12336), .A2(n11390), .ZN(n11338) );
  INHSV2 U13298 ( .I(n11369), .ZN(n12335) );
  NOR2HSV1 U13299 ( .A1(n12335), .A2(n12317), .ZN(n11339) );
  OR2HSV1 U13300 ( .A1(n15178), .A2(n14704), .Z(n11341) );
  NAND2HSV0 U13301 ( .A1(\pe15/got [6]), .A2(n11390), .ZN(n11360) );
  NAND2HSV0 U13302 ( .A1(\pe15/aot [6]), .A2(\pe15/bq[6] ), .ZN(n11345) );
  NAND2HSV0 U13303 ( .A1(\pe15/got [4]), .A2(\pe15/ti_1 ), .ZN(n11344) );
  XOR2HSV0 U13304 ( .A1(n11345), .A2(n11344), .Z(n11349) );
  NAND2HSV0 U13305 ( .A1(\pe15/aot [4]), .A2(\pe15/bq[8] ), .ZN(n11346) );
  XOR2HSV0 U13306 ( .A1(n11347), .A2(n11346), .Z(n11348) );
  XOR2HSV0 U13307 ( .A1(n11349), .A2(n11348), .Z(n11356) );
  NAND2HSV0 U13308 ( .A1(\pe15/aot [7]), .A2(\pe15/bq[5] ), .ZN(n11351) );
  NAND2HSV0 U13309 ( .A1(\pe15/bq[4] ), .A2(\pe15/aot [8]), .ZN(n11350) );
  XOR2HSV0 U13310 ( .A1(n11351), .A2(n11350), .Z(n11354) );
  NAND2HSV0 U13311 ( .A1(\pe15/pvq [5]), .A2(\pe15/ctrq ), .ZN(n11352) );
  XOR2HSV0 U13312 ( .A1(n11352), .A2(\pe15/phq [5]), .Z(n11353) );
  XOR2HSV0 U13313 ( .A1(n11354), .A2(n11353), .Z(n11355) );
  XOR2HSV0 U13314 ( .A1(n11356), .A2(n11355), .Z(n11358) );
  NAND2HSV2 U13315 ( .A1(n11387), .A2(\pe15/got [5]), .ZN(n11357) );
  XNOR2HSV4 U13316 ( .A1(n11358), .A2(n11357), .ZN(n11359) );
  NOR2HSV2 U13317 ( .A1(n11361), .A2(n12317), .ZN(n11364) );
  CLKNHSV0 U13318 ( .I(n11362), .ZN(n11363) );
  NAND3HSV2 U13319 ( .A1(n13865), .A2(n11364), .A3(n11363), .ZN(n11365) );
  OAI21HSV2 U13320 ( .A1(n11366), .A2(n12317), .B(n11365), .ZN(n11399) );
  CLKNHSV0 U13321 ( .I(n11367), .ZN(n11368) );
  CLKNAND2HSV2 U13322 ( .A1(n11368), .A2(n14864), .ZN(n11400) );
  INAND2HSV2 U13323 ( .A1(n11399), .B1(n11400), .ZN(n11398) );
  AND2HSV2 U13324 ( .A1(n11369), .A2(\pe15/got [6]), .Z(n11370) );
  CLKNAND2HSV1 U13325 ( .A1(n11371), .A2(n11370), .ZN(n11372) );
  NOR2HSV2 U13326 ( .A1(n11373), .A2(n11372), .ZN(n11396) );
  NAND2HSV0 U13327 ( .A1(\pe15/aot [7]), .A2(\pe15/bq[4] ), .ZN(n11375) );
  NAND2HSV0 U13328 ( .A1(\pe15/aot [5]), .A2(\pe15/bq[6] ), .ZN(n11374) );
  XOR2HSV0 U13329 ( .A1(n11375), .A2(n11374), .Z(n11379) );
  NAND2HSV0 U13330 ( .A1(\pe15/aot [4]), .A2(\pe15/bq[7] ), .ZN(n11377) );
  NAND2HSV0 U13331 ( .A1(\pe15/bq[3] ), .A2(\pe15/aot [8]), .ZN(n11376) );
  XOR2HSV0 U13332 ( .A1(n11377), .A2(n11376), .Z(n11378) );
  XOR2HSV0 U13333 ( .A1(n11379), .A2(n11378), .Z(n11386) );
  NAND2HSV0 U13334 ( .A1(\pe15/pvq [6]), .A2(\pe15/ctrq ), .ZN(n11384) );
  XOR2HSV0 U13335 ( .A1(n11381), .A2(n11380), .Z(n11382) );
  XOR3HSV2 U13336 ( .A1(n11384), .A2(n11383), .A3(n11382), .Z(n11385) );
  XNOR2HSV4 U13337 ( .A1(n11386), .A2(n11385), .ZN(n11389) );
  NAND2HSV2 U13338 ( .A1(n11387), .A2(\pe15/got [4]), .ZN(n11388) );
  XNOR2HSV4 U13339 ( .A1(n11389), .A2(n11388), .ZN(n11393) );
  NAND2HSV2 U13340 ( .A1(n11390), .A2(\pe15/got [5]), .ZN(n11391) );
  MUX2NHSV2 U13341 ( .I0(n11391), .I1(\pe15/got [5]), .S(n11393), .ZN(n11392)
         );
  XNOR2HSV4 U13342 ( .A1(n11396), .A2(n11395), .ZN(n11401) );
  INHSV3 U13343 ( .I(n11401), .ZN(n11397) );
  INHSV2 U13344 ( .I(n11399), .ZN(n11402) );
  NAND3HSV4 U13345 ( .A1(n11402), .A2(n11401), .A3(n11400), .ZN(n11403) );
  NOR2HSV1 U13346 ( .A1(n10521), .A2(\pe15/ti_7t [5]), .ZN(n12318) );
  NOR2HSV2 U13347 ( .A1(n12318), .A2(n11405), .ZN(n11698) );
  INHSV2 U13348 ( .I(n11698), .ZN(n11409) );
  BUFHSV2 U13349 ( .I(ctro15), .Z(n12829) );
  OR2HSV1 U13350 ( .A1(n11409), .A2(n12829), .Z(n11406) );
  NAND2HSV2 U13351 ( .A1(n11410), .A2(n11698), .ZN(n11411) );
  INHSV2 U13352 ( .I(n11411), .ZN(n11412) );
  NAND2HSV2 U13353 ( .A1(n10522), .A2(\pe15/ti_7t [6]), .ZN(n11413) );
  INHSV2 U13354 ( .I(ctro12), .ZN(n11448) );
  AOI21HSV1 U13355 ( .A1(n11415), .A2(n11447), .B(n11414), .ZN(n11416) );
  NAND2HSV0 U13356 ( .A1(\pe12/ti_7[1] ), .A2(\pe12/got [4]), .ZN(n11433) );
  NAND2HSV0 U13357 ( .A1(\pe12/bq[3] ), .A2(n14876), .ZN(n11419) );
  NAND2HSV0 U13358 ( .A1(\pe12/got [3]), .A2(\pe12/ti_1 ), .ZN(n11418) );
  XOR2HSV0 U13359 ( .A1(n11419), .A2(n11418), .Z(n11430) );
  NAND2HSV2 U13360 ( .A1(\pe12/ctrq ), .A2(\pe12/pvq [6]), .ZN(n11420) );
  XNOR2HSV1 U13361 ( .A1(n11420), .A2(\pe12/phq [6]), .ZN(n11421) );
  NAND2HSV0 U13362 ( .A1(\pe12/bq[7] ), .A2(\pe12/aot [4]), .ZN(n14243) );
  NAND2HSV0 U13363 ( .A1(\pe12/aot [3]), .A2(\pe12/bq[8] ), .ZN(n11422) );
  XOR2HSV0 U13364 ( .A1(n11423), .A2(n11422), .Z(n11427) );
  NAND2HSV0 U13365 ( .A1(\pe12/aot [5]), .A2(\pe12/bq[6] ), .ZN(n11425) );
  NAND2HSV0 U13366 ( .A1(\pe12/aot [6]), .A2(\pe12/bq[5] ), .ZN(n11424) );
  XOR2HSV0 U13367 ( .A1(n11425), .A2(n11424), .Z(n11426) );
  XOR2HSV0 U13368 ( .A1(n11427), .A2(n11426), .Z(n11428) );
  XOR3HSV2 U13369 ( .A1(n11430), .A2(n11429), .A3(n11428), .Z(n11432) );
  NAND2HSV0 U13370 ( .A1(\pe12/got [5]), .A2(n15192), .ZN(n11431) );
  XOR3HSV2 U13371 ( .A1(n11433), .A2(n11432), .A3(n11431), .Z(n11441) );
  INHSV2 U13372 ( .I(n11434), .ZN(n11437) );
  INHSV2 U13373 ( .I(n11435), .ZN(n11439) );
  CLKNHSV0 U13374 ( .I(\pe12/got [6]), .ZN(n12683) );
  NOR2HSV1 U13375 ( .A1(n11438), .A2(n12683), .ZN(n11440) );
  NOR2HSV1 U13376 ( .A1(n11446), .A2(\pe12/ti_7t [5]), .ZN(n11450) );
  NOR2HSV1 U13377 ( .A1(n11450), .A2(n11442), .ZN(n11443) );
  OR2HSV1 U13378 ( .A1(n11447), .A2(\pe12/got [8]), .Z(n11468) );
  CLKNAND2HSV0 U13379 ( .A1(n7206), .A2(n11448), .ZN(n11453) );
  CLKNHSV0 U13380 ( .I(n11450), .ZN(n11451) );
  CLKAND2HSV1 U13381 ( .A1(n11451), .A2(\pe12/got [7]), .Z(n11452) );
  CLKNAND2HSV1 U13382 ( .A1(\pe12/aot [5]), .A2(\pe12/bq[5] ), .ZN(n12667) );
  NAND2HSV0 U13383 ( .A1(\pe12/aot [3]), .A2(\pe12/bq[7] ), .ZN(n11454) );
  NAND2HSV0 U13384 ( .A1(\pe12/aot [6]), .A2(\pe12/bq[4] ), .ZN(n11456) );
  CLKNAND2HSV0 U13385 ( .A1(n14578), .A2(\pe12/pvq [7]), .ZN(n11457) );
  XOR2HSV0 U13386 ( .A1(n11457), .A2(\pe12/phq [7]), .Z(n11458) );
  BUFHSV2 U13387 ( .I(\pe12/ti_1 ), .Z(n13830) );
  NAND2HSV0 U13388 ( .A1(\pe12/got [2]), .A2(n13830), .ZN(n11461) );
  NAND2HSV0 U13389 ( .A1(\pe12/aot [4]), .A2(\pe12/bq[6] ), .ZN(n11460) );
  XOR2HSV0 U13390 ( .A1(n11461), .A2(n11460), .Z(n11465) );
  NAND2HSV0 U13391 ( .A1(\pe12/aot [8]), .A2(\pe12/bq[2] ), .ZN(n11463) );
  NAND2HSV0 U13392 ( .A1(n14507), .A2(\pe12/aot [2]), .ZN(n11462) );
  XOR2HSV0 U13393 ( .A1(n11463), .A2(n11462), .Z(n11464) );
  NOR2HSV2 U13394 ( .A1(n11467), .A2(n11466), .ZN(n13891) );
  CLKNHSV0 U13395 ( .I(n11469), .ZN(n11470) );
  NAND2HSV0 U13396 ( .A1(\pe5/aot [3]), .A2(\pe5/bq[8] ), .ZN(n11482) );
  NAND2HSV2 U13397 ( .A1(\pe5/bq[3] ), .A2(\pe5/aot [4]), .ZN(n13290) );
  NAND2HSV0 U13398 ( .A1(\pe5/aot [6]), .A2(\pe5/bq[5] ), .ZN(n11479) );
  NAND2HSV0 U13399 ( .A1(\pe5/bq[4] ), .A2(\pe5/aot [7]), .ZN(n11478) );
  XOR2HSV0 U13400 ( .A1(n11479), .A2(n11478), .Z(n11480) );
  XOR3HSV2 U13401 ( .A1(n11482), .A2(n11481), .A3(n11480), .Z(n11489) );
  CLKNAND2HSV0 U13402 ( .A1(\pe5/aot [5]), .A2(\pe5/bq[6] ), .ZN(n11484) );
  NAND2HSV0 U13403 ( .A1(\pe5/got [3]), .A2(\pe5/ti_1 ), .ZN(n11483) );
  XOR2HSV0 U13404 ( .A1(n11484), .A2(n11483), .Z(n11487) );
  NAND2HSV0 U13405 ( .A1(\pe5/ctrq ), .A2(\pe5/pvq [6]), .ZN(n11485) );
  XOR2HSV0 U13406 ( .A1(n11485), .A2(\pe5/phq [6]), .Z(n11486) );
  XOR2HSV0 U13407 ( .A1(n11487), .A2(n11486), .Z(n11488) );
  NAND2HSV0 U13408 ( .A1(n10346), .A2(\pe5/got [4]), .ZN(n11490) );
  INHSV2 U13409 ( .I(n11494), .ZN(n11493) );
  AOI21HSV2 U13410 ( .A1(n6922), .A2(\pe5/got [7]), .B(n11493), .ZN(n12777) );
  INHSV2 U13411 ( .I(n12777), .ZN(n12776) );
  INHSV2 U13412 ( .I(n10307), .ZN(n13283) );
  NOR2HSV4 U13413 ( .A1(n11495), .A2(n13283), .ZN(n12821) );
  CLKNAND2HSV2 U13414 ( .A1(n12780), .A2(n12821), .ZN(n12786) );
  NOR2HSV2 U13415 ( .A1(n10307), .A2(\pe5/ti_7t [5]), .ZN(n12817) );
  INHSV2 U13416 ( .I(n15067), .ZN(n12790) );
  OR2HSV1 U13417 ( .A1(n12817), .A2(n12790), .Z(n12784) );
  INHSV2 U13418 ( .I(n12784), .ZN(n12773) );
  NAND3HSV2 U13419 ( .A1(n12787), .A2(n12786), .A3(n12773), .ZN(n13013) );
  NAND2HSV0 U13420 ( .A1(\pe8/aot [7]), .A2(\pe8/bq[5] ), .ZN(n11497) );
  CLKNAND2HSV0 U13421 ( .A1(n14950), .A2(\pe8/bq[4] ), .ZN(n11496) );
  XOR2HSV0 U13422 ( .A1(n11497), .A2(n11496), .Z(n11500) );
  NAND2HSV2 U13423 ( .A1(\pe8/aot [5]), .A2(\pe8/bq[7] ), .ZN(n11565) );
  NAND2HSV0 U13424 ( .A1(\pe8/aot [4]), .A2(\pe8/bq[8] ), .ZN(n11498) );
  XOR2HSV0 U13425 ( .A1(n11565), .A2(n11498), .Z(n11499) );
  XOR2HSV0 U13426 ( .A1(n11500), .A2(n11499), .Z(n11507) );
  NAND2HSV0 U13427 ( .A1(\pe8/got [4]), .A2(\pe8/ti_1 ), .ZN(n11502) );
  NAND2HSV0 U13428 ( .A1(\pe8/aot [6]), .A2(\pe8/bq[6] ), .ZN(n11501) );
  XOR2HSV0 U13429 ( .A1(n11502), .A2(n11501), .Z(n11505) );
  NAND2HSV2 U13430 ( .A1(n11574), .A2(\pe8/pvq [5]), .ZN(n11503) );
  XOR2HSV0 U13431 ( .A1(n11503), .A2(\pe8/phq [5]), .Z(n11504) );
  XOR2HSV0 U13432 ( .A1(n11505), .A2(n11504), .Z(n11506) );
  CLKXOR2HSV4 U13433 ( .A1(n11507), .A2(n11506), .Z(n11509) );
  CLKNAND2HSV1 U13434 ( .A1(n11580), .A2(n13488), .ZN(n11510) );
  NAND2HSV2 U13435 ( .A1(n11517), .A2(n11518), .ZN(n11520) );
  NOR2HSV2 U13436 ( .A1(n11596), .A2(n11521), .ZN(n11592) );
  NAND2HSV2 U13437 ( .A1(n11596), .A2(n11602), .ZN(n11522) );
  INHSV2 U13438 ( .I(n11522), .ZN(n11537) );
  CLKNAND2HSV1 U13439 ( .A1(\pe8/ctrq ), .A2(\pe8/pvq [4]), .ZN(n11524) );
  XNOR2HSV1 U13440 ( .A1(n11524), .A2(\pe8/phq [4]), .ZN(n11526) );
  BUFHSV2 U13441 ( .I(\pe8/bq[8] ), .Z(n11845) );
  NAND2HSV0 U13442 ( .A1(n11845), .A2(\pe8/aot [5]), .ZN(n11525) );
  XNOR2HSV1 U13443 ( .A1(n11526), .A2(n11525), .ZN(n11534) );
  NAND2HSV2 U13444 ( .A1(\pe8/bq[7] ), .A2(\pe8/aot [6]), .ZN(n11528) );
  CLKNAND2HSV0 U13445 ( .A1(\pe8/bq[5] ), .A2(\pe8/aot [8]), .ZN(n11527) );
  XOR2HSV2 U13446 ( .A1(n11528), .A2(n11527), .Z(n11532) );
  CLKNAND2HSV1 U13447 ( .A1(\pe8/ti_1 ), .A2(\pe8/got [5]), .ZN(n11530) );
  NAND2HSV2 U13448 ( .A1(\pe8/aot [7]), .A2(\pe8/bq[6] ), .ZN(n11529) );
  XNOR2HSV4 U13449 ( .A1(n11530), .A2(n11529), .ZN(n11531) );
  XNOR2HSV4 U13450 ( .A1(n11532), .A2(n11531), .ZN(n11533) );
  XNOR2HSV1 U13451 ( .A1(n11534), .A2(n11533), .ZN(n11535) );
  NAND2HSV2 U13452 ( .A1(n11580), .A2(\pe8/got [7]), .ZN(n11536) );
  NOR2HSV4 U13453 ( .A1(n15267), .A2(n14190), .ZN(n11586) );
  NAND2HSV4 U13454 ( .A1(n11586), .A2(n6703), .ZN(n11595) );
  NAND2HSV4 U13455 ( .A1(n11594), .A2(n11595), .ZN(n13877) );
  MUX2NHSV2 U13456 ( .I0(n11592), .I1(n11537), .S(n13877), .ZN(n11711) );
  INHSV2 U13457 ( .I(n11538), .ZN(n11560) );
  NAND2HSV0 U13458 ( .A1(n11580), .A2(\pe8/got [4]), .ZN(n11541) );
  NAND2HSV0 U13459 ( .A1(\pe8/ti_7[1] ), .A2(\pe8/got [3]), .ZN(n11540) );
  XNOR2HSV1 U13460 ( .A1(n11541), .A2(n11540), .ZN(n11557) );
  NAND2HSV0 U13461 ( .A1(n5948), .A2(\pe8/bq[5] ), .ZN(n11543) );
  NAND2HSV0 U13462 ( .A1(n11845), .A2(\pe8/aot [2]), .ZN(n11542) );
  XOR2HSV0 U13463 ( .A1(n11543), .A2(n11542), .Z(n11555) );
  CLKNHSV2 U13464 ( .I(\pe8/aot [4]), .ZN(n14207) );
  NOR2HSV2 U13465 ( .A1(n14207), .A2(n14199), .ZN(n11564) );
  CLKNHSV0 U13466 ( .I(\pe8/aot [3]), .ZN(n11567) );
  NOR2HSV0 U13467 ( .A1(n11567), .A2(n15132), .ZN(n11544) );
  CLKNAND2HSV1 U13468 ( .A1(n8941), .A2(\pe8/aot [3]), .ZN(n14202) );
  CLKNAND2HSV1 U13469 ( .A1(\pe8/aot [4]), .A2(\pe8/bq[7] ), .ZN(n11566) );
  OAI22HSV2 U13470 ( .A1(n11564), .A2(n11544), .B1(n14202), .B2(n11566), .ZN(
        n11545) );
  XNOR2HSV1 U13471 ( .A1(n11546), .A2(n11545), .ZN(n11554) );
  CLKNAND2HSV0 U13472 ( .A1(n14950), .A2(\pe8/bq[2] ), .ZN(n11548) );
  NAND2HSV0 U13473 ( .A1(n14947), .A2(\pe8/bq[4] ), .ZN(n11547) );
  XOR2HSV0 U13474 ( .A1(n11548), .A2(n11547), .Z(n11552) );
  NAND2HSV0 U13475 ( .A1(\pe8/aot [7]), .A2(\pe8/bq[3] ), .ZN(n11550) );
  INHSV2 U13476 ( .I(n15127), .ZN(n11571) );
  NAND2HSV0 U13477 ( .A1(\pe8/got [2]), .A2(n11571), .ZN(n11549) );
  XOR2HSV0 U13478 ( .A1(n11550), .A2(n11549), .Z(n11551) );
  XOR2HSV0 U13479 ( .A1(n11552), .A2(n11551), .Z(n11553) );
  XOR3HSV2 U13480 ( .A1(n11555), .A2(n11554), .A3(n11553), .Z(n11556) );
  XNOR2HSV1 U13481 ( .A1(n11557), .A2(n11556), .ZN(n11559) );
  NAND2HSV0 U13482 ( .A1(n14857), .A2(\pe8/got [5]), .ZN(n11558) );
  NAND2HSV2 U13483 ( .A1(n14189), .A2(\pe8/ti_7t [4]), .ZN(n13876) );
  CLKNAND2HSV2 U13484 ( .A1(n13862), .A2(n13876), .ZN(n11587) );
  NAND2HSV2 U13485 ( .A1(n11560), .A2(n13876), .ZN(n11585) );
  INHSV2 U13486 ( .I(n11589), .ZN(n11561) );
  OAI21HSV4 U13487 ( .A1(n13877), .A2(n11561), .B(n13488), .ZN(n11562) );
  NAND2HSV0 U13488 ( .A1(\pe8/ti_7[1] ), .A2(\pe8/got [4]), .ZN(n11584) );
  NAND2HSV0 U13489 ( .A1(\pe8/bq[4] ), .A2(\pe8/aot [7]), .ZN(n11570) );
  XOR3HSV2 U13490 ( .A1(n11570), .A2(n11569), .A3(n11568), .Z(n11579) );
  NAND2HSV0 U13491 ( .A1(\pe8/got [3]), .A2(n11571), .ZN(n11573) );
  NAND2HSV0 U13492 ( .A1(\pe8/aot [6]), .A2(\pe8/bq[5] ), .ZN(n11572) );
  XOR2HSV0 U13493 ( .A1(n11573), .A2(n11572), .Z(n11577) );
  CLKNAND2HSV1 U13494 ( .A1(n11574), .A2(\pe8/pvq [6]), .ZN(n11575) );
  XOR2HSV0 U13495 ( .A1(n11575), .A2(\pe8/phq [6]), .Z(n11576) );
  XOR2HSV0 U13496 ( .A1(n11577), .A2(n11576), .Z(n11578) );
  CLKXOR2HSV4 U13497 ( .A1(n11579), .A2(n11578), .Z(n11583) );
  NAND2HSV0 U13498 ( .A1(n11580), .A2(\pe8/got [5]), .ZN(n11581) );
  INHSV2 U13499 ( .I(n11581), .ZN(n11582) );
  OAI21HSV1 U13500 ( .A1(n11591), .A2(\pe8/ti_7t [5]), .B(\pe8/got [8]), .ZN(
        n11590) );
  NAND3HSV2 U13501 ( .A1(n11594), .A2(n12316), .A3(n11595), .ZN(n11593) );
  INHSV2 U13502 ( .I(n11596), .ZN(n13878) );
  CLKNHSV0 U13503 ( .I(n11594), .ZN(n11600) );
  CLKNAND2HSV1 U13504 ( .A1(n11595), .A2(n11597), .ZN(n11599) );
  NOR2HSV2 U13505 ( .A1(n11596), .A2(n14190), .ZN(n11598) );
  OAI22HSV4 U13506 ( .A1(n11600), .A2(n11599), .B1(n11598), .B2(n11590), .ZN(
        n11601) );
  NAND2HSV2 U13507 ( .A1(n14190), .A2(\pe8/ti_7t [6]), .ZN(n11605) );
  NAND2HSV2 U13508 ( .A1(ctro12), .A2(\pe12/ti_7t [6]), .ZN(n11609) );
  CLKNAND2HSV1 U13509 ( .A1(n14896), .A2(\pe9/got [3]), .ZN(n11614) );
  NAND2HSV0 U13510 ( .A1(\pe9/ti_7[1] ), .A2(\pe9/got [2]), .ZN(n11613) );
  XNOR2HSV1 U13511 ( .A1(n11614), .A2(n11613), .ZN(n11634) );
  CLKNAND2HSV0 U13512 ( .A1(n13826), .A2(\pe9/pq ), .ZN(n11616) );
  NAND2HSV0 U13513 ( .A1(\pe9/aot [4]), .A2(\pe9/bq[5] ), .ZN(n11615) );
  XOR2HSV0 U13514 ( .A1(n11616), .A2(n11615), .Z(n11620) );
  NAND2HSV0 U13515 ( .A1(\pe9/aot [1]), .A2(\pe9/bq[8] ), .ZN(n11618) );
  NAND2HSV0 U13516 ( .A1(\pe9/aot [2]), .A2(n5976), .ZN(n11617) );
  XOR2HSV0 U13517 ( .A1(n11618), .A2(n11617), .Z(n11619) );
  XOR2HSV0 U13518 ( .A1(n11620), .A2(n11619), .Z(n11624) );
  NAND2HSV0 U13519 ( .A1(\pe9/aot [5]), .A2(\pe9/bq[4] ), .ZN(n11622) );
  NAND2HSV0 U13520 ( .A1(\pe9/bq[2] ), .A2(\pe9/aot [7]), .ZN(n11621) );
  XOR2HSV0 U13521 ( .A1(n11622), .A2(n11621), .Z(n11623) );
  XNOR2HSV1 U13522 ( .A1(n11624), .A2(n11623), .ZN(n11632) );
  NAND2HSV0 U13523 ( .A1(n8944), .A2(\pe9/got [1]), .ZN(n11626) );
  NAND2HSV0 U13524 ( .A1(n11647), .A2(\pe9/aot [3]), .ZN(n11625) );
  XOR2HSV0 U13525 ( .A1(n11626), .A2(n11625), .Z(n11630) );
  NAND2HSV2 U13526 ( .A1(n14942), .A2(\pe9/bq[1] ), .ZN(n11628) );
  NAND2HSV0 U13527 ( .A1(\pe9/aot [6]), .A2(\pe9/bq[3] ), .ZN(n11627) );
  XOR2HSV0 U13528 ( .A1(n11628), .A2(n11627), .Z(n11629) );
  XOR2HSV0 U13529 ( .A1(n11630), .A2(n11629), .Z(n11631) );
  XNOR2HSV1 U13530 ( .A1(n11632), .A2(n11631), .ZN(n11633) );
  XNOR2HSV1 U13531 ( .A1(n11634), .A2(n11633), .ZN(n11635) );
  NAND2HSV0 U13532 ( .A1(n14963), .A2(\pe9/got [1]), .ZN(n11641) );
  CLKNAND2HSV0 U13533 ( .A1(\pe9/aot [3]), .A2(\pe9/bq[1] ), .ZN(n11637) );
  NAND2HSV0 U13534 ( .A1(\pe9/aot [1]), .A2(\pe9/bq[3] ), .ZN(n11636) );
  XOR2HSV0 U13535 ( .A1(n11637), .A2(n11636), .Z(n11639) );
  NAND2HSV0 U13536 ( .A1(\pe9/aot [2]), .A2(\pe9/bq[2] ), .ZN(n11638) );
  XNOR2HSV1 U13537 ( .A1(n11639), .A2(n11638), .ZN(n11640) );
  XOR2HSV0 U13538 ( .A1(n11641), .A2(n11640), .Z(n11642) );
  NAND2HSV2 U13539 ( .A1(n6209), .A2(\pe9/got [3]), .ZN(n11661) );
  CLKNAND2HSV1 U13540 ( .A1(n10443), .A2(\pe9/got [2]), .ZN(n11659) );
  NAND2HSV0 U13541 ( .A1(n14896), .A2(\pe9/got [1]), .ZN(n11657) );
  NAND2HSV0 U13542 ( .A1(\pe9/aot [4]), .A2(\pe9/bq[3] ), .ZN(n11646) );
  NAND2HSV0 U13543 ( .A1(\pe9/bq[4] ), .A2(\pe9/aot [3]), .ZN(n11645) );
  XOR2HSV0 U13544 ( .A1(n11646), .A2(n11645), .Z(n11651) );
  NAND2HSV0 U13545 ( .A1(\pe9/aot [2]), .A2(\pe9/bq[5] ), .ZN(n11649) );
  NAND2HSV0 U13546 ( .A1(n11647), .A2(\pe9/aot [1]), .ZN(n11648) );
  XOR2HSV0 U13547 ( .A1(n11649), .A2(n11648), .Z(n11650) );
  XOR2HSV0 U13548 ( .A1(n11651), .A2(n11650), .Z(n11655) );
  NAND2HSV0 U13549 ( .A1(\pe9/bq[1] ), .A2(\pe9/aot [6]), .ZN(n11653) );
  NAND2HSV0 U13550 ( .A1(n8950), .A2(\pe9/bq[2] ), .ZN(n11652) );
  XOR2HSV0 U13551 ( .A1(n11653), .A2(n11652), .Z(n11654) );
  XNOR2HSV1 U13552 ( .A1(n11655), .A2(n11654), .ZN(n11656) );
  XOR2HSV0 U13553 ( .A1(n11657), .A2(n11656), .Z(n11658) );
  XOR2HSV0 U13554 ( .A1(n11659), .A2(n11658), .Z(n11660) );
  XOR2HSV0 U13555 ( .A1(n11661), .A2(n11660), .Z(n11663) );
  XOR2HSV0 U13556 ( .A1(n11663), .A2(n11662), .Z(n11664) );
  CLKNHSV0 U13557 ( .I(\pe9/got [1]), .ZN(n11667) );
  NAND2HSV0 U13558 ( .A1(\pe9/aot [1]), .A2(\pe9/bq[2] ), .ZN(n11670) );
  NAND2HSV0 U13559 ( .A1(\pe9/aot [2]), .A2(\pe9/bq[1] ), .ZN(n11669) );
  XOR2HSV0 U13560 ( .A1(n11670), .A2(n11669), .Z(n11671) );
  NAND2HSV2 U13561 ( .A1(n6209), .A2(\pe9/got [2]), .ZN(n11686) );
  CLKNAND2HSV0 U13562 ( .A1(n10443), .A2(\pe9/got [1]), .ZN(n11684) );
  NAND2HSV0 U13563 ( .A1(n8950), .A2(\pe9/bq[1] ), .ZN(n11676) );
  NAND2HSV0 U13564 ( .A1(\pe9/aot [3]), .A2(\pe9/bq[3] ), .ZN(n11675) );
  XOR2HSV0 U13565 ( .A1(n11676), .A2(n11675), .Z(n11678) );
  NAND2HSV0 U13566 ( .A1(\pe9/aot [1]), .A2(\pe9/bq[5] ), .ZN(n11677) );
  XNOR2HSV1 U13567 ( .A1(n11678), .A2(n11677), .ZN(n11682) );
  NAND2HSV0 U13568 ( .A1(\pe9/aot [4]), .A2(\pe9/bq[2] ), .ZN(n11680) );
  NAND2HSV0 U13569 ( .A1(\pe9/aot [2]), .A2(\pe9/bq[4] ), .ZN(n11679) );
  XOR2HSV0 U13570 ( .A1(n11680), .A2(n11679), .Z(n11681) );
  XNOR2HSV1 U13571 ( .A1(n11682), .A2(n11681), .ZN(n11683) );
  XNOR2HSV1 U13572 ( .A1(n11684), .A2(n11683), .ZN(n11685) );
  XNOR2HSV1 U13573 ( .A1(n11686), .A2(n11685), .ZN(n11687) );
  CLKNAND2HSV1 U13574 ( .A1(n14583), .A2(n11690), .ZN(n11695) );
  OAI21HSV0 U13575 ( .A1(n15074), .A2(\pe9/ti_7t [7]), .B(\pe9/got [5]), .ZN(
        n11693) );
  CLKNAND2HSV1 U13576 ( .A1(n11695), .A2(n11694), .ZN(n11696) );
  CLKNHSV0 U13577 ( .I(\pe15/ti_7t [5]), .ZN(n11703) );
  NOR2HSV0 U13578 ( .A1(n12337), .A2(n11703), .ZN(n11704) );
  INHSV2 U13579 ( .I(n12614), .ZN(n12514) );
  INHSV2 U13580 ( .I(n12514), .ZN(\pe15/ti_7[5] ) );
  NOR2HSV0 U13581 ( .A1(n13801), .A2(n11705), .ZN(n11706) );
  CLKBUFHSV4 U13582 ( .I(n14196), .Z(n14893) );
  CLKNHSV0 U13583 ( .I(n14219), .ZN(n14222) );
  CLKNHSV0 U13584 ( .I(n14222), .ZN(n11713) );
  INHSV2 U13585 ( .I(n11721), .ZN(n11764) );
  INHSV2 U13586 ( .I(\pe11/got [7]), .ZN(n11745) );
  NOR2HSV2 U13587 ( .A1(n11764), .A2(n11745), .ZN(n11714) );
  CLKBUFHSV4 U13588 ( .I(\pe11/bq[5] ), .Z(n11797) );
  BUFHSV8 U13589 ( .I(\pe11/aot [8]), .Z(n12424) );
  NAND2HSV2 U13590 ( .A1(n12424), .A2(\pe11/bq[4] ), .ZN(n11718) );
  CLKBUFHSV4 U13591 ( .I(\pe11/bq[6] ), .Z(n12562) );
  NAND2HSV0 U13592 ( .A1(\pe11/aot [6]), .A2(\pe11/bq[6] ), .ZN(n11717) );
  NAND2HSV0 U13593 ( .A1(\pe11/aot [5]), .A2(\pe11/bq[7] ), .ZN(n11719) );
  INHSV2 U13594 ( .I(n9609), .ZN(n11944) );
  BUFHSV4 U13595 ( .I(\pe11/got [8]), .Z(n15179) );
  CLKAND2HSV2 U13596 ( .A1(n11721), .A2(n15179), .Z(n11739) );
  NAND2HSV0 U13597 ( .A1(\pe11/got [5]), .A2(\pe11/ti_1 ), .ZN(n11723) );
  NAND2HSV0 U13598 ( .A1(\pe11/bq[5] ), .A2(\pe11/aot [8]), .ZN(n11722) );
  XOR2HSV0 U13599 ( .A1(n11723), .A2(n11722), .Z(n11727) );
  CLKNAND2HSV1 U13600 ( .A1(\pe11/bq[6] ), .A2(\pe11/aot [7]), .ZN(n11725) );
  NAND2HSV2 U13601 ( .A1(\pe11/aot [5]), .A2(\pe11/bq[8] ), .ZN(n11724) );
  XOR2HSV0 U13602 ( .A1(n11725), .A2(n11724), .Z(n11726) );
  CLKXOR2HSV4 U13603 ( .A1(n11727), .A2(n11726), .Z(n11731) );
  CLKNAND2HSV0 U13604 ( .A1(\pe11/aot [6]), .A2(\pe11/bq[7] ), .ZN(n11729) );
  NAND2HSV2 U13605 ( .A1(n14791), .A2(\pe11/pvq [4]), .ZN(n11728) );
  XOR3HSV2 U13606 ( .A1(\pe11/phq [4]), .A2(n11729), .A3(n11728), .Z(n11730)
         );
  XNOR2HSV4 U13607 ( .A1(n11731), .A2(n11730), .ZN(n11736) );
  CLKNAND2HSV1 U13608 ( .A1(n11732), .A2(\pe11/got [6]), .ZN(n11733) );
  NOR2HSV4 U13609 ( .A1(n11734), .A2(n11733), .ZN(n11735) );
  XOR2HSV2 U13610 ( .A1(n11736), .A2(n11735), .Z(n11737) );
  NAND2HSV2 U13611 ( .A1(n11948), .A2(\pe11/ti_7t [4]), .ZN(n11897) );
  INHSV2 U13612 ( .I(n11897), .ZN(n11895) );
  INHSV2 U13613 ( .I(n14365), .ZN(n11776) );
  INHSV3 U13614 ( .I(n11738), .ZN(n11743) );
  NAND3HSV4 U13615 ( .A1(n11741), .A2(n11740), .A3(n11739), .ZN(n11742) );
  NOR2HSV1 U13616 ( .A1(n11944), .A2(\pe11/ti_7t [5]), .ZN(n11903) );
  NOR2HSV1 U13617 ( .A1(n11903), .A2(n11896), .ZN(n11744) );
  BUFHSV2 U13618 ( .I(n14381), .Z(n12561) );
  CLKNAND2HSV1 U13619 ( .A1(n12561), .A2(\pe11/got [5]), .ZN(n11763) );
  NAND2HSV2 U13620 ( .A1(\pe11/ctrq ), .A2(\pe11/pvq [6]), .ZN(n11747) );
  CLKNAND2HSV1 U13621 ( .A1(\pe11/bq[4] ), .A2(n14837), .ZN(n11746) );
  XOR3HSV2 U13622 ( .A1(\pe11/phq [6]), .A2(n11747), .A3(n11746), .Z(n11751)
         );
  CLKBUFHSV4 U13623 ( .I(\pe11/bq[7] ), .Z(n14519) );
  CLKNAND2HSV1 U13624 ( .A1(\pe11/aot [4]), .A2(n14519), .ZN(n11749) );
  NAND2HSV0 U13625 ( .A1(\pe11/got [3]), .A2(\pe11/ti_1 ), .ZN(n11748) );
  XNOR2HSV1 U13626 ( .A1(n11749), .A2(n11748), .ZN(n11750) );
  CLKNAND2HSV0 U13627 ( .A1(\pe11/aot [5]), .A2(\pe11/bq[6] ), .ZN(n11753) );
  NAND2HSV0 U13628 ( .A1(n11924), .A2(\pe11/aot [3]), .ZN(n11752) );
  XOR2HSV0 U13629 ( .A1(n11753), .A2(n11752), .Z(n11757) );
  CLKNAND2HSV1 U13630 ( .A1(n12424), .A2(\pe11/bq[3] ), .ZN(n11755) );
  NAND2HSV0 U13631 ( .A1(\pe11/aot [6]), .A2(\pe11/bq[5] ), .ZN(n11754) );
  XOR2HSV0 U13632 ( .A1(n11755), .A2(n11754), .Z(n11756) );
  XNOR2HSV1 U13633 ( .A1(n11757), .A2(n11756), .ZN(n11758) );
  XNOR2HSV2 U13634 ( .A1(n11759), .A2(n11758), .ZN(n11761) );
  CLKNAND2HSV1 U13635 ( .A1(\pe11/ti_7[1] ), .A2(\pe11/got [4]), .ZN(n11760)
         );
  XNOR2HSV2 U13636 ( .A1(n11761), .A2(n11760), .ZN(n11762) );
  XNOR2HSV4 U13637 ( .A1(n11763), .A2(n11762), .ZN(n11772) );
  NOR2HSV2 U13638 ( .A1(n11764), .A2(n15146), .ZN(n11768) );
  INAND2HSV2 U13639 ( .A1(n7684), .B1(n11766), .ZN(n11769) );
  NAND3HSV2 U13640 ( .A1(n11770), .A2(n11769), .A3(n11768), .ZN(n11771) );
  INHSV1 U13641 ( .I(n11773), .ZN(n14825) );
  INHSV1 U13642 ( .I(n13476), .ZN(n15191) );
  NAND2HSV4 U13643 ( .A1(n13177), .A2(n13176), .ZN(n15168) );
  CLKNHSV0 U13644 ( .I(n11954), .ZN(n14728) );
  CLKNHSV0 U13645 ( .I(n14817), .ZN(n11959) );
  CLKNHSV0 U13646 ( .I(n11959), .ZN(n14801) );
  CLKBUFHSV4 U13647 ( .I(n11775), .Z(n15066) );
  INHSV2 U13648 ( .I(n11776), .ZN(n14737) );
  CLKNHSV0 U13649 ( .I(n11953), .ZN(n14748) );
  NAND2HSV0 U13650 ( .A1(\pe2/ti_7[1] ), .A2(n14818), .ZN(n11779) );
  XNOR2HSV0 U13651 ( .A1(n11779), .A2(n11778), .ZN(n15294) );
  INHSV2 U13652 ( .I(n14005), .ZN(\pe1/ti_7[3] ) );
  AO21HSV1 U13653 ( .A1(n8948), .A2(n9103), .B(n11784), .Z(n14964) );
  CLKNHSV0 U13654 ( .I(rst), .ZN(n11894) );
  CLKNHSV0 U13655 ( .I(\pe21/bq[5] ), .ZN(n11785) );
  INHSV2 U13656 ( .I(n11785), .ZN(n11787) );
  MUX2HSV2 U13657 ( .I0(bo21[5]), .I1(n11787), .S(n11786), .Z(n15172) );
  BUFHSV2 U13658 ( .I(n14578), .Z(n14938) );
  INHSV2 U13659 ( .I(\pe3/pq ), .ZN(n11789) );
  CLKNHSV0 U13660 ( .I(n12357), .ZN(n11788) );
  MUX2HSV2 U13661 ( .I0(n8924), .I1(n11789), .S(n11788), .Z(\pe3/ti_1t ) );
  MUX2HSV2 U13662 ( .I0(bo3[2]), .I1(\pe3/bq[2] ), .S(n12357), .Z(n15102) );
  BUFHSV2 U13663 ( .I(n11790), .Z(n12474) );
  CLKNHSV0 U13664 ( .I(\pe3/bq[6] ), .ZN(n11791) );
  INHSV2 U13665 ( .I(n11791), .ZN(n11792) );
  MUX2HSV2 U13666 ( .I0(bo3[6]), .I1(n11792), .S(n11790), .Z(n15100) );
  INHSV2 U13667 ( .I(\pe10/pq ), .ZN(n11794) );
  INHSV2 U13668 ( .I(n14554), .ZN(n11793) );
  MUX2HSV2 U13669 ( .I0(n15139), .I1(n11794), .S(n11793), .Z(\pe10/ti_1t ) );
  INHSV2 U13670 ( .I(n11796), .ZN(n14925) );
  INHSV2 U13671 ( .I(n11838), .ZN(n14553) );
  MUX2HSV1 U13672 ( .I0(bo11[5]), .I1(n11797), .S(n14553), .Z(n15141) );
  CLKNHSV0 U13673 ( .I(\pe4/bq[3] ), .ZN(n11798) );
  INHSV2 U13674 ( .I(n11798), .ZN(n11799) );
  MUX2HSV2 U13675 ( .I0(bo4[3]), .I1(n11799), .S(n10562), .Z(n15106) );
  BUFHSV2 U13676 ( .I(\pe4/bq[4] ), .Z(n11800) );
  MUX2HSV2 U13677 ( .I0(bo4[4]), .I1(n11800), .S(n10562), .Z(n15107) );
  MUX2HSV1 U13678 ( .I0(bo4[5]), .I1(\pe4/bq[5] ), .S(n10562), .Z(n15105) );
  MUX2HSV2 U13679 ( .I0(bo7[6]), .I1(n8930), .S(n12067), .Z(n15124) );
  MUX2HSV1 U13680 ( .I0(bo4[6]), .I1(n12581), .S(n13822), .Z(n15104) );
  CLKNHSV0 U13681 ( .I(bo5[2]), .ZN(n11803) );
  CLKNHSV0 U13682 ( .I(\pe5/bq[2] ), .ZN(n11802) );
  CLKNHSV0 U13683 ( .I(\pe5/ctrq ), .ZN(n11812) );
  MUX2NHSV1 U13684 ( .I0(n11803), .I1(n11802), .S(n11818), .ZN(n15038) );
  CLKNHSV0 U13685 ( .I(\pe5/bq[8] ), .ZN(n11804) );
  INHSV2 U13686 ( .I(n11804), .ZN(n13419) );
  MUX2HSV2 U13687 ( .I0(bo5[8]), .I1(n13419), .S(n11818), .Z(n15108) );
  BUFHSV2 U13688 ( .I(\pe20/bq[7] ), .Z(n13737) );
  MUX2HSV2 U13689 ( .I0(bo20[7]), .I1(n13737), .S(n12362), .Z(n15169) );
  CLKNHSV0 U13690 ( .I(\pe20/bq[4] ), .ZN(n11805) );
  INHSV2 U13691 ( .I(n11805), .ZN(n11806) );
  MUX2HSV2 U13692 ( .I0(bo20[4]), .I1(n11806), .S(n12362), .Z(n15170) );
  CLKNHSV0 U13693 ( .I(\pe20/bq[3] ), .ZN(n11807) );
  INHSV2 U13694 ( .I(n11807), .ZN(n11808) );
  MUX2HSV2 U13695 ( .I0(bo20[3]), .I1(n11808), .S(n12362), .Z(n15171) );
  INHSV2 U13696 ( .I(\pe8/pq ), .ZN(n11810) );
  INHSV2 U13697 ( .I(n14572), .ZN(n11809) );
  MUX2HSV2 U13698 ( .I0(n15127), .I1(n11810), .S(n11809), .Z(\pe8/ti_1t ) );
  MUX2NHSV1 U13699 ( .I0(bo11[8]), .I1(n11924), .S(n14553), .ZN(n14980) );
  CLKNHSV0 U13700 ( .I(\pe5/bq[6] ), .ZN(n11811) );
  INHSV1 U13701 ( .I(n11811), .ZN(n11813) );
  MUX2HSV1 U13702 ( .I0(bo5[6]), .I1(n11813), .S(n11818), .Z(n15111) );
  CLKNHSV0 U13703 ( .I(\pe5/bq[3] ), .ZN(n11814) );
  INHSV1 U13704 ( .I(n11814), .ZN(n11815) );
  MUX2HSV1 U13705 ( .I0(bo5[3]), .I1(n11815), .S(n11818), .Z(n15112) );
  BUFHSV2 U13706 ( .I(\pe5/bq[4] ), .Z(n11816) );
  MUX2HSV1 U13707 ( .I0(bo5[4]), .I1(n11816), .S(n11818), .Z(n15113) );
  BUFHSV2 U13708 ( .I(\pe18/aot [6]), .Z(n14894) );
  CLKNHSV0 U13709 ( .I(\pe5/bq[5] ), .ZN(n11817) );
  INHSV1 U13710 ( .I(n11817), .ZN(n11819) );
  MUX2HSV1 U13711 ( .I0(bo5[5]), .I1(n11819), .S(n11818), .Z(n15109) );
  CLKNHSV0 U13712 ( .I(\pe6/bq[4] ), .ZN(n11820) );
  INHSV1 U13713 ( .I(n11820), .ZN(n11821) );
  INHSV2 U13714 ( .I(n14869), .ZN(n13828) );
  MUX2HSV1 U13715 ( .I0(bo6[4]), .I1(n11821), .S(n13828), .Z(n15117) );
  CLKNHSV0 U13716 ( .I(\pe6/bq[5] ), .ZN(n11822) );
  INHSV1 U13717 ( .I(n11822), .ZN(n11823) );
  MUX2HSV1 U13718 ( .I0(bo6[5]), .I1(n11823), .S(n13041), .Z(n15116) );
  CLKNHSV0 U13719 ( .I(\pe7/bq[7] ), .ZN(n11824) );
  INHSV2 U13720 ( .I(n11824), .ZN(n11825) );
  MUX2HSV2 U13721 ( .I0(bo7[7]), .I1(n11825), .S(n12067), .Z(n15123) );
  MUX2HSV2 U13722 ( .I0(bo7[3]), .I1(\pe7/bq[3] ), .S(n12067), .Z(n15125) );
  CLKNHSV0 U13723 ( .I(\pe15/aot [6]), .ZN(n11826) );
  INHSV2 U13724 ( .I(n11826), .ZN(n14739) );
  INHSV2 U13725 ( .I(n11827), .ZN(n14743) );
  CLKNHSV0 U13726 ( .I(\pe16/bq[3] ), .ZN(n11828) );
  INHSV1 U13727 ( .I(n11828), .ZN(n11829) );
  MUX2HSV1 U13728 ( .I0(bo16[3]), .I1(n11829), .S(n14570), .Z(n15163) );
  INHSV2 U13729 ( .I(n11834), .ZN(n13820) );
  MUX2HSV1 U13730 ( .I0(bo13[3]), .I1(\pe13/bq[3] ), .S(n13820), .Z(n15152) );
  INHSV2 U13731 ( .I(n11834), .ZN(n14795) );
  MUX2HSV2 U13732 ( .I0(bo13[4]), .I1(\pe13/bq[4] ), .S(n14795), .Z(n15149) );
  CLKNHSV0 U13733 ( .I(\pe9/bq[1] ), .ZN(n11830) );
  INHSV1 U13734 ( .I(n11830), .ZN(n11831) );
  MUX2HSV1 U13735 ( .I0(bo9[1]), .I1(n11831), .S(n13826), .Z(n15138) );
  CLKNHSV0 U13736 ( .I(\pe13/bq[6] ), .ZN(n11833) );
  INHSV2 U13737 ( .I(n11833), .ZN(n11835) );
  MUX2HSV2 U13738 ( .I0(bo13[6]), .I1(n11835), .S(n13820), .Z(n15150) );
  MUX2HSV2 U13739 ( .I0(bo13[7]), .I1(n13591), .S(n13820), .Z(n15148) );
  CLKNHSV0 U13740 ( .I(\pe3/aot [7]), .ZN(n11836) );
  INHSV2 U13741 ( .I(n11836), .ZN(n14738) );
  CLKNHSV0 U13742 ( .I(\pe11/bq[3] ), .ZN(n11837) );
  INHSV1 U13743 ( .I(n11837), .ZN(n11839) );
  INHSV2 U13744 ( .I(n11838), .ZN(n13812) );
  MUX2HSV1 U13745 ( .I0(bo11[3]), .I1(n11839), .S(n13812), .Z(n15144) );
  MUX2HSV1 U13746 ( .I0(bo11[2]), .I1(\pe11/bq[2] ), .S(n13812), .Z(n15143) );
  MUX2HSV1 U13747 ( .I0(bo11[1]), .I1(\pe11/bq[1] ), .S(n13812), .Z(n15145) );
  MUX2HSV1 U13748 ( .I0(bo11[6]), .I1(n12562), .S(n13812), .Z(n15142) );
  BUFHSV2 U13749 ( .I(\pe17/ctrq ), .Z(n14892) );
  MUX2HSV1 U13750 ( .I0(bo17[2]), .I1(\pe17/bq[2] ), .S(n14892), .Z(n15166) );
  CLKNHSV0 U13751 ( .I(\pe17/bq[5] ), .ZN(n11840) );
  INHSV1 U13752 ( .I(n11840), .ZN(n11841) );
  MUX2HSV1 U13753 ( .I0(bo17[5]), .I1(n11841), .S(n14892), .Z(n15165) );
  CLKNHSV0 U13754 ( .I(\pe14/bq[4] ), .ZN(n11842) );
  INHSV2 U13755 ( .I(n11842), .ZN(n11843) );
  INHSV2 U13756 ( .I(n13067), .ZN(n14535) );
  MUX2HSV2 U13757 ( .I0(bo14[4]), .I1(n11843), .S(n14535), .Z(n15153) );
  MUX2HSV2 U13758 ( .I0(bo15[1]), .I1(\pe15/bq[1] ), .S(n13815), .Z(n15159) );
  CLKBUFHSV4 U13759 ( .I(\pe15/bq[5] ), .Z(n12616) );
  INHSV2 U13760 ( .I(n11844), .ZN(n14586) );
  MUX2HSV2 U13761 ( .I0(bo15[5]), .I1(n12616), .S(n14586), .Z(n15158) );
  MUX2HSV2 U13762 ( .I0(bo8[8]), .I1(n11845), .S(n14758), .Z(n15128) );
  CLKNHSV0 U13763 ( .I(\pe15/bq[6] ), .ZN(n11846) );
  INHSV2 U13764 ( .I(n11846), .ZN(n11847) );
  BUFHSV2 U13765 ( .I(\pe15/ctrq ), .Z(n12343) );
  MUX2HSV2 U13766 ( .I0(bo15[6]), .I1(n11847), .S(n12343), .Z(n15156) );
  MUX2HSV2 U13767 ( .I0(bo8[6]), .I1(n8941), .S(n14758), .Z(n15130) );
  CLKNHSV0 U13768 ( .I(\pe15/bq[7] ), .ZN(n11849) );
  INHSV2 U13769 ( .I(n11849), .ZN(n11850) );
  MUX2HSV2 U13770 ( .I0(bo15[7]), .I1(n11850), .S(n12343), .Z(n15157) );
  MUX2HSV2 U13771 ( .I0(bo8[1]), .I1(\pe8/bq[1] ), .S(n14572), .Z(n15131) );
  CLKNHSV0 U13772 ( .I(\pe14/bq[1] ), .ZN(n11851) );
  INHSV2 U13773 ( .I(n11851), .ZN(n11852) );
  MUX2HSV2 U13774 ( .I0(bo14[1]), .I1(n11852), .S(n14535), .Z(n15154) );
  INHSV2 U13775 ( .I(\pe17/got [1]), .ZN(n14319) );
  MUX2HSV1 U13776 ( .I0(bo15[3]), .I1(\pe15/bq[3] ), .S(n15160), .Z(n15161) );
  BUFHSV8 U13777 ( .I(\pe17/bq[7] ), .Z(n14412) );
  MUX2HSV1 U13778 ( .I0(bo17[7]), .I1(n14412), .S(n14892), .Z(n15164) );
  MUX2HSV1 U13779 ( .I0(bo6[3]), .I1(\pe6/bq[3] ), .S(n14870), .Z(n15119) );
  MUX2HSV1 U13780 ( .I0(bo6[2]), .I1(\pe6/bq[2] ), .S(n14870), .Z(n15120) );
  MUX2HSV1 U13781 ( .I0(bo6[1]), .I1(\pe6/bq[1] ), .S(n13041), .Z(n15118) );
  CLKNHSV0 U13782 ( .I(n11957), .ZN(n14833) );
  BUFHSV2 U13783 ( .I(\pe19/aot [7]), .Z(n14945) );
  BUFHSV2 U13784 ( .I(\pe7/got [7]), .Z(n14829) );
  INHSV2 U13785 ( .I(n14848), .ZN(n14849) );
  CLKNHSV0 U13786 ( .I(\pe14/aot [7]), .ZN(n11853) );
  INHSV2 U13787 ( .I(n11853), .ZN(n14706) );
  NAND2HSV2 U13788 ( .A1(n15184), .A2(\pe20/got [6]), .ZN(n11876) );
  CLKNAND2HSV0 U13789 ( .A1(\pe20/aot [3]), .A2(n13737), .ZN(n11857) );
  NAND2HSV0 U13790 ( .A1(\pe20/aot [5]), .A2(\pe20/bq[5] ), .ZN(n11856) );
  XOR2HSV0 U13791 ( .A1(n11857), .A2(n11856), .Z(n11870) );
  NAND2HSV0 U13792 ( .A1(n14946), .A2(\pe20/bq[4] ), .ZN(n11859) );
  NAND2HSV0 U13793 ( .A1(\pe20/got [2]), .A2(n13738), .ZN(n11858) );
  XOR2HSV0 U13794 ( .A1(n11859), .A2(n11858), .Z(n11861) );
  XNOR2HSV1 U13795 ( .A1(n11861), .A2(n11860), .ZN(n11869) );
  NAND2HSV0 U13796 ( .A1(\pe20/aot [4]), .A2(\pe20/bq[6] ), .ZN(n11863) );
  NAND2HSV0 U13797 ( .A1(\pe20/aot [7]), .A2(\pe20/bq[3] ), .ZN(n11862) );
  XOR2HSV0 U13798 ( .A1(n11863), .A2(n11862), .Z(n11867) );
  CLKNAND2HSV0 U13799 ( .A1(\pe20/bq[2] ), .A2(n13733), .ZN(n11865) );
  NAND2HSV0 U13800 ( .A1(\pe20/aot [2]), .A2(\pe20/bq[8] ), .ZN(n11864) );
  XOR2HSV0 U13801 ( .A1(n11865), .A2(n11864), .Z(n11866) );
  XOR2HSV0 U13802 ( .A1(n11867), .A2(n11866), .Z(n11868) );
  XOR3HSV2 U13803 ( .A1(n11870), .A2(n11869), .A3(n11868), .Z(n11871) );
  XNOR2HSV1 U13804 ( .A1(n11872), .A2(n11871), .ZN(n11873) );
  XNOR2HSV4 U13805 ( .A1(n11876), .A2(n11875), .ZN(n11891) );
  INHSV2 U13806 ( .I(n15184), .ZN(n13640) );
  INHSV4 U13807 ( .I(n13640), .ZN(n13695) );
  NOR2HSV2 U13808 ( .A1(n9459), .A2(n15177), .ZN(n13647) );
  INHSV2 U13809 ( .I(n13647), .ZN(n11877) );
  CLKNAND2HSV0 U13810 ( .A1(n11888), .A2(n14821), .ZN(n11878) );
  CLKNHSV0 U13811 ( .I(n11878), .ZN(n11879) );
  NAND2HSV0 U13812 ( .A1(n11879), .A2(n9459), .ZN(n11884) );
  NOR2HSV1 U13813 ( .A1(n15177), .A2(n11880), .ZN(n11892) );
  CLKNHSV0 U13814 ( .I(n11892), .ZN(n11882) );
  CLKNAND2HSV0 U13815 ( .A1(n13641), .A2(n13718), .ZN(n11881) );
  IAO21HSV4 U13816 ( .A1(n9459), .A2(n11882), .B(n11881), .ZN(n11883) );
  CLKNAND2HSV2 U13817 ( .A1(n11883), .A2(n11884), .ZN(n11885) );
  NOR2HSV4 U13818 ( .A1(n11886), .A2(n11885), .ZN(n11890) );
  XNOR2HSV4 U13819 ( .A1(n11891), .A2(n11890), .ZN(n13794) );
  NAND2HSV0 U13820 ( .A1(n13749), .A2(n11888), .ZN(n11889) );
  INHSV2 U13821 ( .I(n11889), .ZN(n11893) );
  CLKNHSV0 U13822 ( .I(n11956), .ZN(n14710) );
  CLKNHSV0 U13823 ( .I(n11953), .ZN(n14711) );
  CLKNHSV0 U13824 ( .I(n11956), .ZN(n14712) );
  CLKNHSV0 U13825 ( .I(n11959), .ZN(n14713) );
  CLKNHSV0 U13826 ( .I(n11954), .ZN(n14714) );
  CLKNHSV0 U13827 ( .I(n8938), .ZN(n11954) );
  CLKNHSV0 U13828 ( .I(n11954), .ZN(n14715) );
  CLKNHSV0 U13829 ( .I(n11954), .ZN(n14716) );
  CLKNHSV0 U13830 ( .I(n11956), .ZN(n14717) );
  CLKNHSV0 U13831 ( .I(n14811), .ZN(n11957) );
  CLKNHSV0 U13832 ( .I(n11957), .ZN(n14718) );
  CLKNHSV0 U13833 ( .I(n11957), .ZN(n14719) );
  CLKNHSV0 U13834 ( .I(n11959), .ZN(n14720) );
  CLKNHSV0 U13835 ( .I(n14713), .ZN(n11952) );
  CLKNHSV0 U13836 ( .I(n11952), .ZN(n14722) );
  CLKNHSV0 U13837 ( .I(n11952), .ZN(n14723) );
  CLKNHSV0 U13838 ( .I(n11957), .ZN(n14724) );
  CLKNHSV0 U13839 ( .I(n14833), .ZN(n11960) );
  CLKNHSV0 U13840 ( .I(n11958), .ZN(n14725) );
  CLKNHSV0 U13841 ( .I(n11953), .ZN(n14726) );
  CLKNHSV0 U13842 ( .I(n12346), .ZN(n14727) );
  CLKNHSV0 U13843 ( .I(n11957), .ZN(n14749) );
  CLKNHSV0 U13844 ( .I(n11957), .ZN(n14729) );
  CLKNHSV0 U13845 ( .I(n11954), .ZN(n14730) );
  CLKNHSV0 U13846 ( .I(n11957), .ZN(n14731) );
  CLKNHSV0 U13847 ( .I(n11952), .ZN(n14732) );
  AOI21HSV1 U13848 ( .A1(ctro11), .A2(n11897), .B(n11896), .ZN(n11900) );
  INHSV2 U13849 ( .I(n11900), .ZN(n11898) );
  INAND2HSV2 U13850 ( .A1(n12348), .B1(n11899), .ZN(n11908) );
  INAND2HSV0 U13851 ( .A1(n11948), .B1(n11900), .ZN(n11901) );
  CLKNHSV0 U13852 ( .I(n11903), .ZN(n11904) );
  CLKNAND2HSV1 U13853 ( .A1(n11904), .A2(\pe11/got [7]), .ZN(n11905) );
  NAND2HSV2 U13854 ( .A1(n11908), .A2(n11907), .ZN(n11941) );
  CLKNAND2HSV1 U13855 ( .A1(n15090), .A2(\pe11/ti_7t [3]), .ZN(n12354) );
  CLKNHSV0 U13856 ( .I(n12354), .ZN(n11911) );
  INHSV1 U13857 ( .I(\pe11/got [5]), .ZN(n11909) );
  AOI21HSV1 U13858 ( .A1(n11948), .A2(n12354), .B(n11909), .ZN(n11910) );
  OAI21HSV2 U13859 ( .A1(n15258), .A2(n11911), .B(n11910), .ZN(n11939) );
  NAND2HSV0 U13860 ( .A1(n12424), .A2(\pe11/bq[2] ), .ZN(n11913) );
  INHSV2 U13861 ( .I(\pe11/phq [7]), .ZN(n11912) );
  XNOR2HSV1 U13862 ( .A1(n11913), .A2(n11912), .ZN(n11915) );
  CLKNAND2HSV0 U13863 ( .A1(n11915), .A2(\pe11/got [3]), .ZN(n11920) );
  NOR2HSV0 U13864 ( .A1(n11915), .A2(n11914), .ZN(n11918) );
  OAI22HSV0 U13865 ( .A1(n11920), .A2(n11916), .B1(\pe11/got [3]), .B2(n11915), 
        .ZN(n11917) );
  AOI21HSV2 U13866 ( .A1(n11921), .A2(n11918), .B(n11917), .ZN(n11919) );
  OAI21HSV2 U13867 ( .A1(n11921), .A2(n11920), .B(n11919), .ZN(n11937) );
  NAND2HSV0 U13868 ( .A1(\pe11/aot [6]), .A2(\pe11/bq[4] ), .ZN(n11923) );
  NAND2HSV0 U13869 ( .A1(\pe11/aot [4]), .A2(n12562), .ZN(n11922) );
  XOR2HSV0 U13870 ( .A1(n11923), .A2(n11922), .Z(n11927) );
  NAND2HSV0 U13871 ( .A1(n11924), .A2(\pe11/aot [2]), .ZN(n12429) );
  NAND2HSV0 U13872 ( .A1(\pe11/aot [5]), .A2(\pe11/bq[5] ), .ZN(n11925) );
  CLKNAND2HSV0 U13873 ( .A1(n14519), .A2(\pe11/aot [3]), .ZN(n11929) );
  CLKNAND2HSV0 U13874 ( .A1(n14837), .A2(\pe11/bq[3] ), .ZN(n11928) );
  XOR2HSV0 U13875 ( .A1(n11929), .A2(n11928), .Z(n11933) );
  NAND2HSV2 U13876 ( .A1(\pe11/got [2]), .A2(n13811), .ZN(n11931) );
  CLKNAND2HSV1 U13877 ( .A1(n14791), .A2(\pe11/pvq [7]), .ZN(n11930) );
  XOR2HSV0 U13878 ( .A1(n11931), .A2(n11930), .Z(n11932) );
  XOR2HSV0 U13879 ( .A1(n11933), .A2(n11932), .Z(n11934) );
  XOR2HSV0 U13880 ( .A1(n11935), .A2(n11934), .Z(n11936) );
  NAND2HSV2 U13881 ( .A1(n12561), .A2(\pe11/got [4]), .ZN(n11938) );
  XNOR2HSV4 U13882 ( .A1(n11941), .A2(n11940), .ZN(n11946) );
  NAND2HSV2 U13883 ( .A1(n9609), .A2(\pe11/ti_7t [6]), .ZN(n12192) );
  MUX2NHSV4 U13884 ( .I0(n11945), .I1(n8909), .S(n14388), .ZN(n12453) );
  INHSV2 U13885 ( .I(n11946), .ZN(n13889) );
  NOR2HSV1 U13886 ( .A1(n15179), .A2(n15090), .ZN(n11947) );
  AOI22HSV4 U13887 ( .A1(n11948), .A2(\pe11/ti_7t [7]), .B1(n13889), .B2(
        n11947), .ZN(n12452) );
  XOR2HSV0 U13888 ( .A1(n11950), .A2(n11949), .Z(n14734) );
  CLKNHSV0 U13889 ( .I(n11951), .ZN(n14887) );
  CLKNHSV0 U13890 ( .I(\pe19/ctrq ), .ZN(n14543) );
  CLKNHSV0 U13891 ( .I(n11954), .ZN(n14744) );
  CLKNHSV0 U13892 ( .I(n11954), .ZN(n14745) );
  CLKNHSV0 U13893 ( .I(n14723), .ZN(n11956) );
  CLKNHSV0 U13894 ( .I(n11956), .ZN(n14746) );
  CLKNHSV0 U13895 ( .I(n11956), .ZN(n14747) );
  CLKNHSV0 U13896 ( .I(n11959), .ZN(n14751) );
  CLKNHSV0 U13897 ( .I(n11957), .ZN(n14752) );
  CLKNHSV0 U13898 ( .I(n14728), .ZN(n11955) );
  CLKNHSV0 U13899 ( .I(n14771), .ZN(n11953) );
  CLKNHSV0 U13900 ( .I(n11953), .ZN(n14753) );
  CLKNHSV0 U13901 ( .I(n11953), .ZN(n14754) );
  CLKNHSV0 U13902 ( .I(n11956), .ZN(n14755) );
  CLKNHSV0 U13903 ( .I(n11957), .ZN(n14756) );
  CLKNHSV0 U13904 ( .I(n11953), .ZN(n14757) );
  CLKNHSV0 U13905 ( .I(n11952), .ZN(n14759) );
  CLKNHSV0 U13906 ( .I(n12346), .ZN(n14760) );
  CLKNHSV0 U13907 ( .I(n11959), .ZN(n14762) );
  CLKNHSV0 U13908 ( .I(n12346), .ZN(n14763) );
  CLKNHSV0 U13909 ( .I(n11952), .ZN(n14764) );
  CLKNHSV0 U13910 ( .I(n11953), .ZN(n14765) );
  CLKNHSV0 U13911 ( .I(n11957), .ZN(n14766) );
  CLKNHSV0 U13912 ( .I(n11952), .ZN(n14767) );
  CLKNHSV0 U13913 ( .I(n14767), .ZN(n11958) );
  CLKNHSV0 U13914 ( .I(n11958), .ZN(n14768) );
  CLKNHSV0 U13915 ( .I(n11956), .ZN(n14769) );
  CLKNHSV0 U13916 ( .I(n11953), .ZN(n14770) );
  CLKNHSV0 U13917 ( .I(n11952), .ZN(n14771) );
  CLKNHSV0 U13918 ( .I(n11960), .ZN(n14772) );
  CLKNHSV0 U13919 ( .I(n11958), .ZN(n14773) );
  CLKNHSV0 U13920 ( .I(n11952), .ZN(n14774) );
  CLKNHSV0 U13921 ( .I(n12346), .ZN(n14775) );
  CLKNHSV0 U13922 ( .I(n11952), .ZN(n14776) );
  CLKNHSV0 U13923 ( .I(n11954), .ZN(n14777) );
  CLKNHSV0 U13924 ( .I(n11953), .ZN(n14778) );
  CLKNHSV0 U13925 ( .I(n12346), .ZN(n14779) );
  CLKNHSV0 U13926 ( .I(n11954), .ZN(n14780) );
  CLKNHSV0 U13927 ( .I(n11952), .ZN(n14781) );
  CLKNHSV0 U13928 ( .I(n11954), .ZN(n14782) );
  CLKNHSV0 U13929 ( .I(n11959), .ZN(n14783) );
  CLKNHSV0 U13930 ( .I(n11953), .ZN(n14784) );
  CLKNHSV0 U13931 ( .I(n11956), .ZN(n14785) );
  CLKNHSV0 U13932 ( .I(n11956), .ZN(n14786) );
  CLKNHSV0 U13933 ( .I(n11957), .ZN(n14787) );
  CLKNHSV0 U13934 ( .I(n12346), .ZN(n14789) );
  CLKNHSV0 U13935 ( .I(n11958), .ZN(n14792) );
  CLKNHSV0 U13936 ( .I(n11958), .ZN(n14793) );
  CLKNHSV0 U13937 ( .I(n11958), .ZN(n14794) );
  CLKNHSV0 U13938 ( .I(n12346), .ZN(n14796) );
  CLKNHSV0 U13939 ( .I(n11959), .ZN(n14797) );
  CLKNHSV0 U13940 ( .I(n11956), .ZN(n14798) );
  CLKNHSV0 U13941 ( .I(n12346), .ZN(n14799) );
  CLKNHSV0 U13942 ( .I(n11953), .ZN(n14800) );
  CLKNHSV0 U13943 ( .I(n11956), .ZN(n14802) );
  CLKNHSV0 U13944 ( .I(n11959), .ZN(n14803) );
  CLKNHSV0 U13945 ( .I(n12346), .ZN(n14804) );
  CLKNHSV0 U13946 ( .I(n11959), .ZN(n14806) );
  CLKNHSV0 U13947 ( .I(n11959), .ZN(n14807) );
  CLKNHSV0 U13948 ( .I(n11953), .ZN(n14808) );
  CLKNHSV0 U13949 ( .I(n11958), .ZN(n14809) );
  CLKNHSV0 U13950 ( .I(n11958), .ZN(n14810) );
  CLKNHSV0 U13951 ( .I(n11959), .ZN(n14811) );
  CLKNHSV0 U13952 ( .I(n11957), .ZN(n14812) );
  CLKNHSV0 U13953 ( .I(n11955), .ZN(n14813) );
  CLKNHSV0 U13954 ( .I(n11954), .ZN(n14814) );
  CLKNHSV0 U13955 ( .I(n11958), .ZN(n14815) );
  CLKNHSV0 U13956 ( .I(n11958), .ZN(n14816) );
  CLKNHSV0 U13957 ( .I(n11894), .ZN(n14817) );
  NAND2HSV0 U13958 ( .A1(\pe13/aot [1]), .A2(\pe13/bq[3] ), .ZN(n11962) );
  NAND2HSV0 U13959 ( .A1(\pe13/aot [3]), .A2(\pe13/bq[1] ), .ZN(n11961) );
  XOR2HSV0 U13960 ( .A1(n11962), .A2(n11961), .Z(n11963) );
  XNOR2HSV1 U13961 ( .A1(n11963), .A2(n13592), .ZN(n11967) );
  CLKNHSV1 U13962 ( .I(\pe13/got [1]), .ZN(n11964) );
  NAND2HSV2 U13963 ( .A1(n12997), .A2(\pe13/got [2]), .ZN(n11965) );
  XOR3HSV2 U13964 ( .A1(n11967), .A2(n11966), .A3(n11965), .Z(n11971) );
  NOR2HSV2 U13965 ( .A1(n13143), .A2(\pe18/got [8]), .ZN(n12006) );
  CLKNHSV0 U13966 ( .I(n13346), .ZN(n11973) );
  AOI21HSV0 U13967 ( .A1(n13139), .A2(n12006), .B(n11974), .ZN(n11975) );
  NOR2HSV2 U13968 ( .A1(n13139), .A2(n12010), .ZN(n11978) );
  NAND2HSV0 U13969 ( .A1(\pe18/aot [2]), .A2(n14511), .ZN(n13154) );
  CLKNAND2HSV0 U13970 ( .A1(n14513), .A2(\pe18/aot [3]), .ZN(n11980) );
  XOR2HSV0 U13971 ( .A1(n13154), .A2(n11980), .Z(n11995) );
  NAND2HSV0 U13972 ( .A1(\pe18/aot [6]), .A2(\pe18/bq[4] ), .ZN(n11982) );
  CLKNAND2HSV0 U13973 ( .A1(\pe18/got [2]), .A2(n13818), .ZN(n11981) );
  XOR2HSV0 U13974 ( .A1(n11982), .A2(n11981), .Z(n11985) );
  XNOR2HSV1 U13975 ( .A1(n11983), .A2(\pe18/phq [7]), .ZN(n11984) );
  XNOR2HSV1 U13976 ( .A1(n11985), .A2(n11984), .ZN(n11994) );
  NAND2HSV0 U13977 ( .A1(\pe18/aot [5]), .A2(\pe18/bq[5] ), .ZN(n11987) );
  NAND2HSV0 U13978 ( .A1(\pe18/aot [7]), .A2(\pe18/bq[3] ), .ZN(n11986) );
  XOR2HSV0 U13979 ( .A1(n11987), .A2(n11986), .Z(n11992) );
  NAND2HSV0 U13980 ( .A1(\pe18/aot [4]), .A2(\pe18/bq[6] ), .ZN(n11990) );
  NAND2HSV0 U13981 ( .A1(n11988), .A2(\pe18/bq[2] ), .ZN(n11989) );
  XOR2HSV0 U13982 ( .A1(n11990), .A2(n11989), .Z(n11991) );
  XOR2HSV0 U13983 ( .A1(n11992), .A2(n11991), .Z(n11993) );
  XOR3HSV2 U13984 ( .A1(n11995), .A2(n11994), .A3(n11993), .Z(n11998) );
  XNOR2HSV4 U13985 ( .A1(n12000), .A2(n11999), .ZN(n12003) );
  AOI21HSV1 U13986 ( .A1(n13143), .A2(n13142), .B(n13147), .ZN(n12001) );
  OAI21HSV2 U13987 ( .A1(n13140), .A2(n15217), .B(n12001), .ZN(n12002) );
  XNOR2HSV4 U13988 ( .A1(n12003), .A2(n12002), .ZN(n12004) );
  INHSV2 U13989 ( .I(\pe18/ti_7t [7]), .ZN(n12007) );
  OR2HSV1 U13990 ( .A1(n13145), .A2(n12007), .Z(n12008) );
  CLKNAND2HSV4 U13991 ( .A1(n12009), .A2(n12008), .ZN(n13184) );
  AOI21HSV4 U13992 ( .A1(n13185), .A2(n13255), .B(n13184), .ZN(n14682) );
  INHSV4 U13993 ( .I(n12102), .ZN(n12038) );
  NAND2HSV2 U13994 ( .A1(n14740), .A2(n8928), .ZN(n12011) );
  NOR2HSV4 U13995 ( .A1(n12038), .A2(n12011), .ZN(n13873) );
  CLKNAND2HSV1 U13996 ( .A1(n12104), .A2(n12103), .ZN(n13872) );
  NOR2HSV4 U13997 ( .A1(n13873), .A2(n12012), .ZN(n12039) );
  AND2HSV2 U13998 ( .A1(n12015), .A2(n12014), .Z(n12016) );
  OAI21HSV0 U13999 ( .A1(n13268), .A2(\pe17/ti_7t [4]), .B(n14429), .ZN(n12018) );
  NAND2HSV2 U14000 ( .A1(n12109), .A2(\pe17/got [6]), .ZN(n12032) );
  NAND2HSV2 U14001 ( .A1(\pe17/ctrq ), .A2(\pe17/pvq [6]), .ZN(n12023) );
  XNOR2HSV1 U14002 ( .A1(n12023), .A2(\pe17/phq [6]), .ZN(n12026) );
  NAND2HSV0 U14003 ( .A1(\pe17/aot [7]), .A2(\pe17/bq[4] ), .ZN(n12024) );
  NAND2HSV0 U14004 ( .A1(\pe17/aot [6]), .A2(\pe17/bq[5] ), .ZN(n12025) );
  XNOR2HSV4 U14005 ( .A1(n12028), .A2(n12027), .ZN(n12030) );
  NOR2HSV3 U14006 ( .A1(n12037), .A2(n12031), .ZN(n12034) );
  INHSV2 U14007 ( .I(n12032), .ZN(n12035) );
  CLKNAND2HSV3 U14008 ( .A1(n12034), .A2(n12033), .ZN(n12041) );
  NAND4HSV2 U14009 ( .A1(n12039), .A2(n12041), .A3(n12040), .A4(n13874), .ZN(
        n12047) );
  NAND3HSV4 U14010 ( .A1(n13875), .A2(n12044), .A3(n12043), .ZN(n12046) );
  NAND2HSV2 U14011 ( .A1(n13269), .A2(\pe17/ti_7t [6]), .ZN(n12045) );
  CLKNHSV0 U14012 ( .I(\pe4/got [1]), .ZN(n12049) );
  NAND2HSV0 U14013 ( .A1(\pe4/aot [1]), .A2(\pe4/bq[5] ), .ZN(n12051) );
  NAND2HSV0 U14014 ( .A1(\pe4/bq[1] ), .A2(\pe4/aot [5]), .ZN(n12050) );
  XOR2HSV0 U14015 ( .A1(n12051), .A2(n12050), .Z(n12052) );
  NAND2HSV0 U14016 ( .A1(\pe4/aot [3]), .A2(\pe4/bq[3] ), .ZN(n12632) );
  XNOR2HSV1 U14017 ( .A1(n12052), .A2(n12632), .ZN(n12056) );
  NAND2HSV0 U14018 ( .A1(\pe4/aot [2]), .A2(\pe4/bq[4] ), .ZN(n12054) );
  NAND2HSV0 U14019 ( .A1(\pe4/aot [4]), .A2(\pe4/bq[2] ), .ZN(n12053) );
  XOR2HSV0 U14020 ( .A1(n12054), .A2(n12053), .Z(n12055) );
  XNOR2HSV4 U14021 ( .A1(n12058), .A2(n12057), .ZN(n12202) );
  NAND2HSV4 U14022 ( .A1(n12060), .A2(n12059), .ZN(n14860) );
  CLKNAND2HSV0 U14023 ( .A1(\pe7/bq[7] ), .A2(\pe7/aot [6]), .ZN(n12235) );
  NAND2HSV0 U14024 ( .A1(\pe7/got [5]), .A2(\pe7/ti_1 ), .ZN(n12061) );
  XOR2HSV0 U14025 ( .A1(n12235), .A2(n12061), .Z(n12065) );
  NAND2HSV0 U14026 ( .A1(\pe7/bq[6] ), .A2(\pe7/aot [7]), .ZN(n12062) );
  XNOR2HSV2 U14027 ( .A1(n12063), .A2(n12062), .ZN(n12064) );
  XNOR2HSV4 U14028 ( .A1(n12065), .A2(n12064), .ZN(n12071) );
  NAND2HSV0 U14029 ( .A1(\pe7/aot [5]), .A2(\pe7/bq[8] ), .ZN(n12066) );
  CLKXOR2HSV2 U14030 ( .A1(n12066), .A2(\pe7/phq [4]), .Z(n12069) );
  NAND2HSV2 U14031 ( .A1(n12067), .A2(\pe7/pvq [4]), .ZN(n12068) );
  XNOR2HSV4 U14032 ( .A1(n12069), .A2(n12068), .ZN(n12070) );
  XNOR2HSV4 U14033 ( .A1(n12071), .A2(n12070), .ZN(n12076) );
  CLKNAND2HSV0 U14034 ( .A1(n12072), .A2(\pe7/got [6]), .ZN(n12073) );
  NOR2HSV3 U14035 ( .A1(n12074), .A2(n12073), .ZN(n12075) );
  XNOR2HSV4 U14036 ( .A1(n12076), .A2(n12075), .ZN(n12077) );
  CLKNAND2HSV2 U14037 ( .A1(n12232), .A2(\pe7/got [7]), .ZN(n12078) );
  XNOR2HSV4 U14038 ( .A1(n12077), .A2(n12078), .ZN(n12247) );
  NAND3HSV4 U14039 ( .A1(n12248), .A2(n12247), .A3(n8905), .ZN(n12264) );
  BUFHSV2 U14040 ( .I(n12276), .Z(n14823) );
  NAND2HSV2 U14041 ( .A1(n12079), .A2(\pe4/got [1]), .ZN(n12085) );
  CLKNAND2HSV0 U14042 ( .A1(\pe4/aot [3]), .A2(\pe4/bq[1] ), .ZN(n12081) );
  NAND2HSV0 U14043 ( .A1(\pe4/aot [2]), .A2(\pe4/bq[2] ), .ZN(n12080) );
  XOR2HSV0 U14044 ( .A1(n12081), .A2(n12080), .Z(n12083) );
  NAND2HSV0 U14045 ( .A1(\pe4/aot [1]), .A2(\pe4/bq[3] ), .ZN(n12082) );
  XNOR2HSV1 U14046 ( .A1(n12083), .A2(n12082), .ZN(n12084) );
  XNOR2HSV1 U14047 ( .A1(n12085), .A2(n12084), .ZN(n12087) );
  NAND2HSV2 U14048 ( .A1(n7519), .A2(\pe21/got [6]), .ZN(n12099) );
  CLKNAND2HSV1 U14049 ( .A1(\pe21/aot [5]), .A2(\pe21/bq[1] ), .ZN(n12552) );
  CLKNAND2HSV0 U14050 ( .A1(\pe21/bq[5] ), .A2(\pe21/aot [3]), .ZN(n12546) );
  XOR2HSV0 U14051 ( .A1(n12092), .A2(n12546), .Z(n12096) );
  NAND2HSV0 U14052 ( .A1(\pe21/bq[4] ), .A2(\pe21/aot [4]), .ZN(n12094) );
  NAND2HSV0 U14053 ( .A1(\pe21/bq[7] ), .A2(\pe21/aot [1]), .ZN(n12093) );
  XOR2HSV0 U14054 ( .A1(n12094), .A2(n12093), .Z(n12095) );
  XNOR2HSV2 U14055 ( .A1(n12099), .A2(n12098), .ZN(n12101) );
  XOR2HSV2 U14056 ( .A1(n12101), .A2(n12100), .Z(\pe21/poht [1]) );
  NOR2HSV0 U14057 ( .A1(n12103), .A2(n13269), .ZN(n12106) );
  CLKNAND2HSV1 U14058 ( .A1(n12104), .A2(n14429), .ZN(n12105) );
  CLKNAND2HSV0 U14059 ( .A1(n12109), .A2(\pe17/got [5]), .ZN(n12110) );
  NAND2HSV0 U14060 ( .A1(\pe17/aot [5]), .A2(\pe17/bq[5] ), .ZN(n13238) );
  NAND2HSV0 U14061 ( .A1(\pe17/aot [4]), .A2(\pe17/bq[6] ), .ZN(n12112) );
  XOR2HSV0 U14062 ( .A1(n13238), .A2(n12112), .Z(n12126) );
  NAND2HSV0 U14063 ( .A1(\pe17/aot [7]), .A2(\pe17/bq[3] ), .ZN(n12113) );
  XOR2HSV0 U14064 ( .A1(n12114), .A2(n12113), .Z(n12117) );
  NAND2HSV2 U14065 ( .A1(\pe17/ctrq ), .A2(\pe17/pvq [7]), .ZN(n12115) );
  XOR2HSV0 U14066 ( .A1(n12115), .A2(\pe17/phq [7]), .Z(n12116) );
  XNOR2HSV4 U14067 ( .A1(n12117), .A2(n12116), .ZN(n12125) );
  NAND2HSV0 U14068 ( .A1(\pe17/aot [6]), .A2(\pe17/bq[4] ), .ZN(n12118) );
  XOR2HSV0 U14069 ( .A1(n12119), .A2(n12118), .Z(n12123) );
  CLKNAND2HSV0 U14070 ( .A1(n14412), .A2(\pe17/aot [3]), .ZN(n12121) );
  NAND2HSV0 U14071 ( .A1(\pe17/got [2]), .A2(n14415), .ZN(n12120) );
  XOR2HSV0 U14072 ( .A1(n12121), .A2(n12120), .Z(n12122) );
  XOR3HSV2 U14073 ( .A1(n12126), .A2(n12125), .A3(n12124), .Z(n12128) );
  INHSV2 U14074 ( .I(\pe17/got [3]), .ZN(n14309) );
  NOR2HSV2 U14075 ( .A1(n14401), .A2(n14309), .ZN(n12127) );
  CLKNAND2HSV0 U14076 ( .A1(n14399), .A2(\pe17/got [4]), .ZN(n12129) );
  INHSV2 U14077 ( .I(\pe17/got [6]), .ZN(n14008) );
  INAND2HSV0 U14078 ( .A1(n12135), .B1(n9541), .ZN(n12136) );
  INHSV2 U14079 ( .I(n12136), .ZN(n12137) );
  NOR2HSV1 U14080 ( .A1(n12140), .A2(n12143), .ZN(n12142) );
  CLKNAND2HSV1 U14081 ( .A1(n12142), .A2(n12141), .ZN(n12147) );
  CLKNHSV0 U14082 ( .I(n12143), .ZN(n12145) );
  NOR2HSV1 U14083 ( .A1(n12143), .A2(n9541), .ZN(n12144) );
  NAND2HSV0 U14084 ( .A1(\pe19/ti_7[1] ), .A2(\pe19/got [3]), .ZN(n12167) );
  NAND2HSV0 U14085 ( .A1(\pe19/aot [6]), .A2(\pe19/bq[4] ), .ZN(n12150) );
  NAND2HSV0 U14086 ( .A1(\pe19/aot [2]), .A2(n14506), .ZN(n12149) );
  XOR2HSV0 U14087 ( .A1(n12150), .A2(n12149), .Z(n12164) );
  NAND2HSV2 U14088 ( .A1(n14501), .A2(\pe19/pvq [7]), .ZN(n12151) );
  XOR2HSV0 U14089 ( .A1(n12151), .A2(\pe19/phq [7]), .Z(n12154) );
  CLKNAND2HSV1 U14090 ( .A1(n13317), .A2(\pe19/bq[2] ), .ZN(n14224) );
  XNOR2HSV1 U14091 ( .A1(n12154), .A2(n12153), .ZN(n12163) );
  CLKNHSV0 U14092 ( .I(\pe19/ti_1 ), .ZN(n12155) );
  NAND2HSV0 U14093 ( .A1(\pe19/got [2]), .A2(n13821), .ZN(n12157) );
  NAND2HSV0 U14094 ( .A1(n14945), .A2(\pe19/bq[3] ), .ZN(n12156) );
  XOR2HSV0 U14095 ( .A1(n12157), .A2(n12156), .Z(n12161) );
  CLKNAND2HSV0 U14096 ( .A1(n14576), .A2(\pe19/aot [3]), .ZN(n12159) );
  NAND2HSV0 U14097 ( .A1(\pe19/aot [4]), .A2(\pe19/bq[6] ), .ZN(n12158) );
  XOR2HSV0 U14098 ( .A1(n12159), .A2(n12158), .Z(n12160) );
  XOR2HSV0 U14099 ( .A1(n12161), .A2(n12160), .Z(n12162) );
  XOR3HSV2 U14100 ( .A1(n12164), .A2(n12163), .A3(n12162), .Z(n12165) );
  XOR3HSV2 U14101 ( .A1(n12167), .A2(n12166), .A3(n12165), .Z(n12168) );
  INHSV2 U14102 ( .I(\pe19/ti_7t [7]), .ZN(n12170) );
  NOR2HSV2 U14103 ( .A1(n9541), .A2(n12170), .ZN(n12171) );
  NAND2HSV2 U14104 ( .A1(n14862), .A2(\pe19/got [4]), .ZN(n12181) );
  NAND2HSV2 U14105 ( .A1(n12172), .A2(\pe19/ti_7t [6]), .ZN(n12340) );
  NAND2HSV0 U14106 ( .A1(n14219), .A2(\pe19/got [1]), .ZN(n12180) );
  NAND2HSV0 U14107 ( .A1(\pe19/aot [2]), .A2(\pe19/bq[3] ), .ZN(n12174) );
  NAND2HSV0 U14108 ( .A1(\pe19/aot [1]), .A2(\pe19/bq[4] ), .ZN(n12173) );
  XOR2HSV0 U14109 ( .A1(n12174), .A2(n12173), .Z(n12178) );
  NAND2HSV0 U14110 ( .A1(\pe19/aot [3]), .A2(\pe19/bq[2] ), .ZN(n12176) );
  NAND2HSV0 U14111 ( .A1(\pe19/bq[1] ), .A2(\pe19/aot [4]), .ZN(n12175) );
  XOR2HSV0 U14112 ( .A1(n12176), .A2(n12175), .Z(n12177) );
  XOR2HSV0 U14113 ( .A1(n12178), .A2(n12177), .Z(n12179) );
  NAND2HSV0 U14114 ( .A1(n12181), .A2(n12182), .ZN(n12186) );
  CLKNHSV2 U14115 ( .I(n12181), .ZN(n12184) );
  CLKNAND2HSV1 U14116 ( .A1(n12184), .A2(n12183), .ZN(n12185) );
  NAND2HSV0 U14117 ( .A1(n12186), .A2(n12185), .ZN(\pe19/poht [4]) );
  INHSV1 U14118 ( .I(bo10[3]), .ZN(n12189) );
  MUX2NHSV1 U14119 ( .I0(n12189), .I1(n12188), .S(n14554), .ZN(n15031) );
  CLKNHSV0 U14120 ( .I(bo4[2]), .ZN(n12191) );
  MUX2NHSV1 U14121 ( .I0(n12191), .I1(n12190), .S(n13822), .ZN(n15040) );
  NAND2HSV4 U14122 ( .A1(n12193), .A2(n12192), .ZN(n14830) );
  CLKNAND2HSV1 U14123 ( .A1(\pe16/ti_7[1] ), .A2(n12194), .ZN(n12197) );
  INHSV2 U14124 ( .I(n10682), .ZN(n12196) );
  XNOR2HSV1 U14125 ( .A1(n12197), .A2(n12196), .ZN(n15230) );
  NAND2HSV2 U14126 ( .A1(ctro7), .A2(\pe7/ti_7t [4]), .ZN(n12277) );
  BUFHSV2 U14127 ( .I(n12277), .Z(n12263) );
  CLKNAND2HSV2 U14128 ( .A1(n12265), .A2(n12263), .ZN(n12200) );
  INHSV2 U14129 ( .I(\pe7/got [7]), .ZN(n12274) );
  AOI21HSV1 U14130 ( .A1(n12277), .A2(n12311), .B(n12274), .ZN(n12198) );
  NAND3HSV2 U14131 ( .A1(n12201), .A2(n12202), .A3(n12252), .ZN(n12230) );
  INHSV2 U14132 ( .I(n12230), .ZN(n12225) );
  INHSV2 U14133 ( .I(n12203), .ZN(n12205) );
  INHSV1 U14134 ( .I(n12206), .ZN(n12228) );
  CLKNHSV0 U14135 ( .I(\pe7/got [6]), .ZN(n12207) );
  NOR2HSV1 U14136 ( .A1(n12228), .A2(n12207), .ZN(n12208) );
  NOR2HSV1 U14137 ( .A1(n12225), .A2(n12223), .ZN(n12224) );
  NAND2HSV0 U14138 ( .A1(\pe7/ti_7[1] ), .A2(\pe7/got [4]), .ZN(n12222) );
  NAND2HSV0 U14139 ( .A1(\pe7/aot [6]), .A2(\pe7/bq[5] ), .ZN(n12210) );
  NAND2HSV0 U14140 ( .A1(\pe7/got [3]), .A2(\pe7/ti_1 ), .ZN(n12209) );
  XOR2HSV0 U14141 ( .A1(n12210), .A2(n12209), .Z(n12219) );
  NAND2HSV0 U14142 ( .A1(\pe7/aot [8]), .A2(\pe7/bq[3] ), .ZN(n12212) );
  NAND2HSV0 U14143 ( .A1(\pe7/aot [7]), .A2(\pe7/bq[4] ), .ZN(n12211) );
  XOR2HSV0 U14144 ( .A1(n12212), .A2(n12211), .Z(n12216) );
  NAND2HSV0 U14145 ( .A1(\pe7/aot [4]), .A2(\pe7/bq[7] ), .ZN(n12214) );
  NAND2HSV0 U14146 ( .A1(\pe7/aot [3]), .A2(\pe7/bq[8] ), .ZN(n12213) );
  XOR2HSV0 U14147 ( .A1(n12214), .A2(n12213), .Z(n12215) );
  XOR2HSV2 U14148 ( .A1(n12216), .A2(n12215), .Z(n12217) );
  XOR3HSV2 U14149 ( .A1(n12219), .A2(n12218), .A3(n12217), .Z(n12221) );
  NAND2HSV0 U14150 ( .A1(n14860), .A2(\pe7/got [5]), .ZN(n12220) );
  NAND2HSV2 U14151 ( .A1(n8902), .A2(n12225), .ZN(n12226) );
  NOR2HSV1 U14152 ( .A1(n12228), .A2(n12274), .ZN(n12229) );
  NAND2HSV0 U14153 ( .A1(n12232), .A2(\pe7/got [6]), .ZN(n12245) );
  NAND2HSV0 U14154 ( .A1(\pe7/ctrq ), .A2(\pe7/pvq [5]), .ZN(n12233) );
  XNOR2HSV1 U14155 ( .A1(n12233), .A2(\pe7/phq [5]), .ZN(n12239) );
  NOR2HSV1 U14156 ( .A1(n12235), .A2(n12234), .ZN(n12237) );
  AOI22HSV0 U14157 ( .A1(\pe7/aot [6]), .A2(\pe7/bq[6] ), .B1(\pe7/aot [5]), 
        .B2(\pe7/bq[7] ), .ZN(n12236) );
  NOR2HSV2 U14158 ( .A1(n12237), .A2(n12236), .ZN(n12238) );
  XNOR2HSV1 U14159 ( .A1(n12239), .A2(n12238), .ZN(n12240) );
  XNOR2HSV4 U14160 ( .A1(n12243), .A2(n12242), .ZN(n12244) );
  AOI21HSV0 U14161 ( .A1(n12248), .A2(n12247), .B(n12309), .ZN(n12249) );
  CLKNAND2HSV0 U14162 ( .A1(n12249), .A2(n12265), .ZN(n12250) );
  CLKAND2HSV2 U14163 ( .A1(n12309), .A2(\pe7/ti_7t [6]), .Z(n12254) );
  AOI31HSV2 U14164 ( .A1(n13882), .A2(n12255), .A3(n12256), .B(n12254), .ZN(
        n12259) );
  CLKNHSV0 U14165 ( .I(n12260), .ZN(n14927) );
  CLKNHSV0 U14166 ( .I(bo10[4]), .ZN(n12262) );
  CLKNHSV0 U14167 ( .I(\pe10/bq[4] ), .ZN(n12261) );
  MUX2NHSV1 U14168 ( .I0(n12262), .I1(n12261), .S(n14554), .ZN(n15030) );
  CLKNHSV2 U14169 ( .I(n12265), .ZN(n12269) );
  AOI21HSV1 U14170 ( .A1(n12267), .A2(n12277), .B(n12266), .ZN(n12268) );
  OAI21HSV4 U14171 ( .A1(n12270), .A2(n12269), .B(n12268), .ZN(n13621) );
  NAND2HSV2 U14172 ( .A1(n12311), .A2(\pe7/ti_7t [5]), .ZN(n13620) );
  CLKNHSV0 U14173 ( .I(n12271), .ZN(n14902) );
  AND2HSV2 U14174 ( .A1(n15189), .A2(n12273), .Z(n12307) );
  INHSV1 U14175 ( .I(n13620), .ZN(n13623) );
  INOR2HSV1 U14176 ( .A1(n13620), .B1(n12308), .ZN(n13627) );
  NOR2HSV2 U14177 ( .A1(n13627), .A2(n12274), .ZN(n12275) );
  OAI21HSV4 U14178 ( .A1(\pov7[5] ), .A2(n13623), .B(n12275), .ZN(n12306) );
  INHSV2 U14179 ( .I(\pe7/got [5]), .ZN(n12279) );
  INAND2HSV0 U14180 ( .A1(n12279), .B1(n12308), .ZN(n12278) );
  CLKNHSV0 U14181 ( .I(n12278), .ZN(n12282) );
  OR2HSV1 U14182 ( .A1(n12280), .A2(n12279), .Z(n12281) );
  IOA21HSV2 U14183 ( .A1(n15271), .A2(n12282), .B(n12281), .ZN(n12303) );
  NAND2HSV2 U14184 ( .A1(n14860), .A2(\pe7/got [4]), .ZN(n12284) );
  NAND2HSV0 U14185 ( .A1(\pe7/ti_7[1] ), .A2(\pe7/got [3]), .ZN(n12283) );
  XNOR2HSV1 U14186 ( .A1(n12284), .A2(n12283), .ZN(n12301) );
  NAND2HSV0 U14187 ( .A1(\pe7/bq[3] ), .A2(\pe7/aot [7]), .ZN(n13609) );
  NAND2HSV0 U14188 ( .A1(\pe7/bq[2] ), .A2(\pe7/aot [8]), .ZN(n12285) );
  XOR2HSV0 U14189 ( .A1(n13609), .A2(n12285), .Z(n12299) );
  NAND2HSV0 U14190 ( .A1(\pe7/aot [4]), .A2(\pe7/bq[6] ), .ZN(n12287) );
  NAND2HSV0 U14191 ( .A1(\pe7/aot [6]), .A2(\pe7/bq[4] ), .ZN(n12286) );
  XOR2HSV0 U14192 ( .A1(n12287), .A2(n12286), .Z(n12290) );
  NAND2HSV2 U14193 ( .A1(n12067), .A2(\pe7/pvq [7]), .ZN(n12288) );
  XNOR2HSV1 U14194 ( .A1(n12288), .A2(\pe7/phq [7]), .ZN(n12289) );
  XNOR2HSV1 U14195 ( .A1(n12290), .A2(n12289), .ZN(n12298) );
  NAND2HSV0 U14196 ( .A1(\pe7/aot [2]), .A2(\pe7/bq[8] ), .ZN(n12292) );
  NAND2HSV0 U14197 ( .A1(\pe7/aot [3]), .A2(\pe7/bq[7] ), .ZN(n12291) );
  XOR2HSV0 U14198 ( .A1(n12292), .A2(n12291), .Z(n12296) );
  CLKNAND2HSV0 U14199 ( .A1(\pe7/aot [5]), .A2(\pe7/bq[5] ), .ZN(n12294) );
  NAND2HSV0 U14200 ( .A1(\pe7/got [2]), .A2(n14480), .ZN(n12293) );
  XOR2HSV0 U14201 ( .A1(n12294), .A2(n12293), .Z(n12295) );
  XOR2HSV0 U14202 ( .A1(n12296), .A2(n12295), .Z(n12297) );
  XOR3HSV2 U14203 ( .A1(n12299), .A2(n12298), .A3(n12297), .Z(n12300) );
  XNOR2HSV1 U14204 ( .A1(n12301), .A2(n12300), .ZN(n12302) );
  XOR2HSV0 U14205 ( .A1(n12303), .A2(n12302), .Z(n12304) );
  BUFHSV8 U14206 ( .I(n12310), .Z(n14055) );
  CLKNAND2HSV3 U14207 ( .A1(n12307), .A2(n14055), .ZN(n12941) );
  INHSV2 U14208 ( .I(n14054), .ZN(n14049) );
  OAI21HSV4 U14209 ( .A1(n12310), .A2(n12309), .B(n14049), .ZN(n12315) );
  INAND2HSV2 U14210 ( .A1(n14054), .B1(n8921), .ZN(n12312) );
  INHSV2 U14211 ( .I(n12312), .ZN(n12313) );
  CLKNAND2HSV3 U14212 ( .A1(n14487), .A2(n12313), .ZN(n12314) );
  CLKNAND2HSV4 U14213 ( .A1(n12315), .A2(n12314), .ZN(n12940) );
  NAND2HSV2 U14214 ( .A1(n12941), .A2(n12940), .ZN(n14852) );
  NAND2HSV2 U14215 ( .A1(n14189), .A2(\pe8/ti_7t [7]), .ZN(n12371) );
  NOR2HSV2 U14216 ( .A1(n12318), .A2(n12317), .ZN(n12319) );
  NAND2HSV0 U14217 ( .A1(n15072), .A2(\pe15/got [3]), .ZN(n12334) );
  NAND2HSV2 U14218 ( .A1(n14735), .A2(\pe15/got [4]), .ZN(n12333) );
  NAND2HSV0 U14219 ( .A1(\pe15/aot [4]), .A2(\pe15/bq[6] ), .ZN(n12322) );
  NAND2HSV0 U14220 ( .A1(n14936), .A2(\pe15/bq[3] ), .ZN(n12321) );
  XOR2HSV0 U14221 ( .A1(n12322), .A2(n12321), .Z(n12331) );
  BUFHSV2 U14222 ( .I(\pe15/ti_1 ), .Z(n14587) );
  NAND2HSV0 U14223 ( .A1(n14937), .A2(\pe15/bq[2] ), .ZN(n12324) );
  NAND2HSV0 U14224 ( .A1(\pe15/aot [5]), .A2(\pe15/bq[5] ), .ZN(n12323) );
  XOR2HSV0 U14225 ( .A1(n12324), .A2(n12323), .Z(n12328) );
  NAND2HSV0 U14226 ( .A1(\pe15/aot [6]), .A2(\pe15/bq[4] ), .ZN(n12326) );
  NAND2HSV0 U14227 ( .A1(\pe15/aot [3]), .A2(\pe15/bq[7] ), .ZN(n12325) );
  XOR2HSV0 U14228 ( .A1(n12326), .A2(n12325), .Z(n12327) );
  XOR2HSV0 U14229 ( .A1(n12328), .A2(n12327), .Z(n12329) );
  XOR3HSV2 U14230 ( .A1(n12331), .A2(n12330), .A3(n12329), .Z(n12332) );
  INHSV2 U14231 ( .I(\pe15/got [5]), .ZN(n12513) );
  CLKNHSV0 U14232 ( .I(n12135), .ZN(n14859) );
  CLKNHSV0 U14233 ( .I(bo10[1]), .ZN(n12339) );
  MUX2NHSV1 U14234 ( .I0(n12339), .I1(n12338), .S(n14554), .ZN(n15033) );
  CLKNHSV0 U14235 ( .I(bo5[1]), .ZN(n12342) );
  CLKNHSV0 U14236 ( .I(\pe5/bq[1] ), .ZN(n12341) );
  MUX2NHSV1 U14237 ( .I0(n12342), .I1(n12341), .S(n11818), .ZN(n15039) );
  INHSV1 U14238 ( .I(bo15[2]), .ZN(n12345) );
  MUX2NHSV1 U14239 ( .I0(n12345), .I1(n12344), .S(n14586), .ZN(n15023) );
  CLKNHSV0 U14240 ( .I(n12346), .ZN(n14871) );
  INHSV1 U14241 ( .I(\pe11/ti_7t [5]), .ZN(n12349) );
  NAND2HSV2 U14242 ( .A1(n9609), .A2(n12349), .ZN(n12350) );
  OAI21HSV4 U14243 ( .A1(n15256), .A2(n15090), .B(n12350), .ZN(n14396) );
  CLKNHSV0 U14244 ( .I(n14396), .ZN(\pe11/ti_7[5] ) );
  CLKNHSV0 U14245 ( .I(n12351), .ZN(n14900) );
  CLKNHSV0 U14246 ( .I(n12352), .ZN(n14909) );
  CLKNHSV0 U14247 ( .I(bo3[3]), .ZN(n12356) );
  MUX2NHSV1 U14248 ( .I0(n12356), .I1(n12355), .S(n10979), .ZN(n15045) );
  CLKNHSV0 U14249 ( .I(bo3[4]), .ZN(n12359) );
  CLKNHSV0 U14250 ( .I(\pe3/bq[4] ), .ZN(n12358) );
  MUX2NHSV1 U14251 ( .I0(n12359), .I1(n12358), .S(n12357), .ZN(n15044) );
  CLKNHSV0 U14252 ( .I(bo3[7]), .ZN(n12361) );
  CLKNHSV0 U14253 ( .I(\pe3/bq[7] ), .ZN(n12360) );
  MUX2NHSV1 U14254 ( .I0(n12361), .I1(n12360), .S(n10979), .ZN(n15042) );
  INHSV1 U14255 ( .I(bo20[5]), .ZN(n12364) );
  CLKNHSV0 U14256 ( .I(\pe20/bq[5] ), .ZN(n12363) );
  MUX2NHSV1 U14257 ( .I0(n12364), .I1(n12363), .S(n12362), .ZN(n15011) );
  INHSV2 U14258 ( .I(bo20[2]), .ZN(n12366) );
  CLKNHSV0 U14259 ( .I(\pe20/bq[2] ), .ZN(n12365) );
  MUX2NHSV1 U14260 ( .I0(n12366), .I1(n12365), .S(n12362), .ZN(n15012) );
  INHSV2 U14261 ( .I(bo20[6]), .ZN(n12368) );
  CLKNHSV0 U14262 ( .I(\pe20/bq[6] ), .ZN(n12367) );
  MUX2NHSV1 U14263 ( .I0(n12368), .I1(n12367), .S(n12362), .ZN(n15010) );
  INHSV2 U14264 ( .I(ao4[8]), .ZN(n14878) );
  INHSV2 U14265 ( .I(go5[8]), .ZN(n14882) );
  INHSV2 U14266 ( .I(ao5[6]), .ZN(n14883) );
  CLKNHSV0 U14267 ( .I(n12369), .ZN(n14886) );
  INHSV2 U14268 ( .I(ao2[8]), .ZN(n14888) );
  CLKNHSV0 U14269 ( .I(n12371), .ZN(n12374) );
  CLKNHSV0 U14270 ( .I(\pe8/got [2]), .ZN(n12370) );
  AOI21HSV1 U14271 ( .A1(n12372), .A2(n12371), .B(n12370), .ZN(n12373) );
  CLKNAND2HSV1 U14272 ( .A1(\pe8/aot [1]), .A2(\pe8/bq[2] ), .ZN(n12376) );
  NAND2HSV0 U14273 ( .A1(\pe8/aot [2]), .A2(\pe8/bq[1] ), .ZN(n12375) );
  XNOR2HSV1 U14274 ( .A1(n12376), .A2(n12375), .ZN(n12377) );
  NAND2HSV0 U14275 ( .A1(\pe19/aot [2]), .A2(\pe19/bq[4] ), .ZN(n12384) );
  NAND2HSV0 U14276 ( .A1(n13317), .A2(\pe19/bq[1] ), .ZN(n12379) );
  NAND2HSV0 U14277 ( .A1(\pe19/bq[2] ), .A2(\pe19/aot [4]), .ZN(n12378) );
  XOR2HSV0 U14278 ( .A1(n12379), .A2(n12378), .Z(n12383) );
  NAND2HSV0 U14279 ( .A1(\pe19/aot [3]), .A2(\pe19/bq[3] ), .ZN(n12381) );
  NAND2HSV0 U14280 ( .A1(\pe19/aot [1]), .A2(\pe19/bq[5] ), .ZN(n12380) );
  XOR2HSV0 U14281 ( .A1(n12381), .A2(n12380), .Z(n12382) );
  CLKNAND2HSV1 U14282 ( .A1(n11777), .A2(\pe19/got [3]), .ZN(n12389) );
  NAND2HSV0 U14283 ( .A1(\pe19/ti_7[1] ), .A2(\pe19/got [2]), .ZN(n12388) );
  XNOR2HSV1 U14284 ( .A1(n12389), .A2(n12388), .ZN(n12409) );
  CLKNAND2HSV0 U14285 ( .A1(n14501), .A2(\pe19/pq ), .ZN(n12391) );
  NAND2HSV0 U14286 ( .A1(\pe19/got [1]), .A2(n13821), .ZN(n12390) );
  XOR2HSV0 U14287 ( .A1(n12391), .A2(n12390), .Z(n12395) );
  NAND2HSV0 U14288 ( .A1(\pe19/aot [6]), .A2(\pe19/bq[3] ), .ZN(n12393) );
  NAND2HSV0 U14289 ( .A1(n14945), .A2(\pe19/bq[2] ), .ZN(n12392) );
  XOR2HSV0 U14290 ( .A1(n12393), .A2(n12392), .Z(n12394) );
  XOR2HSV0 U14291 ( .A1(n12395), .A2(n12394), .Z(n12399) );
  NAND2HSV0 U14292 ( .A1(n14506), .A2(\pe19/aot [1]), .ZN(n12397) );
  NAND2HSV0 U14293 ( .A1(\pe19/bq[7] ), .A2(\pe19/aot [2]), .ZN(n12396) );
  XOR2HSV0 U14294 ( .A1(n12397), .A2(n12396), .Z(n12398) );
  XNOR2HSV1 U14295 ( .A1(n12399), .A2(n12398), .ZN(n12407) );
  NAND2HSV0 U14296 ( .A1(\pe19/aot [3]), .A2(\pe19/bq[6] ), .ZN(n12401) );
  NAND2HSV0 U14297 ( .A1(n13317), .A2(\pe19/bq[4] ), .ZN(n12400) );
  XOR2HSV0 U14298 ( .A1(n12401), .A2(n12400), .Z(n12405) );
  NAND2HSV0 U14299 ( .A1(n14915), .A2(\pe19/bq[1] ), .ZN(n12403) );
  NAND2HSV0 U14300 ( .A1(\pe19/aot [4]), .A2(\pe19/bq[5] ), .ZN(n12402) );
  XOR2HSV0 U14301 ( .A1(n12403), .A2(n12402), .Z(n12404) );
  XOR2HSV0 U14302 ( .A1(n12405), .A2(n12404), .Z(n12406) );
  XNOR2HSV1 U14303 ( .A1(n12407), .A2(n12406), .ZN(n12408) );
  NAND2HSV0 U14304 ( .A1(\pe6/aot [3]), .A2(\pe6/bq[5] ), .ZN(n12413) );
  NAND2HSV0 U14305 ( .A1(\pe6/aot [2]), .A2(\pe6/bq[6] ), .ZN(n12412) );
  NAND2HSV0 U14306 ( .A1(\pe6/aot [7]), .A2(\pe6/bq[1] ), .ZN(n12415) );
  NAND2HSV0 U14307 ( .A1(\pe6/aot [6]), .A2(\pe6/bq[2] ), .ZN(n12414) );
  NOR2HSV0 U14308 ( .A1(n12416), .A2(n13000), .ZN(n12417) );
  NAND2HSV0 U14309 ( .A1(n13057), .A2(\pe6/got [3]), .ZN(n12419) );
  XOR2HSV2 U14310 ( .A1(n12420), .A2(n12419), .Z(n12422) );
  NAND2HSV0 U14311 ( .A1(n15077), .A2(\pe6/got [4]), .ZN(n12421) );
  XNOR2HSV1 U14312 ( .A1(n12422), .A2(n12421), .ZN(n12423) );
  NAND2HSV0 U14313 ( .A1(n14366), .A2(\pe11/got [4]), .ZN(n12446) );
  NAND2HSV0 U14314 ( .A1(\pe11/aot [6]), .A2(\pe11/bq[3] ), .ZN(n12426) );
  NAND2HSV0 U14315 ( .A1(n12424), .A2(\pe11/bq[1] ), .ZN(n12425) );
  XOR2HSV0 U14316 ( .A1(n12426), .A2(n12425), .Z(n12442) );
  CLKNAND2HSV0 U14317 ( .A1(n14553), .A2(\pe11/pq ), .ZN(n12428) );
  NAND2HSV0 U14318 ( .A1(n14837), .A2(\pe11/bq[2] ), .ZN(n12427) );
  XOR2HSV0 U14319 ( .A1(n12428), .A2(n12427), .Z(n12433) );
  CLKNAND2HSV0 U14320 ( .A1(\pe11/aot [1]), .A2(n14519), .ZN(n14375) );
  NOR2HSV0 U14321 ( .A1(n14375), .A2(n12429), .ZN(n12431) );
  AOI22HSV0 U14322 ( .A1(n14519), .A2(\pe11/aot [2]), .B1(n11924), .B2(
        \pe11/aot [1]), .ZN(n12430) );
  NOR2HSV2 U14323 ( .A1(n12431), .A2(n12430), .ZN(n12432) );
  XNOR2HSV1 U14324 ( .A1(n12433), .A2(n12432), .ZN(n12441) );
  NAND2HSV0 U14325 ( .A1(\pe11/aot [5]), .A2(\pe11/bq[4] ), .ZN(n12435) );
  NAND2HSV0 U14326 ( .A1(\pe11/aot [4]), .A2(\pe11/bq[5] ), .ZN(n12434) );
  XOR2HSV0 U14327 ( .A1(n12435), .A2(n12434), .Z(n12439) );
  NAND2HSV0 U14328 ( .A1(n12562), .A2(\pe11/aot [3]), .ZN(n12437) );
  NAND2HSV0 U14329 ( .A1(\pe11/got [1]), .A2(n13811), .ZN(n12436) );
  XOR2HSV0 U14330 ( .A1(n12437), .A2(n12436), .Z(n12438) );
  XOR2HSV0 U14331 ( .A1(n12439), .A2(n12438), .Z(n12440) );
  XOR3HSV2 U14332 ( .A1(n12442), .A2(n12441), .A3(n12440), .Z(n12443) );
  XNOR2HSV1 U14333 ( .A1(n12444), .A2(n12443), .ZN(n12445) );
  XOR2HSV0 U14334 ( .A1(n12446), .A2(n12445), .Z(n12447) );
  NAND2HSV0 U14335 ( .A1(n14830), .A2(\pe11/got [7]), .ZN(n12450) );
  NAND2HSV2 U14336 ( .A1(n14366), .A2(\pe11/got [1]), .ZN(n12463) );
  AND2HSV2 U14337 ( .A1(\pe11/aot [1]), .A2(\pe11/bq[5] ), .Z(n12563) );
  NAND2HSV0 U14338 ( .A1(\pe11/bq[2] ), .A2(\pe11/aot [4]), .ZN(n12457) );
  NAND2HSV0 U14339 ( .A1(\pe11/aot [3]), .A2(\pe11/bq[3] ), .ZN(n12456) );
  XOR2HSV0 U14340 ( .A1(n12457), .A2(n12456), .Z(n12461) );
  NAND2HSV0 U14341 ( .A1(\pe11/aot [5]), .A2(\pe11/bq[1] ), .ZN(n12459) );
  NAND2HSV0 U14342 ( .A1(\pe11/aot [2]), .A2(\pe11/bq[4] ), .ZN(n12458) );
  XOR2HSV0 U14343 ( .A1(n12459), .A2(n12458), .Z(n12460) );
  XOR3HSV2 U14344 ( .A1(n12563), .A2(n12461), .A3(n12460), .Z(n12462) );
  AOI21HSV0 U14345 ( .A1(\pe11/got [2]), .A2(n14365), .B(n12465), .ZN(n12464)
         );
  AOI31HSV0 U14346 ( .A1(\pe11/got [2]), .A2(n12465), .A3(n14737), .B(n12464), 
        .ZN(n12466) );
  XNOR2HSV4 U14347 ( .A1(n12467), .A2(n12466), .ZN(n12469) );
  NAND2HSV0 U14348 ( .A1(\pe11/got [4]), .A2(n14830), .ZN(n12468) );
  NAND2HSV0 U14349 ( .A1(\pe3/got [3]), .A2(n14872), .ZN(n12473) );
  NAND2HSV0 U14350 ( .A1(n5949), .A2(\pe3/got [2]), .ZN(n12472) );
  XNOR2HSV1 U14351 ( .A1(n12473), .A2(n12472), .ZN(n12492) );
  CLKNAND2HSV0 U14352 ( .A1(n12476), .A2(\pe3/aot [1]), .ZN(n12478) );
  NAND2HSV0 U14353 ( .A1(\pe3/aot [2]), .A2(\pe3/bq[7] ), .ZN(n12477) );
  XOR2HSV0 U14354 ( .A1(n12478), .A2(n12477), .Z(n12479) );
  XOR2HSV0 U14355 ( .A1(n12480), .A2(n12479), .Z(n12484) );
  NAND2HSV0 U14356 ( .A1(\pe3/aot [3]), .A2(\pe3/bq[6] ), .ZN(n12482) );
  NAND2HSV0 U14357 ( .A1(\pe3/aot [4]), .A2(\pe3/bq[5] ), .ZN(n12481) );
  XOR2HSV0 U14358 ( .A1(n12482), .A2(n12481), .Z(n12483) );
  NAND2HSV0 U14359 ( .A1(n14738), .A2(\pe3/bq[2] ), .ZN(n12486) );
  NAND2HSV0 U14360 ( .A1(\pe3/aot [5]), .A2(\pe3/bq[4] ), .ZN(n12485) );
  XOR2HSV0 U14361 ( .A1(n12486), .A2(n12485), .Z(n12490) );
  NAND2HSV0 U14362 ( .A1(n14953), .A2(\pe3/bq[1] ), .ZN(n12488) );
  NAND2HSV0 U14363 ( .A1(\pe3/aot [6]), .A2(\pe3/bq[3] ), .ZN(n12487) );
  XOR2HSV0 U14364 ( .A1(n12488), .A2(n12487), .Z(n12489) );
  XOR2HSV0 U14365 ( .A1(n12490), .A2(n12489), .Z(n12491) );
  XOR2HSV0 U14366 ( .A1(n12495), .A2(n12494), .Z(n12496) );
  INHSV2 U14367 ( .I(\pe3/ti_7[5] ), .ZN(n12959) );
  CLKNHSV0 U14368 ( .I(\pe3/got [6]), .ZN(n12497) );
  OR2HSV1 U14369 ( .A1(n12959), .A2(n12497), .Z(n12498) );
  XNOR2HSV4 U14370 ( .A1(n12505), .A2(n12504), .ZN(po3) );
  CLKBUFHSV4 U14371 ( .I(n12879), .Z(n13761) );
  INHSV2 U14372 ( .I(\pe2/got [2]), .ZN(n13100) );
  CLKNAND2HSV0 U14373 ( .A1(n14934), .A2(\pe2/got [1]), .ZN(n12510) );
  NAND2HSV0 U14374 ( .A1(\pe2/aot [5]), .A2(\pe2/bq[1] ), .ZN(n13098) );
  NAND2HSV0 U14375 ( .A1(n14741), .A2(\pe2/bq[2] ), .ZN(n12880) );
  CLKNAND2HSV1 U14376 ( .A1(n6535), .A2(\pe15/got [6]), .ZN(n12541) );
  NOR2HSV3 U14377 ( .A1(n14585), .A2(n12513), .ZN(n12536) );
  NAND2HSV0 U14378 ( .A1(\pe15/aot [3]), .A2(n12616), .ZN(n12516) );
  NAND2HSV0 U14379 ( .A1(n14936), .A2(\pe15/bq[1] ), .ZN(n12515) );
  XOR2HSV0 U14380 ( .A1(n12516), .A2(n12515), .Z(n12520) );
  NAND2HSV0 U14381 ( .A1(\pe15/aot [5]), .A2(\pe15/bq[3] ), .ZN(n12518) );
  NAND2HSV0 U14382 ( .A1(\pe15/aot [6]), .A2(\pe15/bq[2] ), .ZN(n12517) );
  XNOR2HSV1 U14383 ( .A1(n12518), .A2(n12517), .ZN(n12519) );
  XNOR2HSV1 U14384 ( .A1(n12520), .A2(n12519), .ZN(n12522) );
  AOI21HSV0 U14385 ( .A1(n5946), .A2(\pe15/got [2]), .B(n12522), .ZN(n12521)
         );
  AOI31HSV1 U14386 ( .A1(\pe15/got [2]), .A2(n12522), .A3(n5946), .B(n12521), 
        .ZN(n12530) );
  CLKNAND2HSV0 U14387 ( .A1(n15072), .A2(\pe15/got [1]), .ZN(n12528) );
  NAND2HSV0 U14388 ( .A1(\pe15/aot [1]), .A2(\pe15/bq[7] ), .ZN(n12524) );
  NAND2HSV0 U14389 ( .A1(\pe15/aot [4]), .A2(\pe15/bq[4] ), .ZN(n12523) );
  XOR2HSV0 U14390 ( .A1(n12524), .A2(n12523), .Z(n12526) );
  NAND2HSV0 U14391 ( .A1(\pe15/aot [2]), .A2(\pe15/bq[6] ), .ZN(n12525) );
  XNOR2HSV1 U14392 ( .A1(n12526), .A2(n12525), .ZN(n12527) );
  XNOR2HSV1 U14393 ( .A1(n12528), .A2(n12527), .ZN(n12529) );
  XOR2HSV0 U14394 ( .A1(n12530), .A2(n12529), .Z(n12531) );
  XNOR2HSV1 U14395 ( .A1(n12532), .A2(n12531), .ZN(n12534) );
  NAND2HSV0 U14396 ( .A1(\pe15/ti_7[3] ), .A2(\pe15/got [3]), .ZN(n12533) );
  XNOR2HSV1 U14397 ( .A1(n12534), .A2(n12533), .ZN(n12535) );
  XOR2HSV2 U14398 ( .A1(n12536), .A2(n12535), .Z(n12540) );
  XOR3HSV2 U14399 ( .A1(n12541), .A2(n12540), .A3(n12539), .Z(\pe15/poht [1])
         );
  CLKNAND2HSV1 U14400 ( .A1(n12542), .A2(\pe21/got [2]), .ZN(n12556) );
  CLKNAND2HSV1 U14401 ( .A1(\pe21/ti_7[3] ), .A2(\pe21/got [1]), .ZN(n12554)
         );
  INHSV2 U14402 ( .I(\pe21/bq[3] ), .ZN(n14560) );
  CLKNHSV0 U14403 ( .I(\pe21/aot [3]), .ZN(n12544) );
  OAI21HSV0 U14404 ( .A1(n14560), .A2(n12544), .B(n12543), .ZN(n12545) );
  OAI21HSV2 U14405 ( .A1(n12547), .A2(n12546), .B(n12545), .ZN(n12551) );
  NAND2HSV0 U14406 ( .A1(\pe21/bq[4] ), .A2(\pe21/aot [2]), .ZN(n12549) );
  NAND2HSV0 U14407 ( .A1(\pe21/bq[2] ), .A2(\pe21/aot [4]), .ZN(n12548) );
  XOR2HSV0 U14408 ( .A1(n12549), .A2(n12548), .Z(n12550) );
  XOR3HSV2 U14409 ( .A1(n12552), .A2(n12551), .A3(n12550), .Z(n12553) );
  XOR2HSV0 U14410 ( .A1(n12554), .A2(n12553), .Z(n12555) );
  XOR2HSV0 U14411 ( .A1(n12556), .A2(n12555), .Z(n12558) );
  XNOR2HSV4 U14412 ( .A1(n12560), .A2(n12559), .ZN(\pe21/poht [3]) );
  NAND2HSV0 U14413 ( .A1(n14365), .A2(\pe11/got [3]), .ZN(n12567) );
  NAND2HSV0 U14414 ( .A1(n14366), .A2(\pe11/got [2]), .ZN(n12565) );
  CLKNAND2HSV0 U14415 ( .A1(n12562), .A2(\pe11/aot [2]), .ZN(n14370) );
  XOR2HSV0 U14416 ( .A1(n12565), .A2(n12564), .Z(n12566) );
  XOR2HSV0 U14417 ( .A1(n12567), .A2(n12566), .Z(n12568) );
  XNOR2HSV4 U14418 ( .A1(n12569), .A2(n12568), .ZN(n12571) );
  NAND2HSV0 U14419 ( .A1(n14830), .A2(\pe11/got [5]), .ZN(n12570) );
  NAND2HSV2 U14420 ( .A1(n14965), .A2(\pe11/got [6]), .ZN(n12572) );
  CLKNHSV0 U14421 ( .I(\pe4/got [2]), .ZN(n12574) );
  NOR2HSV2 U14422 ( .A1(n12645), .A2(n12574), .ZN(n12589) );
  NAND2HSV0 U14423 ( .A1(\pe4/got [1]), .A2(n10537), .ZN(n12587) );
  NAND2HSV0 U14424 ( .A1(\pe4/aot [4]), .A2(\pe4/bq[3] ), .ZN(n12576) );
  NAND2HSV0 U14425 ( .A1(\pe4/aot [3]), .A2(\pe4/bq[4] ), .ZN(n12575) );
  XOR2HSV0 U14426 ( .A1(n12576), .A2(n12575), .Z(n12580) );
  NAND2HSV0 U14427 ( .A1(\pe4/aot [6]), .A2(\pe4/bq[1] ), .ZN(n12578) );
  NAND2HSV0 U14428 ( .A1(\pe4/aot [5]), .A2(\pe4/bq[2] ), .ZN(n12577) );
  XOR2HSV0 U14429 ( .A1(n12578), .A2(n12577), .Z(n12579) );
  XOR2HSV0 U14430 ( .A1(n12580), .A2(n12579), .Z(n12585) );
  NAND2HSV0 U14431 ( .A1(n12581), .A2(\pe4/aot [1]), .ZN(n12583) );
  NAND2HSV0 U14432 ( .A1(\pe4/aot [2]), .A2(\pe4/bq[5] ), .ZN(n12582) );
  XOR2HSV0 U14433 ( .A1(n12583), .A2(n12582), .Z(n12584) );
  XNOR2HSV1 U14434 ( .A1(n12585), .A2(n12584), .ZN(n12586) );
  XOR2HSV0 U14435 ( .A1(n12587), .A2(n12586), .Z(n12588) );
  XOR2HSV0 U14436 ( .A1(n12589), .A2(n12588), .Z(n12613) );
  NOR2HSV2 U14437 ( .A1(n12590), .A2(n15083), .ZN(n12594) );
  NOR2HSV1 U14438 ( .A1(n12594), .A2(n12591), .ZN(n12593) );
  INHSV2 U14439 ( .I(n12595), .ZN(n12592) );
  NAND2HSV2 U14440 ( .A1(n12593), .A2(n12592), .ZN(n12601) );
  NAND2HSV2 U14441 ( .A1(n12595), .A2(n12594), .ZN(n12600) );
  AOI21HSV0 U14442 ( .A1(n12598), .A2(n12597), .B(n12596), .ZN(n12599) );
  NAND2HSV0 U14443 ( .A1(n12602), .A2(\pe4/got [5]), .ZN(n12611) );
  NAND2HSV2 U14444 ( .A1(n12631), .A2(\pe4/got [3]), .ZN(n12609) );
  NOR2HSV0 U14445 ( .A1(n12603), .A2(n12605), .ZN(n12607) );
  OAI22HSV0 U14446 ( .A1(n12605), .A2(n12604), .B1(\pe4/got [4]), .B2(n12609), 
        .ZN(n12606) );
  NOR2HSV1 U14447 ( .A1(n12607), .A2(n12606), .ZN(n12608) );
  OAI21HSV2 U14448 ( .A1(n14850), .A2(n12609), .B(n12608), .ZN(n12610) );
  XOR4HSV2 U14449 ( .A1(n12613), .A2(n12612), .A3(n12611), .A4(n12610), .Z(
        \pe4/poht [2]) );
  INHSV2 U14450 ( .I(ao3[5]), .ZN(n14897) );
  INHSV2 U14451 ( .I(ao3[8]), .ZN(n14899) );
  INHSV2 U14452 ( .I(ao14[8]), .ZN(n14903) );
  INHSV2 U14453 ( .I(ao9[6]), .ZN(n14905) );
  INHSV2 U14454 ( .I(ao19[8]), .ZN(n14907) );
  INHSV2 U14455 ( .I(go9[7]), .ZN(n14910) );
  INHSV2 U14456 ( .I(go9[8]), .ZN(n14911) );
  INHSV2 U14457 ( .I(go9[6]), .ZN(n14912) );
  INHSV2 U14458 ( .I(ao7[8]), .ZN(n14917) );
  INHSV2 U14459 ( .I(go7[6]), .ZN(n14918) );
  INHSV2 U14460 ( .I(ao3[7]), .ZN(n14919) );
  INHSV2 U14461 ( .I(ao10[8]), .ZN(n14921) );
  INHSV2 U14462 ( .I(ao10[7]), .ZN(n14923) );
  CLKNHSV0 U14463 ( .I(n12561), .ZN(n14924) );
  INHSV2 U14464 ( .I(go3[8]), .ZN(n14928) );
  NAND2HSV2 U14465 ( .A1(n14853), .A2(\pe15/got [5]), .ZN(n12628) );
  INHSV4 U14466 ( .I(n12614), .ZN(n14585) );
  CLKNHSV0 U14467 ( .I(\pe15/got [3]), .ZN(n12615) );
  NOR2HSV4 U14468 ( .A1(n14585), .A2(n12615), .ZN(n12624) );
  NAND2HSV0 U14469 ( .A1(\pe15/aot [2]), .A2(\pe15/bq[4] ), .ZN(n12621) );
  NAND2HSV0 U14470 ( .A1(n12616), .A2(\pe15/aot [1]), .ZN(n12618) );
  NAND2HSV0 U14471 ( .A1(\pe15/aot [4]), .A2(\pe15/bq[2] ), .ZN(n12617) );
  XOR2HSV0 U14472 ( .A1(n12618), .A2(n12617), .Z(n12619) );
  XOR3HSV2 U14473 ( .A1(n12621), .A2(n12620), .A3(n12619), .Z(n12622) );
  NAND2HSV0 U14474 ( .A1(\pe15/ti_7[3] ), .A2(\pe15/got [1]), .ZN(n12623) );
  NAND2HSV2 U14475 ( .A1(n6535), .A2(\pe15/got [4]), .ZN(n12625) );
  XNOR2HSV4 U14476 ( .A1(n12626), .A2(n12625), .ZN(n12627) );
  XNOR2HSV4 U14477 ( .A1(n12628), .A2(n12627), .ZN(\pe15/poht [3]) );
  INHSV2 U14478 ( .I(n12629), .ZN(n14930) );
  CLKNHSV0 U14479 ( .I(n12630), .ZN(n15238) );
  NAND2HSV2 U14480 ( .A1(n12941), .A2(n12940), .ZN(n13605) );
  BUFHSV8 U14481 ( .I(n15189), .Z(n14487) );
  NAND2HSV0 U14482 ( .A1(\pe4/aot [2]), .A2(\pe4/bq[6] ), .ZN(n12641) );
  NOR2HSV0 U14483 ( .A1(n12633), .A2(n12632), .ZN(n12635) );
  AOI22HSV0 U14484 ( .A1(\pe4/aot [5]), .A2(\pe4/bq[3] ), .B1(\pe4/bq[5] ), 
        .B2(\pe4/aot [3]), .ZN(n12634) );
  NOR2HSV2 U14485 ( .A1(n12635), .A2(n12634), .ZN(n12640) );
  CLKNAND2HSV0 U14486 ( .A1(n12636), .A2(\pe4/bq[1] ), .ZN(n12638) );
  NAND2HSV0 U14487 ( .A1(\pe4/aot [6]), .A2(\pe4/bq[2] ), .ZN(n12637) );
  XOR2HSV0 U14488 ( .A1(n12638), .A2(n12637), .Z(n12639) );
  XOR3HSV2 U14489 ( .A1(n12641), .A2(n12640), .A3(n12639), .Z(n12643) );
  CLKNHSV0 U14490 ( .I(n12643), .ZN(n12642) );
  NAND2HSV0 U14491 ( .A1(n12642), .A2(\pe4/got [3]), .ZN(n12644) );
  CLKNAND2HSV0 U14492 ( .A1(\pe4/ti_7[1] ), .A2(\pe4/got [1]), .ZN(n12649) );
  NAND2HSV0 U14493 ( .A1(\pe4/aot [1]), .A2(\pe4/bq[7] ), .ZN(n12647) );
  NAND2HSV0 U14494 ( .A1(\pe4/aot [4]), .A2(\pe4/bq[4] ), .ZN(n12646) );
  XOR2HSV0 U14495 ( .A1(n12647), .A2(n12646), .Z(n12648) );
  XNOR2HSV1 U14496 ( .A1(n12649), .A2(n12648), .ZN(n12651) );
  NAND2HSV0 U14497 ( .A1(\pe4/got [2]), .A2(n14733), .ZN(n12650) );
  XNOR2HSV1 U14498 ( .A1(n12651), .A2(n12650), .ZN(n12652) );
  XOR2HSV2 U14499 ( .A1(n12655), .A2(n12654), .Z(n12660) );
  NAND2HSV0 U14500 ( .A1(n12656), .A2(\pe4/got [5]), .ZN(n12657) );
  NOR2HSV0 U14501 ( .A1(n12658), .A2(n12657), .ZN(n12659) );
  CLKXOR2HSV2 U14502 ( .A1(n12660), .A2(n12659), .Z(n12662) );
  NAND2HSV0 U14503 ( .A1(n12602), .A2(\pe4/got [6]), .ZN(n12661) );
  CLKNHSV1 U14504 ( .I(\pe12/got [3]), .ZN(n14245) );
  CLKNAND2HSV0 U14505 ( .A1(n14943), .A2(\pe12/got [2]), .ZN(n12674) );
  NAND2HSV0 U14506 ( .A1(\pe12/bq[3] ), .A2(\pe12/aot [3]), .ZN(n12670) );
  NAND2HSV0 U14507 ( .A1(\pe12/aot [4]), .A2(\pe12/bq[4] ), .ZN(n14240) );
  CLKNAND2HSV1 U14508 ( .A1(\pe12/bq[2] ), .A2(\pe12/aot [2]), .ZN(n14439) );
  NOR2HSV0 U14509 ( .A1(n14240), .A2(n14439), .ZN(n12665) );
  AOI22HSV0 U14510 ( .A1(\pe12/aot [4]), .A2(\pe12/bq[2] ), .B1(\pe12/bq[4] ), 
        .B2(\pe12/aot [2]), .ZN(n12664) );
  NOR2HSV2 U14511 ( .A1(n12665), .A2(n12664), .ZN(n12669) );
  NAND2HSV2 U14512 ( .A1(\pe12/aot [1]), .A2(\pe12/bq[1] ), .ZN(n13939) );
  AO22HSV2 U14513 ( .A1(\pe12/aot [5]), .A2(\pe12/bq[1] ), .B1(\pe12/bq[5] ), 
        .B2(\pe12/aot [1]), .Z(n12666) );
  OAI21HSV0 U14514 ( .A1(n13939), .A2(n12667), .B(n12666), .ZN(n12668) );
  XOR3HSV2 U14515 ( .A1(n12670), .A2(n12669), .A3(n12668), .Z(n12671) );
  XNOR2HSV1 U14516 ( .A1(n12672), .A2(n12671), .ZN(n12673) );
  XNOR2HSV1 U14517 ( .A1(n12674), .A2(n12673), .ZN(n12675) );
  XNOR2HSV4 U14518 ( .A1(n12676), .A2(n12675), .ZN(n12678) );
  NAND2HSV0 U14519 ( .A1(n15190), .A2(\pe12/got [4]), .ZN(n12677) );
  XNOR2HSV4 U14520 ( .A1(n12678), .A2(n12677), .ZN(n12682) );
  NAND2HSV0 U14521 ( .A1(n14446), .A2(\pe12/got [5]), .ZN(n12681) );
  XOR2HSV0 U14522 ( .A1(n12682), .A2(n12681), .Z(\pe12/poht [3]) );
  NOR2HSV2 U14523 ( .A1(n12713), .A2(n12683), .ZN(n12707) );
  NAND2HSV0 U14524 ( .A1(n14943), .A2(\pe12/got [5]), .ZN(n12705) );
  CLKNAND2HSV0 U14525 ( .A1(n14578), .A2(\pe12/pq ), .ZN(n12685) );
  NAND2HSV0 U14526 ( .A1(n14948), .A2(\pe12/bq[2] ), .ZN(n12684) );
  XOR2HSV0 U14527 ( .A1(n12685), .A2(n12684), .Z(n12689) );
  NAND2HSV0 U14528 ( .A1(\pe12/aot [5]), .A2(\pe12/bq[4] ), .ZN(n12687) );
  NAND2HSV0 U14529 ( .A1(\pe12/got [1]), .A2(n13830), .ZN(n12686) );
  XOR2HSV0 U14530 ( .A1(n12687), .A2(n12686), .Z(n12688) );
  XOR2HSV0 U14531 ( .A1(n12689), .A2(n12688), .Z(n12691) );
  NAND2HSV0 U14532 ( .A1(\pe12/aot [3]), .A2(\pe12/bq[6] ), .ZN(n12725) );
  NAND2HSV0 U14533 ( .A1(\pe12/aot [6]), .A2(\pe12/bq[3] ), .ZN(n12730) );
  XOR2HSV0 U14534 ( .A1(n12725), .A2(n12730), .Z(n12690) );
  XNOR2HSV1 U14535 ( .A1(n12691), .A2(n12690), .ZN(n12699) );
  CLKNHSV0 U14536 ( .I(\pe12/aot [1]), .ZN(n14241) );
  NAND2HSV0 U14537 ( .A1(\pe12/aot [1]), .A2(n14507), .ZN(n12693) );
  NAND2HSV0 U14538 ( .A1(n14876), .A2(\pe12/bq[1] ), .ZN(n12692) );
  XOR2HSV0 U14539 ( .A1(n12693), .A2(n12692), .Z(n12697) );
  NAND2HSV0 U14540 ( .A1(\pe12/aot [2]), .A2(\pe12/bq[7] ), .ZN(n12695) );
  NAND2HSV0 U14541 ( .A1(\pe12/aot [4]), .A2(\pe12/bq[5] ), .ZN(n12694) );
  XOR2HSV0 U14542 ( .A1(n12695), .A2(n12694), .Z(n12696) );
  XOR2HSV0 U14543 ( .A1(n12697), .A2(n12696), .Z(n12698) );
  XNOR2HSV1 U14544 ( .A1(n12699), .A2(n12698), .ZN(n12700) );
  XNOR2HSV1 U14545 ( .A1(n12701), .A2(n12700), .ZN(n12702) );
  XOR2HSV0 U14546 ( .A1(n12703), .A2(n12702), .Z(n12704) );
  XOR2HSV0 U14547 ( .A1(n12704), .A2(n12705), .Z(n12706) );
  XNOR2HSV4 U14548 ( .A1(n12707), .A2(n12706), .ZN(n12709) );
  NAND2HSV0 U14549 ( .A1(n15190), .A2(\pe12/got [7]), .ZN(n12708) );
  XNOR2HSV4 U14550 ( .A1(n12709), .A2(n12708), .ZN(n12711) );
  NAND2HSV0 U14551 ( .A1(n14446), .A2(n5958), .ZN(n12710) );
  XOR2HSV0 U14552 ( .A1(n12711), .A2(n12710), .Z(po12) );
  CLKNHSV0 U14553 ( .I(\pe12/got [2]), .ZN(n12712) );
  NOR2HSV2 U14554 ( .A1(n14442), .A2(n12712), .ZN(n12721) );
  NAND2HSV0 U14555 ( .A1(n14943), .A2(\pe12/got [1]), .ZN(n12719) );
  CLKNAND2HSV0 U14556 ( .A1(\pe12/aot [1]), .A2(\pe12/bq[4] ), .ZN(n14244) );
  NAND2HSV0 U14557 ( .A1(\pe12/aot [4]), .A2(\pe12/bq[1] ), .ZN(n12729) );
  XOR2HSV0 U14558 ( .A1(n14244), .A2(n12729), .Z(n12717) );
  NAND2HSV0 U14559 ( .A1(\pe12/aot [3]), .A2(\pe12/bq[2] ), .ZN(n12715) );
  NAND2HSV0 U14560 ( .A1(\pe12/aot [2]), .A2(\pe12/bq[3] ), .ZN(n12714) );
  XOR2HSV0 U14561 ( .A1(n12715), .A2(n12714), .Z(n12716) );
  XOR2HSV0 U14562 ( .A1(n12717), .A2(n12716), .Z(n12718) );
  XOR2HSV0 U14563 ( .A1(n12719), .A2(n12718), .Z(n12720) );
  XNOR2HSV4 U14564 ( .A1(n12721), .A2(n12720), .ZN(n12722) );
  CLKNHSV1 U14565 ( .I(\pe12/got [4]), .ZN(n14248) );
  NOR2HSV2 U14566 ( .A1(n14442), .A2(n14248), .ZN(n12744) );
  CLKNAND2HSV1 U14567 ( .A1(n14943), .A2(\pe12/got [3]), .ZN(n12742) );
  NAND2HSV0 U14568 ( .A1(\pe12/aot [5]), .A2(\pe12/bq[2] ), .ZN(n12724) );
  NAND2HSV0 U14569 ( .A1(\pe12/aot [2]), .A2(\pe12/bq[5] ), .ZN(n12723) );
  XOR2HSV0 U14570 ( .A1(n12724), .A2(n12723), .Z(n12738) );
  CLKNHSV0 U14571 ( .I(n12725), .ZN(n12728) );
  CLKNHSV0 U14572 ( .I(n14244), .ZN(n12727) );
  AOI22HSV0 U14573 ( .A1(\pe12/aot [3]), .A2(\pe12/bq[4] ), .B1(\pe12/bq[6] ), 
        .B2(\pe12/aot [1]), .ZN(n12726) );
  AOI21HSV2 U14574 ( .A1(n12728), .A2(n12727), .B(n12726), .ZN(n12735) );
  CLKNHSV0 U14575 ( .I(n12729), .ZN(n12733) );
  CLKNHSV0 U14576 ( .I(n12730), .ZN(n12732) );
  AOI22HSV0 U14577 ( .A1(\pe12/aot [6]), .A2(\pe12/bq[1] ), .B1(\pe12/aot [4]), 
        .B2(\pe12/bq[3] ), .ZN(n12731) );
  AOI21HSV2 U14578 ( .A1(n12733), .A2(n12732), .B(n12731), .ZN(n12734) );
  XOR2HSV0 U14579 ( .A1(n12735), .A2(n12734), .Z(n12737) );
  NAND2HSV0 U14580 ( .A1(n14255), .A2(\pe12/got [1]), .ZN(n12736) );
  XOR3HSV2 U14581 ( .A1(n12738), .A2(n12737), .A3(n12736), .Z(n12739) );
  XOR2HSV0 U14582 ( .A1(n12740), .A2(n12739), .Z(n12741) );
  XOR2HSV0 U14583 ( .A1(n12742), .A2(n12741), .Z(n12743) );
  XNOR2HSV4 U14584 ( .A1(n12744), .A2(n12743), .ZN(n12746) );
  NAND2HSV2 U14585 ( .A1(n14446), .A2(\pe12/got [6]), .ZN(n12745) );
  NAND2HSV0 U14586 ( .A1(n14820), .A2(\pe3/got [3]), .ZN(n12764) );
  NAND2HSV0 U14587 ( .A1(\pe3/aot [5]), .A2(\pe3/bq[3] ), .ZN(n12747) );
  XOR2HSV0 U14588 ( .A1(n12748), .A2(n12747), .Z(n12752) );
  NAND2HSV0 U14589 ( .A1(\pe3/aot [1]), .A2(\pe3/bq[7] ), .ZN(n12749) );
  XOR2HSV0 U14590 ( .A1(n12750), .A2(n12749), .Z(n12751) );
  XOR2HSV0 U14591 ( .A1(n12752), .A2(n12751), .Z(n12758) );
  NAND2HSV0 U14592 ( .A1(\pe3/aot [7]), .A2(\pe3/bq[1] ), .ZN(n12754) );
  NAND2HSV0 U14593 ( .A1(\pe3/aot [4]), .A2(\pe3/bq[4] ), .ZN(n12753) );
  XOR2HSV0 U14594 ( .A1(n12754), .A2(n12753), .Z(n12756) );
  NAND2HSV0 U14595 ( .A1(\pe3/bq[2] ), .A2(\pe3/aot [6]), .ZN(n12755) );
  XNOR2HSV1 U14596 ( .A1(n12756), .A2(n12755), .ZN(n12757) );
  XNOR2HSV1 U14597 ( .A1(n12758), .A2(n12757), .ZN(n12760) );
  NAND2HSV0 U14598 ( .A1(n5949), .A2(\pe3/got [1]), .ZN(n12759) );
  XOR2HSV0 U14599 ( .A1(n12760), .A2(n12759), .Z(n12762) );
  CLKNAND2HSV0 U14600 ( .A1(\pe3/got [2]), .A2(n14872), .ZN(n12761) );
  XNOR2HSV1 U14601 ( .A1(n12762), .A2(n12761), .ZN(n12763) );
  XOR2HSV0 U14602 ( .A1(n12764), .A2(n12763), .Z(n12765) );
  XOR2HSV0 U14603 ( .A1(n12766), .A2(n12765), .Z(n12767) );
  NAND2HSV0 U14604 ( .A1(\pe3/got [5]), .A2(\pe3/ti_7[5] ), .ZN(n12768) );
  XNOR2HSV1 U14605 ( .A1(n12770), .A2(n12769), .ZN(n15203) );
  CLKNHSV0 U14606 ( .I(bo4[1]), .ZN(n12772) );
  MUX2NHSV0 U14607 ( .I0(n12772), .I1(n12771), .S(n10562), .ZN(n15041) );
  AND2HSV2 U14608 ( .A1(n12773), .A2(n10307), .Z(n12774) );
  INHSV2 U14609 ( .I(\pe5/ti_7t [6]), .ZN(n12778) );
  AND2HSV2 U14610 ( .A1(n13015), .A2(n12778), .Z(n12783) );
  AOI31HSV1 U14611 ( .A1(n6922), .A2(n10307), .A3(n12779), .B(n12783), .ZN(
        n12781) );
  CLKNAND2HSV1 U14612 ( .A1(n12782), .A2(n12781), .ZN(n12789) );
  NOR2HSV1 U14613 ( .A1(n12784), .A2(n12783), .ZN(n12785) );
  INAND2HSV2 U14614 ( .A1(n12791), .B1(\pe5/got [6]), .ZN(n12815) );
  NAND2HSV0 U14615 ( .A1(n10346), .A2(\pe5/got [3]), .ZN(n12810) );
  NAND2HSV2 U14616 ( .A1(n14952), .A2(\pe5/got [4]), .ZN(n12809) );
  NAND2HSV0 U14617 ( .A1(\pe5/got [2]), .A2(\pe5/ti_1 ), .ZN(n12793) );
  NAND2HSV0 U14618 ( .A1(\pe5/aot [2]), .A2(\pe5/bq[8] ), .ZN(n12792) );
  XOR2HSV0 U14619 ( .A1(n12793), .A2(n12792), .Z(n12807) );
  NAND2HSV0 U14620 ( .A1(\pe5/aot [7]), .A2(\pe5/bq[3] ), .ZN(n12795) );
  NAND2HSV0 U14621 ( .A1(\pe5/aot [8]), .A2(\pe5/bq[2] ), .ZN(n12794) );
  XOR2HSV0 U14622 ( .A1(n12795), .A2(n12794), .Z(n12798) );
  NAND2HSV0 U14623 ( .A1(\pe5/ctrq ), .A2(\pe5/pvq [7]), .ZN(n12796) );
  XOR2HSV0 U14624 ( .A1(n12796), .A2(\pe5/phq [7]), .Z(n12797) );
  XNOR2HSV1 U14625 ( .A1(n12798), .A2(n12797), .ZN(n12806) );
  NAND2HSV0 U14626 ( .A1(\pe5/bq[5] ), .A2(\pe5/aot [5]), .ZN(n12800) );
  NAND2HSV0 U14627 ( .A1(\pe5/aot [6]), .A2(\pe5/bq[4] ), .ZN(n12799) );
  XOR2HSV0 U14628 ( .A1(n12800), .A2(n12799), .Z(n12804) );
  NAND2HSV0 U14629 ( .A1(\pe5/aot [4]), .A2(\pe5/bq[6] ), .ZN(n12802) );
  NAND2HSV0 U14630 ( .A1(\pe5/aot [3]), .A2(\pe5/bq[7] ), .ZN(n12801) );
  XOR2HSV0 U14631 ( .A1(n12802), .A2(n12801), .Z(n12803) );
  XOR2HSV0 U14632 ( .A1(n12804), .A2(n12803), .Z(n12805) );
  XOR3HSV2 U14633 ( .A1(n12807), .A2(n12806), .A3(n12805), .Z(n12808) );
  XOR3HSV2 U14634 ( .A1(n12810), .A2(n12808), .A3(n12809), .Z(n12813) );
  NAND2HSV0 U14635 ( .A1(n6710), .A2(\pe5/got [5]), .ZN(n12812) );
  XOR2HSV2 U14636 ( .A1(n12815), .A2(n12814), .Z(n12826) );
  CLKNAND2HSV2 U14637 ( .A1(n12816), .A2(n15067), .ZN(n12820) );
  INAND2HSV0 U14638 ( .A1(n12817), .B1(\pe5/got [7]), .ZN(n12818) );
  AOI21HSV2 U14639 ( .A1(n12819), .A2(n12820), .B(n12818), .ZN(n12824) );
  INHSV2 U14640 ( .I(n12820), .ZN(n12822) );
  CLKNAND2HSV1 U14641 ( .A1(n12822), .A2(n12821), .ZN(n12823) );
  CLKNHSV0 U14642 ( .I(\pe15/ti_7t [7]), .ZN(n12827) );
  AOI21HSV2 U14643 ( .A1(n12827), .A2(n12829), .B(n14584), .ZN(n12828) );
  OAI21HSV4 U14644 ( .A1(n15231), .A2(n12829), .B(n12828), .ZN(n12849) );
  NAND2HSV0 U14645 ( .A1(\pe15/ti_7[3] ), .A2(\pe15/got [2]), .ZN(n12845) );
  CLKNAND2HSV0 U14646 ( .A1(n5946), .A2(\pe15/got [1]), .ZN(n12842) );
  NAND2HSV0 U14647 ( .A1(\pe15/aot [2]), .A2(\pe15/bq[5] ), .ZN(n12832) );
  NAND2HSV0 U14648 ( .A1(\pe15/aot [5]), .A2(\pe15/bq[2] ), .ZN(n12831) );
  XOR2HSV0 U14649 ( .A1(n12832), .A2(n12831), .Z(n12836) );
  NAND2HSV0 U14650 ( .A1(\pe15/aot [3]), .A2(\pe15/bq[4] ), .ZN(n12834) );
  NAND2HSV0 U14651 ( .A1(\pe15/aot [6]), .A2(\pe15/bq[1] ), .ZN(n12833) );
  XOR2HSV0 U14652 ( .A1(n12834), .A2(n12833), .Z(n12835) );
  XOR2HSV0 U14653 ( .A1(n12836), .A2(n12835), .Z(n12840) );
  NAND2HSV0 U14654 ( .A1(\pe15/aot [4]), .A2(\pe15/bq[3] ), .ZN(n12838) );
  NAND2HSV0 U14655 ( .A1(\pe15/aot [1]), .A2(\pe15/bq[6] ), .ZN(n12837) );
  XOR2HSV0 U14656 ( .A1(n12838), .A2(n12837), .Z(n12839) );
  XNOR2HSV1 U14657 ( .A1(n12840), .A2(n12839), .ZN(n12841) );
  XOR2HSV0 U14658 ( .A1(n12842), .A2(n12841), .Z(n12843) );
  CLKNHSV0 U14659 ( .I(\pe15/got [4]), .ZN(n12844) );
  NAND2HSV2 U14660 ( .A1(n6535), .A2(\pe15/got [5]), .ZN(n12846) );
  XNOR2HSV4 U14661 ( .A1(n12849), .A2(n12848), .ZN(\pe15/poht [2]) );
  NAND2HSV0 U14662 ( .A1(n14847), .A2(\pe1/got [1]), .ZN(n12856) );
  NAND2HSV0 U14663 ( .A1(\pe1/aot [2]), .A2(\pe1/bq[3] ), .ZN(n12851) );
  NAND2HSV0 U14664 ( .A1(\pe1/bq[2] ), .A2(\pe1/aot [3]), .ZN(n12850) );
  XOR2HSV0 U14665 ( .A1(n12851), .A2(n12850), .Z(n12854) );
  CLKNAND2HSV0 U14666 ( .A1(\pe1/aot [1]), .A2(\pe1/bq[4] ), .ZN(n12864) );
  NAND2HSV0 U14667 ( .A1(\pe1/aot [4]), .A2(\pe1/bq[1] ), .ZN(n12852) );
  XOR2HSV0 U14668 ( .A1(n12864), .A2(n12852), .Z(n12853) );
  XOR2HSV0 U14669 ( .A1(n12854), .A2(n12853), .Z(n12855) );
  XNOR2HSV1 U14670 ( .A1(n12856), .A2(n12855), .ZN(n12859) );
  CLKBUFHSV4 U14671 ( .I(\pe1/ti_7[5] ), .Z(n14006) );
  NAND2HSV2 U14672 ( .A1(n14006), .A2(\pe1/got [2]), .ZN(n12858) );
  CLKNAND2HSV0 U14673 ( .A1(\pe1/ti_7[6] ), .A2(\pe1/got [3]), .ZN(n12857) );
  XNOR3HSV1 U14674 ( .A1(n12859), .A2(n12858), .A3(n12857), .ZN(n12861) );
  XOR2HSV0 U14675 ( .A1(n12861), .A2(n12860), .Z(\pe1/poht [4]) );
  NAND2HSV0 U14676 ( .A1(\pe1/aot [4]), .A2(\pe1/bq[2] ), .ZN(n13998) );
  NAND2HSV0 U14677 ( .A1(\pe1/aot [2]), .A2(\pe1/bq[5] ), .ZN(n13945) );
  NAND2HSV0 U14678 ( .A1(\pe1/aot [1]), .A2(\pe1/bq[5] ), .ZN(n13970) );
  NAND2HSV0 U14679 ( .A1(\pe1/aot [2]), .A2(\pe1/bq[4] ), .ZN(n12862) );
  CLKNAND2HSV1 U14680 ( .A1(n13970), .A2(n12862), .ZN(n12863) );
  OAI21HSV2 U14681 ( .A1(n13945), .A2(n12864), .B(n12863), .ZN(n12868) );
  NAND2HSV0 U14682 ( .A1(\pe1/bq[1] ), .A2(\pe1/aot [5]), .ZN(n12865) );
  XOR2HSV0 U14683 ( .A1(n12866), .A2(n12865), .Z(n12867) );
  XOR3HSV2 U14684 ( .A1(n13998), .A2(n12868), .A3(n12867), .Z(n12872) );
  CLKNHSV0 U14685 ( .I(\pe1/got [1]), .ZN(n12869) );
  NOR2HSV1 U14686 ( .A1(n13953), .A2(n12869), .ZN(n12871) );
  NAND2HSV0 U14687 ( .A1(n14847), .A2(\pe1/got [2]), .ZN(n12870) );
  XOR3HSV2 U14688 ( .A1(n12872), .A2(n12871), .A3(n12870), .Z(n12875) );
  NAND2HSV2 U14689 ( .A1(n14006), .A2(\pe1/got [3]), .ZN(n12874) );
  CLKNAND2HSV0 U14690 ( .A1(\pe1/ti_7[6] ), .A2(\pe1/got [4]), .ZN(n12873) );
  XNOR3HSV1 U14691 ( .A1(n12875), .A2(n12874), .A3(n12873), .ZN(n12877) );
  NAND2HSV0 U14692 ( .A1(\pe1/ti_7[7] ), .A2(\pe1/got [5]), .ZN(n12876) );
  XOR2HSV0 U14693 ( .A1(n12877), .A2(n12876), .Z(\pe1/poht [3]) );
  NOR2HSV0 U14694 ( .A1(n13102), .A2(n12878), .ZN(n12906) );
  INHSV1 U14695 ( .I(\pe2/got [3]), .ZN(n13101) );
  NOR2HSV2 U14696 ( .A1(n12879), .A2(n13101), .ZN(n12887) );
  NAND2HSV0 U14697 ( .A1(\pe2/bq[5] ), .A2(\pe2/aot [3]), .ZN(n13093) );
  XOR2HSV0 U14698 ( .A1(n13093), .A2(n12880), .Z(n12885) );
  NAND2HSV2 U14699 ( .A1(\pe2/aot [1]), .A2(\pe2/bq[1] ), .ZN(n14062) );
  NOR2HSV0 U14700 ( .A1(n14062), .A2(n12881), .ZN(n12883) );
  AOI22HSV0 U14701 ( .A1(\pe2/aot [1]), .A2(n14504), .B1(\pe2/aot [7]), .B2(
        \pe2/bq[1] ), .ZN(n12882) );
  NOR2HSV1 U14702 ( .A1(n12883), .A2(n12882), .ZN(n12884) );
  XNOR2HSV1 U14703 ( .A1(n12885), .A2(n12884), .ZN(n12886) );
  CLKNHSV0 U14704 ( .I(n12889), .ZN(n12888) );
  NOR2HSV1 U14705 ( .A1(n12888), .A2(n13760), .ZN(n12891) );
  AOI21HSV0 U14706 ( .A1(\pe2/got [4]), .A2(n12907), .B(n12889), .ZN(n12890)
         );
  AOI21HSV2 U14707 ( .A1(n12891), .A2(n14935), .B(n12890), .ZN(n12901) );
  NAND2HSV0 U14708 ( .A1(\pe2/ti_7[1] ), .A2(\pe2/got [1]), .ZN(n12897) );
  NAND2HSV0 U14709 ( .A1(\pe2/aot [5]), .A2(\pe2/bq[3] ), .ZN(n12893) );
  NAND2HSV0 U14710 ( .A1(\pe2/aot [2]), .A2(n14510), .ZN(n12892) );
  XOR2HSV0 U14711 ( .A1(n12893), .A2(n12892), .Z(n12895) );
  NAND2HSV0 U14712 ( .A1(\pe2/aot [4]), .A2(\pe2/bq[4] ), .ZN(n12894) );
  XNOR2HSV1 U14713 ( .A1(n12895), .A2(n12894), .ZN(n12896) );
  XNOR2HSV1 U14714 ( .A1(n12897), .A2(n12896), .ZN(n12899) );
  NAND2HSV0 U14715 ( .A1(n14934), .A2(\pe2/got [2]), .ZN(n12898) );
  XOR2HSV0 U14716 ( .A1(n12899), .A2(n12898), .Z(n12900) );
  XOR2HSV0 U14717 ( .A1(n12901), .A2(n12900), .Z(n12902) );
  XNOR2HSV4 U14718 ( .A1(n12903), .A2(n12902), .ZN(n12905) );
  NAND2HSV2 U14719 ( .A1(n14061), .A2(\pe2/got [7]), .ZN(n12904) );
  XOR3HSV2 U14720 ( .A1(n12906), .A2(n12905), .A3(n12904), .Z(\pe2/poht [1])
         );
  CLKNAND2HSV0 U14721 ( .A1(n12907), .A2(\pe2/got [1]), .ZN(n12915) );
  NAND2HSV0 U14722 ( .A1(\pe2/bq[1] ), .A2(\pe2/aot [4]), .ZN(n12909) );
  NAND2HSV0 U14723 ( .A1(\pe2/bq[2] ), .A2(\pe2/aot [3]), .ZN(n12908) );
  XOR2HSV0 U14724 ( .A1(n12909), .A2(n12908), .Z(n12913) );
  NAND2HSV0 U14725 ( .A1(\pe2/aot [1]), .A2(\pe2/bq[4] ), .ZN(n12911) );
  NAND2HSV0 U14726 ( .A1(\pe2/bq[3] ), .A2(\pe2/aot [2]), .ZN(n12910) );
  XOR2HSV0 U14727 ( .A1(n12911), .A2(n12910), .Z(n12912) );
  XOR2HSV0 U14728 ( .A1(n12913), .A2(n12912), .Z(n12914) );
  XOR2HSV0 U14729 ( .A1(n12915), .A2(n12914), .Z(n12918) );
  NOR2HSV0 U14730 ( .A1(n13102), .A2(n13100), .ZN(n12916) );
  XNOR3HSV2 U14731 ( .A1(n12918), .A2(n12917), .A3(n12916), .ZN(n12920) );
  XOR2HSV0 U14732 ( .A1(n12920), .A2(n12919), .Z(\pe2/poht [4]) );
  CLKNHSV0 U14733 ( .I(\pe13/got [3]), .ZN(n12921) );
  NAND2HSV2 U14734 ( .A1(n15065), .A2(\pe13/got [1]), .ZN(n12931) );
  NAND2HSV0 U14735 ( .A1(\pe13/aot [2]), .A2(\pe13/bq[4] ), .ZN(n12929) );
  NAND2HSV0 U14736 ( .A1(\pe13/aot [5]), .A2(\pe13/bq[1] ), .ZN(n12923) );
  AOI22HSV0 U14737 ( .A1(n12924), .A2(n12923), .B1(n12922), .B2(n13337), .ZN(
        n12928) );
  NAND2HSV0 U14738 ( .A1(\pe13/aot [4]), .A2(\pe13/bq[2] ), .ZN(n12926) );
  NAND2HSV0 U14739 ( .A1(\pe13/bq[3] ), .A2(\pe13/aot [3]), .ZN(n12925) );
  XOR2HSV0 U14740 ( .A1(n12926), .A2(n12925), .Z(n12927) );
  XOR3HSV1 U14741 ( .A1(n12929), .A2(n12928), .A3(n12927), .Z(n12930) );
  XNOR2HSV1 U14742 ( .A1(n12931), .A2(n12930), .ZN(n12933) );
  AOI21HSV0 U14743 ( .A1(\pe13/got [2]), .A2(\pe13/ti_7[4] ), .B(n12933), .ZN(
        n12932) );
  NAND2HSV2 U14744 ( .A1(n14961), .A2(\pe13/got [5]), .ZN(n12934) );
  XOR2HSV0 U14745 ( .A1(n12935), .A2(n12934), .Z(\pe13/poht [3]) );
  CLKAND2HSV2 U14746 ( .A1(n13034), .A2(\pe6/got [1]), .Z(n12938) );
  CLKNAND2HSV0 U14747 ( .A1(\pe6/aot [2]), .A2(\pe6/bq[3] ), .ZN(n12999) );
  NAND2HSV2 U14748 ( .A1(\pe6/aot [4]), .A2(\pe6/bq[5] ), .ZN(n13048) );
  NAND2HSV2 U14749 ( .A1(\pe6/aot [3]), .A2(\pe6/bq[6] ), .ZN(n13049) );
  INHSV2 U14750 ( .I(n14845), .ZN(n13827) );
  NAND2HSV0 U14751 ( .A1(n13057), .A2(\pe6/got [2]), .ZN(n12939) );
  CLKNHSV0 U14752 ( .I(\pe7/got [1]), .ZN(n12943) );
  NAND2HSV0 U14753 ( .A1(\pe7/aot [4]), .A2(\pe7/bq[2] ), .ZN(n12945) );
  NAND2HSV0 U14754 ( .A1(\pe7/aot [2]), .A2(\pe7/bq[4] ), .ZN(n12944) );
  XOR2HSV0 U14755 ( .A1(n12945), .A2(n12944), .Z(n12946) );
  NAND2HSV0 U14756 ( .A1(\pe7/aot [5]), .A2(\pe7/bq[1] ), .ZN(n13610) );
  NAND2HSV0 U14757 ( .A1(\pe7/aot [3]), .A2(\pe7/bq[3] ), .ZN(n12948) );
  NAND2HSV0 U14758 ( .A1(\pe7/aot [1]), .A2(\pe7/bq[5] ), .ZN(n12947) );
  NAND2HSV0 U14759 ( .A1(\pe3/aot [2]), .A2(\pe3/bq[3] ), .ZN(n12950) );
  NAND2HSV0 U14760 ( .A1(\pe3/aot [1]), .A2(\pe3/bq[4] ), .ZN(n12949) );
  XOR2HSV0 U14761 ( .A1(n12950), .A2(n12949), .Z(n12954) );
  NAND2HSV0 U14762 ( .A1(\pe3/aot [3]), .A2(\pe3/bq[2] ), .ZN(n12952) );
  NAND2HSV0 U14763 ( .A1(\pe3/aot [4]), .A2(\pe3/bq[1] ), .ZN(n12951) );
  XOR2HSV0 U14764 ( .A1(n12952), .A2(n12951), .Z(n12953) );
  XOR2HSV0 U14765 ( .A1(n12954), .A2(n12953), .Z(n12955) );
  XNOR2HSV1 U14766 ( .A1(n12956), .A2(n12955), .ZN(n12962) );
  CLKNHSV0 U14767 ( .I(\pe3/got [2]), .ZN(n12958) );
  NOR2HSV2 U14768 ( .A1(n12959), .A2(n12958), .ZN(n12960) );
  XOR3HSV2 U14769 ( .A1(n12962), .A2(n12961), .A3(n12960), .Z(n12964) );
  NAND2HSV0 U14770 ( .A1(\pe3/aot [2]), .A2(\pe3/bq[2] ), .ZN(n12966) );
  NAND2HSV0 U14771 ( .A1(\pe3/aot [1]), .A2(\pe3/bq[3] ), .ZN(n12965) );
  XOR2HSV0 U14772 ( .A1(n12966), .A2(n12965), .Z(n12968) );
  NAND2HSV0 U14773 ( .A1(\pe3/aot [3]), .A2(\pe3/bq[1] ), .ZN(n12967) );
  XNOR2HSV1 U14774 ( .A1(n12968), .A2(n12967), .ZN(n12972) );
  INHSV2 U14775 ( .I(n12969), .ZN(n12971) );
  NAND2HSV0 U14776 ( .A1(n12981), .A2(\pe3/got [2]), .ZN(n12970) );
  XOR3HSV2 U14777 ( .A1(n12972), .A2(n12971), .A3(n12970), .Z(n12974) );
  NAND2HSV0 U14778 ( .A1(\pe3/aot [4]), .A2(\pe3/bq[2] ), .ZN(n12976) );
  NAND2HSV0 U14779 ( .A1(\pe3/aot [2]), .A2(\pe3/bq[4] ), .ZN(n12975) );
  XNOR2HSV1 U14780 ( .A1(n12976), .A2(n12975), .ZN(n12980) );
  NAND2HSV0 U14781 ( .A1(\pe3/aot [5]), .A2(\pe3/bq[1] ), .ZN(n12978) );
  NAND2HSV0 U14782 ( .A1(\pe3/aot [1]), .A2(\pe3/bq[5] ), .ZN(n12977) );
  XOR2HSV0 U14783 ( .A1(n12978), .A2(n12977), .Z(n12979) );
  NAND2HSV0 U14784 ( .A1(\pe6/aot [1]), .A2(\pe6/bq[3] ), .ZN(n12983) );
  NAND2HSV0 U14785 ( .A1(\pe6/aot [2]), .A2(\pe6/bq[2] ), .ZN(n12982) );
  XOR2HSV0 U14786 ( .A1(n12983), .A2(n12982), .Z(n12985) );
  XOR2HSV0 U14787 ( .A1(n12985), .A2(n12984), .Z(n12986) );
  XOR2HSV0 U14788 ( .A1(n12987), .A2(n12986), .Z(n12988) );
  NAND2HSV0 U14789 ( .A1(\pe13/aot [4]), .A2(\pe13/bq[1] ), .ZN(n12993) );
  NAND2HSV0 U14790 ( .A1(\pe13/aot [2]), .A2(\pe13/bq[3] ), .ZN(n12992) );
  NAND2HSV0 U14791 ( .A1(\pe13/aot [3]), .A2(\pe13/bq[2] ), .ZN(n12995) );
  NAND2HSV0 U14792 ( .A1(\pe13/aot [1]), .A2(\pe13/bq[4] ), .ZN(n12994) );
  XOR2HSV0 U14793 ( .A1(n12995), .A2(n12994), .Z(n12996) );
  CLKNAND2HSV2 U14794 ( .A1(\pe6/ti_7[5] ), .A2(\pe6/got [2]), .ZN(n13006) );
  NAND2HSV0 U14795 ( .A1(n15077), .A2(\pe6/got [1]), .ZN(n13004) );
  XOR2HSV0 U14796 ( .A1(n13000), .A2(n12999), .Z(n13002) );
  XNOR2HSV1 U14797 ( .A1(n13002), .A2(n13001), .ZN(n13003) );
  XNOR2HSV1 U14798 ( .A1(n13004), .A2(n13003), .ZN(n13005) );
  XNOR2HSV1 U14799 ( .A1(n13006), .A2(n13005), .ZN(n13007) );
  XNOR2HSV4 U14800 ( .A1(n13008), .A2(n13007), .ZN(n13009) );
  XNOR2HSV4 U14801 ( .A1(n13010), .A2(n13009), .ZN(\pe6/poht [4]) );
  NAND2HSV0 U14802 ( .A1(n10307), .A2(n13861), .ZN(n13011) );
  AOI21HSV2 U14803 ( .A1(n13013), .A2(n13012), .B(n13011), .ZN(n13017) );
  CLKAND2HSV2 U14804 ( .A1(n13015), .A2(\pe5/ti_7t [7]), .Z(n13016) );
  CLKNAND2HSV0 U14805 ( .A1(n10346), .A2(\pe5/got [1]), .ZN(n13033) );
  NAND2HSV0 U14806 ( .A1(\pe5/aot [6]), .A2(\pe5/bq[2] ), .ZN(n13021) );
  NAND2HSV0 U14807 ( .A1(\pe5/aot [4]), .A2(\pe5/bq[4] ), .ZN(n13020) );
  XOR2HSV0 U14808 ( .A1(n13021), .A2(n13020), .Z(n13025) );
  NAND2HSV0 U14809 ( .A1(\pe5/aot [5]), .A2(\pe5/bq[3] ), .ZN(n13023) );
  NAND2HSV0 U14810 ( .A1(\pe5/aot [3]), .A2(\pe5/bq[5] ), .ZN(n13022) );
  XOR2HSV0 U14811 ( .A1(n13023), .A2(n13022), .Z(n13024) );
  XOR2HSV0 U14812 ( .A1(n13025), .A2(n13024), .Z(n13031) );
  NAND2HSV0 U14813 ( .A1(\pe5/aot [1]), .A2(\pe5/bq[6] ), .ZN(n13293) );
  NAND2HSV0 U14814 ( .A1(\pe5/aot [2]), .A2(\pe5/bq[7] ), .ZN(n13413) );
  NOR2HSV0 U14815 ( .A1(n13293), .A2(n13413), .ZN(n13027) );
  AOI22HSV0 U14816 ( .A1(\pe5/aot [2]), .A2(\pe5/bq[6] ), .B1(\pe5/bq[7] ), 
        .B2(\pe5/aot [1]), .ZN(n13026) );
  NOR2HSV2 U14817 ( .A1(n13027), .A2(n13026), .ZN(n13029) );
  NAND2HSV0 U14818 ( .A1(\pe5/aot [7]), .A2(\pe5/bq[1] ), .ZN(n13028) );
  XOR2HSV0 U14819 ( .A1(n13029), .A2(n13028), .Z(n13030) );
  XNOR2HSV1 U14820 ( .A1(n13031), .A2(n13030), .ZN(n13032) );
  INHSV1 U14821 ( .I(\pe5/got [6]), .ZN(n13280) );
  CLKAND2HSV2 U14822 ( .A1(n13034), .A2(\pe6/got [3]), .Z(n13056) );
  NAND2HSV0 U14823 ( .A1(\pe6/bq[1] ), .A2(\pe6/aot [8]), .ZN(n13036) );
  NAND2HSV0 U14824 ( .A1(\pe6/aot [5]), .A2(\pe6/bq[4] ), .ZN(n13035) );
  XOR2HSV0 U14825 ( .A1(n13036), .A2(n13035), .Z(n13040) );
  NAND2HSV0 U14826 ( .A1(\pe6/aot [6]), .A2(\pe6/bq[3] ), .ZN(n13038) );
  NAND2HSV0 U14827 ( .A1(\pe6/aot [7]), .A2(\pe6/bq[2] ), .ZN(n13037) );
  XOR2HSV0 U14828 ( .A1(n13038), .A2(n13037), .Z(n13039) );
  XOR2HSV0 U14829 ( .A1(n13040), .A2(n13039), .Z(n13054) );
  CLKNAND2HSV1 U14830 ( .A1(n13041), .A2(\pe6/pq ), .ZN(n13043) );
  XOR2HSV0 U14831 ( .A1(n13043), .A2(n13042), .Z(n13047) );
  NAND2HSV0 U14832 ( .A1(\pe6/aot [1]), .A2(\pe6/bq[8] ), .ZN(n13045) );
  NAND2HSV0 U14833 ( .A1(\pe6/aot [2]), .A2(\pe6/bq[7] ), .ZN(n13044) );
  XOR2HSV0 U14834 ( .A1(n13045), .A2(n13044), .Z(n13046) );
  XOR2HSV0 U14835 ( .A1(n13047), .A2(n13046), .Z(n13051) );
  XOR2HSV0 U14836 ( .A1(n13049), .A2(n13048), .Z(n13050) );
  XNOR2HSV1 U14837 ( .A1(n13051), .A2(n13050), .ZN(n13053) );
  CLKNAND2HSV0 U14838 ( .A1(n14895), .A2(\pe6/got [2]), .ZN(n13052) );
  XOR3HSV2 U14839 ( .A1(n13054), .A2(n13053), .A3(n13052), .Z(n13055) );
  NAND2HSV0 U14840 ( .A1(n13057), .A2(\pe6/got [4]), .ZN(n13058) );
  NOR2HSV2 U14841 ( .A1(n14489), .A2(n13059), .ZN(n13084) );
  NAND2HSV0 U14842 ( .A1(n15195), .A2(\pe14/got [5]), .ZN(n13082) );
  NAND2HSV1 U14843 ( .A1(\pe14/bq[7] ), .A2(\pe14/aot [2]), .ZN(n13555) );
  NAND2HSV0 U14844 ( .A1(n14518), .A2(\pe14/aot [3]), .ZN(n13060) );
  XOR2HSV0 U14845 ( .A1(n13555), .A2(n13060), .Z(n13076) );
  NAND2HSV0 U14846 ( .A1(\pe14/got [1]), .A2(n5968), .ZN(n13062) );
  NAND2HSV0 U14847 ( .A1(\pe14/aot [1]), .A2(n14505), .ZN(n13061) );
  XOR2HSV0 U14848 ( .A1(n13062), .A2(n13061), .Z(n13066) );
  CLKNAND2HSV0 U14849 ( .A1(n14891), .A2(\pe14/bq[1] ), .ZN(n13064) );
  NAND2HSV0 U14850 ( .A1(\pe14/aot [4]), .A2(\pe14/bq[5] ), .ZN(n13063) );
  XOR2HSV0 U14851 ( .A1(n13064), .A2(n13063), .Z(n13065) );
  XNOR2HSV1 U14852 ( .A1(n13066), .A2(n13065), .ZN(n13075) );
  CLKNHSV0 U14853 ( .I(n13067), .ZN(n14566) );
  NAND2HSV0 U14854 ( .A1(n14566), .A2(\pe14/pq ), .ZN(n13069) );
  NAND2HSV0 U14855 ( .A1(\pe14/bq[2] ), .A2(n14706), .ZN(n13068) );
  XOR2HSV0 U14856 ( .A1(n13069), .A2(n13068), .Z(n13073) );
  NAND2HSV0 U14857 ( .A1(n14889), .A2(\pe14/bq[3] ), .ZN(n13071) );
  NAND2HSV0 U14858 ( .A1(\pe14/bq[4] ), .A2(\pe14/aot [5]), .ZN(n13070) );
  XOR2HSV0 U14859 ( .A1(n13071), .A2(n13070), .Z(n13072) );
  XOR2HSV0 U14860 ( .A1(n13073), .A2(n13072), .Z(n13074) );
  XOR3HSV2 U14861 ( .A1(n13076), .A2(n13075), .A3(n13074), .Z(n13077) );
  XNOR2HSV1 U14862 ( .A1(n13078), .A2(n13077), .ZN(n13079) );
  XNOR2HSV1 U14863 ( .A1(n13080), .A2(n13079), .ZN(n13081) );
  XOR2HSV0 U14864 ( .A1(n13082), .A2(n13081), .Z(n13083) );
  XOR2HSV0 U14865 ( .A1(n13084), .A2(n13083), .Z(n13088) );
  XNOR2HSV4 U14866 ( .A1(n13091), .A2(n13090), .ZN(po14) );
  NOR2HSV2 U14867 ( .A1(n13761), .A2(n13776), .ZN(n13099) );
  NAND2HSV0 U14868 ( .A1(\pe2/aot [2]), .A2(\pe2/bq[4] ), .ZN(n13095) );
  NAND2HSV0 U14869 ( .A1(\pe2/aot [4]), .A2(\pe2/bq[2] ), .ZN(n13094) );
  XNOR2HSV1 U14870 ( .A1(n13095), .A2(n13094), .ZN(n13096) );
  AOI21HSV1 U14871 ( .A1(n13104), .A2(n13897), .B(n13103), .ZN(n13106) );
  NAND2HSV0 U14872 ( .A1(n15175), .A2(\pe21/got [5]), .ZN(n13133) );
  CLKNAND2HSV1 U14873 ( .A1(\pe21/ti_7[3] ), .A2(\pe21/got [4]), .ZN(n13131)
         );
  NAND2HSV0 U14874 ( .A1(n14538), .A2(\pe21/aot [3]), .ZN(n13109) );
  NAND2HSV0 U14875 ( .A1(\pe21/bq[7] ), .A2(\pe21/aot [2]), .ZN(n13108) );
  XOR2HSV0 U14876 ( .A1(n13109), .A2(n13108), .Z(n13113) );
  NAND2HSV0 U14877 ( .A1(\pe21/bq[3] ), .A2(\pe21/aot [6]), .ZN(n13111) );
  NAND2HSV0 U14878 ( .A1(n13834), .A2(\pe21/got [1]), .ZN(n13110) );
  XOR2HSV0 U14879 ( .A1(n13111), .A2(n13110), .Z(n13112) );
  XOR2HSV0 U14880 ( .A1(n13113), .A2(n13112), .Z(n13117) );
  CLKNAND2HSV0 U14881 ( .A1(n11786), .A2(\pe21/pq ), .ZN(n13115) );
  NAND2HSV0 U14882 ( .A1(\pe21/bq[5] ), .A2(\pe21/aot [4]), .ZN(n13114) );
  XOR2HSV0 U14883 ( .A1(n13115), .A2(n13114), .Z(n13116) );
  XNOR2HSV1 U14884 ( .A1(n13117), .A2(n13116), .ZN(n13118) );
  XNOR2HSV1 U14885 ( .A1(n13119), .A2(n13118), .ZN(n13129) );
  NAND2HSV0 U14886 ( .A1(\pe21/ti_7[1] ), .A2(\pe21/got [2]), .ZN(n13127) );
  NAND2HSV0 U14887 ( .A1(\pe21/bq[1] ), .A2(\pe21/aot [8]), .ZN(n13121) );
  NAND2HSV0 U14888 ( .A1(\pe21/bq[8] ), .A2(\pe21/aot [1]), .ZN(n13120) );
  XOR2HSV0 U14889 ( .A1(n13121), .A2(n13120), .Z(n13125) );
  NAND2HSV0 U14890 ( .A1(\pe21/bq[2] ), .A2(\pe21/aot [7]), .ZN(n13123) );
  NAND2HSV0 U14891 ( .A1(\pe21/bq[4] ), .A2(\pe21/aot [5]), .ZN(n13122) );
  XOR2HSV0 U14892 ( .A1(n13123), .A2(n13122), .Z(n13124) );
  XOR2HSV0 U14893 ( .A1(n13125), .A2(n13124), .Z(n13126) );
  XOR2HSV0 U14894 ( .A1(n13127), .A2(n13126), .Z(n13128) );
  XOR2HSV0 U14895 ( .A1(n13129), .A2(n13128), .Z(n13130) );
  XOR2HSV0 U14896 ( .A1(n13131), .A2(n13130), .Z(n13132) );
  XOR2HSV0 U14897 ( .A1(n13133), .A2(n13132), .Z(n13134) );
  INHSV4 U14898 ( .I(n13139), .ZN(n13804) );
  AO21HSV1 U14899 ( .A1(n13143), .A2(n13142), .B(n13141), .Z(n13144) );
  NAND2HSV0 U14900 ( .A1(\pe18/ti_7[1] ), .A2(\pe18/got [2]), .ZN(n13148) );
  XNOR2HSV1 U14901 ( .A1(n13149), .A2(n13148), .ZN(n13169) );
  NAND2HSV0 U14902 ( .A1(\pe18/got [1]), .A2(n13818), .ZN(n13151) );
  INHSV2 U14903 ( .I(\pe18/bq[1] ), .ZN(n14624) );
  NAND2HSV0 U14904 ( .A1(n11988), .A2(\pe18/bq[1] ), .ZN(n13150) );
  XOR2HSV0 U14905 ( .A1(n13151), .A2(n13150), .Z(n13167) );
  NAND2HSV0 U14906 ( .A1(\pe18/aot [7]), .A2(\pe18/bq[2] ), .ZN(n13152) );
  XOR2HSV0 U14907 ( .A1(n13153), .A2(n13152), .Z(n13158) );
  NAND2HSV0 U14908 ( .A1(\pe18/aot [1]), .A2(n14513), .ZN(n14632) );
  NOR2HSV0 U14909 ( .A1(n13154), .A2(n14632), .ZN(n13156) );
  AOI22HSV0 U14910 ( .A1(\pe18/aot [2]), .A2(n14513), .B1(n14511), .B2(
        \pe18/aot [1]), .ZN(n13155) );
  NOR2HSV2 U14911 ( .A1(n13156), .A2(n13155), .ZN(n13157) );
  XNOR2HSV1 U14912 ( .A1(n13158), .A2(n13157), .ZN(n13166) );
  NAND2HSV0 U14913 ( .A1(n14894), .A2(\pe18/bq[3] ), .ZN(n13160) );
  NAND2HSV0 U14914 ( .A1(\pe18/aot [5]), .A2(\pe18/bq[4] ), .ZN(n13159) );
  XOR2HSV0 U14915 ( .A1(n13160), .A2(n13159), .Z(n13164) );
  NAND2HSV0 U14916 ( .A1(\pe18/bq[5] ), .A2(\pe18/aot [4]), .ZN(n13162) );
  NAND2HSV0 U14917 ( .A1(\pe18/aot [3]), .A2(\pe18/bq[6] ), .ZN(n13161) );
  XOR2HSV0 U14918 ( .A1(n13162), .A2(n13161), .Z(n13163) );
  XOR2HSV0 U14919 ( .A1(n13164), .A2(n13163), .Z(n13165) );
  XOR3HSV2 U14920 ( .A1(n13167), .A2(n13166), .A3(n13165), .Z(n13168) );
  XNOR2HSV1 U14921 ( .A1(n13169), .A2(n13168), .ZN(n13170) );
  XNOR2HSV1 U14922 ( .A1(n13171), .A2(n13170), .ZN(n13172) );
  XNOR2HSV1 U14923 ( .A1(n13173), .A2(n13172), .ZN(n13174) );
  XOR2HSV0 U14924 ( .A1(n13175), .A2(n13174), .Z(n13179) );
  NAND2HSV4 U14925 ( .A1(n13177), .A2(n13176), .ZN(n14669) );
  NAND2HSV0 U14926 ( .A1(n14669), .A2(\pe18/got [7]), .ZN(n13180) );
  CLKNHSV0 U14927 ( .I(n13180), .ZN(n13178) );
  CLKNAND2HSV1 U14928 ( .A1(n13179), .A2(n13178), .ZN(n13183) );
  INHSV1 U14929 ( .I(n13179), .ZN(n13181) );
  CLKNAND2HSV1 U14930 ( .A1(n13181), .A2(n13180), .ZN(n13182) );
  CLKNAND2HSV1 U14931 ( .A1(n13183), .A2(n13182), .ZN(n13187) );
  AOI21HSV4 U14932 ( .A1(n13185), .A2(n13255), .B(n13184), .ZN(n13186) );
  OAI21HSV4 U14933 ( .A1(n15226), .A2(n8956), .B(n13188), .ZN(n14298) );
  CLKNHSV0 U14934 ( .I(n14298), .ZN(\pe16/ti_7[7] ) );
  NOR2HSV2 U14935 ( .A1(n14364), .A2(n13189), .ZN(n13204) );
  INHSV3 U14936 ( .I(n13191), .ZN(n14350) );
  INHSV2 U14937 ( .I(\pe16/got [1]), .ZN(n13378) );
  NOR2HSV2 U14938 ( .A1(n14350), .A2(n13378), .ZN(n13198) );
  NAND2HSV0 U14939 ( .A1(\pe16/aot [4]), .A2(\pe16/bq[1] ), .ZN(n13193) );
  NAND2HSV0 U14940 ( .A1(\pe16/aot [1]), .A2(\pe16/bq[4] ), .ZN(n13192) );
  XOR2HSV0 U14941 ( .A1(n13193), .A2(n13192), .Z(n13196) );
  CLKNAND2HSV0 U14942 ( .A1(\pe16/aot [3]), .A2(\pe16/bq[2] ), .ZN(n14351) );
  NAND2HSV0 U14943 ( .A1(\pe16/aot [2]), .A2(\pe16/bq[3] ), .ZN(n13194) );
  XOR2HSV0 U14944 ( .A1(n14351), .A2(n13194), .Z(n13195) );
  XOR2HSV0 U14945 ( .A1(n13196), .A2(n13195), .Z(n13197) );
  XOR2HSV0 U14946 ( .A1(n13198), .A2(n13197), .Z(n13199) );
  CLKNAND2HSV1 U14947 ( .A1(n14835), .A2(\pe16/got [2]), .ZN(n13201) );
  XNOR2HSV4 U14948 ( .A1(n13202), .A2(n13201), .ZN(n13203) );
  XNOR2HSV4 U14949 ( .A1(n13204), .A2(n13203), .ZN(\pe16/poht [4]) );
  CLKAND2HSV1 U14950 ( .A1(n14827), .A2(\pe16/got [4]), .Z(n13225) );
  CLKNAND2HSV0 U14951 ( .A1(\pe16/ti_7[3] ), .A2(\pe16/got [3]), .ZN(n13223)
         );
  NAND2HSV0 U14952 ( .A1(\pe16/aot [7]), .A2(\pe16/bq[1] ), .ZN(n13206) );
  NAND2HSV0 U14953 ( .A1(n14932), .A2(\pe16/bq[2] ), .ZN(n13205) );
  XOR2HSV0 U14954 ( .A1(n13206), .A2(n13205), .Z(n13210) );
  NAND2HSV0 U14955 ( .A1(\pe16/bq[3] ), .A2(\pe16/aot [5]), .ZN(n13208) );
  NAND2HSV0 U14956 ( .A1(\pe16/aot [4]), .A2(\pe16/bq[4] ), .ZN(n13207) );
  XOR2HSV0 U14957 ( .A1(n13208), .A2(n13207), .Z(n13209) );
  XOR2HSV0 U14958 ( .A1(n13210), .A2(n13209), .Z(n13216) );
  NAND2HSV0 U14959 ( .A1(\pe16/aot [1]), .A2(n6004), .ZN(n14274) );
  NAND2HSV0 U14960 ( .A1(\pe16/aot [3]), .A2(\pe16/bq[5] ), .ZN(n13213) );
  CLKNAND2HSV1 U14961 ( .A1(\pe16/aot [1]), .A2(\pe16/bq[5] ), .ZN(n14353) );
  NOR2HSV0 U14962 ( .A1(n13211), .A2(n14353), .ZN(n13212) );
  AOI21HSV2 U14963 ( .A1(n14274), .A2(n13213), .B(n13212), .ZN(n13214) );
  XOR2HSV0 U14964 ( .A1(n13214), .A2(n14083), .Z(n13215) );
  XNOR2HSV1 U14965 ( .A1(n13216), .A2(n13215), .ZN(n13218) );
  NAND2HSV0 U14966 ( .A1(\pe16/ti_7[1] ), .A2(\pe16/got [1]), .ZN(n13217) );
  XOR2HSV0 U14967 ( .A1(n13218), .A2(n13217), .Z(n13221) );
  NAND2HSV0 U14968 ( .A1(n13219), .A2(\pe16/got [2]), .ZN(n13220) );
  XNOR2HSV1 U14969 ( .A1(n13221), .A2(n13220), .ZN(n13222) );
  XNOR2HSV1 U14970 ( .A1(n13223), .A2(n13222), .ZN(n13224) );
  XOR2HSV0 U14971 ( .A1(n13225), .A2(n13224), .Z(n13228) );
  NAND2HSV0 U14972 ( .A1(n14293), .A2(\pe16/got [5]), .ZN(n13226) );
  NOR2HSV2 U14973 ( .A1(n14298), .A2(n13229), .ZN(n13230) );
  XOR2HSV0 U14974 ( .A1(n13231), .A2(n13230), .Z(\pe16/poht [1]) );
  NAND2HSV0 U14975 ( .A1(\pe15/aot [4]), .A2(\pe15/bq[1] ), .ZN(n13233) );
  NAND2HSV0 U14976 ( .A1(\pe15/aot [2]), .A2(\pe15/bq[3] ), .ZN(n13232) );
  NAND2HSV0 U14977 ( .A1(\pe15/aot [3]), .A2(\pe15/bq[2] ), .ZN(n13235) );
  NAND2HSV0 U14978 ( .A1(\pe15/aot [1]), .A2(\pe15/bq[4] ), .ZN(n13234) );
  CLKNAND2HSV0 U14979 ( .A1(\pe17/ti_7[3] ), .A2(\pe17/got [1]), .ZN(n13245)
         );
  NAND2HSV0 U14980 ( .A1(\pe17/aot [2]), .A2(\pe17/bq[4] ), .ZN(n13243) );
  NAND2HSV0 U14981 ( .A1(\pe17/aot [1]), .A2(\pe17/bq[5] ), .ZN(n14017) );
  NAND2HSV2 U14982 ( .A1(\pe17/aot [1]), .A2(\pe17/bq[1] ), .ZN(n13270) );
  NAND2HSV0 U14983 ( .A1(\pe17/aot [4]), .A2(\pe17/bq[2] ), .ZN(n13240) );
  NAND2HSV0 U14984 ( .A1(\pe17/aot [3]), .A2(\pe17/bq[3] ), .ZN(n13239) );
  XOR2HSV0 U14985 ( .A1(n13240), .A2(n13239), .Z(n13241) );
  XOR3HSV2 U14986 ( .A1(n13243), .A2(n13242), .A3(n13241), .Z(n13244) );
  XNOR2HSV1 U14987 ( .A1(n13245), .A2(n13244), .ZN(n13247) );
  XOR2HSV0 U14988 ( .A1(n13247), .A2(n13246), .Z(n13248) );
  XNOR2HSV4 U14989 ( .A1(n13249), .A2(n13248), .ZN(n13251) );
  CLKNAND2HSV1 U14990 ( .A1(n14824), .A2(\pe17/got [3]), .ZN(n13250) );
  XNOR2HSV4 U14991 ( .A1(n13251), .A2(n13250), .ZN(n13254) );
  INHSV2 U14992 ( .I(\pe17/got [5]), .ZN(n14398) );
  NOR2HSV2 U14993 ( .A1(n13261), .A2(n14398), .ZN(n13253) );
  XNOR2HSV4 U14994 ( .A1(n13254), .A2(n13253), .ZN(\pe17/poht [3]) );
  INHSV2 U14995 ( .I(n13761), .ZN(\pe2/ti_7[3] ) );
  NOR2HSV2 U14996 ( .A1(n13261), .A2(n14400), .ZN(n13267) );
  NAND2HSV0 U14997 ( .A1(\pe17/aot [1]), .A2(\pe17/bq[2] ), .ZN(n13263) );
  NAND2HSV0 U14998 ( .A1(\pe17/bq[1] ), .A2(\pe17/aot [2]), .ZN(n13262) );
  XOR2HSV0 U14999 ( .A1(n13263), .A2(n13262), .Z(n13264) );
  XOR2HSV0 U15000 ( .A1(n13265), .A2(n13264), .Z(n13266) );
  XNOR2HSV1 U15001 ( .A1(n13267), .A2(n13266), .ZN(\pe17/poht [6]) );
  XNOR2HSV1 U15002 ( .A1(n13271), .A2(n13270), .ZN(\pe17/poht [7]) );
  NAND2HSV0 U15003 ( .A1(\pe1/aot [3]), .A2(\pe1/bq[1] ), .ZN(n13273) );
  NAND2HSV0 U15004 ( .A1(\pe1/aot [2]), .A2(\pe1/bq[2] ), .ZN(n13272) );
  XOR2HSV0 U15005 ( .A1(n13273), .A2(n13272), .Z(n13274) );
  CLKNAND2HSV1 U15006 ( .A1(\pe1/aot [1]), .A2(\pe1/bq[3] ), .ZN(n13992) );
  XNOR2HSV1 U15007 ( .A1(n13274), .A2(n13992), .ZN(n13277) );
  CLKNAND2HSV1 U15008 ( .A1(n14006), .A2(\pe1/got [1]), .ZN(n13276) );
  CLKNAND2HSV0 U15009 ( .A1(\pe1/ti_7[6] ), .A2(\pe1/got [2]), .ZN(n13275) );
  XOR3HSV2 U15010 ( .A1(n13277), .A2(n13276), .A3(n13275), .Z(n13279) );
  CLKNAND2HSV1 U15011 ( .A1(n8947), .A2(\pe1/got [3]), .ZN(n13278) );
  XNOR2HSV1 U15012 ( .A1(n13279), .A2(n13278), .ZN(\pe1/poht [5]) );
  CLKNHSV0 U15013 ( .I(\pe5/ti_7t [7]), .ZN(n13281) );
  AOI21HSV2 U15014 ( .A1(n13281), .A2(n13283), .B(n13280), .ZN(n13282) );
  OAI21HSV4 U15015 ( .A1(n15275), .A2(n13283), .B(n13282), .ZN(n13311) );
  CLKNAND2HSV1 U15016 ( .A1(n13406), .A2(\pe5/got [4]), .ZN(n13303) );
  NAND2HSV0 U15017 ( .A1(n14916), .A2(\pe5/got [2]), .ZN(n13299) );
  NAND2HSV0 U15018 ( .A1(n14952), .A2(\pe5/got [1]), .ZN(n13297) );
  NAND2HSV0 U15019 ( .A1(\pe5/aot [5]), .A2(\pe5/bq[2] ), .ZN(n13287) );
  NAND2HSV0 U15020 ( .A1(\pe5/aot [6]), .A2(\pe5/bq[1] ), .ZN(n13286) );
  XOR2HSV0 U15021 ( .A1(n13287), .A2(n13286), .Z(n13292) );
  NAND2HSV0 U15022 ( .A1(\pe5/aot [2]), .A2(\pe5/bq[5] ), .ZN(n13289) );
  CLKNAND2HSV0 U15023 ( .A1(\pe5/aot [2]), .A2(\pe5/bq[3] ), .ZN(n13385) );
  NAND2HSV0 U15024 ( .A1(\pe5/bq[5] ), .A2(\pe5/aot [4]), .ZN(n13414) );
  NOR2HSV0 U15025 ( .A1(n13385), .A2(n13414), .ZN(n13288) );
  AOI21HSV1 U15026 ( .A1(n13290), .A2(n13289), .B(n13288), .ZN(n13291) );
  XNOR2HSV1 U15027 ( .A1(n13292), .A2(n13291), .ZN(n13295) );
  NAND2HSV0 U15028 ( .A1(\pe5/aot [3]), .A2(\pe5/bq[4] ), .ZN(n13386) );
  XOR2HSV0 U15029 ( .A1(n13386), .A2(n13293), .Z(n13294) );
  XNOR2HSV1 U15030 ( .A1(n13295), .A2(n13294), .ZN(n13296) );
  XOR2HSV0 U15031 ( .A1(n13297), .A2(n13296), .Z(n13298) );
  XNOR2HSV1 U15032 ( .A1(n13299), .A2(n13298), .ZN(n13301) );
  AOI21HSV0 U15033 ( .A1(n12780), .A2(\pe5/got [3]), .B(n13301), .ZN(n13300)
         );
  AOI31HSV0 U15034 ( .A1(\pe5/got [3]), .A2(n6922), .A3(n13301), .B(n13300), 
        .ZN(n13302) );
  OAI21HSV4 U15035 ( .A1(n13306), .A2(n13305), .B(n13304), .ZN(n13401) );
  CLKNHSV0 U15036 ( .I(\pe5/got [5]), .ZN(n13307) );
  CLKNAND2HSV0 U15037 ( .A1(\pe19/aot [3]), .A2(\pe19/bq[1] ), .ZN(n13313) );
  NAND2HSV0 U15038 ( .A1(\pe19/aot [2]), .A2(\pe19/bq[2] ), .ZN(n13312) );
  XNOR2HSV1 U15039 ( .A1(n13313), .A2(n13312), .ZN(n13314) );
  CLKNAND2HSV1 U15040 ( .A1(n12148), .A2(\pe19/got [3]), .ZN(n13335) );
  NAND2HSV0 U15041 ( .A1(n13317), .A2(\pe19/bq[3] ), .ZN(n13319) );
  NAND2HSV0 U15042 ( .A1(n14576), .A2(\pe19/aot [1]), .ZN(n13318) );
  XOR2HSV0 U15043 ( .A1(n13319), .A2(n13318), .Z(n13323) );
  NAND2HSV0 U15044 ( .A1(\pe19/aot [4]), .A2(\pe19/bq[4] ), .ZN(n13321) );
  NAND2HSV0 U15045 ( .A1(n14542), .A2(\pe19/aot [2]), .ZN(n13320) );
  XOR2HSV0 U15046 ( .A1(n13321), .A2(n13320), .Z(n13322) );
  XOR2HSV0 U15047 ( .A1(n13323), .A2(n13322), .Z(n13329) );
  NAND2HSV0 U15048 ( .A1(n14945), .A2(\pe19/bq[1] ), .ZN(n13325) );
  NAND2HSV0 U15049 ( .A1(\pe19/aot [3]), .A2(\pe19/bq[5] ), .ZN(n13324) );
  XOR2HSV0 U15050 ( .A1(n13325), .A2(n13324), .Z(n13327) );
  NAND2HSV0 U15051 ( .A1(\pe19/aot [6]), .A2(\pe19/bq[2] ), .ZN(n13326) );
  XNOR2HSV1 U15052 ( .A1(n13327), .A2(n13326), .ZN(n13328) );
  XNOR2HSV1 U15053 ( .A1(n13329), .A2(n13328), .ZN(n13331) );
  NAND2HSV0 U15054 ( .A1(\pe19/ti_7[1] ), .A2(\pe19/got [1]), .ZN(n13330) );
  XOR2HSV0 U15055 ( .A1(n13331), .A2(n13330), .Z(n13333) );
  NAND2HSV0 U15056 ( .A1(n11777), .A2(\pe19/got [2]), .ZN(n13332) );
  XNOR2HSV1 U15057 ( .A1(n13333), .A2(n13332), .ZN(n13334) );
  NAND2HSV2 U15058 ( .A1(\pe5/ti_7[7] ), .A2(\pe5/got [1]), .ZN(n13340) );
  AND2HSV2 U15059 ( .A1(\pe5/aot [1]), .A2(\pe5/bq[1] ), .Z(n13339) );
  XNOR2HSV1 U15060 ( .A1(n13340), .A2(n13339), .ZN(\pe5/poht [7]) );
  NAND2HSV2 U15061 ( .A1(n15168), .A2(\pe18/got [5]), .ZN(n13369) );
  NOR2HSV4 U15062 ( .A1(n13344), .A2(n13341), .ZN(n13347) );
  CLKNHSV0 U15063 ( .I(\pe18/got [4]), .ZN(n13345) );
  CLKNAND2HSV1 U15064 ( .A1(n14851), .A2(\pe18/got [3]), .ZN(n13350) );
  AOI21HSV2 U15065 ( .A1(n13351), .A2(n13350), .B(n13349), .ZN(n13367) );
  NAND2HSV0 U15066 ( .A1(n14894), .A2(\pe18/bq[1] ), .ZN(n13353) );
  NAND2HSV0 U15067 ( .A1(\pe18/aot [5]), .A2(\pe18/bq[2] ), .ZN(n13352) );
  XOR2HSV0 U15068 ( .A1(n13353), .A2(n13352), .Z(n13357) );
  NAND2HSV0 U15069 ( .A1(\pe18/aot [4]), .A2(\pe18/bq[3] ), .ZN(n13355) );
  NAND2HSV0 U15070 ( .A1(\pe18/aot [3]), .A2(\pe18/bq[4] ), .ZN(n13354) );
  XOR2HSV0 U15071 ( .A1(n13355), .A2(n13354), .Z(n13356) );
  XOR2HSV0 U15072 ( .A1(n13357), .A2(n13356), .Z(n13361) );
  NAND2HSV0 U15073 ( .A1(\pe18/aot [1]), .A2(\pe18/bq[6] ), .ZN(n13359) );
  NAND2HSV0 U15074 ( .A1(\pe18/aot [2]), .A2(\pe18/bq[5] ), .ZN(n13358) );
  XOR2HSV0 U15075 ( .A1(n13359), .A2(n13358), .Z(n13360) );
  XNOR2HSV1 U15076 ( .A1(n13361), .A2(n13360), .ZN(n13362) );
  XOR2HSV0 U15077 ( .A1(n13363), .A2(n13362), .Z(n13364) );
  XOR2HSV0 U15078 ( .A1(n13365), .A2(n13364), .Z(n13366) );
  CLKXOR2HSV2 U15079 ( .A1(n13367), .A2(n13366), .Z(n13368) );
  INHSV2 U15080 ( .I(\pe16/got [2]), .ZN(n14349) );
  NAND2HSV1 U15081 ( .A1(n14069), .A2(\pe16/got [1]), .ZN(n13375) );
  CLKNAND2HSV1 U15082 ( .A1(\pe16/aot [1]), .A2(\pe16/bq[2] ), .ZN(n13373) );
  NAND2HSV0 U15083 ( .A1(\pe16/aot [2]), .A2(\pe16/bq[1] ), .ZN(n13372) );
  XOR2HSV0 U15084 ( .A1(n13373), .A2(n13372), .Z(n13374) );
  XOR2HSV0 U15085 ( .A1(n13375), .A2(n13374), .Z(n13376) );
  XNOR2HSV1 U15086 ( .A1(n13377), .A2(n13376), .ZN(\pe16/poht [6]) );
  NOR2HSV2 U15087 ( .A1(n14298), .A2(n13378), .ZN(n13380) );
  NAND2HSV0 U15088 ( .A1(\pe16/aot [1]), .A2(\pe16/bq[1] ), .ZN(n13379) );
  XNOR2HSV1 U15089 ( .A1(n13380), .A2(n13379), .ZN(\pe16/poht [7]) );
  NAND2HSV0 U15090 ( .A1(\pe5/aot [1]), .A2(\pe5/bq[4] ), .ZN(n13382) );
  NAND2HSV0 U15091 ( .A1(\pe5/aot [3]), .A2(\pe5/bq[2] ), .ZN(n13381) );
  NAND2HSV0 U15092 ( .A1(\pe5/aot [4]), .A2(\pe5/bq[1] ), .ZN(n13383) );
  XOR2HSV0 U15093 ( .A1(n13385), .A2(n13383), .Z(n13384) );
  NAND2HSV0 U15094 ( .A1(\pe5/aot [4]), .A2(\pe5/bq[2] ), .ZN(n13393) );
  NOR2HSV0 U15095 ( .A1(n13386), .A2(n13385), .ZN(n13388) );
  AOI22HSV0 U15096 ( .A1(\pe5/aot [3]), .A2(\pe5/bq[3] ), .B1(\pe5/bq[4] ), 
        .B2(\pe5/aot [2]), .ZN(n13387) );
  NOR2HSV2 U15097 ( .A1(n13388), .A2(n13387), .ZN(n13392) );
  NAND2HSV0 U15098 ( .A1(\pe5/aot [5]), .A2(\pe5/bq[1] ), .ZN(n13390) );
  NAND2HSV0 U15099 ( .A1(\pe5/aot [1]), .A2(\pe5/bq[5] ), .ZN(n13389) );
  XOR2HSV0 U15100 ( .A1(n13390), .A2(n13389), .Z(n13391) );
  NAND2HSV2 U15101 ( .A1(\pe5/ti_7[7] ), .A2(\pe5/got [3]), .ZN(n13405) );
  CLKNAND2HSV1 U15102 ( .A1(n14846), .A2(\pe5/got [1]), .ZN(n13399) );
  NAND2HSV0 U15103 ( .A1(\pe5/aot [3]), .A2(\pe5/bq[1] ), .ZN(n13395) );
  NAND2HSV0 U15104 ( .A1(\pe5/aot [1]), .A2(\pe5/bq[3] ), .ZN(n13394) );
  XOR2HSV0 U15105 ( .A1(n13395), .A2(n13394), .Z(n13397) );
  NAND2HSV0 U15106 ( .A1(\pe5/aot [2]), .A2(\pe5/bq[2] ), .ZN(n13396) );
  XNOR2HSV1 U15107 ( .A1(n13397), .A2(n13396), .ZN(n13398) );
  XOR2HSV0 U15108 ( .A1(n13399), .A2(n13398), .Z(n13403) );
  CLKNHSV0 U15109 ( .I(\pe5/got [2]), .ZN(n13400) );
  NOR2HSV2 U15110 ( .A1(n13401), .A2(n13400), .ZN(n13402) );
  XNOR2HSV1 U15111 ( .A1(n13405), .A2(n13404), .ZN(\pe5/poht [5]) );
  NAND2HSV0 U15112 ( .A1(n10346), .A2(\pe5/got [2]), .ZN(n13428) );
  NAND2HSV2 U15113 ( .A1(n14952), .A2(\pe5/got [3]), .ZN(n13427) );
  NAND2HSV0 U15114 ( .A1(\pe5/pq ), .A2(\pe5/ctrq ), .ZN(n13408) );
  NAND2HSV0 U15115 ( .A1(\pe5/aot [8]), .A2(\pe5/bq[1] ), .ZN(n13407) );
  XOR2HSV0 U15116 ( .A1(n13408), .A2(n13407), .Z(n13412) );
  NAND2HSV0 U15117 ( .A1(\pe5/aot [7]), .A2(\pe5/bq[2] ), .ZN(n13410) );
  NAND2HSV0 U15118 ( .A1(\pe5/aot [6]), .A2(\pe5/bq[3] ), .ZN(n13409) );
  XOR2HSV0 U15119 ( .A1(n13410), .A2(n13409), .Z(n13411) );
  XOR2HSV0 U15120 ( .A1(n13412), .A2(n13411), .Z(n13416) );
  XOR2HSV0 U15121 ( .A1(n13414), .A2(n13413), .Z(n13415) );
  XNOR2HSV1 U15122 ( .A1(n13416), .A2(n13415), .ZN(n13425) );
  NAND2HSV0 U15123 ( .A1(\pe5/aot [3]), .A2(\pe5/bq[6] ), .ZN(n13418) );
  NAND2HSV0 U15124 ( .A1(\pe5/got [1]), .A2(\pe5/ti_1 ), .ZN(n13417) );
  XOR2HSV0 U15125 ( .A1(n13418), .A2(n13417), .Z(n13423) );
  NAND2HSV0 U15126 ( .A1(n13419), .A2(\pe5/aot [1]), .ZN(n13421) );
  NAND2HSV0 U15127 ( .A1(\pe5/bq[4] ), .A2(\pe5/aot [5]), .ZN(n13420) );
  XOR2HSV0 U15128 ( .A1(n13421), .A2(n13420), .Z(n13422) );
  XOR2HSV0 U15129 ( .A1(n13423), .A2(n13422), .Z(n13424) );
  XNOR2HSV1 U15130 ( .A1(n13425), .A2(n13424), .ZN(n13426) );
  NAND2HSV2 U15131 ( .A1(n14957), .A2(\pe2/got [2]), .ZN(n13435) );
  CLKNAND2HSV1 U15132 ( .A1(\pe2/aot [1]), .A2(\pe2/bq[2] ), .ZN(n13431) );
  NAND2HSV0 U15133 ( .A1(\pe2/aot [2]), .A2(\pe2/bq[1] ), .ZN(n13430) );
  XOR2HSV0 U15134 ( .A1(n13431), .A2(n13430), .Z(n13432) );
  XNOR2HSV1 U15135 ( .A1(n13435), .A2(n13434), .ZN(\pe2/poht [6]) );
  NOR2HSV2 U15136 ( .A1(n13476), .A2(n13899), .ZN(n13443) );
  NAND2HSV0 U15137 ( .A1(\pe10/bq[2] ), .A2(\pe10/aot [3]), .ZN(n13437) );
  NAND2HSV0 U15138 ( .A1(\pe10/aot [2]), .A2(\pe10/bq[3] ), .ZN(n13436) );
  XOR2HSV0 U15139 ( .A1(n13437), .A2(n13436), .Z(n13441) );
  NAND2HSV0 U15140 ( .A1(\pe10/aot [4]), .A2(\pe10/bq[1] ), .ZN(n13439) );
  NAND2HSV0 U15141 ( .A1(\pe10/aot [1]), .A2(\pe10/bq[4] ), .ZN(n13438) );
  XOR2HSV0 U15142 ( .A1(n13439), .A2(n13438), .Z(n13440) );
  XOR2HSV0 U15143 ( .A1(n13441), .A2(n13440), .Z(n13442) );
  NAND2HSV0 U15144 ( .A1(\pe10/ti_7[5] ), .A2(\pe10/got [2]), .ZN(n13444) );
  XOR2HSV0 U15145 ( .A1(n13445), .A2(n13444), .Z(n13447) );
  NAND2HSV0 U15146 ( .A1(\pe10/ti_7[6] ), .A2(\pe10/got [3]), .ZN(n13446) );
  XOR2HSV0 U15147 ( .A1(n13447), .A2(n13446), .Z(n13448) );
  CLKNHSV0 U15148 ( .I(\pe10/got [3]), .ZN(n13449) );
  NOR2HSV2 U15149 ( .A1(n13476), .A2(n13449), .ZN(n13465) );
  NAND2HSV0 U15150 ( .A1(n14132), .A2(\pe10/got [2]), .ZN(n13463) );
  NAND2HSV0 U15151 ( .A1(\pe10/aot [2]), .A2(\pe10/bq[5] ), .ZN(n13451) );
  NAND2HSV0 U15152 ( .A1(\pe10/aot [1]), .A2(\pe10/bq[6] ), .ZN(n13450) );
  XOR2HSV0 U15153 ( .A1(n13451), .A2(n13450), .Z(n13455) );
  NAND2HSV0 U15154 ( .A1(n14133), .A2(\pe10/bq[1] ), .ZN(n13453) );
  NAND2HSV0 U15155 ( .A1(\pe10/aot [5]), .A2(\pe10/bq[2] ), .ZN(n13452) );
  XOR2HSV0 U15156 ( .A1(n13453), .A2(n13452), .Z(n13454) );
  XOR2HSV0 U15157 ( .A1(n13455), .A2(n13454), .Z(n13459) );
  NAND2HSV0 U15158 ( .A1(\pe10/aot [3]), .A2(\pe10/bq[4] ), .ZN(n13457) );
  NAND2HSV0 U15159 ( .A1(\pe10/aot [4]), .A2(\pe10/bq[3] ), .ZN(n13456) );
  XOR2HSV0 U15160 ( .A1(n13457), .A2(n13456), .Z(n13458) );
  XNOR2HSV1 U15161 ( .A1(n13459), .A2(n13458), .ZN(n13460) );
  XOR2HSV0 U15162 ( .A1(n13461), .A2(n13460), .Z(n13462) );
  XOR2HSV0 U15163 ( .A1(n13463), .A2(n13462), .Z(n13464) );
  NAND2HSV0 U15164 ( .A1(\pe10/aot [2]), .A2(\pe10/bq[4] ), .ZN(n13475) );
  NAND2HSV0 U15165 ( .A1(\pe10/aot [3]), .A2(\pe10/bq[3] ), .ZN(n13470) );
  NAND2HSV0 U15166 ( .A1(\pe10/aot [1]), .A2(\pe10/bq[5] ), .ZN(n13469) );
  XOR2HSV0 U15167 ( .A1(n13470), .A2(n13469), .Z(n13474) );
  NAND2HSV0 U15168 ( .A1(\pe10/aot [5]), .A2(\pe10/bq[1] ), .ZN(n13472) );
  NAND2HSV0 U15169 ( .A1(\pe10/aot [4]), .A2(\pe10/bq[2] ), .ZN(n13471) );
  XOR2HSV0 U15170 ( .A1(n13472), .A2(n13471), .Z(n13473) );
  NAND2HSV2 U15171 ( .A1(n15091), .A2(\pe8/got [3]), .ZN(n13485) );
  NAND2HSV0 U15172 ( .A1(n14196), .A2(\pe8/got [1]), .ZN(n13481) );
  CLKNAND2HSV0 U15173 ( .A1(\pe8/aot [2]), .A2(\pe8/bq[2] ), .ZN(n13478) );
  NAND2HSV0 U15174 ( .A1(\pe8/aot [3]), .A2(\pe8/bq[1] ), .ZN(n13477) );
  XNOR2HSV1 U15175 ( .A1(n13478), .A2(n13477), .ZN(n13479) );
  CLKNAND2HSV1 U15176 ( .A1(\pe8/aot [1]), .A2(\pe8/bq[3] ), .ZN(n13519) );
  XOR2HSV0 U15177 ( .A1(n13479), .A2(n13519), .Z(n13480) );
  XNOR2HSV1 U15178 ( .A1(n13481), .A2(n13480), .ZN(n13483) );
  AOI21HSV0 U15179 ( .A1(n15182), .A2(\pe8/got [2]), .B(n13483), .ZN(n13482)
         );
  AOI31HSV0 U15180 ( .A1(\pe8/got [2]), .A2(n13483), .A3(n15182), .B(n13482), 
        .ZN(n13484) );
  XNOR2HSV1 U15181 ( .A1(n13485), .A2(n13484), .ZN(\pe8/poht [5]) );
  CLKNAND2HSV0 U15182 ( .A1(\pe8/aot [1]), .A2(\pe8/bq[4] ), .ZN(n14203) );
  CLKNAND2HSV0 U15183 ( .A1(\pe8/aot [2]), .A2(\pe8/bq[3] ), .ZN(n14208) );
  CLKNAND2HSV0 U15184 ( .A1(\pe8/aot [3]), .A2(\pe8/bq[2] ), .ZN(n13487) );
  NAND2HSV0 U15185 ( .A1(\pe8/aot [4]), .A2(\pe8/bq[1] ), .ZN(n13486) );
  NAND2HSV2 U15186 ( .A1(n15091), .A2(\pe8/got [7]), .ZN(n13511) );
  CLKNAND2HSV1 U15187 ( .A1(n15182), .A2(n13488), .ZN(n13509) );
  NAND2HSV2 U15188 ( .A1(n15066), .A2(\pe8/got [4]), .ZN(n13505) );
  NAND2HSV0 U15189 ( .A1(n14857), .A2(\pe8/got [3]), .ZN(n13503) );
  NAND2HSV0 U15190 ( .A1(\pe8/ti_7[1] ), .A2(\pe8/got [1]), .ZN(n13499) );
  NAND2HSV0 U15191 ( .A1(\pe8/bq[1] ), .A2(\pe8/aot [7]), .ZN(n13497) );
  NAND2HSV0 U15192 ( .A1(\pe8/aot [4]), .A2(\pe8/bq[4] ), .ZN(n13490) );
  NAND2HSV0 U15193 ( .A1(n14947), .A2(\pe8/bq[2] ), .ZN(n13489) );
  XOR2HSV0 U15194 ( .A1(n13490), .A2(n13489), .Z(n13496) );
  CLKNAND2HSV0 U15195 ( .A1(\pe8/aot [2]), .A2(\pe8/bq[5] ), .ZN(n14206) );
  AO22HSV1 U15196 ( .A1(\pe8/aot [3]), .A2(\pe8/bq[5] ), .B1(n8941), .B2(
        \pe8/aot [2]), .Z(n13491) );
  OAI21HSV0 U15197 ( .A1(n14202), .A2(n14206), .B(n13491), .ZN(n13495) );
  NAND2HSV0 U15198 ( .A1(\pe8/aot [1]), .A2(\pe8/bq[7] ), .ZN(n13493) );
  NAND2HSV0 U15199 ( .A1(n5948), .A2(\pe8/bq[3] ), .ZN(n13492) );
  XOR2HSV0 U15200 ( .A1(n13493), .A2(n13492), .Z(n13494) );
  XOR4HSV1 U15201 ( .A1(n13497), .A2(n13496), .A3(n13495), .A4(n13494), .Z(
        n13498) );
  XNOR2HSV1 U15202 ( .A1(n13499), .A2(n13498), .ZN(n13501) );
  CLKNHSV0 U15203 ( .I(n15079), .ZN(n14191) );
  NAND2HSV0 U15204 ( .A1(\pe8/got [2]), .A2(n14191), .ZN(n13500) );
  XNOR2HSV1 U15205 ( .A1(n13501), .A2(n13500), .ZN(n13502) );
  XNOR2HSV1 U15206 ( .A1(n13503), .A2(n13502), .ZN(n13504) );
  XNOR2HSV1 U15207 ( .A1(n13505), .A2(n13504), .ZN(n13507) );
  NAND2HSV0 U15208 ( .A1(n14196), .A2(\pe8/got [5]), .ZN(n13506) );
  XOR2HSV0 U15209 ( .A1(n13507), .A2(n13506), .Z(n13508) );
  XNOR2HSV1 U15210 ( .A1(n13511), .A2(n13510), .ZN(\pe8/poht [1]) );
  NAND2HSV2 U15211 ( .A1(n15091), .A2(\pe8/got [1]), .ZN(n13513) );
  AND2HSV1 U15212 ( .A1(\pe8/aot [1]), .A2(\pe8/bq[1] ), .Z(n13512) );
  XNOR2HSV1 U15213 ( .A1(n13513), .A2(n13512), .ZN(\pe8/poht [7]) );
  NAND2HSV0 U15214 ( .A1(\pe8/aot [4]), .A2(\pe8/bq[5] ), .ZN(n14209) );
  XOR2HSV0 U15215 ( .A1(n14202), .A2(n14209), .Z(n13530) );
  CLKNAND2HSV0 U15216 ( .A1(n14572), .A2(\pe8/pq ), .ZN(n13515) );
  NAND2HSV0 U15217 ( .A1(n14950), .A2(\pe8/bq[1] ), .ZN(n13514) );
  XOR2HSV0 U15218 ( .A1(n13515), .A2(n13514), .Z(n13521) );
  CLKNHSV0 U15219 ( .I(\pe8/aot [1]), .ZN(n14200) );
  IOA22HSV0 U15220 ( .B1(n14200), .B2(n13516), .A1(n14947), .A2(\pe8/bq[3] ), 
        .ZN(n13517) );
  OAI21HSV0 U15221 ( .A1(n13519), .A2(n13518), .B(n13517), .ZN(n13520) );
  XNOR2HSV1 U15222 ( .A1(n13521), .A2(n13520), .ZN(n13529) );
  NAND2HSV0 U15223 ( .A1(n11571), .A2(\pe8/got [1]), .ZN(n13523) );
  NAND2HSV0 U15224 ( .A1(\pe8/aot [2]), .A2(\pe8/bq[7] ), .ZN(n13522) );
  XOR2HSV0 U15225 ( .A1(n13523), .A2(n13522), .Z(n13527) );
  NAND2HSV0 U15226 ( .A1(\pe8/bq[2] ), .A2(\pe8/aot [7]), .ZN(n13525) );
  NAND2HSV0 U15227 ( .A1(n5948), .A2(\pe8/bq[4] ), .ZN(n13524) );
  XOR2HSV0 U15228 ( .A1(n13525), .A2(n13524), .Z(n13526) );
  XOR2HSV0 U15229 ( .A1(n13527), .A2(n13526), .Z(n13528) );
  NAND2HSV0 U15230 ( .A1(\pe8/ti_7[1] ), .A2(\pe8/got [2]), .ZN(n13531) );
  NAND2HSV2 U15231 ( .A1(n15091), .A2(\pe8/got [5]), .ZN(n13551) );
  INHSV2 U15232 ( .I(n13532), .ZN(n13534) );
  NAND2HSV2 U15233 ( .A1(n13534), .A2(n14197), .ZN(n13537) );
  NAND3HSV2 U15234 ( .A1(n13535), .A2(n13534), .A3(n13533), .ZN(n13536) );
  NAND3HSV2 U15235 ( .A1(n13538), .A2(n13537), .A3(n13536), .ZN(n13549) );
  NAND2HSV0 U15236 ( .A1(n15066), .A2(\pe8/got [2]), .ZN(n13547) );
  NAND2HSV0 U15237 ( .A1(n14857), .A2(\pe8/got [1]), .ZN(n13545) );
  NAND2HSV0 U15238 ( .A1(n5948), .A2(\pe8/bq[1] ), .ZN(n13543) );
  NAND2HSV0 U15239 ( .A1(\pe8/aot [4]), .A2(\pe8/bq[2] ), .ZN(n13540) );
  NAND2HSV0 U15240 ( .A1(\pe8/aot [3]), .A2(\pe8/bq[3] ), .ZN(n13539) );
  XOR2HSV0 U15241 ( .A1(n13540), .A2(n13539), .Z(n13541) );
  XOR3HSV2 U15242 ( .A1(n13543), .A2(n13542), .A3(n13541), .Z(n13544) );
  XNOR2HSV1 U15243 ( .A1(n13545), .A2(n13544), .ZN(n13546) );
  XNOR2HSV1 U15244 ( .A1(n13547), .A2(n13546), .ZN(n13548) );
  XNOR2HSV1 U15245 ( .A1(n13551), .A2(n13550), .ZN(\pe8/poht [3]) );
  NAND2HSV2 U15246 ( .A1(n14855), .A2(\pe14/got [6]), .ZN(n13579) );
  MUX2NHSV1 U15247 ( .I0(n15236), .I1(\pe14/ti_7t [5]), .S(n14702), .ZN(n13806) );
  NAND2HSV0 U15248 ( .A1(n15195), .A2(\pe14/got [4]), .ZN(n13576) );
  NOR2HSV0 U15249 ( .A1(n13555), .A2(n13554), .ZN(n13557) );
  AOI22HSV0 U15250 ( .A1(\pe14/aot [2]), .A2(\pe14/bq[6] ), .B1(\pe14/bq[7] ), 
        .B2(\pe14/aot [1]), .ZN(n13556) );
  NOR2HSV2 U15251 ( .A1(n13557), .A2(n13556), .ZN(n13559) );
  NAND2HSV0 U15252 ( .A1(\pe14/aot [4]), .A2(\pe14/bq[4] ), .ZN(n13558) );
  XOR2HSV0 U15253 ( .A1(n13559), .A2(n13558), .Z(n13570) );
  NAND2HSV0 U15254 ( .A1(\pe14/bq[3] ), .A2(\pe14/aot [5]), .ZN(n13562) );
  NAND2HSV0 U15255 ( .A1(\pe14/bq[1] ), .A2(\pe14/aot [7]), .ZN(n13561) );
  XOR2HSV0 U15256 ( .A1(n13562), .A2(n13561), .Z(n13566) );
  NAND2HSV0 U15257 ( .A1(\pe14/aot [3]), .A2(\pe14/bq[5] ), .ZN(n13564) );
  NAND2HSV0 U15258 ( .A1(n14889), .A2(\pe14/bq[2] ), .ZN(n13563) );
  XOR2HSV0 U15259 ( .A1(n13564), .A2(n13563), .Z(n13565) );
  XOR2HSV0 U15260 ( .A1(n13566), .A2(n13565), .Z(n13569) );
  NOR2HSV1 U15261 ( .A1(n13853), .A2(n13567), .ZN(n13568) );
  XOR3HSV2 U15262 ( .A1(n13570), .A2(n13569), .A3(n13568), .Z(n13572) );
  NAND2HSV0 U15263 ( .A1(n14944), .A2(\pe14/got [2]), .ZN(n13571) );
  XOR2HSV0 U15264 ( .A1(n13572), .A2(n13571), .Z(n13573) );
  XOR2HSV0 U15265 ( .A1(n13574), .A2(n13573), .Z(n13575) );
  XOR2HSV0 U15266 ( .A1(n13576), .A2(n13575), .Z(n13577) );
  AOI21HSV2 U15267 ( .A1(n13581), .A2(n13582), .B(n13580), .ZN(n13585) );
  AOI22HSV0 U15268 ( .A1(n13585), .A2(n13584), .B1(n13583), .B2(\pe14/got [7]), 
        .ZN(n13586) );
  NAND2HSV2 U15269 ( .A1(\pe13/aot [4]), .A2(\pe13/bq[5] ), .ZN(n13589) );
  NAND2HSV0 U15270 ( .A1(\pe13/aot [3]), .A2(\pe13/bq[6] ), .ZN(n13588) );
  XOR2HSV0 U15271 ( .A1(n13589), .A2(n13588), .Z(n13601) );
  NAND2HSV0 U15272 ( .A1(\pe13/aot [5]), .A2(\pe13/bq[4] ), .ZN(n13594) );
  NAND2HSV0 U15273 ( .A1(\pe13/got [1]), .A2(n13819), .ZN(n13593) );
  XOR2HSV0 U15274 ( .A1(n13594), .A2(n13593), .Z(n13598) );
  NAND2HSV0 U15275 ( .A1(\pe13/aot [6]), .A2(\pe13/bq[3] ), .ZN(n13596) );
  NAND2HSV0 U15276 ( .A1(\pe13/aot [1]), .A2(\pe13/bq[8] ), .ZN(n13595) );
  XOR2HSV0 U15277 ( .A1(n13596), .A2(n13595), .Z(n13597) );
  XOR2HSV0 U15278 ( .A1(n13598), .A2(n13597), .Z(n13599) );
  CLKNHSV0 U15279 ( .I(\pe7/got [3]), .ZN(n13617) );
  NAND2HSV0 U15280 ( .A1(\pe7/bq[1] ), .A2(\pe7/aot [7]), .ZN(n13607) );
  NAND2HSV0 U15281 ( .A1(\pe7/aot [5]), .A2(\pe7/bq[3] ), .ZN(n13606) );
  CLKNAND2HSV0 U15282 ( .A1(n13607), .A2(n13606), .ZN(n13608) );
  OAI21HSV0 U15283 ( .A1(n13610), .A2(n13609), .B(n13608), .ZN(n13612) );
  NAND2HSV0 U15284 ( .A1(\pe7/bq[2] ), .A2(\pe7/aot [6]), .ZN(n13611) );
  XNOR2HSV1 U15285 ( .A1(n13612), .A2(n13611), .ZN(n13616) );
  NAND2HSV0 U15286 ( .A1(\pe7/aot [4]), .A2(\pe7/bq[4] ), .ZN(n13614) );
  NAND2HSV0 U15287 ( .A1(\pe7/aot [1]), .A2(\pe7/bq[7] ), .ZN(n13613) );
  XNOR2HSV1 U15288 ( .A1(n13614), .A2(n13613), .ZN(n13615) );
  NAND2HSV0 U15289 ( .A1(\pe7/aot [2]), .A2(n8930), .ZN(n13618) );
  NAND2HSV0 U15290 ( .A1(n13624), .A2(n13620), .ZN(n13622) );
  BUFHSV2 U15291 ( .I(n13621), .Z(n13625) );
  NOR2HSV2 U15292 ( .A1(n13622), .A2(n13625), .ZN(n13633) );
  CLKNHSV0 U15293 ( .I(n13633), .ZN(n13631) );
  NOR2HSV0 U15294 ( .A1(n13624), .A2(n13623), .ZN(n13626) );
  CLKAND2HSV2 U15295 ( .A1(n13626), .A2(n13625), .Z(n13634) );
  CLKNHSV1 U15296 ( .I(n13634), .ZN(n13630) );
  CLKNHSV0 U15297 ( .I(n13627), .ZN(n13628) );
  NAND2HSV0 U15298 ( .A1(n13628), .A2(\pe7/got [5]), .ZN(n13632) );
  CLKNHSV0 U15299 ( .I(n13632), .ZN(n13629) );
  NAND3HSV2 U15300 ( .A1(n13631), .A2(n13630), .A3(n13629), .ZN(n13636) );
  NOR3HSV2 U15301 ( .A1(n13634), .A2(n13633), .A3(n13632), .ZN(n13635) );
  NAND2HSV0 U15302 ( .A1(n15189), .A2(\pe7/got [6]), .ZN(n13637) );
  CLKNHSV0 U15303 ( .I(\pe20/got [3]), .ZN(n13639) );
  NOR2HSV2 U15304 ( .A1(n13640), .A2(n13639), .ZN(n13651) );
  CLKNHSV1 U15305 ( .I(n13651), .ZN(n13644) );
  CLKNHSV0 U15306 ( .I(n13641), .ZN(n13643) );
  CLKNHSV0 U15307 ( .I(\pe20/got [4]), .ZN(n13642) );
  NOR2HSV2 U15308 ( .A1(n13643), .A2(n13642), .ZN(n13649) );
  NAND2HSV2 U15309 ( .A1(n13644), .A2(n13649), .ZN(n13653) );
  NAND2HSV0 U15310 ( .A1(n9459), .A2(n13645), .ZN(n13646) );
  CLKNHSV1 U15311 ( .I(n13646), .ZN(n13648) );
  INHSV2 U15312 ( .I(n13650), .ZN(n13652) );
  CLKNAND2HSV0 U15313 ( .A1(n11854), .A2(\pe20/got [2]), .ZN(n13666) );
  NAND2HSV0 U15314 ( .A1(n6026), .A2(\pe20/got [1]), .ZN(n13665) );
  NAND2HSV0 U15315 ( .A1(\pe20/aot [3]), .A2(\pe20/bq[4] ), .ZN(n13655) );
  NAND2HSV0 U15316 ( .A1(\pe20/aot [1]), .A2(\pe20/bq[6] ), .ZN(n13654) );
  XOR2HSV0 U15317 ( .A1(n13655), .A2(n13654), .Z(n13659) );
  NAND2HSV0 U15318 ( .A1(\pe20/aot [4]), .A2(\pe20/bq[3] ), .ZN(n13657) );
  NAND2HSV0 U15319 ( .A1(\pe20/aot [2]), .A2(\pe20/bq[5] ), .ZN(n13656) );
  XOR2HSV0 U15320 ( .A1(n13657), .A2(n13656), .Z(n13658) );
  XOR2HSV0 U15321 ( .A1(n13659), .A2(n13658), .Z(n13663) );
  NAND2HSV0 U15322 ( .A1(n14946), .A2(\pe20/bq[1] ), .ZN(n13661) );
  NAND2HSV0 U15323 ( .A1(\pe20/aot [5]), .A2(\pe20/bq[2] ), .ZN(n13660) );
  XOR2HSV0 U15324 ( .A1(n13661), .A2(n13660), .Z(n13662) );
  XNOR2HSV1 U15325 ( .A1(n13663), .A2(n13662), .ZN(n13664) );
  NAND2HSV0 U15326 ( .A1(n15184), .A2(\pe20/got [1]), .ZN(n13674) );
  NAND2HSV0 U15327 ( .A1(\pe20/aot [2]), .A2(\pe20/bq[3] ), .ZN(n13668) );
  NAND2HSV0 U15328 ( .A1(\pe20/aot [1]), .A2(\pe20/bq[4] ), .ZN(n13667) );
  XOR2HSV0 U15329 ( .A1(n13668), .A2(n13667), .Z(n13672) );
  NAND2HSV0 U15330 ( .A1(\pe20/aot [3]), .A2(\pe20/bq[2] ), .ZN(n13670) );
  NAND2HSV0 U15331 ( .A1(\pe20/aot [4]), .A2(\pe20/bq[1] ), .ZN(n13669) );
  XOR2HSV0 U15332 ( .A1(n13670), .A2(n13669), .Z(n13671) );
  XOR2HSV0 U15333 ( .A1(n13672), .A2(n13671), .Z(n13673) );
  XOR2HSV0 U15334 ( .A1(n13674), .A2(n13673), .Z(n13675) );
  INHSV1 U15335 ( .I(\pe20/got [2]), .ZN(n13692) );
  NOR2HSV4 U15336 ( .A1(n13751), .A2(n13692), .ZN(n13678) );
  NAND2HSV0 U15337 ( .A1(\pe20/aot [2]), .A2(\pe20/bq[2] ), .ZN(n13680) );
  NAND2HSV0 U15338 ( .A1(\pe20/aot [1]), .A2(\pe20/bq[3] ), .ZN(n13679) );
  NAND2HSV0 U15339 ( .A1(\pe20/aot [2]), .A2(\pe20/bq[4] ), .ZN(n13689) );
  NAND2HSV0 U15340 ( .A1(\pe20/aot [4]), .A2(\pe20/bq[2] ), .ZN(n13684) );
  NAND2HSV0 U15341 ( .A1(\pe20/aot [1]), .A2(\pe20/bq[5] ), .ZN(n13683) );
  XNOR2HSV1 U15342 ( .A1(n13684), .A2(n13683), .ZN(n13688) );
  NAND2HSV0 U15343 ( .A1(\pe20/aot [5]), .A2(\pe20/bq[1] ), .ZN(n13686) );
  NAND2HSV0 U15344 ( .A1(\pe20/aot [3]), .A2(\pe20/bq[3] ), .ZN(n13685) );
  XOR2HSV0 U15345 ( .A1(n13686), .A2(n13685), .Z(n13687) );
  XOR3HSV2 U15346 ( .A1(n13689), .A2(n13688), .A3(n13687), .Z(n13690) );
  XNOR2HSV1 U15347 ( .A1(n13691), .A2(n13690), .ZN(n13694) );
  CLKNHSV0 U15348 ( .I(n13694), .ZN(n13693) );
  NAND2HSV0 U15349 ( .A1(n13695), .A2(\pe20/got [4]), .ZN(n13715) );
  CLKNAND2HSV0 U15350 ( .A1(n11854), .A2(\pe20/got [3]), .ZN(n13713) );
  CLKNAND2HSV0 U15351 ( .A1(n13737), .A2(\pe20/aot [1]), .ZN(n13697) );
  NAND2HSV0 U15352 ( .A1(\pe20/bq[1] ), .A2(n8937), .ZN(n13696) );
  XOR2HSV0 U15353 ( .A1(n13697), .A2(n13696), .Z(n13701) );
  CLKNAND2HSV0 U15354 ( .A1(n14946), .A2(\pe20/bq[2] ), .ZN(n13699) );
  NAND2HSV0 U15355 ( .A1(\pe20/aot [5]), .A2(\pe20/bq[3] ), .ZN(n13698) );
  XOR2HSV0 U15356 ( .A1(n13699), .A2(n13698), .Z(n13700) );
  XOR2HSV0 U15357 ( .A1(n13701), .A2(n13700), .Z(n13707) );
  NAND2HSV0 U15358 ( .A1(\pe20/aot [4]), .A2(\pe20/bq[4] ), .ZN(n13703) );
  NAND2HSV0 U15359 ( .A1(\pe20/aot [2]), .A2(\pe20/bq[6] ), .ZN(n13702) );
  XOR2HSV0 U15360 ( .A1(n13703), .A2(n13702), .Z(n13705) );
  NAND2HSV0 U15361 ( .A1(\pe20/aot [3]), .A2(\pe20/bq[5] ), .ZN(n13704) );
  XNOR2HSV1 U15362 ( .A1(n13705), .A2(n13704), .ZN(n13706) );
  XNOR2HSV1 U15363 ( .A1(n13707), .A2(n13706), .ZN(n13709) );
  XOR2HSV0 U15364 ( .A1(n13709), .A2(n13708), .Z(n13711) );
  NAND2HSV0 U15365 ( .A1(n6026), .A2(\pe20/got [2]), .ZN(n13710) );
  XNOR2HSV1 U15366 ( .A1(n13711), .A2(n13710), .ZN(n13712) );
  XOR2HSV0 U15367 ( .A1(n13713), .A2(n13712), .Z(n13714) );
  XOR2HSV0 U15368 ( .A1(n13715), .A2(n13714), .Z(n13716) );
  CLKNAND2HSV1 U15369 ( .A1(\pe20/ti_7[5] ), .A2(\pe20/got [5]), .ZN(n13717)
         );
  CLKNAND2HSV0 U15370 ( .A1(n11854), .A2(\pe20/got [4]), .ZN(n13748) );
  NAND2HSV0 U15371 ( .A1(n6026), .A2(\pe20/got [3]), .ZN(n13722) );
  XNOR2HSV1 U15372 ( .A1(n13722), .A2(n13721), .ZN(n13746) );
  CLKNAND2HSV0 U15373 ( .A1(\pe20/pq ), .A2(n12362), .ZN(n13724) );
  NAND2HSV0 U15374 ( .A1(\pe20/aot [7]), .A2(\pe20/bq[2] ), .ZN(n13723) );
  XOR2HSV0 U15375 ( .A1(n13724), .A2(n13723), .Z(n13728) );
  NAND2HSV0 U15376 ( .A1(\pe20/aot [5]), .A2(\pe20/bq[4] ), .ZN(n13726) );
  NAND2HSV0 U15377 ( .A1(\pe20/aot [4]), .A2(\pe20/bq[5] ), .ZN(n13725) );
  XOR2HSV0 U15378 ( .A1(n13726), .A2(n13725), .Z(n13727) );
  XOR2HSV0 U15379 ( .A1(n13728), .A2(n13727), .Z(n13732) );
  NAND2HSV0 U15380 ( .A1(\pe20/aot [3]), .A2(\pe20/bq[6] ), .ZN(n13730) );
  NAND2HSV0 U15381 ( .A1(n14946), .A2(\pe20/bq[3] ), .ZN(n13729) );
  XOR2HSV0 U15382 ( .A1(n13730), .A2(n13729), .Z(n13731) );
  XNOR2HSV1 U15383 ( .A1(n13732), .A2(n13731), .ZN(n13744) );
  CLKNAND2HSV0 U15384 ( .A1(n13733), .A2(\pe20/bq[1] ), .ZN(n13736) );
  NAND2HSV0 U15385 ( .A1(\pe20/aot [1]), .A2(n13734), .ZN(n13735) );
  XOR2HSV0 U15386 ( .A1(n13736), .A2(n13735), .Z(n13742) );
  NAND2HSV0 U15387 ( .A1(n13737), .A2(\pe20/aot [2]), .ZN(n13740) );
  NAND2HSV0 U15388 ( .A1(\pe20/got [1]), .A2(n13738), .ZN(n13739) );
  XOR2HSV0 U15389 ( .A1(n13740), .A2(n13739), .Z(n13741) );
  XOR2HSV0 U15390 ( .A1(n13742), .A2(n13741), .Z(n13743) );
  XNOR2HSV1 U15391 ( .A1(n13744), .A2(n13743), .ZN(n13745) );
  XOR2HSV0 U15392 ( .A1(n13746), .A2(n13745), .Z(n13747) );
  CLKNHSV0 U15393 ( .I(\pe20/got [6]), .ZN(n13750) );
  NAND2HSV0 U15394 ( .A1(\pe11/aot [2]), .A2(\pe11/bq[3] ), .ZN(n13754) );
  NAND2HSV0 U15395 ( .A1(\pe11/aot [1]), .A2(\pe11/bq[4] ), .ZN(n13753) );
  XOR2HSV0 U15396 ( .A1(n13754), .A2(n13753), .Z(n13758) );
  NAND2HSV0 U15397 ( .A1(\pe11/aot [3]), .A2(\pe11/bq[2] ), .ZN(n13756) );
  NAND2HSV0 U15398 ( .A1(\pe11/aot [4]), .A2(\pe11/bq[1] ), .ZN(n13755) );
  XOR2HSV0 U15399 ( .A1(n13756), .A2(n13755), .Z(n13757) );
  CLKNHSV0 U15400 ( .I(\pe2/bq[8] ), .ZN(n13763) );
  INHSV2 U15401 ( .I(n13763), .ZN(n14559) );
  NAND2HSV0 U15402 ( .A1(\pe2/aot [1]), .A2(n14559), .ZN(n13765) );
  NAND2HSV0 U15403 ( .A1(\pe2/aot [7]), .A2(\pe2/bq[2] ), .ZN(n13764) );
  XOR2HSV0 U15404 ( .A1(n13765), .A2(n13764), .Z(n13783) );
  INHSV2 U15405 ( .I(n13766), .ZN(n14523) );
  NAND2HSV0 U15406 ( .A1(n14858), .A2(\pe2/bq[1] ), .ZN(n13767) );
  XOR2HSV0 U15407 ( .A1(n13768), .A2(n13767), .Z(n13772) );
  NAND2HSV0 U15408 ( .A1(\pe2/aot [4]), .A2(\pe2/bq[5] ), .ZN(n13770) );
  NAND2HSV0 U15409 ( .A1(\pe2/aot [3]), .A2(n14510), .ZN(n13769) );
  XOR2HSV0 U15410 ( .A1(n13770), .A2(n13769), .Z(n13771) );
  XNOR2HSV1 U15411 ( .A1(n13772), .A2(n13771), .ZN(n13782) );
  NAND2HSV0 U15412 ( .A1(\pe2/aot [6]), .A2(\pe2/bq[3] ), .ZN(n13774) );
  NAND2HSV0 U15413 ( .A1(\pe2/aot [5]), .A2(\pe2/bq[4] ), .ZN(n13773) );
  XOR2HSV0 U15414 ( .A1(n13774), .A2(n13773), .Z(n13780) );
  NOR2HSV0 U15415 ( .A1(n13776), .A2(n13775), .ZN(n13778) );
  NAND2HSV0 U15416 ( .A1(\pe2/aot [2]), .A2(n14504), .ZN(n13777) );
  XOR2HSV0 U15417 ( .A1(n13778), .A2(n13777), .Z(n13779) );
  XOR2HSV0 U15418 ( .A1(n13780), .A2(n13779), .Z(n13781) );
  XOR3HSV2 U15419 ( .A1(n13783), .A2(n13782), .A3(n13781), .Z(n13784) );
  NAND2HSV2 U15420 ( .A1(n14487), .A2(n10459), .ZN(n13787) );
  INHSV2 U15421 ( .I(n14055), .ZN(n13786) );
  CLKNAND2HSV1 U15422 ( .A1(n8947), .A2(\pe1/got [2]), .ZN(n13793) );
  CLKNAND2HSV1 U15423 ( .A1(\pe1/ti_7[6] ), .A2(\pe1/got [1]), .ZN(n13791) );
  CLKNAND2HSV1 U15424 ( .A1(\pe1/aot [2]), .A2(\pe1/bq[1] ), .ZN(n13789) );
  NAND2HSV0 U15425 ( .A1(\pe1/aot [1]), .A2(\pe1/bq[2] ), .ZN(n13788) );
  XOR2HSV0 U15426 ( .A1(n13789), .A2(n13788), .Z(n13790) );
  XNOR2HSV1 U15427 ( .A1(n13791), .A2(n13790), .ZN(n13792) );
  XNOR2HSV1 U15428 ( .A1(n13793), .A2(n13792), .ZN(\pe1/poht [6]) );
  NAND2HSV0 U15429 ( .A1(\pe21/ti_7[1] ), .A2(n13797), .ZN(n13798) );
  NOR2HSV2 U15430 ( .A1(n13799), .A2(n13801), .ZN(n13800) );
  XOR2HSV0 U15431 ( .A1(n13800), .A2(poh21[2]), .Z(po[3]) );
  XOR2HSV0 U15432 ( .A1(n13802), .A2(poh21[3]), .Z(po[4]) );
  OAI21HSV0 U15433 ( .A1(n13805), .A2(n13804), .B(n13803), .ZN(n15216) );
  CLKNHSV0 U15434 ( .I(n13806), .ZN(\pe14/ti_7[5] ) );
  NOR2HSV2 U15435 ( .A1(n13808), .A2(n13807), .ZN(n14688) );
  CLKNHSV0 U15436 ( .I(n14688), .ZN(\pe18/ti_7[5] ) );
  CLKNHSV0 U15437 ( .I(n13809), .ZN(n15193) );
  CLKNHSV0 U15438 ( .I(n14310), .ZN(\pe17/ti_7[7] ) );
  BUFHSV2 U15439 ( .I(n14812), .Z(n15173) );
  BUFHSV2 U15440 ( .I(n14721), .Z(n15094) );
  BUFHSV2 U15441 ( .I(n15094), .Z(n15174) );
  INHSV2 U15442 ( .I(\pe5/pq ), .ZN(n13814) );
  MUX2NHSV1 U15443 ( .I0(n13814), .I1(n10316), .S(n11818), .ZN(\pe5/ti_1t ) );
  INHSV2 U15444 ( .I(\pe14/pq ), .ZN(n13817) );
  CLKNHSV0 U15445 ( .I(n5968), .ZN(n13816) );
  MUX2NHSV1 U15446 ( .I0(n13817), .I1(n13816), .S(n14742), .ZN(\pe14/ti_1t )
         );
  MUX2NHSV1 U15447 ( .I0(bo4[8]), .I1(n13823), .S(n13822), .ZN(n15103) );
  MUX2NHSV1 U15448 ( .I0(bo8[7]), .I1(n13825), .S(n14758), .ZN(n15129) );
  MUX2NHSV1 U15449 ( .I0(bo6[6]), .I1(n13827), .S(n13828), .ZN(n15115) );
  MUX2NHSV1 U15450 ( .I0(bo6[8]), .I1(n13829), .S(n13828), .ZN(n15114) );
  INHSV2 U15451 ( .I(n14415), .ZN(n13837) );
  INHSV2 U15452 ( .I(\pe17/pq ), .ZN(n13836) );
  CLKNHSV0 U15453 ( .I(\pe17/ctrq ), .ZN(n14404) );
  INHSV2 U15454 ( .I(n14571), .ZN(n13835) );
  MUX2NHSV1 U15455 ( .I0(n13837), .I1(n13836), .S(n13835), .ZN(\pe17/ti_1t )
         );
  NAND2HSV0 U15456 ( .A1(n10242), .A2(\pe1/got [8]), .ZN(n13839) );
  XOR2HSV0 U15457 ( .A1(n13839), .A2(n13838), .Z(pov1[2]) );
  NAND2HSV0 U15458 ( .A1(n5949), .A2(n15180), .ZN(n13843) );
  XOR2HSV0 U15459 ( .A1(n13843), .A2(n13842), .Z(n15289) );
  NAND2HSV0 U15460 ( .A1(\pe19/ti_7[1] ), .A2(n13844), .ZN(n13846) );
  XNOR2HSV1 U15461 ( .A1(n13846), .A2(n13845), .ZN(n15213) );
  NAND2HSV0 U15462 ( .A1(\pe12/ti_7[1] ), .A2(n5958), .ZN(n13850) );
  XNOR2HSV1 U15463 ( .A1(n13850), .A2(n13849), .ZN(n15252) );
  CLKNAND2HSV0 U15464 ( .A1(n15072), .A2(n15178), .ZN(n13858) );
  XOR2HSV0 U15465 ( .A1(n13858), .A2(n13857), .Z(n15234) );
  XNOR2HSV1 U15466 ( .A1(n13860), .A2(n6702), .ZN(n15295) );
  CLKNAND2HSV0 U15467 ( .A1(n14857), .A2(\pe8/got [8]), .ZN(n13863) );
  XOR2HSV0 U15468 ( .A1(n13863), .A2(n13862), .Z(n15266) );
  BUFHSV2 U15469 ( .I(n13865), .Z(n13866) );
  XNOR2HSV1 U15470 ( .A1(n13867), .A2(n13866), .ZN(\pov15[4] ) );
  MUX2NHSV1 U15471 ( .I0(n6730), .I1(n13881), .S(n13880), .ZN(n15281) );
  XOR2HSV0 U15472 ( .A1(n13883), .A2(n6714), .Z(n15270) );
  NAND2HSV0 U15473 ( .A1(\pe1/ti_7[5] ), .A2(\pe1/got [8]), .ZN(n13885) );
  XOR2HSV0 U15474 ( .A1(n13885), .A2(n13884), .Z(pov1[6]) );
  XOR2HSV0 U15475 ( .A1(n13887), .A2(n13886), .Z(n15290) );
  CLKNAND2HSV1 U15476 ( .A1(n15190), .A2(n5958), .ZN(n13896) );
  CLKNHSV0 U15477 ( .I(n13891), .ZN(n13894) );
  CLKNHSV0 U15478 ( .I(n13893), .ZN(n13892) );
  OA22HSV2 U15479 ( .A1(n13894), .A2(n13893), .B1(n13892), .B2(n13890), .Z(
        n13895) );
  XOR2HSV0 U15480 ( .A1(n13896), .A2(n13895), .Z(n15247) );
  AOI21HSV0 U15481 ( .A1(n10058), .A2(n13900), .B(n13899), .ZN(n13901) );
  NAND2HSV2 U15482 ( .A1(\pe10/bq[1] ), .A2(\pe10/aot [1]), .ZN(n13903) );
  XOR2HSV0 U15483 ( .A1(n13903), .A2(n13904), .Z(\pe10/poht [7]) );
  CLKNAND2HSV1 U15484 ( .A1(n8947), .A2(\pe1/got [1]), .ZN(n13906) );
  NAND2HSV0 U15485 ( .A1(\pe1/aot [1]), .A2(\pe1/bq[1] ), .ZN(n13905) );
  XOR2HSV0 U15486 ( .A1(n13906), .A2(n13905), .Z(\pe1/poht [7]) );
  NAND2HSV0 U15487 ( .A1(\pe4/aot [1]), .A2(\pe4/bq[1] ), .ZN(n13907) );
  NAND2HSV0 U15488 ( .A1(\pe9/aot [1]), .A2(\pe9/bq[1] ), .ZN(n13908) );
  XOR2HSV0 U15489 ( .A1(n13909), .A2(n13908), .Z(\pe9/poht [7]) );
  NAND2HSV2 U15490 ( .A1(\pe9/aot [5]), .A2(\pe9/bq[3] ), .ZN(n13913) );
  NAND2HSV0 U15491 ( .A1(n5976), .A2(\pe9/aot [1]), .ZN(n13912) );
  XOR2HSV0 U15492 ( .A1(n13913), .A2(n13912), .Z(n13917) );
  NAND2HSV0 U15493 ( .A1(\pe9/aot [3]), .A2(\pe9/bq[5] ), .ZN(n13914) );
  XOR2HSV0 U15494 ( .A1(n13915), .A2(n13914), .Z(n13916) );
  XOR2HSV0 U15495 ( .A1(n13917), .A2(n13916), .Z(n13925) );
  CLKNHSV0 U15496 ( .I(n13918), .ZN(n13921) );
  AOI22HSV0 U15497 ( .A1(\pe9/bq[1] ), .A2(\pe9/aot [7]), .B1(\pe9/bq[4] ), 
        .B2(\pe9/aot [4]), .ZN(n13919) );
  AOI21HSV0 U15498 ( .A1(n13921), .A2(n7021), .B(n13919), .ZN(n13923) );
  XOR2HSV0 U15499 ( .A1(n13923), .A2(n13922), .Z(n13924) );
  XNOR2HSV1 U15500 ( .A1(n13925), .A2(n13924), .ZN(n13927) );
  NAND2HSV0 U15501 ( .A1(\pe9/ti_7[1] ), .A2(\pe9/got [1]), .ZN(n13926) );
  XOR2HSV0 U15502 ( .A1(n13927), .A2(n13926), .Z(n13929) );
  NAND2HSV0 U15503 ( .A1(n14896), .A2(\pe9/got [2]), .ZN(n13928) );
  CLKNHSV0 U15504 ( .I(\pe9/got [6]), .ZN(n13930) );
  CLKNAND2HSV1 U15505 ( .A1(\pe6/aot [1]), .A2(\pe6/bq[2] ), .ZN(n13933) );
  NAND2HSV0 U15506 ( .A1(\pe6/aot [2]), .A2(\pe6/bq[1] ), .ZN(n13932) );
  XOR2HSV0 U15507 ( .A1(n13933), .A2(n13932), .Z(n13934) );
  NAND2HSV2 U15508 ( .A1(n14862), .A2(\pe19/got [1]), .ZN(n13936) );
  CLKNAND2HSV0 U15509 ( .A1(\pe19/bq[1] ), .A2(\pe19/aot [1]), .ZN(n13935) );
  XOR2HSV0 U15510 ( .A1(n13936), .A2(n13935), .Z(\pe19/poht [7]) );
  NAND2HSV2 U15511 ( .A1(n14965), .A2(\pe11/got [1]), .ZN(n13938) );
  NAND2HSV0 U15512 ( .A1(\pe11/aot [1]), .A2(\pe11/bq[1] ), .ZN(n13937) );
  XOR2HSV0 U15513 ( .A1(n13938), .A2(n13937), .Z(\pe11/poht [7]) );
  CLKNAND2HSV1 U15514 ( .A1(n14959), .A2(\pe12/got [1]), .ZN(n13940) );
  XOR2HSV0 U15515 ( .A1(n13940), .A2(n13939), .Z(\pe12/poht [7]) );
  NAND2HSV0 U15516 ( .A1(n6027), .A2(\pe1/got [1]), .ZN(n13942) );
  XNOR2HSV1 U15517 ( .A1(n13942), .A2(n13941), .ZN(n13951) );
  NAND2HSV0 U15518 ( .A1(\pe1/aot [6]), .A2(\pe1/bq[1] ), .ZN(n13944) );
  NAND2HSV0 U15519 ( .A1(\pe1/aot [5]), .A2(\pe1/bq[2] ), .ZN(n13943) );
  XOR2HSV0 U15520 ( .A1(n13944), .A2(n13943), .Z(n13949) );
  INHSV2 U15521 ( .I(n13968), .ZN(n14581) );
  NAND2HSV0 U15522 ( .A1(n14581), .A2(\pe1/aot [2]), .ZN(n14002) );
  CLKNHSV0 U15523 ( .I(\pe1/aot [1]), .ZN(n13946) );
  OAI21HSV0 U15524 ( .A1(n13946), .A2(n13968), .B(n13945), .ZN(n13947) );
  OAI21HSV1 U15525 ( .A1(n13970), .A2(n14002), .B(n13947), .ZN(n13948) );
  XNOR2HSV1 U15526 ( .A1(n13949), .A2(n13948), .ZN(n13950) );
  XNOR2HSV1 U15527 ( .A1(n13951), .A2(n13950), .ZN(n13956) );
  CLKNHSV0 U15528 ( .I(\pe1/got [2]), .ZN(n13952) );
  NOR2HSV1 U15529 ( .A1(n13953), .A2(n13952), .ZN(n13955) );
  NAND2HSV0 U15530 ( .A1(n14847), .A2(\pe1/got [3]), .ZN(n13954) );
  XOR3HSV2 U15531 ( .A1(n13956), .A2(n13955), .A3(n13954), .Z(n13959) );
  NAND2HSV2 U15532 ( .A1(n14006), .A2(\pe1/got [4]), .ZN(n13958) );
  NAND2HSV0 U15533 ( .A1(\pe1/ti_7[6] ), .A2(\pe1/got [5]), .ZN(n13957) );
  XOR3HSV2 U15534 ( .A1(n13959), .A2(n13958), .A3(n13957), .Z(n13961) );
  NAND2HSV0 U15535 ( .A1(\pe1/ti_7[7] ), .A2(\pe1/got [6]), .ZN(n13960) );
  XOR2HSV0 U15536 ( .A1(n13961), .A2(n13960), .Z(\pe1/poht [2]) );
  NAND2HSV0 U15537 ( .A1(\pe1/aot [5]), .A2(\pe1/bq[4] ), .ZN(n13963) );
  NAND2HSV0 U15538 ( .A1(\pe1/aot [8]), .A2(\pe1/bq[1] ), .ZN(n13962) );
  XOR2HSV0 U15539 ( .A1(n13963), .A2(n13962), .Z(n13967) );
  NAND2HSV0 U15540 ( .A1(\pe1/aot [2]), .A2(n8945), .ZN(n13964) );
  XOR2HSV0 U15541 ( .A1(n13965), .A2(n13964), .Z(n13966) );
  XOR2HSV0 U15542 ( .A1(n13967), .A2(n13966), .Z(n13975) );
  XNOR2HSV1 U15543 ( .A1(n13973), .A2(n13972), .ZN(n13974) );
  XNOR2HSV1 U15544 ( .A1(n13975), .A2(n13974), .ZN(n13979) );
  NAND2HSV0 U15545 ( .A1(n6027), .A2(\pe1/got [3]), .ZN(n13977) );
  NAND2HSV0 U15546 ( .A1(n10242), .A2(\pe1/got [2]), .ZN(n13976) );
  XOR2HSV0 U15547 ( .A1(n13977), .A2(n13976), .Z(n13978) );
  XNOR2HSV1 U15548 ( .A1(n13979), .A2(n13978), .ZN(n13983) );
  CLKNHSV0 U15549 ( .I(\pe1/got [4]), .ZN(n13980) );
  NOR2HSV1 U15550 ( .A1(n14005), .A2(n13980), .ZN(n13982) );
  NAND2HSV0 U15551 ( .A1(n14847), .A2(\pe1/got [5]), .ZN(n13981) );
  XOR3HSV2 U15552 ( .A1(n13983), .A2(n13982), .A3(n13981), .Z(n13986) );
  NAND2HSV2 U15553 ( .A1(n14006), .A2(\pe1/got [6]), .ZN(n13985) );
  NAND2HSV0 U15554 ( .A1(\pe1/ti_7[6] ), .A2(n14703), .ZN(n13984) );
  XOR3HSV2 U15555 ( .A1(n13986), .A2(n13985), .A3(n13984), .Z(n13988) );
  NAND2HSV0 U15556 ( .A1(\pe1/ti_7[7] ), .A2(\pe1/got [8]), .ZN(n13987) );
  XOR2HSV0 U15557 ( .A1(n13988), .A2(n13987), .Z(po1) );
  NAND2HSV0 U15558 ( .A1(\pe1/bq[5] ), .A2(\pe1/aot [3]), .ZN(n13990) );
  NAND2HSV0 U15559 ( .A1(\pe1/aot [7]), .A2(\pe1/bq[1] ), .ZN(n13989) );
  XOR2HSV0 U15560 ( .A1(n13990), .A2(n13989), .Z(n13995) );
  AO22HSV1 U15561 ( .A1(\pe1/bq[3] ), .A2(\pe1/aot [5]), .B1(n8945), .B2(
        \pe1/aot [1]), .Z(n13991) );
  OAI21HSV0 U15562 ( .A1(n13993), .A2(n13992), .B(n13991), .ZN(n13994) );
  XNOR2HSV1 U15563 ( .A1(n13995), .A2(n13994), .ZN(n13997) );
  NAND2HSV0 U15564 ( .A1(n6027), .A2(\pe1/got [2]), .ZN(n13996) );
  CLKNHSV0 U15565 ( .I(n13998), .ZN(n14001) );
  AOI22HSV0 U15566 ( .A1(\pe1/aot [6]), .A2(\pe1/bq[2] ), .B1(\pe1/bq[4] ), 
        .B2(\pe1/aot [4]), .ZN(n13999) );
  AOI21HSV0 U15567 ( .A1(n14001), .A2(n14000), .B(n13999), .ZN(n14003) );
  XOR2HSV0 U15568 ( .A1(n14003), .A2(n14002), .Z(n14004) );
  CLKNHSV0 U15569 ( .I(\pe17/ti_7t [7]), .ZN(n14009) );
  AOI21HSV0 U15570 ( .A1(n14010), .A2(n14009), .B(n14008), .ZN(n14014) );
  CLKNAND2HSV0 U15571 ( .A1(\pe17/ti_7[3] ), .A2(\pe17/got [2]), .ZN(n14028)
         );
  NAND2HSV0 U15572 ( .A1(n14399), .A2(\pe17/got [1]), .ZN(n14026) );
  NAND2HSV0 U15573 ( .A1(\pe17/aot [5]), .A2(\pe17/bq[2] ), .ZN(n14016) );
  NAND2HSV0 U15574 ( .A1(\pe17/bq[4] ), .A2(\pe17/aot [3]), .ZN(n14015) );
  XOR2HSV0 U15575 ( .A1(n14016), .A2(n14015), .Z(n14021) );
  NAND2HSV0 U15576 ( .A1(\pe17/aot [2]), .A2(\pe17/bq[6] ), .ZN(n14336) );
  NOR2HSV0 U15577 ( .A1(n14336), .A2(n14017), .ZN(n14019) );
  AOI22HSV0 U15578 ( .A1(\pe17/aot [2]), .A2(\pe17/bq[5] ), .B1(n14525), .B2(
        \pe17/aot [1]), .ZN(n14018) );
  NOR2HSV2 U15579 ( .A1(n14019), .A2(n14018), .ZN(n14020) );
  XNOR2HSV1 U15580 ( .A1(n14021), .A2(n14020), .ZN(n14024) );
  NAND2HSV0 U15581 ( .A1(\pe17/aot [4]), .A2(\pe17/bq[3] ), .ZN(n14022) );
  XOR2HSV0 U15582 ( .A1(n14409), .A2(n14022), .Z(n14023) );
  XNOR2HSV1 U15583 ( .A1(n14024), .A2(n14023), .ZN(n14025) );
  XOR2HSV0 U15584 ( .A1(n14026), .A2(n14025), .Z(n14027) );
  CLKNHSV0 U15585 ( .I(\pe7/got [2]), .ZN(n14029) );
  NAND2HSV0 U15586 ( .A1(\pe7/got [1]), .A2(n14860), .ZN(n14041) );
  NAND2HSV0 U15587 ( .A1(\pe7/aot [5]), .A2(\pe7/bq[2] ), .ZN(n14031) );
  NAND2HSV0 U15588 ( .A1(\pe7/aot [4]), .A2(\pe7/bq[3] ), .ZN(n14030) );
  XOR2HSV0 U15589 ( .A1(n14031), .A2(n14030), .Z(n14035) );
  NAND2HSV0 U15590 ( .A1(\pe7/aot [3]), .A2(\pe7/bq[4] ), .ZN(n14033) );
  NAND2HSV0 U15591 ( .A1(\pe7/aot [2]), .A2(\pe7/bq[5] ), .ZN(n14032) );
  XOR2HSV0 U15592 ( .A1(n14033), .A2(n14032), .Z(n14034) );
  XOR2HSV0 U15593 ( .A1(n14035), .A2(n14034), .Z(n14039) );
  NAND2HSV0 U15594 ( .A1(\pe7/bq[1] ), .A2(n14705), .ZN(n14037) );
  NAND2HSV0 U15595 ( .A1(\pe7/aot [1]), .A2(\pe7/bq[6] ), .ZN(n14036) );
  XOR2HSV0 U15596 ( .A1(n14037), .A2(n14036), .Z(n14038) );
  XNOR2HSV1 U15597 ( .A1(n14039), .A2(n14038), .ZN(n14040) );
  XNOR2HSV1 U15598 ( .A1(n14041), .A2(n14040), .ZN(n14042) );
  CLKNHSV0 U15599 ( .I(\pe7/got [4]), .ZN(n14464) );
  NOR2HSV2 U15600 ( .A1(n14043), .A2(n14464), .ZN(n14046) );
  AOI21HSV0 U15601 ( .A1(\pe7/ti_7[5] ), .A2(n6038), .B(n14044), .ZN(n14045)
         );
  AOI21HSV2 U15602 ( .A1(n14046), .A2(\pe7/ti_7[5] ), .B(n14045), .ZN(n14048)
         );
  NAND2HSV0 U15603 ( .A1(n14487), .A2(\pe7/got [5]), .ZN(n14047) );
  NOR2HSV0 U15604 ( .A1(n14054), .A2(n10459), .ZN(n14053) );
  NAND3HSV0 U15605 ( .A1(n15189), .A2(n5967), .A3(n14049), .ZN(n14051) );
  OA21HSV2 U15606 ( .A1(n14054), .A2(n12252), .B(\pe7/got [6]), .Z(n14050) );
  OAI21HSV2 U15607 ( .A1(n14055), .A2(n14051), .B(n14050), .ZN(n14052) );
  AOI21HSV2 U15608 ( .A1(n14055), .A2(n14053), .B(n14052), .ZN(n14058) );
  NOR2HSV2 U15609 ( .A1(n14487), .A2(n14054), .ZN(n14056) );
  CLKNAND2HSV0 U15610 ( .A1(n14056), .A2(n14055), .ZN(n14057) );
  CLKNAND2HSV1 U15611 ( .A1(n14058), .A2(n14057), .ZN(n14059) );
  XOR2HSV0 U15612 ( .A1(n14060), .A2(n14059), .Z(\pe7/poht [2]) );
  XOR2HSV0 U15613 ( .A1(n14063), .A2(n14062), .Z(\pe2/poht [7]) );
  NAND3HSV2 U15614 ( .A1(n14069), .A2(n6654), .A3(n14064), .ZN(n14077) );
  CLKNHSV0 U15615 ( .I(n6654), .ZN(n14068) );
  NAND2HSV2 U15616 ( .A1(n14069), .A2(\pe16/got [5]), .ZN(n14075) );
  AOI21HSV0 U15617 ( .A1(n14071), .A2(n8957), .B(n14070), .ZN(n14076) );
  CLKNAND2HSV0 U15618 ( .A1(n14075), .A2(n14076), .ZN(n14073) );
  AOI21HSV2 U15619 ( .A1(n14077), .A2(n14076), .B(n14075), .ZN(n14078) );
  CLKNAND2HSV1 U15620 ( .A1(n14835), .A2(\pe16/got [4]), .ZN(n14100) );
  NAND2HSV0 U15621 ( .A1(\pe16/ti_7[3] ), .A2(\pe16/got [2]), .ZN(n14095) );
  NAND2HSV0 U15622 ( .A1(n14080), .A2(\pe16/got [1]), .ZN(n14093) );
  NAND2HSV0 U15623 ( .A1(n14932), .A2(\pe16/bq[1] ), .ZN(n14082) );
  NAND2HSV0 U15624 ( .A1(\pe16/aot [5]), .A2(\pe16/bq[2] ), .ZN(n14081) );
  XOR2HSV0 U15625 ( .A1(n14082), .A2(n14081), .Z(n14088) );
  CLKNHSV0 U15626 ( .I(n14353), .ZN(n14086) );
  CLKNHSV0 U15627 ( .I(n14083), .ZN(n14085) );
  AOI22HSV0 U15628 ( .A1(\pe16/aot [2]), .A2(\pe16/bq[5] ), .B1(\pe16/bq[6] ), 
        .B2(\pe16/aot [1]), .ZN(n14084) );
  AOI21HSV2 U15629 ( .A1(n14086), .A2(n14085), .B(n14084), .ZN(n14087) );
  XNOR2HSV1 U15630 ( .A1(n14088), .A2(n14087), .ZN(n14091) );
  NAND2HSV0 U15631 ( .A1(\pe16/bq[3] ), .A2(\pe16/aot [4]), .ZN(n14352) );
  NAND2HSV0 U15632 ( .A1(\pe16/aot [3]), .A2(\pe16/bq[4] ), .ZN(n14089) );
  XOR2HSV0 U15633 ( .A1(n14352), .A2(n14089), .Z(n14090) );
  XNOR2HSV1 U15634 ( .A1(n14091), .A2(n14090), .ZN(n14092) );
  XOR2HSV0 U15635 ( .A1(n14093), .A2(n14092), .Z(n14094) );
  XOR2HSV0 U15636 ( .A1(n14095), .A2(n14094), .Z(n14098) );
  NOR2HSV2 U15637 ( .A1(n14350), .A2(n14096), .ZN(n14097) );
  XOR2HSV0 U15638 ( .A1(n14098), .A2(n14097), .Z(n14099) );
  XOR2HSV0 U15639 ( .A1(n14100), .A2(n14099), .Z(n14101) );
  XOR2HSV0 U15640 ( .A1(n14102), .A2(n14101), .Z(\pe16/poht [2]) );
  NAND2HSV0 U15641 ( .A1(\pe10/ti_7[6] ), .A2(\pe10/got [1]), .ZN(n14106) );
  CLKNAND2HSV1 U15642 ( .A1(\pe10/aot [1]), .A2(\pe10/bq[2] ), .ZN(n14104) );
  CLKNAND2HSV0 U15643 ( .A1(\pe10/bq[1] ), .A2(\pe10/aot [2]), .ZN(n14103) );
  XOR2HSV0 U15644 ( .A1(n14104), .A2(n14103), .Z(n14105) );
  XOR2HSV0 U15645 ( .A1(n14106), .A2(n14105), .Z(n14107) );
  XOR2HSV0 U15646 ( .A1(n14108), .A2(n14107), .Z(\pe10/poht [6]) );
  CLKNAND2HSV0 U15647 ( .A1(\pe10/aot [3]), .A2(\pe10/bq[1] ), .ZN(n14110) );
  NAND2HSV0 U15648 ( .A1(\pe10/aot [1]), .A2(\pe10/bq[3] ), .ZN(n14109) );
  XOR2HSV0 U15649 ( .A1(n14110), .A2(n14109), .Z(n14112) );
  NAND2HSV0 U15650 ( .A1(\pe10/aot [2]), .A2(\pe10/bq[2] ), .ZN(n14111) );
  XNOR2HSV1 U15651 ( .A1(n14112), .A2(n14111), .ZN(n14113) );
  XNOR2HSV1 U15652 ( .A1(n14114), .A2(n14113), .ZN(n14115) );
  NAND3HSV0 U15653 ( .A1(n10040), .A2(\pe10/got [5]), .A3(n15262), .ZN(n14131)
         );
  CLKNHSV0 U15654 ( .I(\pe10/got [4]), .ZN(n14118) );
  INAND2HSV0 U15655 ( .A1(n14118), .B1(n10925), .ZN(n14116) );
  CLKNHSV0 U15656 ( .I(n14116), .ZN(n14117) );
  CLKNAND2HSV0 U15657 ( .A1(n15200), .A2(n14117), .ZN(n14121) );
  NAND2HSV0 U15658 ( .A1(n14119), .A2(\pe10/got [4]), .ZN(n14120) );
  NAND2HSV2 U15659 ( .A1(n14121), .A2(n14120), .ZN(n14127) );
  NAND2HSV0 U15660 ( .A1(n14122), .A2(\pe10/got [5]), .ZN(n14123) );
  CLKNHSV1 U15661 ( .I(n14123), .ZN(n14124) );
  NOR2HSV2 U15662 ( .A1(n14127), .A2(n14124), .ZN(n14130) );
  AND2HSV2 U15663 ( .A1(n14125), .A2(\pe10/got [5]), .Z(n14126) );
  CLKNAND2HSV1 U15664 ( .A1(n14127), .A2(n14126), .ZN(n14128) );
  NAND2HSV0 U15665 ( .A1(n14132), .A2(\pe10/got [3]), .ZN(n14151) );
  NAND2HSV0 U15666 ( .A1(n14844), .A2(\pe10/bq[1] ), .ZN(n14135) );
  NAND2HSV0 U15667 ( .A1(n14133), .A2(\pe10/bq[2] ), .ZN(n14134) );
  XOR2HSV0 U15668 ( .A1(n14135), .A2(n14134), .Z(n14139) );
  NAND2HSV0 U15669 ( .A1(n14567), .A2(\pe10/aot [1]), .ZN(n14137) );
  NAND2HSV0 U15670 ( .A1(\pe10/aot [5]), .A2(\pe10/bq[3] ), .ZN(n14136) );
  XOR2HSV0 U15671 ( .A1(n14137), .A2(n14136), .Z(n14138) );
  XOR2HSV0 U15672 ( .A1(n14139), .A2(n14138), .Z(n14145) );
  NAND2HSV0 U15673 ( .A1(\pe10/bq[4] ), .A2(\pe10/aot [4]), .ZN(n14141) );
  NAND2HSV0 U15674 ( .A1(\pe10/bq[6] ), .A2(\pe10/aot [2]), .ZN(n14140) );
  XOR2HSV0 U15675 ( .A1(n14141), .A2(n14140), .Z(n14143) );
  NAND2HSV0 U15676 ( .A1(\pe10/aot [3]), .A2(\pe10/bq[5] ), .ZN(n14142) );
  XNOR2HSV1 U15677 ( .A1(n14143), .A2(n14142), .ZN(n14144) );
  XNOR2HSV1 U15678 ( .A1(n14145), .A2(n14144), .ZN(n14147) );
  NAND2HSV0 U15679 ( .A1(n6033), .A2(\pe10/got [1]), .ZN(n14146) );
  XOR2HSV0 U15680 ( .A1(n14147), .A2(n14146), .Z(n14149) );
  NAND2HSV0 U15681 ( .A1(n14940), .A2(\pe10/got [2]), .ZN(n14148) );
  XNOR2HSV1 U15682 ( .A1(n14149), .A2(n14148), .ZN(n14150) );
  XOR2HSV0 U15683 ( .A1(n14151), .A2(n14150), .Z(n14152) );
  XOR2HSV0 U15684 ( .A1(n14153), .A2(n14152), .Z(n14155) );
  XOR2HSV0 U15685 ( .A1(n14156), .A2(n14157), .Z(\pe10/poht [1]) );
  NAND2HSV0 U15686 ( .A1(n14819), .A2(\pe3/got [1]), .ZN(n14159) );
  NAND2HSV0 U15687 ( .A1(\pe3/aot [1]), .A2(\pe3/bq[1] ), .ZN(n14158) );
  XOR2HSV0 U15688 ( .A1(n14159), .A2(n14158), .Z(\pe3/poht [7]) );
  CLKNAND2HSV0 U15689 ( .A1(n14959), .A2(\pe12/got [2]), .ZN(n14165) );
  NAND2HSV0 U15690 ( .A1(n15190), .A2(\pe12/got [1]), .ZN(n14163) );
  CLKNAND2HSV1 U15691 ( .A1(\pe12/aot [1]), .A2(\pe12/bq[2] ), .ZN(n14161) );
  NAND2HSV0 U15692 ( .A1(\pe12/aot [2]), .A2(\pe12/bq[1] ), .ZN(n14160) );
  XOR2HSV0 U15693 ( .A1(n14161), .A2(n14160), .Z(n14162) );
  XOR2HSV0 U15694 ( .A1(n14163), .A2(n14162), .Z(n14164) );
  XOR2HSV0 U15695 ( .A1(n14165), .A2(n14164), .Z(\pe12/poht [6]) );
  NAND2HSV0 U15696 ( .A1(n14819), .A2(\pe3/got [2]), .ZN(n14171) );
  NAND2HSV2 U15697 ( .A1(n14941), .A2(\pe3/got [1]), .ZN(n14169) );
  CLKNAND2HSV1 U15698 ( .A1(\pe3/aot [1]), .A2(\pe3/bq[2] ), .ZN(n14167) );
  CLKNAND2HSV0 U15699 ( .A1(\pe3/bq[1] ), .A2(\pe3/aot [2]), .ZN(n14166) );
  XOR2HSV0 U15700 ( .A1(n14167), .A2(n14166), .Z(n14168) );
  XOR2HSV0 U15701 ( .A1(n14169), .A2(n14168), .Z(n14170) );
  XOR2HSV0 U15702 ( .A1(n14171), .A2(n14170), .Z(\pe3/poht [6]) );
  NAND2HSV0 U15703 ( .A1(\pe20/aot [1]), .A2(\pe20/bq[1] ), .ZN(n14172) );
  CLKNAND2HSV1 U15704 ( .A1(\pe20/aot [1]), .A2(\pe20/bq[2] ), .ZN(n14174) );
  NAND2HSV0 U15705 ( .A1(\pe20/aot [2]), .A2(\pe20/bq[1] ), .ZN(n14173) );
  XOR2HSV0 U15706 ( .A1(n14174), .A2(n14173), .Z(n14175) );
  XOR2HSV0 U15707 ( .A1(n14176), .A2(n14175), .Z(n14177) );
  XOR2HSV0 U15708 ( .A1(n14178), .A2(n14177), .Z(\pe20/poht [6]) );
  NAND2HSV0 U15709 ( .A1(\pe6/aot [1]), .A2(\pe6/bq[1] ), .ZN(n14180) );
  NAND2HSV2 U15710 ( .A1(n14683), .A2(\pe18/got [1]), .ZN(n14182) );
  NAND2HSV0 U15711 ( .A1(\pe18/aot [1]), .A2(\pe18/bq[1] ), .ZN(n14181) );
  XOR2HSV0 U15712 ( .A1(n14182), .A2(n14181), .Z(\pe18/poht [7]) );
  NAND2HSV2 U15713 ( .A1(n14683), .A2(\pe18/got [2]), .ZN(n14188) );
  NAND2HSV2 U15714 ( .A1(n14669), .A2(\pe18/got [1]), .ZN(n14186) );
  CLKNAND2HSV1 U15715 ( .A1(\pe18/aot [1]), .A2(\pe18/bq[2] ), .ZN(n14184) );
  NAND2HSV0 U15716 ( .A1(\pe18/aot [2]), .A2(\pe18/bq[1] ), .ZN(n14183) );
  XOR2HSV0 U15717 ( .A1(n14184), .A2(n14183), .Z(n14185) );
  XOR2HSV0 U15718 ( .A1(n14186), .A2(n14185), .Z(n14187) );
  XOR2HSV0 U15719 ( .A1(n14188), .A2(n14187), .Z(\pe18/poht [6]) );
  NAND2HSV0 U15720 ( .A1(n14857), .A2(\pe8/got [2]), .ZN(n14195) );
  NAND2HSV0 U15721 ( .A1(n14191), .A2(\pe8/got [1]), .ZN(n14193) );
  NAND2HSV0 U15722 ( .A1(n5948), .A2(\pe8/bq[2] ), .ZN(n14192) );
  XOR2HSV0 U15723 ( .A1(n14193), .A2(n14192), .Z(n14194) );
  CLKNHSV0 U15724 ( .I(\pe8/got [4]), .ZN(n14197) );
  INAND2HSV2 U15725 ( .A1(n14197), .B1(n14196), .ZN(n14212) );
  NAND2HSV0 U15726 ( .A1(\pe8/aot [3]), .A2(\pe8/bq[4] ), .ZN(n14198) );
  OAI21HSV1 U15727 ( .A1(n14200), .A2(n14199), .B(n14198), .ZN(n14201) );
  OAI21HSV2 U15728 ( .A1(n14203), .A2(n14202), .B(n14201), .ZN(n14205) );
  NAND2HSV0 U15729 ( .A1(n14947), .A2(\pe8/bq[1] ), .ZN(n14204) );
  XNOR2HSV1 U15730 ( .A1(n14205), .A2(n14204), .ZN(n14211) );
  NAND2HSV0 U15731 ( .A1(\pe19/aot [2]), .A2(\pe19/bq[5] ), .ZN(n14214) );
  NAND2HSV0 U15732 ( .A1(\pe19/aot [1]), .A2(\pe19/bq[6] ), .ZN(n14213) );
  XOR2HSV0 U15733 ( .A1(n14214), .A2(n14213), .Z(n14218) );
  NAND2HSV0 U15734 ( .A1(\pe19/aot [3]), .A2(\pe19/bq[4] ), .ZN(n14216) );
  NAND2HSV0 U15735 ( .A1(\pe19/aot [4]), .A2(\pe19/bq[3] ), .ZN(n14215) );
  XNOR2HSV1 U15736 ( .A1(n14216), .A2(n14215), .ZN(n14217) );
  XNOR2HSV1 U15737 ( .A1(n14218), .A2(n14217), .ZN(n14220) );
  NAND2HSV0 U15738 ( .A1(n14220), .A2(\pe19/got [3]), .ZN(n14221) );
  NAND2HSV0 U15739 ( .A1(n11777), .A2(\pe19/got [1]), .ZN(n14226) );
  NAND2HSV0 U15740 ( .A1(\pe19/aot [6]), .A2(\pe19/bq[1] ), .ZN(n14223) );
  XOR2HSV0 U15741 ( .A1(n14224), .A2(n14223), .Z(n14225) );
  NAND2HSV2 U15742 ( .A1(\pe21/got [1]), .A2(n15085), .ZN(n14228) );
  CLKNAND2HSV0 U15743 ( .A1(\pe21/bq[1] ), .A2(\pe21/aot [1]), .ZN(n14227) );
  XOR2HSV0 U15744 ( .A1(n14228), .A2(n14227), .Z(\pe21/poht [7]) );
  NAND2HSV2 U15745 ( .A1(n14852), .A2(\pe7/got [1]), .ZN(n14230) );
  NAND2HSV0 U15746 ( .A1(\pe7/aot [1]), .A2(\pe7/bq[1] ), .ZN(n14229) );
  XOR2HSV0 U15747 ( .A1(n14230), .A2(n14229), .Z(\pe7/poht [7]) );
  NAND2HSV2 U15748 ( .A1(n14449), .A2(\pe7/got [2]), .ZN(n14236) );
  NAND2HSV0 U15749 ( .A1(n14487), .A2(\pe7/got [1]), .ZN(n14234) );
  CLKNAND2HSV1 U15750 ( .A1(\pe7/aot [1]), .A2(\pe7/bq[2] ), .ZN(n14232) );
  NAND2HSV0 U15751 ( .A1(\pe7/aot [2]), .A2(\pe7/bq[1] ), .ZN(n14231) );
  XOR2HSV0 U15752 ( .A1(n14232), .A2(n14231), .Z(n14233) );
  XOR2HSV0 U15753 ( .A1(n14234), .A2(n14233), .Z(n14235) );
  XOR2HSV0 U15754 ( .A1(n14236), .A2(n14235), .Z(\pe7/poht [6]) );
  NAND2HSV0 U15755 ( .A1(\pe12/aot [6]), .A2(\pe12/bq[2] ), .ZN(n14239) );
  NAND2HSV0 U15756 ( .A1(\pe12/bq[5] ), .A2(\pe12/aot [3]), .ZN(n14238) );
  OAI21HSV0 U15757 ( .A1(n14241), .A2(n14577), .B(n14240), .ZN(n14242) );
  NAND2HSV0 U15758 ( .A1(\pe12/ti_7[1] ), .A2(\pe12/got [1]), .ZN(n14254) );
  NAND2HSV0 U15759 ( .A1(\pe12/aot [5]), .A2(\pe12/bq[3] ), .ZN(n14250) );
  NAND2HSV0 U15760 ( .A1(n14948), .A2(\pe12/bq[1] ), .ZN(n14249) );
  XOR2HSV0 U15761 ( .A1(n14250), .A2(n14249), .Z(n14252) );
  NAND2HSV0 U15762 ( .A1(\pe12/aot [2]), .A2(\pe12/bq[6] ), .ZN(n14251) );
  XNOR2HSV1 U15763 ( .A1(n14252), .A2(n14251), .ZN(n14253) );
  XNOR2HSV1 U15764 ( .A1(n14254), .A2(n14253), .ZN(n14256) );
  NAND2HSV2 U15765 ( .A1(n14830), .A2(\pe11/got [1]), .ZN(n14261) );
  NAND2HSV0 U15766 ( .A1(\pe11/aot [1]), .A2(\pe11/bq[2] ), .ZN(n14259) );
  NAND2HSV0 U15767 ( .A1(\pe11/aot [2]), .A2(\pe11/bq[1] ), .ZN(n14258) );
  XOR2HSV0 U15768 ( .A1(n14259), .A2(n14258), .Z(n14260) );
  XOR2HSV0 U15769 ( .A1(n14261), .A2(n14260), .Z(n14262) );
  XOR2HSV0 U15770 ( .A1(n14263), .A2(n14262), .Z(\pe11/poht [6]) );
  NOR2HSV2 U15771 ( .A1(n14350), .A2(n14363), .ZN(n14291) );
  CLKNAND2HSV0 U15772 ( .A1(\pe16/ti_7[3] ), .A2(\pe16/got [4]), .ZN(n14289)
         );
  NAND2HSV0 U15773 ( .A1(\pe16/ti_7[1] ), .A2(\pe16/got [2]), .ZN(n14264) );
  XNOR2HSV1 U15774 ( .A1(n14265), .A2(n14264), .ZN(n14287) );
  NAND2HSV0 U15775 ( .A1(\pe16/bq[2] ), .A2(\pe16/aot [7]), .ZN(n14268) );
  NAND2HSV0 U15776 ( .A1(\pe16/got [1]), .A2(n14266), .ZN(n14267) );
  XOR2HSV0 U15777 ( .A1(n14268), .A2(n14267), .Z(n14285) );
  CLKNAND2HSV0 U15778 ( .A1(n14743), .A2(\pe16/pq ), .ZN(n14270) );
  NAND2HSV0 U15779 ( .A1(\pe16/aot [4]), .A2(\pe16/bq[5] ), .ZN(n14269) );
  XOR2HSV0 U15780 ( .A1(n14270), .A2(n14269), .Z(n14276) );
  INHSV2 U15781 ( .I(n6004), .ZN(n14565) );
  IOA22HSV1 U15782 ( .B1(n14271), .B2(n14565), .A1(n5947), .A2(\pe16/aot [1]), 
        .ZN(n14272) );
  OAI21HSV0 U15783 ( .A1(n14274), .A2(n14273), .B(n14272), .ZN(n14275) );
  XNOR2HSV1 U15784 ( .A1(n14276), .A2(n14275), .ZN(n14284) );
  NAND2HSV0 U15785 ( .A1(\pe16/aot [3]), .A2(\pe16/bq[6] ), .ZN(n14278) );
  NAND2HSV0 U15786 ( .A1(\pe16/aot [5]), .A2(\pe16/bq[4] ), .ZN(n14277) );
  XOR2HSV0 U15787 ( .A1(n14278), .A2(n14277), .Z(n14282) );
  NAND2HSV0 U15788 ( .A1(n14932), .A2(\pe16/bq[3] ), .ZN(n14280) );
  NAND2HSV0 U15789 ( .A1(\pe16/aot [8]), .A2(\pe16/bq[1] ), .ZN(n14279) );
  XOR2HSV0 U15790 ( .A1(n14280), .A2(n14279), .Z(n14281) );
  XOR2HSV0 U15791 ( .A1(n14282), .A2(n14281), .Z(n14283) );
  XOR3HSV2 U15792 ( .A1(n14285), .A2(n14284), .A3(n14283), .Z(n14286) );
  XNOR2HSV1 U15793 ( .A1(n14287), .A2(n14286), .ZN(n14288) );
  XNOR2HSV1 U15794 ( .A1(n14289), .A2(n14288), .ZN(n14290) );
  XOR2HSV0 U15795 ( .A1(n14291), .A2(n14290), .Z(n14296) );
  NAND2HSV0 U15796 ( .A1(n14293), .A2(\pe16/got [6]), .ZN(n14294) );
  NOR2HSV2 U15797 ( .A1(n14298), .A2(n14297), .ZN(n14299) );
  XOR2HSV0 U15798 ( .A1(n14300), .A2(n14299), .Z(po16) );
  NAND2HSV2 U15799 ( .A1(n14853), .A2(\pe15/got [2]), .ZN(n14306) );
  NAND2HSV2 U15800 ( .A1(n6535), .A2(\pe15/got [1]), .ZN(n14304) );
  CLKNAND2HSV1 U15801 ( .A1(\pe15/aot [1]), .A2(\pe15/bq[2] ), .ZN(n14302) );
  NAND2HSV0 U15802 ( .A1(\pe15/aot [2]), .A2(\pe15/bq[1] ), .ZN(n14301) );
  XOR2HSV0 U15803 ( .A1(n14302), .A2(n14301), .Z(n14303) );
  XOR2HSV0 U15804 ( .A1(n14304), .A2(n14303), .Z(n14305) );
  XOR2HSV0 U15805 ( .A1(n14306), .A2(n14305), .Z(\pe15/poht [6]) );
  NAND2HSV2 U15806 ( .A1(n14853), .A2(\pe15/got [1]), .ZN(n14308) );
  NAND2HSV0 U15807 ( .A1(\pe15/aot [1]), .A2(\pe15/bq[1] ), .ZN(n14307) );
  XOR2HSV0 U15808 ( .A1(n14308), .A2(n14307), .Z(\pe15/poht [7]) );
  NOR2HSV2 U15809 ( .A1(n14310), .A2(n14309), .ZN(n14318) );
  NAND2HSV0 U15810 ( .A1(\pe17/aot [2]), .A2(\pe17/bq[2] ), .ZN(n14312) );
  NAND2HSV0 U15811 ( .A1(\pe17/aot [3]), .A2(\pe17/bq[1] ), .ZN(n14311) );
  XOR2HSV0 U15812 ( .A1(n14312), .A2(n14311), .Z(n14313) );
  CLKNAND2HSV1 U15813 ( .A1(\pe17/aot [1]), .A2(\pe17/bq[3] ), .ZN(n14334) );
  XNOR2HSV1 U15814 ( .A1(n14313), .A2(n14334), .ZN(n14316) );
  NAND2HSV2 U15815 ( .A1(n14824), .A2(\pe17/got [1]), .ZN(n14314) );
  XOR3HSV2 U15816 ( .A1(n14316), .A2(n14315), .A3(n14314), .Z(n14317) );
  XOR2HSV0 U15817 ( .A1(n14318), .A2(n14317), .Z(\pe17/poht [5]) );
  INHSV2 U15818 ( .I(\pe17/got [4]), .ZN(n14347) );
  NOR2HSV2 U15819 ( .A1(n14310), .A2(n14347), .ZN(n14332) );
  NAND2HSV0 U15820 ( .A1(\pe17/aot [2]), .A2(\pe17/bq[3] ), .ZN(n14321) );
  NAND2HSV0 U15821 ( .A1(\pe17/aot [1]), .A2(\pe17/bq[4] ), .ZN(n14320) );
  XOR2HSV0 U15822 ( .A1(n14321), .A2(n14320), .Z(n14325) );
  NAND2HSV0 U15823 ( .A1(\pe17/bq[2] ), .A2(\pe17/aot [3]), .ZN(n14323) );
  NAND2HSV0 U15824 ( .A1(\pe17/aot [4]), .A2(\pe17/bq[1] ), .ZN(n14322) );
  XOR2HSV0 U15825 ( .A1(n14323), .A2(n14322), .Z(n14324) );
  XOR2HSV0 U15826 ( .A1(n14325), .A2(n14324), .Z(n14326) );
  NAND2HSV2 U15827 ( .A1(n14824), .A2(\pe17/got [2]), .ZN(n14328) );
  XOR3HSV2 U15828 ( .A1(n14330), .A2(n14329), .A3(n14328), .Z(n14331) );
  XOR2HSV0 U15829 ( .A1(n14332), .A2(n14331), .Z(\pe17/poht [4]) );
  NAND2HSV0 U15830 ( .A1(\pe17/aot [4]), .A2(\pe17/bq[4] ), .ZN(n14338) );
  NAND2HSV0 U15831 ( .A1(\pe17/bq[1] ), .A2(\pe17/aot [7]), .ZN(n14337) );
  XOR2HSV0 U15832 ( .A1(n14338), .A2(n14337), .Z(n14342) );
  NAND2HSV0 U15833 ( .A1(n5973), .A2(\pe17/bq[2] ), .ZN(n14340) );
  NAND2HSV0 U15834 ( .A1(\pe17/bq[5] ), .A2(\pe17/aot [3]), .ZN(n14339) );
  XOR2HSV0 U15835 ( .A1(n14340), .A2(n14339), .Z(n14341) );
  XOR2HSV0 U15836 ( .A1(n14342), .A2(n14341), .Z(n14344) );
  NAND2HSV0 U15837 ( .A1(\pe17/got [2]), .A2(n14962), .ZN(n14346) );
  NOR2HSV2 U15838 ( .A1(n14350), .A2(n14349), .ZN(n14361) );
  NAND2HSV0 U15839 ( .A1(\pe16/ti_7[3] ), .A2(\pe16/got [1]), .ZN(n14359) );
  NAND2HSV0 U15840 ( .A1(\pe16/aot [2]), .A2(\pe16/bq[4] ), .ZN(n14355) );
  NAND2HSV0 U15841 ( .A1(\pe16/aot [5]), .A2(\pe16/bq[1] ), .ZN(n14354) );
  XOR2HSV0 U15842 ( .A1(n14355), .A2(n14354), .Z(n14356) );
  XOR2HSV0 U15843 ( .A1(n14357), .A2(n14356), .Z(n14358) );
  XOR2HSV0 U15844 ( .A1(n14359), .A2(n14358), .Z(n14360) );
  CLKNAND2HSV0 U15845 ( .A1(n14835), .A2(\pe16/got [3]), .ZN(n14362) );
  NAND2HSV0 U15846 ( .A1(n14365), .A2(\pe11/got [4]), .ZN(n14387) );
  NAND2HSV0 U15847 ( .A1(n14366), .A2(\pe11/got [3]), .ZN(n14385) );
  NAND2HSV0 U15848 ( .A1(\pe11/aot [5]), .A2(\pe11/bq[3] ), .ZN(n14368) );
  NAND2HSV0 U15849 ( .A1(\pe11/aot [3]), .A2(\pe11/bq[5] ), .ZN(n14367) );
  XOR2HSV0 U15850 ( .A1(n14368), .A2(n14367), .Z(n14372) );
  NAND2HSV0 U15851 ( .A1(\pe11/aot [4]), .A2(\pe11/bq[4] ), .ZN(n14369) );
  XOR2HSV0 U15852 ( .A1(n14370), .A2(n14369), .Z(n14371) );
  XOR2HSV0 U15853 ( .A1(n14372), .A2(n14371), .Z(n14378) );
  NAND2HSV0 U15854 ( .A1(\pe11/aot [6]), .A2(\pe11/bq[2] ), .ZN(n14374) );
  NAND2HSV0 U15855 ( .A1(n14837), .A2(\pe11/bq[1] ), .ZN(n14373) );
  XOR2HSV0 U15856 ( .A1(n14374), .A2(n14373), .Z(n14376) );
  XNOR2HSV1 U15857 ( .A1(n14376), .A2(n14375), .ZN(n14377) );
  XNOR2HSV1 U15858 ( .A1(n14378), .A2(n14377), .ZN(n14380) );
  NAND2HSV0 U15859 ( .A1(\pe11/ti_7[1] ), .A2(\pe11/got [1]), .ZN(n14379) );
  XOR2HSV0 U15860 ( .A1(n14380), .A2(n14379), .Z(n14383) );
  NAND2HSV0 U15861 ( .A1(\pe11/got [2]), .A2(n6713), .ZN(n14382) );
  XNOR2HSV1 U15862 ( .A1(n14383), .A2(n14382), .ZN(n14384) );
  XOR2HSV0 U15863 ( .A1(n14385), .A2(n14384), .Z(n14386) );
  XNOR2HSV1 U15864 ( .A1(n14387), .A2(n14386), .ZN(n14391) );
  NAND2HSV0 U15865 ( .A1(n14388), .A2(\pe11/got [6]), .ZN(n14389) );
  NAND2HSV2 U15866 ( .A1(n14965), .A2(\pe11/got [7]), .ZN(n14392) );
  XOR2HSV0 U15867 ( .A1(n14393), .A2(n14392), .Z(\pe11/poht [1]) );
  NAND2HSV0 U15868 ( .A1(\pe11/aot [2]), .A2(\pe11/bq[2] ), .ZN(n14395) );
  NAND2HSV0 U15869 ( .A1(\pe11/aot [1]), .A2(\pe11/bq[3] ), .ZN(n14394) );
  NOR2HSV2 U15870 ( .A1(n14310), .A2(n14397), .ZN(n14434) );
  CLKNAND2HSV0 U15871 ( .A1(\pe17/ti_7[3] ), .A2(\pe17/got [4]), .ZN(n14426)
         );
  NAND2HSV0 U15872 ( .A1(\pe17/aot [7]), .A2(\pe17/bq[2] ), .ZN(n14403) );
  NAND2HSV0 U15873 ( .A1(\pe17/aot [5]), .A2(\pe17/bq[4] ), .ZN(n14402) );
  XOR2HSV0 U15874 ( .A1(n14403), .A2(n14402), .Z(n14422) );
  CLKNAND2HSV0 U15875 ( .A1(n14571), .A2(\pe17/pq ), .ZN(n14406) );
  NAND2HSV0 U15876 ( .A1(\pe17/aot [4]), .A2(\pe17/bq[5] ), .ZN(n14405) );
  XOR2HSV0 U15877 ( .A1(n14406), .A2(n14405), .Z(n14411) );
  AOI22HSV0 U15878 ( .A1(n14949), .A2(\pe17/bq[1] ), .B1(n5973), .B2(
        \pe17/bq[3] ), .ZN(n14407) );
  AOI21HSV0 U15879 ( .A1(n14409), .A2(n14408), .B(n14407), .ZN(n14410) );
  XNOR2HSV1 U15880 ( .A1(n14411), .A2(n14410), .ZN(n14421) );
  NAND2HSV0 U15881 ( .A1(\pe17/aot [2]), .A2(n14412), .ZN(n14414) );
  XOR2HSV0 U15882 ( .A1(n14414), .A2(n14413), .Z(n14419) );
  NAND2HSV0 U15883 ( .A1(\pe17/aot [3]), .A2(\pe17/bq[6] ), .ZN(n14417) );
  NAND2HSV0 U15884 ( .A1(\pe17/got [1]), .A2(n14415), .ZN(n14416) );
  XOR2HSV0 U15885 ( .A1(n14417), .A2(n14416), .Z(n14418) );
  XOR2HSV0 U15886 ( .A1(n14419), .A2(n14418), .Z(n14420) );
  XOR3HSV2 U15887 ( .A1(n14422), .A2(n14421), .A3(n14420), .Z(n14423) );
  XNOR2HSV1 U15888 ( .A1(n14424), .A2(n14423), .ZN(n14425) );
  XNOR2HSV1 U15889 ( .A1(n14426), .A2(n14425), .ZN(n14427) );
  XOR2HSV0 U15890 ( .A1(n14428), .A2(n14427), .Z(n14432) );
  NAND2HSV0 U15891 ( .A1(n14824), .A2(\pe17/got [6]), .ZN(n14430) );
  XOR3HSV2 U15892 ( .A1(n14432), .A2(n14431), .A3(n14430), .Z(n14433) );
  XOR2HSV0 U15893 ( .A1(n14434), .A2(n14433), .Z(po17) );
  NAND2HSV0 U15894 ( .A1(\pe14/aot [1]), .A2(\pe14/bq[1] ), .ZN(n14435) );
  XOR2HSV0 U15895 ( .A1(n14436), .A2(n14435), .Z(\pe14/poht [7]) );
  NAND2HSV0 U15896 ( .A1(\pe12/aot [3]), .A2(\pe12/bq[1] ), .ZN(n14438) );
  NAND2HSV0 U15897 ( .A1(\pe12/aot [1]), .A2(\pe12/bq[3] ), .ZN(n14437) );
  XOR2HSV0 U15898 ( .A1(n14438), .A2(n14437), .Z(n14440) );
  XNOR2HSV1 U15899 ( .A1(n14440), .A2(n14439), .ZN(n14445) );
  CLKNHSV1 U15900 ( .I(\pe12/got [1]), .ZN(n14441) );
  NOR2HSV4 U15901 ( .A1(n14442), .A2(n14441), .ZN(n14444) );
  XOR3HSV2 U15902 ( .A1(n14445), .A2(n14444), .A3(n14443), .Z(n14448) );
  CLKNAND2HSV1 U15903 ( .A1(n14446), .A2(\pe12/got [3]), .ZN(n14447) );
  XOR2HSV0 U15904 ( .A1(n14448), .A2(n14447), .Z(\pe12/poht [5]) );
  NAND2HSV2 U15905 ( .A1(n14449), .A2(n6038), .ZN(n14463) );
  CLKNAND2HSV1 U15906 ( .A1(n15081), .A2(\pe7/got [1]), .ZN(n14458) );
  NAND2HSV0 U15907 ( .A1(\pe7/aot [2]), .A2(\pe7/bq[3] ), .ZN(n14452) );
  NAND2HSV0 U15908 ( .A1(\pe7/aot [1]), .A2(\pe7/bq[4] ), .ZN(n14451) );
  XOR2HSV0 U15909 ( .A1(n14452), .A2(n14451), .Z(n14456) );
  NAND2HSV0 U15910 ( .A1(\pe7/bq[2] ), .A2(\pe7/aot [3]), .ZN(n14454) );
  NAND2HSV0 U15911 ( .A1(\pe7/aot [4]), .A2(\pe7/bq[1] ), .ZN(n14453) );
  XOR2HSV0 U15912 ( .A1(n14454), .A2(n14453), .Z(n14455) );
  XOR2HSV0 U15913 ( .A1(n14456), .A2(n14455), .Z(n14457) );
  XOR2HSV0 U15914 ( .A1(n14458), .A2(n14457), .Z(n14461) );
  NAND2HSV2 U15915 ( .A1(\pe7/ti_7[5] ), .A2(\pe7/got [2]), .ZN(n14460) );
  NAND2HSV2 U15916 ( .A1(n14487), .A2(\pe7/got [3]), .ZN(n14459) );
  XOR3HSV2 U15917 ( .A1(n14461), .A2(n14460), .A3(n14459), .Z(n14462) );
  XOR2HSV0 U15918 ( .A1(n14463), .A2(n14462), .Z(\pe7/poht [4]) );
  NAND2HSV0 U15919 ( .A1(n14860), .A2(\pe7/got [3]), .ZN(n14467) );
  NAND2HSV0 U15920 ( .A1(\pe7/ti_7[1] ), .A2(\pe7/got [2]), .ZN(n14466) );
  CLKNAND2HSV0 U15921 ( .A1(n12067), .A2(\pe7/pq ), .ZN(n14469) );
  NAND2HSV0 U15922 ( .A1(\pe7/aot [6]), .A2(\pe7/bq[3] ), .ZN(n14468) );
  XOR2HSV0 U15923 ( .A1(n14469), .A2(n14468), .Z(n14473) );
  NAND2HSV0 U15924 ( .A1(\pe7/aot [5]), .A2(\pe7/bq[4] ), .ZN(n14471) );
  NAND2HSV0 U15925 ( .A1(\pe7/aot [7]), .A2(\pe7/bq[2] ), .ZN(n14470) );
  XOR2HSV0 U15926 ( .A1(n14471), .A2(n14470), .Z(n14472) );
  XOR2HSV0 U15927 ( .A1(n14473), .A2(n14472), .Z(n14477) );
  NAND2HSV0 U15928 ( .A1(\pe7/aot [4]), .A2(\pe7/bq[5] ), .ZN(n14475) );
  NAND2HSV0 U15929 ( .A1(\pe7/aot [3]), .A2(\pe7/bq[6] ), .ZN(n14474) );
  XOR2HSV0 U15930 ( .A1(n14475), .A2(n14474), .Z(n14476) );
  XNOR2HSV1 U15931 ( .A1(n14477), .A2(n14476), .ZN(n14486) );
  NAND2HSV0 U15932 ( .A1(\pe7/aot [1]), .A2(\pe7/bq[8] ), .ZN(n14479) );
  NAND2HSV0 U15933 ( .A1(\pe7/bq[1] ), .A2(\pe7/aot [8]), .ZN(n14478) );
  XOR2HSV0 U15934 ( .A1(n14479), .A2(n14478), .Z(n14484) );
  NAND2HSV0 U15935 ( .A1(\pe7/got [1]), .A2(n14480), .ZN(n14482) );
  NAND2HSV0 U15936 ( .A1(\pe7/aot [2]), .A2(\pe7/bq[7] ), .ZN(n14481) );
  XOR2HSV0 U15937 ( .A1(n14482), .A2(n14481), .Z(n14483) );
  XOR2HSV0 U15938 ( .A1(n14484), .A2(n14483), .Z(n14485) );
  NAND2HSV0 U15939 ( .A1(\pe14/aot [5]), .A2(\pe14/bq[1] ), .ZN(n14491) );
  NAND2HSV0 U15940 ( .A1(\pe14/aot [1]), .A2(\pe14/bq[5] ), .ZN(n14490) );
  XOR2HSV0 U15941 ( .A1(n14491), .A2(n14490), .Z(n14493) );
  XNOR2HSV1 U15942 ( .A1(n14493), .A2(n14492), .ZN(n14496) );
  NAND2HSV0 U15943 ( .A1(\pe14/aot [3]), .A2(\pe14/bq[3] ), .ZN(n14495) );
  NAND2HSV0 U15944 ( .A1(\pe14/aot [4]), .A2(\pe14/bq[2] ), .ZN(n14494) );
  MUX2HSV2 U15945 ( .I0(bo2[3]), .I1(\pe2/bq[3] ), .S(n14805), .Z(n14966) );
  BUFHSV2 U15946 ( .I(\pe1/bq[2] ), .Z(n14497) );
  MUX2HSV2 U15947 ( .I0(bo1[2]), .I1(n14497), .S(\pe1/ctrq ), .Z(n14967) );
  MUX2HSV2 U15948 ( .I0(bo19[1]), .I1(\pe19/bq[1] ), .S(n14501), .Z(n14968) );
  CLKBUFHSV1 U15949 ( .I(\pe18/bq[3] ), .Z(n14498) );
  MUX2HSV2 U15950 ( .I0(bo18[3]), .I1(n14498), .S(n14790), .Z(n14969) );
  CLKBUFHSV1 U15951 ( .I(\pe2/bq[4] ), .Z(n14499) );
  MUX2HSV2 U15952 ( .I0(bo2[4]), .I1(n14499), .S(n14558), .Z(n14970) );
  MUX2HSV2 U15953 ( .I0(bo1[4]), .I1(\pe1/bq[4] ), .S(\pe1/ctrq ), .Z(n14971)
         );
  MUX2HSV2 U15954 ( .I0(bo19[2]), .I1(\pe19/bq[2] ), .S(n14501), .Z(n14972) );
  MUX2HSV2 U15955 ( .I0(bo18[1]), .I1(\pe18/bq[1] ), .S(n14790), .Z(n14973) );
  MUX2HSV2 U15956 ( .I0(bo1[8]), .I1(n14502), .S(\pe1/ctrq ), .Z(n14974) );
  MUX2HSV2 U15957 ( .I0(bo2[7]), .I1(n14504), .S(n14523), .Z(n14976) );
  MUX2HSV2 U15958 ( .I0(bo14[8]), .I1(n14505), .S(n14516), .Z(n14977) );
  MUX2HSV2 U15959 ( .I0(bo19[8]), .I1(n14506), .S(n14501), .Z(n14978) );
  BUFHSV2 U15960 ( .I(n14578), .Z(n14521) );
  MUX2HSV2 U15961 ( .I0(bo12[8]), .I1(n14507), .S(n14521), .Z(n14979) );
  MUX2HSV2 U15962 ( .I0(bo13[2]), .I1(\pe13/bq[2] ), .S(n14552), .Z(n14981) );
  CLKNHSV0 U15963 ( .I(\pe12/bq[1] ), .ZN(n14508) );
  INHSV2 U15964 ( .I(n14508), .ZN(n14509) );
  BUFHSV2 U15965 ( .I(n14578), .Z(n14531) );
  MUX2HSV2 U15966 ( .I0(bo12[1]), .I1(n14509), .S(n14531), .Z(n14982) );
  MUX2HSV2 U15967 ( .I0(bo2[1]), .I1(\pe2/bq[1] ), .S(n8946), .Z(n14983) );
  MUX2HSV2 U15968 ( .I0(bo2[6]), .I1(n14510), .S(n14558), .Z(n14984) );
  MUX2HSV2 U15969 ( .I0(bo12[4]), .I1(\pe12/bq[4] ), .S(n14578), .Z(n14985) );
  MUX2HSV2 U15970 ( .I0(bo8[5]), .I1(\pe8/bq[5] ), .S(n14572), .Z(n14986) );
  MUX2HSV2 U15971 ( .I0(bo17[3]), .I1(\pe17/bq[3] ), .S(n14571), .Z(n14987) );
  MUX2HSV2 U15972 ( .I0(bo18[8]), .I1(n14511), .S(n14790), .Z(n14988) );
  MUX2HSV2 U15973 ( .I0(bo18[7]), .I1(n14513), .S(n14790), .Z(n14990) );
  CLKNHSV0 U15974 ( .I(\pe16/bq[5] ), .ZN(n14514) );
  INHSV2 U15975 ( .I(n14514), .ZN(n14515) );
  MUX2HSV2 U15976 ( .I0(bo16[5]), .I1(n14515), .S(n14743), .Z(n14991) );
  CLKNHSV0 U15977 ( .I(n14516), .ZN(n14517) );
  INHSV2 U15978 ( .I(n14517), .ZN(n14551) );
  MUX2HSV2 U15979 ( .I0(bo14[6]), .I1(n14518), .S(n14551), .Z(n14993) );
  MUX2HSV2 U15980 ( .I0(bo12[2]), .I1(\pe12/bq[2] ), .S(n14578), .Z(n14994) );
  MUX2HSV2 U15981 ( .I0(bo11[7]), .I1(n14519), .S(n14553), .Z(n14995) );
  MUX2HSV2 U15982 ( .I0(bo8[4]), .I1(\pe8/bq[4] ), .S(n14572), .Z(n14996) );
  BUFHSV2 U15983 ( .I(\pe1/bq[5] ), .Z(n14520) );
  MUX2HSV2 U15984 ( .I0(bo1[5]), .I1(n14520), .S(\pe1/ctrq ), .Z(n14997) );
  BUFHSV2 U15985 ( .I(\pe12/bq[3] ), .Z(n14522) );
  MUX2HSV2 U15986 ( .I0(bo12[3]), .I1(n14522), .S(n14521), .Z(n14998) );
  MUX2HSV2 U15987 ( .I0(bo2[2]), .I1(\pe2/bq[2] ), .S(n14523), .Z(n14999) );
  CLKNHSV0 U15988 ( .I(\pe17/bq[6] ), .ZN(n14524) );
  INHSV2 U15989 ( .I(n14524), .ZN(n14525) );
  MUX2HSV2 U15990 ( .I0(bo17[6]), .I1(n14525), .S(n14571), .Z(n15000) );
  CLKNHSV0 U15991 ( .I(\pe16/bq[6] ), .ZN(n14526) );
  INHSV2 U15992 ( .I(n14526), .ZN(n14527) );
  CLKNHSV0 U15993 ( .I(\pe12/bq[6] ), .ZN(n14528) );
  INHSV2 U15994 ( .I(n14528), .ZN(n14529) );
  MUX2HSV2 U15995 ( .I0(bo12[6]), .I1(n14529), .S(n14938), .Z(n15002) );
  CLKNHSV0 U15996 ( .I(\pe12/bq[5] ), .ZN(n14530) );
  INHSV2 U15997 ( .I(n14530), .ZN(n14532) );
  MUX2HSV2 U15998 ( .I0(bo12[5]), .I1(n14532), .S(n14531), .Z(n15003) );
  CLKNHSV0 U15999 ( .I(\pe2/bq[5] ), .ZN(n14533) );
  INHSV2 U16000 ( .I(n14533), .ZN(n14534) );
  MUX2HSV2 U16001 ( .I0(bo2[5]), .I1(n14534), .S(n8946), .Z(n15004) );
  MUX2HSV2 U16002 ( .I0(bo17[1]), .I1(\pe17/bq[1] ), .S(n14892), .Z(n15005) );
  MUX2HSV2 U16003 ( .I0(bo14[7]), .I1(\pe14/bq[7] ), .S(n14535), .Z(n15006) );
  CLKNHSV0 U16004 ( .I(\pe21/bq[6] ), .ZN(n14536) );
  INHSV2 U16005 ( .I(n14536), .ZN(n14538) );
  MUX2HSV2 U16006 ( .I0(bo21[6]), .I1(n14538), .S(n6014), .Z(n15007) );
  MUX2HSV2 U16007 ( .I0(bo1[3]), .I1(\pe1/bq[3] ), .S(\pe1/ctrq ), .Z(n15008)
         );
  MUX2HSV2 U16008 ( .I0(bo21[1]), .I1(\pe21/bq[1] ), .S(n14574), .Z(n15009) );
  CLKNHSV0 U16009 ( .I(\pe19/bq[6] ), .ZN(n14541) );
  INHSV2 U16010 ( .I(n14541), .ZN(n14542) );
  MUX2HSV2 U16011 ( .I0(bo19[6]), .I1(n14542), .S(n14501), .Z(n15014) );
  CLKBUFHSV1 U16012 ( .I(\pe19/bq[4] ), .Z(n14544) );
  MUX2HSV2 U16013 ( .I0(bo19[4]), .I1(n14544), .S(n14501), .Z(n15015) );
  CLKBUFHSV1 U16014 ( .I(\pe19/bq[3] ), .Z(n14545) );
  MUX2HSV2 U16015 ( .I0(bo19[3]), .I1(n14545), .S(n14501), .Z(n15016) );
  CLKNHSV0 U16016 ( .I(\pe18/bq[4] ), .ZN(n14547) );
  INHSV2 U16017 ( .I(n14547), .ZN(n14548) );
  MUX2HSV2 U16018 ( .I0(bo18[4]), .I1(n14548), .S(n14564), .Z(n15018) );
  MUX2HSV2 U16019 ( .I0(bo18[2]), .I1(\pe18/bq[2] ), .S(n14564), .Z(n15019) );
  CLKNHSV0 U16020 ( .I(\pe17/bq[4] ), .ZN(n14549) );
  INHSV2 U16021 ( .I(n14549), .ZN(n14550) );
  MUX2HSV2 U16022 ( .I0(bo17[4]), .I1(n14550), .S(n14892), .Z(n15020) );
  MUX2HSV2 U16023 ( .I0(bo16[1]), .I1(\pe16/bq[1] ), .S(n14743), .Z(n15021) );
  MUX2HSV2 U16024 ( .I0(bo14[5]), .I1(\pe14/bq[5] ), .S(n14742), .Z(n15024) );
  MUX2HSV2 U16025 ( .I0(bo14[2]), .I1(\pe14/bq[2] ), .S(n14551), .Z(n15025) );
  MUX2HSV2 U16026 ( .I0(bo13[1]), .I1(\pe13/bq[1] ), .S(n14552), .Z(n15026) );
  MUX2HSV2 U16027 ( .I0(bo11[4]), .I1(\pe11/bq[4] ), .S(n14553), .Z(n15027) );
  MUX2HSV2 U16028 ( .I0(bo10[6]), .I1(\pe10/bq[6] ), .S(n14554), .Z(n15029) );
  BUFHSV2 U16029 ( .I(\pe10/bq[2] ), .Z(n14555) );
  MUX2HSV2 U16030 ( .I0(bo10[2]), .I1(n14555), .S(n14554), .Z(n15032) );
  MUX2HSV2 U16031 ( .I0(bo9[2]), .I1(\pe9/bq[2] ), .S(n13826), .Z(n15034) );
  MUX2HSV2 U16032 ( .I0(bo8[2]), .I1(\pe8/bq[2] ), .S(n14758), .Z(n15035) );
  MUX2HSV2 U16033 ( .I0(bo7[2]), .I1(\pe7/bq[2] ), .S(n12067), .Z(n15036) );
  CLKNHSV0 U16034 ( .I(\pe1/bq[1] ), .ZN(n14556) );
  INHSV2 U16035 ( .I(n14556), .ZN(n14557) );
  MUX2HSV2 U16036 ( .I0(bo1[1]), .I1(n14557), .S(\pe1/ctrq ), .Z(n15046) );
  MUX2HSV2 U16037 ( .I0(bo2[8]), .I1(n14559), .S(n14558), .Z(n15047) );
  CLKNHSV0 U16038 ( .I(\pe21/bq[7] ), .ZN(n14561) );
  INHSV2 U16039 ( .I(n14561), .ZN(n14562) );
  MUX2HSV2 U16040 ( .I0(bo21[7]), .I1(n14562), .S(n14574), .Z(n15049) );
  MUX2HSV2 U16041 ( .I0(bo14[3]), .I1(\pe14/bq[3] ), .S(n14566), .Z(n15052) );
  MUX2HSV2 U16042 ( .I0(bo10[7]), .I1(n14567), .S(n14554), .Z(n15053) );
  CLKNHSV0 U16043 ( .I(\pe19/bq[5] ), .ZN(n14568) );
  INHSV2 U16044 ( .I(n14568), .ZN(n14569) );
  MUX2HSV2 U16045 ( .I0(bo19[5]), .I1(n14569), .S(n14501), .Z(n15055) );
  MUX2HSV2 U16046 ( .I0(bo16[8]), .I1(n5947), .S(n14570), .Z(n15056) );
  MUX2HSV2 U16047 ( .I0(bo8[3]), .I1(\pe8/bq[3] ), .S(n14572), .Z(n15058) );
  MUX2HSV2 U16048 ( .I0(bo9[4]), .I1(\pe9/bq[4] ), .S(n13826), .Z(n15059) );
  CLKNHSV0 U16049 ( .I(\pe21/bq[2] ), .ZN(n14573) );
  INHSV2 U16050 ( .I(n14573), .ZN(n14575) );
  MUX2HSV2 U16051 ( .I0(bo21[2]), .I1(n14575), .S(n14574), .Z(n15060) );
  MUX2HSV2 U16052 ( .I0(bo19[7]), .I1(n14576), .S(n14501), .Z(n15061) );
  CLKNHSV0 U16053 ( .I(\pe21/bq[4] ), .ZN(n14579) );
  INHSV2 U16054 ( .I(n14579), .ZN(n14580) );
  MUX2HSV2 U16055 ( .I0(bo21[4]), .I1(n14580), .S(n14574), .Z(n15063) );
  MUX2HSV2 U16056 ( .I0(bo1[6]), .I1(n14581), .S(\pe1/ctrq ), .Z(n15064) );
  XNOR2HSV1 U16057 ( .A1(n14583), .A2(n6810), .ZN(pov9[7]) );
  CLKNAND2HSV1 U16058 ( .A1(n6535), .A2(n14864), .ZN(n14620) );
  NOR2HSV2 U16059 ( .A1(n12514), .A2(n14584), .ZN(n14617) );
  NAND2HSV0 U16060 ( .A1(n15072), .A2(\pe15/got [2]), .ZN(n14611) );
  CLKNAND2HSV1 U16061 ( .A1(n5946), .A2(\pe15/got [3]), .ZN(n14610) );
  CLKNAND2HSV0 U16062 ( .A1(n14586), .A2(\pe15/pq ), .ZN(n14589) );
  NAND2HSV0 U16063 ( .A1(\pe15/got [1]), .A2(n14587), .ZN(n14588) );
  XOR2HSV0 U16064 ( .A1(n14589), .A2(n14588), .Z(n14593) );
  NAND2HSV0 U16065 ( .A1(n14936), .A2(\pe15/bq[2] ), .ZN(n14591) );
  NAND2HSV0 U16066 ( .A1(n14937), .A2(\pe15/bq[1] ), .ZN(n14590) );
  XOR2HSV0 U16067 ( .A1(n14591), .A2(n14590), .Z(n14592) );
  XOR2HSV0 U16068 ( .A1(n14593), .A2(n14592), .Z(n14597) );
  NAND2HSV0 U16069 ( .A1(\pe15/aot [3]), .A2(\pe15/bq[6] ), .ZN(n14595) );
  NAND2HSV0 U16070 ( .A1(\pe15/aot [4]), .A2(\pe15/bq[5] ), .ZN(n14594) );
  XOR2HSV0 U16071 ( .A1(n14595), .A2(n14594), .Z(n14596) );
  XNOR2HSV1 U16072 ( .A1(n14597), .A2(n14596), .ZN(n14608) );
  NAND2HSV0 U16073 ( .A1(\pe15/aot [5]), .A2(\pe15/bq[4] ), .ZN(n14599) );
  NAND2HSV0 U16074 ( .A1(\pe15/aot [2]), .A2(\pe15/bq[7] ), .ZN(n14598) );
  XOR2HSV0 U16075 ( .A1(n14599), .A2(n14598), .Z(n14606) );
  CLKNHSV0 U16076 ( .I(\pe15/bq[3] ), .ZN(n14600) );
  CLKNHSV0 U16077 ( .I(n14600), .ZN(n14601) );
  NAND2HSV0 U16078 ( .A1(n14739), .A2(n14601), .ZN(n14604) );
  NAND2HSV0 U16079 ( .A1(\pe15/aot [1]), .A2(n14602), .ZN(n14603) );
  XOR2HSV0 U16080 ( .A1(n14604), .A2(n14603), .Z(n14605) );
  XOR2HSV0 U16081 ( .A1(n14606), .A2(n14605), .Z(n14607) );
  XNOR2HSV1 U16082 ( .A1(n14608), .A2(n14607), .ZN(n14609) );
  XOR3HSV2 U16083 ( .A1(n14611), .A2(n14610), .A3(n14609), .Z(n14612) );
  NAND2HSV0 U16084 ( .A1(\pe15/ti_7[3] ), .A2(\pe15/got [4]), .ZN(n14614) );
  CLKXOR2HSV2 U16085 ( .A1(n14617), .A2(n14616), .Z(n14619) );
  CLKNAND2HSV2 U16086 ( .A1(n14853), .A2(n15178), .ZN(n14618) );
  XOR3HSV2 U16087 ( .A1(n14620), .A2(n14619), .A3(n14618), .Z(po15) );
  NOR2HSV2 U16088 ( .A1(n14650), .A2(n14621), .ZN(n14645) );
  NAND2HSV0 U16089 ( .A1(n14851), .A2(\pe18/got [4]), .ZN(n14643) );
  NAND2HSV0 U16090 ( .A1(\pe18/aot [2]), .A2(\pe18/bq[6] ), .ZN(n14623) );
  NAND2HSV0 U16091 ( .A1(\pe18/aot [5]), .A2(\pe18/bq[3] ), .ZN(n14622) );
  XOR2HSV0 U16092 ( .A1(n14623), .A2(n14622), .Z(n14629) );
  NOR2HSV0 U16093 ( .A1(n14625), .A2(n14624), .ZN(n14627) );
  NAND2HSV0 U16094 ( .A1(\pe18/aot [3]), .A2(\pe18/bq[5] ), .ZN(n14626) );
  XOR2HSV0 U16095 ( .A1(n14627), .A2(n14626), .Z(n14628) );
  XOR2HSV0 U16096 ( .A1(n14629), .A2(n14628), .Z(n14635) );
  CLKNAND2HSV0 U16097 ( .A1(n14894), .A2(\pe18/bq[2] ), .ZN(n14631) );
  NAND2HSV0 U16098 ( .A1(\pe18/aot [4]), .A2(\pe18/bq[4] ), .ZN(n14630) );
  XOR2HSV0 U16099 ( .A1(n14631), .A2(n14630), .Z(n14633) );
  XOR2HSV0 U16100 ( .A1(n14633), .A2(n14632), .Z(n14634) );
  XOR2HSV0 U16101 ( .A1(n14635), .A2(n14634), .Z(n14637) );
  NAND2HSV0 U16102 ( .A1(\pe18/ti_7[1] ), .A2(\pe18/got [1]), .ZN(n14636) );
  XNOR2HSV1 U16103 ( .A1(n14637), .A2(n14636), .ZN(n14639) );
  XNOR2HSV1 U16104 ( .A1(n14639), .A2(n14638), .ZN(n14640) );
  XNOR2HSV1 U16105 ( .A1(n14641), .A2(n14640), .ZN(n14642) );
  XNOR2HSV1 U16106 ( .A1(n14643), .A2(n14642), .ZN(n14644) );
  XOR2HSV0 U16107 ( .A1(n14645), .A2(n14644), .Z(n14647) );
  NAND2HSV2 U16108 ( .A1(n14695), .A2(\pe18/got [7]), .ZN(n14646) );
  XOR3HSV2 U16109 ( .A1(n14648), .A2(n14647), .A3(n14646), .Z(\pe18/poht [1])
         );
  CLKNAND2HSV1 U16110 ( .A1(n14669), .A2(\pe18/got [4]), .ZN(n14668) );
  CLKNHSV0 U16111 ( .I(\pe18/got [3]), .ZN(n14649) );
  NOR2HSV2 U16112 ( .A1(n14650), .A2(n14649), .ZN(n14665) );
  NAND2HSV0 U16113 ( .A1(\pe18/aot [2]), .A2(\pe18/bq[4] ), .ZN(n14657) );
  NAND2HSV0 U16114 ( .A1(\pe18/bq[2] ), .A2(\pe18/aot [4]), .ZN(n14652) );
  NAND2HSV0 U16115 ( .A1(\pe18/aot [1]), .A2(\pe18/bq[5] ), .ZN(n14651) );
  XNOR2HSV1 U16116 ( .A1(n14652), .A2(n14651), .ZN(n14656) );
  NAND2HSV0 U16117 ( .A1(\pe18/aot [5]), .A2(\pe18/bq[1] ), .ZN(n14654) );
  NAND2HSV0 U16118 ( .A1(\pe18/aot [3]), .A2(\pe18/bq[3] ), .ZN(n14653) );
  XOR2HSV0 U16119 ( .A1(n14654), .A2(n14653), .Z(n14655) );
  XOR3HSV2 U16120 ( .A1(n14657), .A2(n14656), .A3(n14655), .Z(n14658) );
  XNOR2HSV1 U16121 ( .A1(n14659), .A2(n14658), .ZN(n14661) );
  CLKNHSV0 U16122 ( .I(n14661), .ZN(n14660) );
  INHSV1 U16123 ( .I(\pe18/got [2]), .ZN(n14670) );
  NOR2HSV1 U16124 ( .A1(n14660), .A2(n14670), .ZN(n14663) );
  AOI21HSV0 U16125 ( .A1(n14851), .A2(\pe18/got [2]), .B(n14661), .ZN(n14662)
         );
  AOI21HSV1 U16126 ( .A1(n14663), .A2(n14851), .B(n14662), .ZN(n14664) );
  XOR2HSV0 U16127 ( .A1(n14665), .A2(n14664), .Z(n14667) );
  NAND2HSV2 U16128 ( .A1(n14695), .A2(\pe18/got [5]), .ZN(n14666) );
  XOR3HSV2 U16129 ( .A1(n14668), .A2(n14667), .A3(n14666), .Z(\pe18/poht [3])
         );
  CLKNAND2HSV1 U16130 ( .A1(n14669), .A2(\pe18/got [3]), .ZN(n14686) );
  NOR2HSV2 U16131 ( .A1(n14688), .A2(n14670), .ZN(n14680) );
  NAND2HSV0 U16132 ( .A1(n14851), .A2(\pe18/got [1]), .ZN(n14678) );
  NAND2HSV0 U16133 ( .A1(\pe18/aot [3]), .A2(\pe18/bq[2] ), .ZN(n14672) );
  NAND2HSV0 U16134 ( .A1(\pe18/aot [1]), .A2(\pe18/bq[4] ), .ZN(n14671) );
  XOR2HSV0 U16135 ( .A1(n14672), .A2(n14671), .Z(n14676) );
  NAND2HSV0 U16136 ( .A1(\pe18/aot [4]), .A2(\pe18/bq[1] ), .ZN(n14674) );
  NAND2HSV0 U16137 ( .A1(\pe18/aot [2]), .A2(\pe18/bq[3] ), .ZN(n14673) );
  XOR2HSV0 U16138 ( .A1(n14674), .A2(n14673), .Z(n14675) );
  XOR2HSV0 U16139 ( .A1(n14676), .A2(n14675), .Z(n14677) );
  XNOR2HSV1 U16140 ( .A1(n14678), .A2(n14677), .ZN(n14679) );
  XOR2HSV0 U16141 ( .A1(n14680), .A2(n14679), .Z(n14685) );
  CLKNAND2HSV2 U16142 ( .A1(n14681), .A2(n14682), .ZN(n14683) );
  XOR3HSV2 U16143 ( .A1(n14686), .A2(n14685), .A3(n14684), .Z(\pe18/poht [4])
         );
  CLKNHSV0 U16144 ( .I(\pe18/got [1]), .ZN(n14687) );
  NOR2HSV2 U16145 ( .A1(n14688), .A2(n14687), .ZN(n14694) );
  NAND2HSV0 U16146 ( .A1(\pe18/aot [3]), .A2(\pe18/bq[1] ), .ZN(n14690) );
  NAND2HSV0 U16147 ( .A1(\pe18/aot [2]), .A2(\pe18/bq[2] ), .ZN(n14689) );
  XOR2HSV0 U16148 ( .A1(n14690), .A2(n14689), .Z(n14692) );
  NAND2HSV0 U16149 ( .A1(\pe18/aot [1]), .A2(\pe18/bq[3] ), .ZN(n14691) );
  XNOR2HSV1 U16150 ( .A1(n14692), .A2(n14691), .ZN(n14693) );
  XOR2HSV0 U16151 ( .A1(n14694), .A2(n14693), .Z(n14697) );
  NAND2HSV2 U16152 ( .A1(n14695), .A2(\pe18/got [3]), .ZN(n14696) );
  XOR3HSV2 U16153 ( .A1(n14698), .A2(n14697), .A3(n14696), .Z(\pe18/poht [5])
         );
endmodule

