
module topcell ( clk, ctr, rst, ai, gi, bi, po );
  input [16:1] ai;
  input [16:1] gi;
  input [16:1] bi;
  output [1:16] po;
  input clk, ctr, rst;
  wire   po1, ctro1, \pov2[10] , po2, ctro2, po3, ctro3, po4, ctro4, po5,
         ctro5, po6, ctro6, \pov7[10] , po7, ctro7, po8, ctro8, po9, ctro9,
         po10, ctro10, po11, ctro11, \pe1/bq[1] , \pe1/bq[2] , \pe1/bq[3] ,
         \pe1/bq[4] , \pe1/bq[5] , \pe1/bq[6] , \pe1/bq[7] , \pe1/bq[8] ,
         \pe1/bq[9] , \pe1/bq[10] , \pe1/bq[11] , \pe1/bq[12] , \pe1/bq[13] ,
         \pe1/bq[14] , \pe1/bq[15] , \pe1/bq[16] , \pe1/ctrq , \pe2/ti_1 ,
         \pe2/ti_1t , \pe2/bq[1] , \pe2/bq[2] , \pe2/bq[3] , \pe2/bq[4] ,
         \pe2/bq[5] , \pe2/bq[6] , \pe2/bq[7] , \pe2/bq[8] , \pe2/bq[9] ,
         \pe2/bq[10] , \pe2/bq[11] , \pe2/bq[12] , \pe2/bq[13] , \pe2/bq[14] ,
         \pe2/bq[15] , \pe2/bq[16] , \pe2/ctrq , \pe2/pq , \pe3/ti_1 ,
         \pe3/ti_1t , \pe3/bq[1] , \pe3/bq[2] , \pe3/bq[3] , \pe3/bq[4] ,
         \pe3/bq[5] , \pe3/bq[6] , \pe3/bq[7] , \pe3/bq[8] , \pe3/bq[9] ,
         \pe3/bq[10] , \pe3/bq[11] , \pe3/bq[12] , \pe3/bq[13] , \pe3/bq[14] ,
         \pe3/bq[15] , \pe3/bq[16] , \pe3/ctrq , \pe3/pq , \pe4/ti_7[7] ,
         \pe4/ti_1 , \pe4/ti_1t , \pe4/bq[1] , \pe4/bq[2] , \pe4/bq[3] ,
         \pe4/bq[4] , \pe4/bq[5] , \pe4/bq[6] , \pe4/bq[7] , \pe4/bq[8] ,
         \pe4/bq[9] , \pe4/bq[10] , \pe4/bq[11] , \pe4/bq[12] , \pe4/bq[13] ,
         \pe4/bq[14] , \pe4/bq[15] , \pe4/bq[16] , \pe4/ctrq , \pe4/pq ,
         \pe5/ti_7[10] , \pe5/ti_1 , \pe5/ti_1t , \pe5/bq[1] , \pe5/bq[2] ,
         \pe5/bq[3] , \pe5/bq[4] , \pe5/bq[5] , \pe5/bq[6] , \pe5/bq[7] ,
         \pe5/bq[8] , \pe5/bq[9] , \pe5/bq[10] , \pe5/bq[11] , \pe5/bq[12] ,
         \pe5/bq[13] , \pe5/bq[14] , \pe5/bq[15] , \pe5/bq[16] , \pe5/ctrq ,
         \pe5/pq , \pe6/ti_7[7] , \pe6/ti_7[1] , \pe6/ti_1 , \pe6/ti_1t ,
         \pe6/bq[1] , \pe6/bq[2] , \pe6/bq[3] , \pe6/bq[4] , \pe6/bq[5] ,
         \pe6/bq[6] , \pe6/bq[7] , \pe6/bq[8] , \pe6/bq[9] , \pe6/bq[10] ,
         \pe6/bq[11] , \pe6/bq[12] , \pe6/bq[13] , \pe6/bq[14] , \pe6/bq[15] ,
         \pe6/bq[16] , \pe6/ctrq , \pe6/pq , \pe7/ti_7[1] , \pe7/ti_1 ,
         \pe7/ti_1t , \pe7/bq[1] , \pe7/bq[2] , \pe7/bq[3] , \pe7/bq[4] ,
         \pe7/bq[5] , \pe7/bq[6] , \pe7/bq[7] , \pe7/bq[8] , \pe7/bq[9] ,
         \pe7/bq[10] , \pe7/bq[11] , \pe7/bq[12] , \pe7/bq[13] , \pe7/bq[14] ,
         \pe7/bq[15] , \pe7/bq[16] , \pe7/ctrq , \pe7/pq , \pe8/ti_1 ,
         \pe8/ti_1t , \pe8/bq[1] , \pe8/bq[2] , \pe8/bq[3] , \pe8/bq[4] ,
         \pe8/bq[5] , \pe8/bq[6] , \pe8/bq[7] , \pe8/bq[8] , \pe8/bq[9] ,
         \pe8/bq[10] , \pe8/bq[11] , \pe8/bq[12] , \pe8/bq[13] , \pe8/bq[14] ,
         \pe8/bq[15] , \pe8/ctrq , \pe8/pq , \pe9/ti_7[14] , \pe9/ti_1 ,
         \pe9/ti_1t , \pe9/bq[1] , \pe9/bq[2] , \pe9/bq[3] , \pe9/bq[4] ,
         \pe9/bq[5] , \pe9/bq[6] , \pe9/bq[7] , \pe9/bq[8] , \pe9/bq[9] ,
         \pe9/bq[10] , \pe9/bq[11] , \pe9/bq[12] , \pe9/bq[13] , \pe9/bq[14] ,
         \pe9/bq[15] , \pe9/bq[16] , \pe9/ctrq , \pe9/pq , \pe10/ti_1 ,
         \pe10/ti_1t , \pe10/bq[1] , \pe10/bq[2] , \pe10/bq[3] , \pe10/bq[4] ,
         \pe10/bq[5] , \pe10/bq[6] , \pe10/bq[7] , \pe10/bq[8] , \pe10/bq[9] ,
         \pe10/bq[10] , \pe10/bq[11] , \pe10/bq[12] , \pe10/bq[13] ,
         \pe10/bq[14] , \pe10/bq[15] , \pe10/bq[16] , \pe10/ctrq , \pe10/pq ,
         \pe11/ti_1 , \pe11/ti_1t , \pe11/bq[1] , \pe11/bq[2] , \pe11/bq[3] ,
         \pe11/bq[4] , \pe11/bq[5] , \pe11/bq[6] , \pe11/bq[7] , \pe11/bq[8] ,
         \pe11/bq[9] , \pe11/bq[10] , \pe11/bq[11] , \pe11/bq[12] ,
         \pe11/bq[13] , \pe11/bq[14] , \pe11/bq[15] , \pe11/bq[16] ,
         \pe11/ctrq , \pe11/pq , n11800, n11801, n11802, n11803, n11804,
         n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812,
         n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820,
         n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828,
         n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
         n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844,
         n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852,
         n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860,
         n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868,
         n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
         n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
         n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
         n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900,
         n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908,
         n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916,
         n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924,
         n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932,
         n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940,
         n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
         n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956,
         n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964,
         n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972,
         n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
         n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988,
         n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
         n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004,
         n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012,
         n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
         n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028,
         n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036,
         n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044,
         n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052,
         n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060,
         n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
         n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
         n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
         n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
         n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100,
         n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108,
         n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116,
         n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124,
         n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132,
         n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140,
         n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148,
         n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156,
         n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
         n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172,
         n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180,
         n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
         n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
         n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204,
         n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
         n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
         n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
         n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236,
         n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
         n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252,
         n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
         n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268,
         n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
         n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
         n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292,
         n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
         n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
         n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
         n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324,
         n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
         n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340,
         n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348,
         n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
         n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
         n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
         n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380,
         n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
         n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396,
         n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404,
         n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
         n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420,
         n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
         n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
         n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
         n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452,
         n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460,
         n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468,
         n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
         n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484,
         n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492,
         n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
         n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
         n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
         n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
         n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
         n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540,
         n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
         n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
         n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564,
         n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
         n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
         n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588,
         n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596,
         n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604,
         n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612,
         n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620,
         n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628,
         n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636,
         n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
         n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652,
         n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660,
         n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668,
         n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676,
         n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684,
         n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692,
         n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
         n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708,
         n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
         n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
         n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732,
         n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740,
         n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
         n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756,
         n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
         n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
         n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
         n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
         n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804,
         n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812,
         n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
         n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828,
         n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
         n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
         n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852,
         n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
         n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868,
         n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876,
         n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884,
         n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892,
         n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900,
         n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908,
         n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
         n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
         n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
         n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
         n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
         n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
         n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
         n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
         n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028,
         n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
         n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
         n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
         n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
         n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
         n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
         n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
         n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212,
         n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
         n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
         n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
         n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
         n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
         n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
         n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
         n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
         n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
         n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476,
         n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
         n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
         n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
         n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508,
         n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
         n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524,
         n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
         n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
         n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
         n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
         n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
         n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
         n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
         n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692,
         n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
         n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
         n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
         n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
         n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
         n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740,
         n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
         n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756,
         n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
         n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772,
         n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780,
         n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
         n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
         n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
         n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812,
         n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
         n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828,
         n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836,
         n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844,
         n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
         n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
         n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
         n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
         n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
         n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
         n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
         n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
         n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
         n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
         n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
         n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
         n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
         n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
         n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
         n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
         n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
         n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
         n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
         n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
         n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
         n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
         n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
         n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
         n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
         n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
         n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
         n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
         n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
         n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
         n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
         n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
         n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
         n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
         n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
         n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
         n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
         n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
         n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
         n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
         n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
         n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,
         n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
         n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
         n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748,
         n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
         n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764,
         n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772,
         n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780,
         n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
         n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796,
         n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
         n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
         n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820,
         n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828,
         n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836,
         n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844,
         n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852,
         n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
         n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868,
         n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
         n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
         n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
         n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908,
         n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916,
         n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
         n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
         n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
         n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
         n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956,
         n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964,
         n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
         n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980,
         n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988,
         n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996,
         n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004,
         n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
         n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
         n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028,
         n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036,
         n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
         n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
         n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
         n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
         n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100,
         n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108,
         n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116,
         n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124,
         n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132,
         n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140,
         n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
         n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
         n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
         n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172,
         n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180,
         n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188,
         n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196,
         n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204,
         n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212,
         n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220,
         n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
         n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
         n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244,
         n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252,
         n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260,
         n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
         n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276,
         n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284,
         n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
         n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300,
         n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
         n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316,
         n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324,
         n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332,
         n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340,
         n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
         n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356,
         n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
         n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372,
         n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
         n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388,
         n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396,
         n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404,
         n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412,
         n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
         n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428,
         n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
         n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444,
         n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
         n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460,
         n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468,
         n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476,
         n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484,
         n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492,
         n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500,
         n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
         n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516,
         n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524,
         n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532,
         n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540,
         n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
         n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
         n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564,
         n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572,
         n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
         n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588,
         n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596,
         n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604,
         n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612,
         n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620,
         n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628,
         n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636,
         n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644,
         n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652,
         n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660,
         n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668,
         n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676,
         n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684,
         n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692,
         n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700,
         n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708,
         n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716,
         n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724,
         n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732,
         n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740,
         n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748,
         n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756,
         n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764,
         n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772,
         n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780,
         n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788,
         n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796,
         n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804,
         n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812,
         n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820,
         n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828,
         n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836,
         n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844,
         n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852,
         n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860,
         n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868,
         n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876,
         n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884,
         n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892,
         n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900,
         n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908,
         n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916,
         n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924,
         n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932,
         n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940,
         n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948,
         n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956,
         n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964,
         n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972,
         n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980,
         n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988,
         n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996,
         n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004,
         n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012,
         n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020,
         n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028,
         n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036,
         n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044,
         n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052,
         n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060,
         n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068,
         n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076,
         n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084,
         n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092,
         n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100,
         n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108,
         n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116,
         n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124,
         n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132,
         n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140,
         n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148,
         n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156,
         n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164,
         n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172,
         n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180,
         n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188,
         n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196,
         n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204,
         n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212,
         n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220,
         n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228,
         n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236,
         n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244,
         n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252,
         n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260,
         n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268,
         n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276,
         n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284,
         n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292,
         n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300,
         n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308,
         n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316,
         n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324,
         n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332,
         n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340,
         n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348,
         n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356,
         n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364,
         n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372,
         n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380,
         n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388,
         n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396,
         n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404,
         n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412,
         n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420,
         n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428,
         n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436,
         n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444,
         n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452,
         n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460,
         n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468,
         n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476,
         n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484,
         n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492,
         n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500,
         n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508,
         n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516,
         n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524,
         n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532,
         n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540,
         n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548,
         n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556,
         n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564,
         n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572,
         n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580,
         n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588,
         n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596,
         n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604,
         n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612,
         n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620,
         n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628,
         n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636,
         n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644,
         n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652,
         n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660,
         n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668,
         n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676,
         n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684,
         n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692,
         n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700,
         n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708,
         n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716,
         n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724,
         n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732,
         n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740,
         n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748,
         n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756,
         n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764,
         n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772,
         n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780,
         n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788,
         n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796,
         n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804,
         n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812,
         n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820,
         n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828,
         n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836,
         n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844,
         n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852,
         n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860,
         n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868,
         n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876,
         n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884,
         n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892,
         n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900,
         n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908,
         n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916,
         n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924,
         n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932,
         n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940,
         n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948,
         n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956,
         n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964,
         n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972,
         n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980,
         n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988,
         n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996,
         n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004,
         n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012,
         n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020,
         n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028,
         n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036,
         n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044,
         n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052,
         n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060,
         n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068,
         n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076,
         n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084,
         n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092,
         n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100,
         n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108,
         n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116,
         n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124,
         n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132,
         n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140,
         n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148,
         n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156,
         n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164,
         n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172,
         n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180,
         n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188,
         n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196,
         n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204,
         n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212,
         n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220,
         n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228,
         n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236,
         n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244,
         n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252,
         n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260,
         n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268,
         n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276,
         n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284,
         n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292,
         n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300,
         n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308,
         n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316,
         n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324,
         n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332,
         n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340,
         n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348,
         n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356,
         n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364,
         n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372,
         n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380,
         n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388,
         n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396,
         n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404,
         n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412,
         n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420,
         n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428,
         n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436,
         n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444,
         n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452,
         n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460,
         n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468,
         n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476,
         n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484,
         n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492,
         n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500,
         n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508,
         n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516,
         n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524,
         n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532,
         n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540,
         n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548,
         n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556,
         n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564,
         n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572,
         n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580,
         n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588,
         n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596,
         n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604,
         n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612,
         n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620,
         n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628,
         n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636,
         n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644,
         n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652,
         n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660,
         n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668,
         n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676,
         n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684,
         n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692,
         n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700,
         n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708,
         n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716,
         n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724,
         n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732,
         n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740,
         n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748,
         n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756,
         n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764,
         n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772,
         n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780,
         n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788,
         n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796,
         n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804,
         n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812,
         n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820,
         n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828,
         n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836,
         n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844,
         n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852,
         n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860,
         n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868,
         n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876,
         n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884,
         n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892,
         n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900,
         n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908,
         n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916,
         n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924,
         n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932,
         n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940,
         n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948,
         n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956,
         n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964,
         n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972,
         n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980,
         n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988,
         n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996,
         n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004,
         n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012,
         n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020,
         n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028,
         n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036,
         n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044,
         n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052,
         n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060,
         n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068,
         n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076,
         n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084,
         n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092,
         n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100,
         n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108,
         n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116,
         n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124,
         n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132,
         n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140,
         n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148,
         n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156,
         n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164,
         n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172,
         n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180,
         n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188,
         n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196,
         n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204,
         n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212,
         n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220,
         n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228,
         n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236,
         n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244,
         n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252,
         n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260,
         n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268,
         n18269, n18270, n18271, n18272, n18273, n18274, n18275, n18276,
         n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284,
         n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292,
         n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300,
         n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308,
         n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316,
         n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324,
         n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332,
         n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340,
         n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348,
         n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356,
         n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364,
         n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372,
         n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380,
         n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388,
         n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396,
         n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404,
         n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412,
         n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420,
         n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428,
         n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436,
         n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444,
         n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452,
         n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460,
         n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468,
         n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476,
         n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484,
         n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492,
         n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500,
         n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508,
         n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516,
         n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524,
         n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532,
         n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540,
         n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548,
         n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556,
         n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564,
         n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572,
         n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580,
         n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588,
         n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596,
         n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604,
         n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612,
         n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620,
         n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628,
         n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636,
         n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644,
         n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652,
         n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660,
         n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668,
         n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676,
         n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684,
         n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692,
         n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700,
         n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708,
         n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716,
         n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724,
         n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732,
         n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740,
         n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748,
         n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756,
         n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764,
         n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772,
         n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780,
         n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788,
         n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796,
         n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804,
         n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812,
         n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820,
         n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828,
         n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836,
         n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844,
         n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852,
         n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860,
         n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868,
         n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876,
         n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884,
         n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892,
         n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900,
         n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908,
         n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916,
         n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924,
         n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932,
         n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940,
         n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948,
         n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956,
         n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964,
         n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972,
         n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980,
         n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988,
         n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996,
         n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004,
         n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012,
         n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020,
         n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028,
         n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036,
         n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044,
         n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052,
         n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060,
         n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068,
         n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076,
         n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084,
         n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092,
         n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100,
         n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108,
         n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116,
         n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124,
         n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132,
         n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140,
         n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148,
         n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156,
         n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164,
         n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172,
         n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180,
         n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188,
         n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196,
         n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204,
         n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212,
         n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220,
         n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228,
         n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236,
         n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244,
         n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252,
         n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260,
         n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268,
         n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276,
         n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284,
         n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292,
         n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300,
         n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308,
         n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316,
         n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324,
         n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332,
         n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340,
         n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348,
         n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356,
         n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364,
         n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372,
         n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380,
         n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388,
         n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396,
         n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404,
         n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412,
         n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420,
         n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428,
         n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436,
         n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444,
         n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452,
         n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460,
         n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468,
         n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476,
         n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484,
         n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492,
         n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500,
         n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508,
         n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516,
         n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524,
         n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532,
         n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540,
         n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548,
         n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556,
         n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564,
         n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572,
         n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580,
         n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588,
         n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596,
         n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604,
         n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612,
         n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620,
         n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628,
         n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636,
         n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644,
         n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652,
         n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660,
         n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668,
         n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676,
         n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684,
         n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692,
         n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700,
         n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708,
         n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716,
         n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724,
         n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732,
         n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740,
         n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748,
         n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756,
         n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764,
         n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772,
         n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780,
         n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788,
         n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796,
         n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804,
         n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812,
         n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820,
         n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828,
         n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836,
         n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844,
         n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852,
         n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860,
         n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868,
         n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876,
         n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884,
         n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892,
         n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900,
         n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908,
         n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916,
         n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924,
         n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932,
         n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940,
         n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948,
         n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956,
         n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964,
         n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972,
         n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980,
         n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988,
         n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996,
         n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004,
         n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012,
         n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020,
         n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028,
         n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036,
         n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044,
         n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052,
         n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060,
         n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068,
         n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076,
         n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084,
         n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092,
         n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100,
         n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108,
         n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116,
         n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124,
         n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132,
         n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140,
         n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148,
         n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156,
         n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164,
         n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172,
         n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180,
         n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188,
         n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196,
         n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204,
         n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212,
         n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220,
         n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228,
         n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236,
         n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244,
         n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252,
         n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260,
         n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268,
         n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276,
         n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284,
         n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292,
         n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300,
         n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308,
         n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316,
         n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324,
         n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332,
         n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340,
         n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348,
         n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356,
         n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364,
         n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372,
         n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380,
         n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388,
         n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396,
         n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404,
         n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412,
         n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420,
         n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428,
         n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436,
         n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444,
         n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452,
         n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460,
         n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468,
         n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476,
         n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484,
         n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492,
         n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500,
         n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508,
         n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516,
         n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524,
         n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532,
         n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540,
         n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548,
         n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556,
         n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564,
         n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572,
         n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580,
         n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588,
         n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596,
         n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604,
         n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612,
         n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620,
         n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628,
         n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636,
         n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644,
         n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652,
         n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660,
         n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668,
         n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676,
         n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684,
         n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692,
         n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700,
         n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708,
         n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716,
         n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724,
         n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732,
         n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740,
         n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748,
         n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756,
         n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764,
         n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772,
         n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780,
         n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788,
         n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796,
         n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804,
         n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812,
         n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820,
         n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828,
         n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836,
         n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844,
         n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852,
         n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860,
         n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868,
         n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876,
         n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884,
         n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892,
         n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900,
         n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908,
         n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916,
         n20917, n20918, n20919, n20920, n20921, n20922, n20923, n20924,
         n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932,
         n20933, n20934, n20935, n20936, n20937, n20938, n20939, n20940,
         n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948,
         n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956,
         n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964,
         n20965, n20966, n20967, n20968, n20969, n20970, n20971, n20972,
         n20973, n20974, n20975, n20976, n20977, n20978, n20979, n20980,
         n20981, n20982, n20983, n20984, n20985, n20986, n20987, n20988,
         n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996,
         n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004,
         n21005, n21006, n21007, n21008, n21009, n21010, n21011, n21012,
         n21013, n21014, n21015, n21016, n21017, n21018, n21019, n21020,
         n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028,
         n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21036,
         n21037, n21038, n21039, n21040, n21041, n21042, n21043, n21044,
         n21045, n21046, n21047, n21048, n21049, n21050, n21051, n21052,
         n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060,
         n21061, n21062, n21063, n21064, n21065, n21066, n21067, n21068,
         n21069, n21070, n21071, n21072, n21073, n21074, n21075, n21076,
         n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084,
         n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092,
         n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21100,
         n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108,
         n21109, n21110, n21111, n21112, n21113, n21114, n21115, n21116,
         n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124,
         n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132,
         n21133, n21134, n21135, n21136, n21137, n21138, n21139, n21140,
         n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148,
         n21149, n21150, n21151, n21152, n21153, n21154, n21155, n21156,
         n21157, n21158, n21159, n21160, n21161, n21162, n21163, n21164,
         n21165, n21166, n21167, n21168, n21169, n21170, n21171, n21172,
         n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180,
         n21181, n21182, n21183, n21184, n21185, n21186, n21187, n21188,
         n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196,
         n21197, n21198, n21199, n21200, n21201, n21202, n21203, n21204,
         n21205, n21206, n21207, n21208, n21209, n21210, n21211, n21212,
         n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220,
         n21221, n21222, n21223, n21224, n21225, n21226, n21227, n21228,
         n21229, n21230, n21231, n21232, n21233, n21234, n21235, n21236,
         n21237, n21238, n21239, n21240, n21241, n21242, n21243, n21244,
         n21245, n21246, n21247, n21248, n21249, n21250, n21251, n21252,
         n21253, n21254, n21255, n21256, n21257, n21258, n21259, n21260,
         n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268,
         n21269, n21270, n21271, n21272, n21273, n21274, n21275, n21276,
         n21277, n21278, n21279, n21280, n21281, n21282, n21283, n21284,
         n21285, n21286, n21287, n21288, n21289, n21290, n21291, n21292,
         n21293, n21294, n21295, n21296, n21297, n21298, n21299, n21300,
         n21301, n21302, n21303, n21304, n21305, n21306, n21307, n21308,
         n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21316,
         n21317, n21318, n21319, n21320, n21321, n21322, n21323, n21324,
         n21325, n21326, n21327, n21328, n21329, n21330, n21331, n21332,
         n21333, n21334, n21335, n21336, n21337, n21338, n21339, n21340,
         n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348,
         n21349, n21350, n21351, n21352, n21353, n21354, n21355, n21356,
         n21357, n21358, n21359, n21360, n21361, n21362, n21363, n21364,
         n21365, n21366, n21367, n21368, n21369, n21370, n21371, n21372,
         n21373, n21374, n21375, n21376, n21377, n21378, n21379, n21380,
         n21381, n21382, n21383, n21384, n21385, n21386, n21387, n21388,
         n21389, n21390, n21391, n21392, n21393, n21394, n21395, n21396,
         n21397, n21398, n21399, n21400, n21401, n21402, n21403, n21404,
         n21405, n21406, n21407, n21408, n21409, n21410, n21411, n21412,
         n21413, n21414, n21415, n21416, n21417, n21418, n21419, n21420,
         n21421, n21422, n21423, n21424, n21425, n21426, n21427, n21428,
         n21429, n21430, n21431, n21432, n21433, n21434, n21435, n21436,
         n21437, n21438, n21439, n21440, n21441, n21442, n21443, n21444,
         n21445, n21446, n21447, n21448, n21449, n21450, n21451, n21452,
         n21453, n21454, n21455, n21456, n21457, n21458, n21459, n21460,
         n21461, n21462, n21463, n21464, n21465, n21466, n21467, n21468,
         n21469, n21470, n21471, n21472, n21473, n21474, n21475, n21476,
         n21477, n21478, n21479, n21480, n21481, n21482, n21483, n21484,
         n21485, n21486, n21487, n21488, n21489, n21490, n21491, n21492,
         n21493, n21494, n21495, n21496, n21497, n21498, n21499, n21500,
         n21501, n21502, n21503, n21504, n21505, n21506, n21507, n21508,
         n21509, n21510, n21511, n21512, n21513, n21514, n21515, n21516,
         n21517, n21518, n21519, n21520, n21521, n21522, n21523, n21524,
         n21525, n21526, n21527, n21528, n21529, n21530, n21531, n21532,
         n21533, n21534, n21535, n21536, n21537, n21538, n21539, n21540,
         n21541, n21542, n21543, n21544, n21545, n21546, n21547, n21548,
         n21549, n21550, n21551, n21552, n21553, n21554, n21555, n21556,
         n21557, n21558, n21559, n21560, n21561, n21562, n21563, n21564,
         n21565, n21566, n21567, n21568, n21569, n21570, n21571, n21572,
         n21573, n21574, n21575, n21576, n21577, n21578, n21579, n21580,
         n21581, n21582, n21583, n21584, n21585, n21586, n21587, n21588,
         n21589, n21590, n21591, n21592, n21593, n21594, n21595, n21596,
         n21597, n21598, n21599, n21600, n21601, n21602, n21603, n21604,
         n21605, n21606, n21607, n21608, n21609, n21610, n21611, n21612,
         n21613, n21614, n21615, n21616, n21617, n21618, n21619, n21620,
         n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21628,
         n21629, n21630, n21631, n21632, n21633, n21634, n21635, n21636,
         n21637, n21638, n21639, n21640, n21641, n21642, n21643, n21644,
         n21645, n21646, n21647, n21648, n21649, n21650, n21651, n21652,
         n21653, n21654, n21655, n21656, n21657, n21658, n21659, n21660,
         n21661, n21662, n21663, n21664, n21665, n21666, n21667, n21668,
         n21669, n21670, n21671, n21672, n21673, n21674, n21675, n21676,
         n21677, n21678, n21679, n21680, n21681, n21682, n21683, n21684,
         n21685, n21686, n21687, n21688, n21689, n21690, n21691, n21692,
         n21693, n21694, n21695, n21696, n21697, n21698, n21699, n21700,
         n21701, n21702, n21703, n21704, n21705, n21706, n21707, n21708,
         n21709, n21710, n21711, n21712, n21713, n21714, n21715, n21716,
         n21717, n21718, n21719, n21720, n21721, n21722, n21723, n21724,
         n21725, n21726, n21727, n21728, n21729, n21730, n21731, n21732,
         n21733, n21734, n21735, n21736, n21737, n21738, n21739, n21740,
         n21741, n21742, n21743, n21744, n21745, n21746, n21747, n21748,
         n21749, n21750, n21751, n21752, n21753, n21754, n21755, n21756,
         n21757, n21758, n21759, n21760, n21761, n21762, n21763, n21764,
         n21765, n21766, n21767, n21768, n21769, n21770, n21771, n21772,
         n21773, n21774, n21775, n21776, n21777, n21778, n21779, n21780,
         n21781, n21782, n21783, n21784, n21785, n21786, n21787, n21788,
         n21789, n21790, n21791, n21792, n21793, n21794, n21795, n21796,
         n21797, n21798, n21799, n21800, n21801, n21802, n21803, n21804,
         n21805, n21806, n21807, n21808, n21809, n21810, n21811, n21812,
         n21813, n21814, n21815, n21816, n21817, n21818, n21819, n21820,
         n21821, n21822, n21823, n21824, n21825, n21826, n21827, n21828,
         n21829, n21830, n21831, n21832, n21833, n21834, n21835, n21836,
         n21837, n21838, n21839, n21840, n21841, n21842, n21843, n21844,
         n21845, n21846, n21847, n21848, n21849, n21850, n21851, n21852,
         n21853, n21854, n21855, n21856, n21857, n21858, n21859, n21860,
         n21861, n21862, n21863, n21864, n21865, n21866, n21867, n21868,
         n21869, n21870, n21871, n21872, n21873, n21874, n21875, n21876,
         n21877, n21878, n21879, n21880, n21881, n21882, n21883, n21884,
         n21885, n21886, n21887, n21888, n21889, n21890, n21891, n21892,
         n21893, n21894, n21895, n21896, n21897, n21898, n21899, n21900,
         n21901, n21902, n21903, n21904, n21905, n21906, n21907, n21908,
         n21909, n21910, n21911, n21912, n21913, n21914, n21915, n21916,
         n21917, n21918, n21919, n21920, n21921, n21922, n21923, n21924,
         n21925, n21926, n21927, n21928, n21929, n21930, n21931, n21932,
         n21933, n21934, n21935, n21936, n21937, n21938, n21939, n21940,
         n21941, n21942, n21943, n21944, n21945, n21946, n21947, n21948,
         n21949, n21950, n21951, n21952, n21953, n21954, n21955, n21956,
         n21957, n21958, n21959, n21960, n21961, n21962, n21963, n21964,
         n21965, n21966, n21967, n21968, n21969, n21970, n21971, n21972,
         n21973, n21974, n21975, n21976, n21977, n21978, n21979, n21980,
         n21981, n21982, n21983, n21984, n21985, n21986, n21987, n21988,
         n21989, n21990, n21991, n21992, n21993, n21994, n21995, n21996,
         n21997, n21998, n21999, n22000, n22001, n22002, n22003, n22004,
         n22005, n22006, n22007, n22008, n22009, n22010, n22011, n22012,
         n22013, n22014, n22015, n22016, n22017, n22018, n22019, n22020,
         n22021, n22022, n22023, n22024, n22025, n22026, n22027, n22028,
         n22029, n22030, n22031, n22032, n22033, n22034, n22035, n22036,
         n22037, n22038, n22039, n22040, n22041, n22042, n22043, n22044,
         n22045, n22046, n22047, n22048, n22049, n22050, n22051, n22052,
         n22053, n22054, n22055, n22056, n22057, n22058, n22059, n22060,
         n22061, n22062, n22063, n22064, n22065, n22066, n22067, n22068,
         n22069, n22070, n22071, n22072, n22073, n22074, n22075, n22076,
         n22077, n22078, n22079, n22080, n22081, n22082, n22083, n22084,
         n22085, n22086, n22087, n22088, n22089, n22090, n22091, n22092,
         n22093, n22094, n22095, n22096, n22097, n22098, n22099, n22100,
         n22101, n22102, n22103, n22104, n22105, n22106, n22107, n22108,
         n22109, n22110, n22111, n22112, n22113, n22114, n22115, n22116,
         n22117, n22118, n22119, n22120, n22121, n22122, n22123, n22124,
         n22125, n22126, n22127, n22128, n22129, n22130, n22131, n22132,
         n22133, n22134, n22135, n22136, n22137, n22138, n22139, n22140,
         n22141, n22142, n22143, n22144, n22145, n22146, n22147, n22148,
         n22149, n22150, n22151, n22152, n22153, n22154, n22155, n22156,
         n22157, n22158, n22159, n22160, n22161, n22162, n22163, n22164,
         n22165, n22166, n22167, n22168, n22169, n22170, n22171, n22172,
         n22173, n22174, n22175, n22176, n22177, n22178, n22179, n22180,
         n22181, n22182, n22183, n22184, n22185, n22186, n22187, n22188,
         n22189, n22190, n22191, n22192, n22193, n22194, n22195, n22196,
         n22197, n22198, n22199, n22200, n22201, n22202, n22203, n22204,
         n22205, n22206, n22207, n22208, n22209, n22210, n22211, n22212,
         n22213, n22214, n22215, n22216, n22217, n22218, n22219, n22220,
         n22221, n22222, n22223, n22224, n22225, n22226, n22227, n22228,
         n22229, n22230, n22231, n22232, n22233, n22234, n22235, n22236,
         n22237, n22238, n22239, n22240, n22241, n22242, n22243, n22244,
         n22245, n22246, n22247, n22248, n22249, n22250, n22251, n22252,
         n22253, n22254, n22255, n22256, n22257, n22258, n22259, n22260,
         n22261, n22262, n22263, n22264, n22265, n22266, n22267, n22268,
         n22269, n22270, n22271, n22272, n22273, n22274, n22275, n22276,
         n22277, n22278, n22279, n22280, n22281, n22282, n22283, n22284,
         n22285, n22286, n22287, n22288, n22289, n22290, n22291, n22292,
         n22293, n22294, n22295, n22296, n22297, n22298, n22299, n22300,
         n22301, n22302, n22303, n22304, n22305, n22306, n22307, n22308,
         n22309, n22310, n22311, n22312, n22313, n22314, n22315, n22316,
         n22317, n22318, n22319, n22320, n22321, n22322, n22323, n22324,
         n22325, n22326, n22327, n22328, n22329, n22330, n22331, n22332,
         n22333, n22334, n22335, n22336, n22337, n22338, n22339, n22340,
         n22341, n22342, n22343, n22344, n22345, n22346, n22347, n22348,
         n22349, n22350, n22351, n22352, n22353, n22354, n22355, n22356,
         n22357, n22358, n22359, n22360, n22361, n22362, n22363, n22364,
         n22365, n22366, n22367, n22368, n22369, n22370, n22371, n22372,
         n22373, n22374, n22375, n22376, n22377, n22378, n22379, n22380,
         n22381, n22382, n22383, n22384, n22385, n22386, n22387, n22388,
         n22389, n22390, n22391, n22392, n22393, n22394, n22395, n22396,
         n22397, n22398, n22399, n22400, n22401, n22402, n22403, n22404,
         n22405, n22406, n22407, n22408, n22409, n22410, n22411, n22412,
         n22413, n22414, n22415, n22416, n22417, n22418, n22419, n22420,
         n22421, n22422, n22423, n22424, n22425, n22426, n22427, n22428,
         n22429, n22430, n22431, n22432, n22433, n22434, n22435, n22436,
         n22437, n22438, n22439, n22440, n22441, n22442, n22443, n22444,
         n22445, n22446, n22447, n22448, n22449, n22450, n22451, n22452,
         n22453, n22454, n22455, n22456, n22457, n22458, n22459, n22460,
         n22461, n22462, n22463, n22464, n22465, n22466, n22467, n22468,
         n22469, n22470, n22471, n22472, n22473, n22474, n22475, n22476,
         n22477, n22478, n22479, n22480, n22481, n22482, n22483, n22484,
         n22485, n22486, n22487, n22488, n22489, n22490, n22491, n22492,
         n22493, n22494, n22495, n22496, n22497, n22498, n22499, n22500,
         n22501, n22502, n22503, n22504, n22505, n22506, n22507, n22508,
         n22509, n22510, n22511, n22512, n22513, n22514, n22515, n22516,
         n22517, n22518, n22519, n22520, n22521, n22522, n22523, n22524,
         n22525, n22526, n22527, n22528, n22529, n22530, n22531, n22532,
         n22533, n22534, n22535, n22536, n22537, n22538, n22539, n22540,
         n22541, n22542, n22543, n22544, n22545, n22546, n22547, n22548,
         n22549, n22550, n22551, n22552, n22553, n22554, n22555, n22556,
         n22557, n22558, n22559, n22560, n22561, n22562, n22563, n22564,
         n22565, n22566, n22567, n22568, n22569, n22570, n22571, n22572,
         n22573, n22574, n22575, n22576, n22577, n22578, n22579, n22580,
         n22581, n22582, n22583, n22584, n22585, n22586, n22587, n22588,
         n22589, n22590, n22591, n22592, n22593, n22594, n22595, n22596,
         n22597, n22598, n22599, n22600, n22601, n22602, n22603, n22604,
         n22605, n22606, n22607, n22608, n22609, n22610, n22611, n22612,
         n22613, n22614, n22615, n22616, n22617, n22618, n22619, n22620,
         n22621, n22622, n22623, n22624, n22625, n22626, n22627, n22628,
         n22629, n22630, n22631, n22632, n22633, n22634, n22635, n22636,
         n22637, n22638, n22639, n22640, n22641, n22642, n22643, n22644,
         n22645, n22646, n22647, n22648, n22649, n22650, n22651, n22652,
         n22653, n22654, n22655, n22656, n22657, n22658, n22659, n22660,
         n22661, n22662, n22663, n22664, n22665, n22666, n22667, n22668,
         n22669, n22670, n22671, n22672, n22673, n22674, n22675, n22676,
         n22677, n22678, n22679, n22680, n22681, n22682, n22683, n22684,
         n22685, n22686, n22687, n22688, n22689, n22690, n22691, n22692,
         n22693, n22694, n22695, n22696, n22697, n22698, n22699, n22700,
         n22701, n22702, n22703, n22704, n22705, n22706, n22707, n22708,
         n22709, n22710, n22711, n22712, n22713, n22714, n22715, n22716,
         n22717, n22718, n22719, n22720, n22721, n22722, n22723, n22724,
         n22725, n22726, n22727, n22728, n22729, n22730, n22731, n22732,
         n22733, n22734, n22735, n22736, n22737, n22738, n22739, n22740,
         n22741, n22742, n22743, n22744, n22745, n22746, n22747, n22748,
         n22749, n22750, n22751, n22752, n22753, n22754, n22755, n22756,
         n22757, n22758, n22759, n22760, n22761, n22762, n22763, n22764,
         n22765, n22766, n22767, n22768, n22769, n22770, n22771, n22772,
         n22773, n22774, n22775, n22776, n22777, n22778, n22779, n22780,
         n22781, n22782, n22783, n22784, n22785, n22786, n22787, n22788,
         n22789, n22790, n22791, n22792, n22793, n22794, n22795, n22796,
         n22797, n22798, n22799, n22800, n22801, n22802, n22803, n22804,
         n22805, n22806, n22807, n22808, n22809, n22810, n22811, n22812,
         n22813, n22814, n22815, n22816, n22817, n22818, n22819, n22820,
         n22821, n22822, n22823, n22824, n22825, n22826, n22827, n22828,
         n22829, n22830, n22831, n22832, n22833, n22834, n22835, n22836,
         n22837, n22838, n22839, n22840, n22841, n22842, n22843, n22844,
         n22845, n22846, n22847, n22848, n22849, n22850, n22851, n22852,
         n22853, n22854, n22855, n22856, n22857, n22858, n22859, n22860,
         n22861, n22862, n22863, n22864, n22865, n22866, n22867, n22868,
         n22869, n22870, n22871, n22872, n22873, n22874, n22875, n22876,
         n22877, n22878, n22879, n22880, n22881, n22882, n22883, n22884,
         n22885, n22886, n22887, n22888, n22889, n22890, n22891, n22892,
         n22893, n22894, n22895, n22896, n22897, n22898, n22899, n22900,
         n22901, n22902, n22903, n22904, n22905, n22906, n22907, n22908,
         n22909, n22910, n22911, n22912, n22913, n22914, n22915, n22916,
         n22917, n22918, n22919, n22920, n22921, n22922, n22923, n22924,
         n22925, n22926, n22927, n22928, n22929, n22930, n22931, n22932,
         n22933, n22934, n22935, n22936, n22937, n22938, n22939, n22940,
         n22941, n22942, n22943, n22944, n22945, n22946, n22947, n22948,
         n22949, n22950, n22951, n22952, n22953, n22954, n22955, n22956,
         n22957, n22958, n22959, n22960, n22961, n22962, n22963, n22964,
         n22965, n22966, n22967, n22968, n22969, n22970, n22971, n22972,
         n22973, n22974, n22975, n22976, n22977, n22978, n22979, n22980,
         n22981, n22982, n22983, n22984, n22985, n22986, n22987, n22988,
         n22989, n22990, n22991, n22992, n22993, n22994, n22995, n22996,
         n22997, n22998, n22999, n23000, n23001, n23002, n23003, n23004,
         n23005, n23006, n23007, n23008, n23009, n23010, n23011, n23012,
         n23013, n23014, n23015, n23016, n23017, n23018, n23019, n23020,
         n23021, n23022, n23023, n23024, n23025, n23026, n23027, n23028,
         n23029, n23030, n23031, n23032, n23033, n23034, n23035, n23036,
         n23037, n23038, n23039, n23040, n23041, n23042, n23043, n23044,
         n23045, n23046, n23047, n23048, n23049, n23050, n23051, n23052,
         n23053, n23054, n23055, n23056, n23057, n23058, n23059, n23060,
         n23061, n23062, n23063, n23064, n23065, n23066, n23067, n23068,
         n23069, n23070, n23071, n23072, n23073, n23074, n23075, n23076,
         n23077, n23078, n23079, n23080, n23081, n23082, n23083, n23084,
         n23085, n23086, n23087, n23088, n23089, n23090, n23091, n23092,
         n23093, n23094, n23095, n23096, n23097, n23098, n23099, n23100,
         n23101, n23102, n23103, n23104, n23105, n23106, n23107, n23108,
         n23109, n23110, n23111, n23112, n23113, n23114, n23115, n23116,
         n23117, n23118, n23119, n23120, n23121, n23122, n23123, n23124,
         n23125, n23126, n23127, n23128, n23129, n23130, n23131, n23132,
         n23133, n23134, n23135, n23136, n23137, n23138, n23139, n23140,
         n23141, n23142, n23143, n23144, n23145, n23146, n23147, n23148,
         n23149, n23150, n23151, n23152, n23153, n23154, n23155, n23156,
         n23157, n23158, n23159, n23160, n23161, n23162, n23163, n23164,
         n23165, n23166, n23167, n23168, n23169, n23170, n23171, n23172,
         n23173, n23174, n23175, n23176, n23177, n23178, n23179, n23180,
         n23181, n23182, n23183, n23184, n23185, n23186, n23187, n23188,
         n23189, n23190, n23191, n23192, n23193, n23194, n23195, n23196,
         n23197, n23198, n23199, n23200, n23201, n23202, n23203, n23204,
         n23205, n23206, n23207, n23208, n23209, n23210, n23211, n23212,
         n23213, n23214, n23215, n23216, n23217, n23218, n23219, n23220,
         n23221, n23222, n23223, n23224, n23225, n23226, n23227, n23228,
         n23229, n23230, n23231, n23232, n23233, n23234, n23235, n23236,
         n23237, n23238, n23239, n23240, n23241, n23242, n23243, n23244,
         n23245, n23246, n23247, n23248, n23249, n23250, n23251, n23252,
         n23253, n23254, n23255, n23256, n23257, n23258, n23259, n23260,
         n23261, n23262, n23263, n23264, n23265, n23266, n23267, n23268,
         n23269, n23270, n23271, n23272, n23273, n23274, n23275, n23276,
         n23277, n23278, n23279, n23280, n23281, n23282, n23283, n23284,
         n23285, n23286, n23287, n23288, n23289, n23290, n23291, n23292,
         n23293, n23294, n23295, n23296, n23297, n23298, n23299, n23300,
         n23301, n23302, n23303, n23304, n23305, n23306, n23307, n23308,
         n23309, n23310, n23311, n23312, n23313, n23314, n23315, n23316,
         n23317, n23318, n23319, n23320, n23321, n23322, n23323, n23324,
         n23325, n23326, n23327, n23328, n23329, n23330, n23331, n23332,
         n23333, n23334, n23335, n23336, n23337, n23338, n23339, n23340,
         n23341, n23342, n23343, n23344, n23345, n23346, n23347, n23348,
         n23349, n23350, n23351, n23352, n23353, n23354, n23355, n23356,
         n23357, n23358, n23359, n23360, n23361, n23362, n23363, n23364,
         n23365, n23366, n23367, n23368, n23369, n23370, n23371, n23372,
         n23373, n23374, n23375, n23376, n23377, n23378, n23379, n23380,
         n23381, n23382, n23383, n23384, n23385, n23386, n23387, n23388,
         n23389, n23390, n23391, n23392, n23393, n23394, n23395, n23396,
         n23397, n23398, n23399, n23400, n23401, n23402, n23403, n23404,
         n23405, n23406, n23407, n23408, n23409, n23410, n23411, n23412,
         n23413, n23414, n23415, n23416, n23417, n23418, n23419, n23420,
         n23421, n23422, n23423, n23424, n23425, n23426, n23427, n23428,
         n23429, n23430, n23431, n23432, n23433, n23434, n23435, n23436,
         n23437, n23438, n23439, n23440, n23441, n23442, n23443, n23444,
         n23445, n23446, n23447, n23448, n23449, n23450, n23451, n23452,
         n23453, n23454, n23455, n23456, n23457, n23458, n23459, n23460,
         n23461, n23462, n23463, n23464, n23465, n23466, n23467, n23468,
         n23469, n23470, n23471, n23472, n23473, n23474, n23475, n23476,
         n23477, n23478, n23479, n23480, n23481, n23482, n23483, n23484,
         n23485, n23486, n23487, n23488, n23489, n23490, n23491, n23492,
         n23493, n23494, n23495, n23496, n23497, n23498, n23499, n23500,
         n23501, n23502, n23503, n23504, n23505, n23506, n23507, n23508,
         n23509, n23510, n23511, n23512, n23513, n23514, n23515, n23516,
         n23517, n23518, n23519, n23520, n23521, n23522, n23523, n23524,
         n23525, n23526, n23527, n23528, n23529, n23530, n23531, n23532,
         n23533, n23534, n23535, n23536, n23537, n23538, n23539, n23540,
         n23541, n23542, n23543, n23544, n23545, n23546, n23547, n23548,
         n23549, n23550, n23551, n23552, n23553, n23554, n23555, n23556,
         n23557, n23558, n23559, n23560, n23561, n23562, n23563, n23564,
         n23565, n23566, n23567, n23568, n23569, n23570, n23571, n23572,
         n23573, n23574, n23575, n23576, n23577, n23578, n23579, n23580,
         n23581, n23582, n23583, n23584, n23585, n23586, n23587, n23588,
         n23589, n23590, n23591, n23592, n23593, n23594, n23595, n23596,
         n23597, n23598, n23599, n23600, n23601, n23602, n23603, n23604,
         n23605, n23606, n23607, n23608, n23609, n23610, n23611, n23612,
         n23613, n23614, n23615, n23616, n23617, n23618, n23619, n23620,
         n23621, n23622, n23623, n23624, n23625, n23626, n23627, n23628,
         n23629, n23630, n23631, n23632, n23633, n23634, n23635, n23636,
         n23637, n23638, n23639, n23640, n23641, n23642, n23643, n23644,
         n23645, n23646, n23647, n23648, n23649, n23650, n23651, n23652,
         n23653, n23654, n23655, n23656, n23657, n23658, n23659, n23660,
         n23661, n23662, n23663, n23664, n23665, n23666, n23667, n23668,
         n23669, n23670, n23671, n23672, n23673, n23674, n23675, n23676,
         n23677, n23678, n23679, n23680, n23681, n23682, n23683, n23684,
         n23685, n23686, n23687, n23688, n23689, n23690, n23691, n23692,
         n23693, n23694, n23695, n23696, n23697, n23698, n23699, n23700,
         n23701, n23702, n23703, n23704, n23705, n23706, n23707, n23708,
         n23709, n23710, n23711, n23712, n23713, n23714, n23715, n23716,
         n23717, n23718, n23719, n23720, n23721, n23722, n23723, n23724,
         n23725, n23726, n23727, n23728, n23729, n23730, n23731, n23732,
         n23733, n23734, n23735, n23736, n23737, n23738, n23739, n23740,
         n23741, n23742, n23743, n23744, n23745, n23746, n23747, n23748,
         n23749, n23750, n23751, n23752, n23753, n23754, n23755, n23756,
         n23757, n23758, n23759, n23760, n23761, n23762, n23763, n23764,
         n23765, n23766, n23767, n23768, n23769, n23770, n23771, n23772,
         n23773, n23774, n23775, n23776, n23777, n23778, n23779, n23780,
         n23781, n23782, n23783, n23784, n23785, n23786, n23787, n23788,
         n23789, n23790, n23791, n23792, n23793, n23794, n23795, n23796,
         n23797, n23798, n23799, n23800, n23801, n23802, n23803, n23804,
         n23805, n23806, n23807, n23808, n23809, n23810, n23811, n23812,
         n23813, n23814, n23815, n23816, n23817, n23818, n23819, n23820,
         n23821, n23822, n23823, n23824, n23825, n23826, n23827, n23828,
         n23829, n23830, n23831, n23832, n23833, n23834, n23835, n23836,
         n23837, n23838, n23839, n23840, n23841, n23842, n23843, n23844,
         n23845, n23846, n23847, n23848, n23849, n23850, n23851, n23852,
         n23853, n23854, n23855, n23856, n23857, n23858, n23859, n23860,
         n23861, n23862, n23863, n23864, n23865, n23866, n23867, n23868,
         n23869, n23870, n23871, n23872, n23873, n23874, n23875, n23876,
         n23877, n23878, n23879, n23880, n23881, n23882, n23883, n23884,
         n23885, n23886, n23887, n23888, n23889, n23890, n23891, n23892,
         n23893, n23894, n23895, n23896, n23897, n23898, n23899, n23900,
         n23901, n23902, n23903, n23904, n23905, n23906, n23907, n23908,
         n23909, n23910, n23911, n23912, n23913, n23914, n23915, n23916,
         n23917, n23918, n23919, n23920, n23921, n23922, n23923, n23924,
         n23925, n23926, n23927, n23928, n23929, n23930, n23931, n23932,
         n23933, n23934, n23935, n23936, n23937, n23938, n23939, n23940,
         n23941, n23942, n23943, n23944, n23945, n23946, n23947, n23948,
         n23949, n23950, n23951, n23952, n23953, n23954, n23955, n23956,
         n23957, n23958, n23959, n23960, n23961, n23962, n23963, n23964,
         n23965, n23966, n23967, n23968, n23969, n23970, n23971, n23972,
         n23973, n23974, n23975, n23976, n23977, n23978, n23979, n23980,
         n23981, n23982, n23983, n23984, n23985, n23986, n23987, n23988,
         n23989, n23990, n23991, n23992, n23993, n23994, n23995, n23996,
         n23997, n23998, n23999, n24000, n24001, n24002, n24003, n24004,
         n24005, n24006, n24007, n24008, n24009, n24010, n24011, n24012,
         n24013, n24014, n24015, n24016, n24017, n24018, n24019, n24020,
         n24021, n24022, n24023, n24024, n24025, n24026, n24027, n24028,
         n24029, n24030, n24031, n24032, n24033, n24034, n24035, n24036,
         n24037, n24038, n24039, n24040, n24041, n24042, n24043, n24044,
         n24045, n24046, n24047, n24048, n24049, n24050, n24051, n24052,
         n24053, n24054, n24055, n24056, n24057, n24058, n24059, n24060,
         n24061, n24062, n24063, n24064, n24065, n24066, n24067, n24068,
         n24069, n24070, n24071, n24072, n24073, n24074, n24075, n24076,
         n24077, n24078, n24079, n24080, n24081, n24082, n24083, n24084,
         n24085, n24086, n24087, n24088, n24089, n24090, n24091, n24092,
         n24093, n24094, n24095, n24096, n24097, n24098, n24099, n24100,
         n24101, n24102, n24103, n24104, n24105, n24106, n24107, n24108,
         n24109, n24110, n24111, n24112, n24113, n24114, n24115, n24116,
         n24117, n24118, n24119, n24120, n24121, n24122, n24123, n24124,
         n24125, n24126, n24127, n24128, n24129, n24130, n24131, n24132,
         n24133, n24134, n24135, n24136, n24137, n24138, n24139, n24140,
         n24141, n24142, n24143, n24144, n24145, n24146, n24147, n24148,
         n24149, n24150, n24151, n24152, n24153, n24154, n24155, n24156,
         n24157, n24158, n24159, n24160, n24161, n24162, n24163, n24164,
         n24165, n24166, n24167, n24168, n24169, n24170, n24171, n24172,
         n24173, n24174, n24175, n24176, n24177, n24178, n24179, n24180,
         n24181, n24182, n24183, n24184, n24185, n24186, n24187, n24188,
         n24189, n24190, n24191, n24192, n24193, n24194, n24195, n24196,
         n24197, n24198, n24199, n24200, n24201, n24202, n24203, n24204,
         n24205, n24206, n24207, n24208, n24209, n24210, n24211, n24212,
         n24213, n24214, n24215, n24216, n24217, n24218, n24219, n24220,
         n24221, n24222, n24223, n24224, n24225, n24226, n24227, n24228,
         n24229, n24230, n24231, n24232, n24233, n24234, n24235, n24236,
         n24237, n24238, n24239, n24240, n24241, n24242, n24243, n24244,
         n24245, n24246, n24247, n24248, n24249, n24250, n24251, n24252,
         n24253, n24254, n24255, n24256, n24257, n24258, n24259, n24260,
         n24261, n24262, n24263, n24264, n24265, n24266, n24267, n24268,
         n24269, n24270, n24271, n24272, n24273, n24274, n24275, n24276,
         n24277, n24278, n24279, n24280, n24281, n24282, n24283, n24284,
         n24285, n24286, n24287, n24288, n24289, n24290, n24291, n24292,
         n24293, n24294, n24295, n24296, n24297, n24298, n24299, n24300,
         n24301, n24302, n24303, n24304, n24305, n24306, n24307, n24308,
         n24309, n24310, n24311, n24312, n24313, n24314, n24315, n24316,
         n24317, n24318, n24319, n24320, n24321, n24322, n24323, n24324,
         n24325, n24326, n24327, n24328, n24329, n24330, n24331, n24332,
         n24333, n24334, n24335, n24336, n24337, n24338, n24339, n24340,
         n24341, n24342, n24343, n24344, n24345, n24346, n24347, n24348,
         n24349, n24350, n24351, n24352, n24353, n24354, n24355, n24356,
         n24357, n24358, n24359, n24360, n24361, n24362, n24363, n24364,
         n24365, n24366, n24367, n24368, n24369, n24370, n24371, n24372,
         n24373, n24374, n24375, n24376, n24377, n24378, n24379, n24380,
         n24381, n24382, n24383, n24384, n24385, n24386, n24387, n24388,
         n24389, n24390, n24391, n24392, n24393, n24394, n24395, n24396,
         n24397, n24398, n24399, n24400, n24401, n24402, n24403, n24404,
         n24405, n24406, n24407, n24408, n24409, n24410, n24411, n24412,
         n24413, n24414, n24415, n24416, n24417, n24418, n24419, n24420,
         n24421, n24422, n24423, n24424, n24425, n24426, n24427, n24428,
         n24429, n24430, n24431, n24432, n24433, n24434, n24435, n24436,
         n24437, n24438, n24439, n24440, n24441, n24442, n24443, n24444,
         n24445, n24446, n24447, n24448, n24449, n24450, n24451, n24452,
         n24453, n24454, n24455, n24456, n24457, n24458, n24459, n24460,
         n24461, n24462, n24463, n24464, n24465, n24466, n24467, n24468,
         n24469, n24470, n24471, n24472, n24473, n24474, n24475, n24476,
         n24477, n24478, n24479, n24480, n24481, n24482, n24483, n24484,
         n24485, n24486, n24487, n24488, n24489, n24490, n24491, n24492,
         n24493, n24494, n24495, n24496, n24497, n24498, n24499, n24500,
         n24501, n24502, n24503, n24504, n24505, n24506, n24507, n24508,
         n24509, n24510, n24511, n24512, n24513, n24514, n24515, n24516,
         n24517, n24518, n24519, n24520, n24521, n24522, n24523, n24524,
         n24525, n24526, n24527, n24528, n24529, n24530, n24531, n24532,
         n24533, n24534, n24535, n24536, n24537, n24538, n24539, n24540,
         n24541, n24542, n24543, n24544, n24545, n24546, n24547, n24548,
         n24549, n24550, n24551, n24552, n24553, n24554, n24555, n24556,
         n24557, n24558, n24559, n24560, n24561, n24562, n24563, n24564,
         n24565, n24566, n24567, n24568, n24569, n24570, n24571, n24572,
         n24573, n24574, n24575, n24576, n24577, n24578, n24579, n24580,
         n24581, n24582, n24583, n24584, n24585, n24586, n24587, n24588,
         n24589, n24590, n24591, n24592, n24593, n24594, n24595, n24596,
         n24597, n24598, n24599, n24600, n24601, n24602, n24603, n24604,
         n24605, n24606, n24607, n24608, n24609, n24610, n24611, n24612,
         n24613, n24614, n24615, n24616, n24617, n24618, n24619, n24620,
         n24621, n24622, n24623, n24624, n24625, n24626, n24627, n24628,
         n24629, n24630, n24631, n24632, n24633, n24634, n24635, n24636,
         n24637, n24638, n24639, n24640, n24641, n24642, n24643, n24644,
         n24645, n24646, n24647, n24648, n24649, n24650, n24651, n24652,
         n24653, n24654, n24655, n24656, n24657, n24658, n24659, n24660,
         n24661, n24662, n24663, n24664, n24665, n24666, n24667, n24668,
         n24669, n24670, n24671, n24672, n24673, n24674, n24675, n24676,
         n24677, n24678, n24679, n24680, n24681, n24682, n24683, n24684,
         n24685, n24686, n24687, n24688, n24689, n24690, n24691, n24692,
         n24693, n24694, n24695, n24696, n24697, n24698, n24699, n24700,
         n24701, n24702, n24703, n24704, n24705, n24706, n24707, n24708,
         n24709, n24710, n24711, n24712, n24713, n24714, n24715, n24716,
         n24717, n24718, n24719, n24720, n24721, n24722, n24723, n24724,
         n24725, n24726, n24727, n24728, n24729, n24730, n24731, n24732,
         n24733, n24734, n24735, n24736, n24737, n24738, n24739, n24740,
         n24741, n24742, n24743, n24744, n24745, n24746, n24747, n24748,
         n24749, n24750, n24751, n24752, n24753, n24754, n24755, n24756,
         n24757, n24758, n24759, n24760, n24761, n24762, n24763, n24764,
         n24765, n24766, n24767, n24768, n24769, n24770, n24771, n24772,
         n24773, n24774, n24775, n24776, n24777, n24778, n24779, n24780,
         n24781, n24782, n24783, n24784, n24785, n24786, n24787, n24788,
         n24789, n24790, n24791, n24792, n24793, n24794, n24795, n24796,
         n24797, n24798, n24799, n24800, n24801, n24802, n24803, n24804,
         n24805, n24806, n24807, n24808, n24809, n24810, n24811, n24812,
         n24813, n24814, n24815, n24816, n24817, n24818, n24819, n24820,
         n24821, n24822, n24823, n24824, n24825, n24826, n24827, n24828,
         n24829, n24830, n24831, n24832, n24833, n24834, n24835, n24836,
         n24837, n24838, n24839, n24840, n24841, n24842, n24843, n24844,
         n24845, n24846, n24847, n24848, n24849, n24850, n24851, n24852,
         n24853, n24854, n24855, n24856, n24857, n24858, n24859, n24860,
         n24861, n24862, n24863, n24864, n24865, n24866, n24867, n24868,
         n24869, n24870, n24871, n24872, n24873, n24874, n24875, n24876,
         n24877, n24878, n24879, n24880, n24881, n24882, n24883, n24884,
         n24885, n24886, n24887, n24888, n24889, n24890, n24891, n24892,
         n24893, n24894, n24895, n24896, n24897, n24898, n24899, n24900,
         n24901, n24902, n24903, n24904, n24905, n24906, n24907, n24908,
         n24909, n24910, n24911, n24912, n24913, n24914, n24915, n24916,
         n24917, n24918, n24919, n24920, n24921, n24922, n24923, n24924,
         n24925, n24926, n24927, n24928, n24929, n24930, n24931, n24932,
         n24933, n24934, n24935, n24936, n24937, n24938, n24939, n24940,
         n24941, n24942, n24943, n24944, n24945, n24946, n24947, n24948,
         n24949, n24950, n24951, n24952, n24953, n24954, n24955, n24956,
         n24957, n24958, n24959, n24960, n24961, n24962, n24963, n24964,
         n24965, n24966, n24967, n24968, n24969, n24970, n24971, n24972,
         n24973, n24974, n24975, n24976, n24977, n24978, n24979, n24980,
         n24981, n24982, n24983, n24984, n24985, n24986, n24987, n24988,
         n24989, n24990, n24991, n24992, n24993, n24994, n24995, n24996,
         n24997, n24998, n24999, n25000, n25001, n25002, n25003, n25004,
         n25005, n25006, n25007, n25008, n25009, n25010, n25011, n25012,
         n25013, n25014, n25015, n25016, n25017, n25018, n25019, n25020,
         n25021, n25022, n25023, n25024, n25025, n25026, n25027, n25028,
         n25029, n25030, n25031, n25032, n25033, n25034, n25035, n25036,
         n25037, n25038, n25039, n25040, n25041, n25042, n25043, n25044,
         n25045, n25046, n25047, n25048, n25049, n25050, n25051, n25052,
         n25053, n25054, n25055, n25056, n25057, n25058, n25059, n25060,
         n25061, n25062, n25063, n25064, n25065, n25066, n25067, n25068,
         n25069, n25070, n25071, n25072, n25073, n25074, n25075, n25076,
         n25077, n25078, n25079, n25080, n25081, n25082, n25083, n25084,
         n25085, n25086, n25087, n25088, n25089, n25090, n25091, n25092,
         n25093, n25094, n25095, n25096, n25097, n25098, n25099, n25100,
         n25101, n25102, n25103, n25104, n25105, n25106, n25107, n25108,
         n25109, n25110, n25111, n25112, n25113, n25114, n25115, n25116,
         n25117, n25118, n25119, n25120, n25121, n25122, n25123, n25124,
         n25125, n25126, n25127, n25128, n25129, n25130, n25131, n25132,
         n25133, n25134, n25135, n25136, n25137, n25138, n25139, n25140,
         n25141, n25142, n25143, n25144, n25145, n25146, n25147, n25148,
         n25149, n25150, n25151, n25152, n25153, n25154, n25155, n25156,
         n25157, n25158, n25159, n25160, n25161, n25162, n25163, n25164,
         n25165, n25166, n25167, n25168, n25169, n25170, n25171, n25172,
         n25173, n25174, n25175, n25176, n25177, n25178, n25179, n25180,
         n25181, n25182, n25183, n25184, n25185, n25186, n25187, n25188,
         n25189, n25190, n25191, n25192, n25193, n25194, n25195, n25196,
         n25197, n25198, n25199, n25200, n25201, n25202, n25203, n25204,
         n25205, n25206, n25207, n25208, n25209, n25210, n25211, n25212,
         n25213, n25214, n25215, n25216, n25217, n25218, n25219, n25220,
         n25221, n25222, n25223, n25224, n25225, n25226, n25227, n25228,
         n25229, n25230, n25231, n25232, n25233, n25234, n25235, n25236,
         n25237, n25238, n25239, n25240, n25241, n25242, n25243, n25244,
         n25245, n25246, n25247, n25248, n25249, n25250, n25251, n25252,
         n25253, n25254, n25255, n25256, n25257, n25258, n25259, n25260,
         n25261, n25262, n25263, n25264, n25265, n25266, n25267, n25268,
         n25269, n25270, n25271, n25272, n25273, n25274, n25275, n25276,
         n25277, n25278, n25279, n25280, n25281, n25282, n25283, n25284,
         n25285, n25286, n25287, n25288, n25289, n25290, n25291, n25292,
         n25293, n25294, n25295, n25296, n25297, n25298, n25299, n25300,
         n25301, n25302, n25303, n25304, n25305, n25306, n25307, n25308,
         n25309, n25310, n25311, n25312, n25313, n25314, n25315, n25316,
         n25317, n25318, n25319, n25320, n25321, n25322, n25323, n25324,
         n25325, n25326, n25327, n25328, n25329, n25330, n25331, n25332,
         n25333, n25334, n25335, n25336, n25337, n25338, n25339, n25340,
         n25341, n25342, n25343, n25344, n25345, n25346, n25347, n25348,
         n25349, n25350, n25351, n25352, n25353, n25354, n25355, n25356,
         n25357, n25358, n25359, n25360, n25361, n25362, n25363, n25364,
         n25365, n25366, n25367, n25368, n25369, n25370, n25371, n25372,
         n25373, n25374, n25375, n25376, n25377, n25378, n25379, n25380,
         n25381, n25382, n25383, n25384, n25385, n25386, n25387, n25388,
         n25389, n25390, n25391, n25392, n25393, n25394, n25395, n25396,
         n25397, n25398, n25399, n25400, n25401, n25402, n25403, n25404,
         n25405, n25406, n25407, n25408, n25409, n25410, n25411, n25412,
         n25413, n25414, n25415, n25416, n25417, n25418, n25419, n25420,
         n25421, n25422, n25423, n25424, n25425, n25426, n25427, n25428,
         n25429, n25430, n25431, n25432, n25433, n25434, n25435, n25436,
         n25437, n25438, n25439, n25440, n25441, n25442, n25443, n25444,
         n25445, n25446, n25447, n25448, n25449, n25450, n25451, n25452,
         n25453, n25454, n25455, n25456, n25457, n25458, n25459, n25460,
         n25461, n25462, n25463, n25464, n25465, n25466, n25467, n25468,
         n25469, n25470, n25471, n25472, n25473, n25474, n25475, n25476,
         n25477, n25478, n25479, n25480, n25481, n25482, n25483, n25484,
         n25485, n25486, n25487, n25488, n25489, n25490, n25491, n25492,
         n25493, n25494, n25495, n25496, n25497, n25498, n25499, n25500,
         n25501, n25502, n25503, n25504, n25505, n25506, n25507, n25508,
         n25509, n25510, n25511, n25512, n25513, n25514, n25515, n25516,
         n25517, n25518, n25519, n25520, n25521, n25522, n25523, n25524,
         n25525, n25526, n25527, n25528, n25529, n25530, n25531, n25532,
         n25533, n25534, n25535, n25536, n25537, n25538, n25539, n25540,
         n25541, n25542, n25543, n25544, n25545, n25546, n25547, n25548,
         n25549, n25550, n25551, n25552, n25553, n25554, n25555, n25556,
         n25557, n25558, n25559, n25560, n25561, n25562, n25563, n25564,
         n25565, n25566, n25567, n25568, n25569, n25570, n25571, n25572,
         n25573, n25574, n25575, n25576, n25577, n25578, n25579, n25580,
         n25581, n25582, n25583, n25584, n25585, n25586, n25587, n25588,
         n25589, n25590, n25591, n25592, n25593, n25594, n25595, n25596,
         n25597, n25598, n25599, n25600, n25601, n25602, n25603, n25604,
         n25605, n25606, n25607, n25608, n25609, n25610, n25611, n25612,
         n25613, n25614, n25615, n25616, n25617, n25618, n25619, n25620,
         n25621, n25622, n25623, n25624, n25625, n25626, n25627, n25628,
         n25629, n25630, n25631, n25632, n25633, n25634, n25635, n25636,
         n25637, n25638, n25639, n25640, n25641, n25642, n25643, n25644,
         n25645, n25646, n25647, n25648, n25649, n25650, n25651, n25652,
         n25653, n25654, n25655, n25656, n25657, n25658, n25659, n25660,
         n25661, n25662, n25663, n25664, n25665, n25666, n25667, n25668,
         n25669, n25670, n25671, n25672, n25673, n25674, n25675, n25676,
         n25677, n25678, n25679, n25680, n25681, n25682, n25683, n25684,
         n25685, n25686, n25687, n25688, n25689, n25690, n25691, n25692,
         n25693, n25694, n25695, n25696, n25697, n25698, n25699, n25700,
         n25701, n25702, n25703, n25704, n25705, n25706, n25707, n25708,
         n25709, n25710, n25711, n25712, n25713, n25714, n25715, n25716,
         n25717, n25718, n25719, n25720, n25721, n25722, n25723, n25724,
         n25725, n25726, n25727, n25728, n25729, n25730, n25731, n25732,
         n25733, n25734, n25735, n25736, n25737, n25738, n25739, n25740,
         n25741, n25742, n25743, n25744, n25745, n25746, n25747, n25748,
         n25749, n25750, n25751, n25752, n25753, n25754, n25755, n25756,
         n25757, n25758, n25759, n25760, n25761, n25762, n25763, n25764,
         n25765, n25766, n25767, n25768, n25769, n25770, n25771, n25772,
         n25773, n25774, n25775, n25776, n25777, n25778, n25779, n25780,
         n25781, n25782, n25783, n25784, n25785, n25786, n25787, n25788,
         n25789, n25790, n25791, n25792, n25793, n25794, n25795, n25796,
         n25797, n25798, n25799, n25800, n25801, n25802, n25803, n25804,
         n25805, n25806, n25807, n25808, n25809, n25810, n25811, n25812,
         n25813, n25814, n25815, n25816, n25817, n25818, n25819, n25820,
         n25821, n25822, n25823, n25824, n25825, n25826, n25827, n25828,
         n25829, n25830, n25831, n25832, n25833, n25834, n25835, n25836,
         n25837, n25838, n25839, n25840, n25841, n25842, n25843, n25844,
         n25845, n25846, n25847, n25848, n25849, n25850, n25851, n25852,
         n25853, n25854, n25855, n25856, n25857, n25858, n25859, n25860,
         n25861, n25862, n25863, n25864, n25865, n25866, n25867, n25868,
         n25869, n25870, n25871, n25872, n25873, n25874, n25875, n25876,
         n25877, n25878, n25879, n25880, n25881, n25882, n25883, n25884,
         n25885, n25886, n25887, n25888, n25889, n25890, n25891, n25892,
         n25893, n25894, n25895, n25896, n25897, n25898, n25899, n25900,
         n25901, n25902, n25903, n25904, n25905, n25906, n25907, n25908,
         n25909, n25910, n25911, n25912, n25913, n25914, n25915, n25916,
         n25917, n25918, n25919, n25920, n25921, n25922, n25923, n25924,
         n25925, n25926, n25927, n25928, n25929, n25930, n25931, n25932,
         n25933, n25934, n25935, n25936, n25937, n25938, n25939, n25940,
         n25941, n25942, n25943, n25944, n25945, n25946, n25947, n25948,
         n25949, n25950, n25951, n25952, n25953, n25954, n25955, n25956,
         n25957, n25958, n25959, n25960, n25961, n25962, n25963, n25964,
         n25965, n25966, n25967, n25968, n25969, n25970, n25971, n25972,
         n25973, n25974, n25975, n25976, n25977, n25978, n25979, n25980,
         n25981, n25982, n25983, n25984, n25985, n25986, n25987, n25988,
         n25989, n25990, n25991, n25992, n25993, n25994, n25995, n25996,
         n25997, n25998, n25999, n26000, n26001, n26002, n26003, n26004,
         n26005, n26006, n26007, n26008, n26009, n26010, n26011, n26012,
         n26013, n26014, n26015, n26016, n26017, n26018, n26019, n26020,
         n26021, n26022, n26023, n26024, n26025, n26026, n26027, n26028,
         n26029, n26030, n26031, n26032, n26033, n26034, n26035, n26036,
         n26037, n26038, n26039, n26040, n26041, n26042, n26043, n26044,
         n26045, n26046, n26047, n26048, n26049, n26050, n26051, n26052,
         n26053, n26054, n26055, n26056, n26057, n26058, n26059, n26060,
         n26061, n26062, n26063, n26064, n26065, n26066, n26067, n26068,
         n26069, n26070, n26071, n26072, n26073, n26074, n26075, n26076,
         n26077, n26078, n26079, n26080, n26081, n26082, n26083, n26084,
         n26085, n26086, n26087, n26088, n26089, n26090, n26091, n26092,
         n26093, n26094, n26095, n26096, n26097, n26098, n26099, n26100,
         n26101, n26102, n26103, n26104, n26105, n26106, n26107, n26108,
         n26109, n26110, n26111, n26112, n26113, n26114, n26115, n26116,
         n26117, n26118, n26119, n26120, n26121, n26122, n26123, n26124,
         n26125, n26126, n26127, n26128, n26129, n26130, n26131, n26132,
         n26133, n26134, n26135, n26136, n26137, n26138, n26139, n26140,
         n26141, n26142, n26143, n26144, n26145, n26146, n26147, n26148,
         n26149, n26150, n26151, n26152, n26153, n26154, n26155, n26156,
         n26157, n26158, n26159, n26160, n26161, n26162, n26163, n26164,
         n26165, n26166, n26167, n26168, n26169, n26170, n26171, n26172,
         n26173, n26174, n26175, n26176, n26177, n26178, n26179, n26180,
         n26181, n26182, n26183, n26184, n26185, n26186, n26187, n26188,
         n26189, n26190, n26191, n26192, n26193, n26194, n26195, n26196,
         n26197, n26198, n26199, n26200, n26201, n26202, n26203, n26204,
         n26205, n26206, n26207, n26208, n26209, n26210, n26211, n26212,
         n26213, n26214, n26215, n26216, n26217, n26218, n26219, n26220,
         n26221, n26222, n26223, n26224, n26225, n26226, n26227, n26228,
         n26229, n26230, n26231, n26232, n26233, n26234, n26235, n26236,
         n26237, n26238, n26239, n26240, n26241, n26242, n26243, n26244,
         n26245, n26246, n26247, n26248, n26249, n26250, n26251, n26252,
         n26253, n26254, n26255, n26256, n26257, n26258, n26259, n26260,
         n26261, n26262, n26263, n26264, n26265, n26266, n26267, n26268,
         n26269, n26270, n26271, n26272, n26273, n26274, n26275, n26276,
         n26277, n26278, n26279, n26280, n26281, n26282, n26283, n26284,
         n26285, n26286, n26287, n26288, n26289, n26290, n26291, n26292,
         n26293, n26294, n26295, n26296, n26297, n26298, n26299, n26300,
         n26301, n26302, n26303, n26304, n26305, n26306, n26307, n26308,
         n26309, n26310, n26311, n26312, n26313, n26314, n26315, n26316,
         n26317, n26318, n26319, n26320, n26321, n26322, n26323, n26324,
         n26325, n26326, n26327, n26328, n26329, n26330, n26331, n26332,
         n26333, n26334, n26335, n26336, n26337, n26338, n26339, n26340,
         n26341, n26342, n26343, n26344, n26345, n26346, n26347, n26348,
         n26349, n26350, n26351, n26352, n26353, n26354, n26355, n26356,
         n26357, n26358, n26359, n26360, n26361, n26362, n26363, n26364,
         n26365, n26366, n26367, n26368, n26369, n26370, n26371, n26372,
         n26373, n26374, n26375, n26376, n26377, n26378, n26379, n26380,
         n26381, n26382, n26383, n26384, n26385, n26386, n26387, n26388,
         n26389, n26390, n26391, n26392, n26393, n26394, n26395, n26396,
         n26397, n26398, n26399, n26400, n26401, n26402, n26403, n26404,
         n26405, n26406, n26407, n26408, n26409, n26410, n26411, n26412,
         n26413, n26414, n26415, n26416, n26417, n26418, n26419, n26420,
         n26421, n26422, n26423, n26424, n26425, n26426, n26427, n26428,
         n26429, n26430, n26431, n26432, n26433, n26434, n26435, n26436,
         n26437, n26438, n26439, n26440, n26441, n26442, n26443, n26444,
         n26445, n26446, n26447, n26448, n26449, n26450, n26451, n26452,
         n26453, n26454, n26455, n26456, n26457, n26458, n26459, n26460,
         n26461, n26462, n26463, n26464, n26465, n26466, n26467, n26468,
         n26469, n26470, n26471, n26472, n26473, n26474, n26475, n26476,
         n26477, n26478, n26479, n26480, n26481, n26482, n26483, n26484,
         n26485, n26486, n26487, n26488, n26489, n26490, n26491, n26492,
         n26493, n26494, n26495, n26496, n26497, n26498, n26499, n26500,
         n26501, n26502, n26503, n26504, n26505, n26506, n26507, n26508,
         n26509, n26510, n26511, n26512, n26513, n26514, n26515, n26516,
         n26517, n26518, n26519, n26520, n26521, n26522, n26523, n26524,
         n26525, n26526, n26527, n26528, n26529, n26530, n26531, n26532,
         n26533, n26534, n26535, n26536, n26537, n26538, n26539, n26540,
         n26541, n26542, n26543, n26544, n26545, n26546, n26547, n26548,
         n26549, n26550, n26551, n26552, n26553, n26554, n26555, n26556,
         n26557, n26558, n26559, n26560, n26561, n26562, n26563, n26564,
         n26565, n26566, n26567, n26568, n26569, n26570, n26571, n26572,
         n26573, n26574, n26575, n26576, n26577, n26578, n26579, n26580,
         n26581, n26582, n26583, n26584, n26585, n26586, n26587, n26588,
         n26589, n26590, n26591, n26592, n26593, n26594, n26595, n26596,
         n26597, n26598, n26599, n26600, n26601, n26602, n26603, n26604,
         n26605, n26606, n26607, n26608, n26609, n26610, n26611, n26612,
         n26613, n26614, n26615, n26616, n26617, n26618, n26619, n26620,
         n26621, n26622, n26623, n26624, n26625, n26626, n26627, n26628,
         n26629, n26630, n26631, n26632, n26633, n26634, n26635, n26636,
         n26637, n26638, n26639, n26640, n26641, n26642, n26643, n26644,
         n26645, n26646, n26647, n26648, n26649, n26650, n26651, n26652,
         n26653, n26654, n26655, n26656, n26657, n26658, n26659, n26660,
         n26661, n26662, n26663, n26664, n26665, n26666, n26667, n26668,
         n26669, n26670, n26671, n26672, n26673, n26674, n26675, n26676,
         n26677, n26678, n26679, n26680, n26681, n26682, n26683, n26684,
         n26685, n26686, n26687, n26688, n26689, n26690, n26691, n26692,
         n26693, n26694, n26695, n26696, n26697, n26698, n26699, n26700,
         n26701, n26702, n26703, n26704, n26705, n26706, n26707, n26708,
         n26709, n26710, n26711, n26712, n26713, n26714, n26715, n26716,
         n26717, n26718, n26719, n26720, n26721, n26722, n26723, n26724,
         n26725, n26726, n26727, n26728, n26729, n26730, n26731, n26732,
         n26733, n26734, n26735, n26736, n26737, n26738, n26739, n26740,
         n26741, n26742, n26743, n26744, n26745, n26746, n26747, n26748,
         n26749, n26750, n26751, n26752, n26753, n26754, n26755, n26756,
         n26757, n26758, n26759, n26760, n26761, n26762, n26763, n26764,
         n26765, n26766, n26767, n26768, n26769, n26770, n26771, n26772,
         n26773, n26774, n26775, n26776, n26777, n26778, n26779, n26780,
         n26781, n26782, n26783, n26784, n26785, n26786, n26787, n26788,
         n26789, n26790, n26791, n26792, n26793, n26794, n26795, n26796,
         n26797, n26798, n26799, n26800, n26801, n26802, n26803, n26804,
         n26805, n26806, n26807, n26808, n26809, n26810, n26811, n26812,
         n26813, n26814, n26815, n26816, n26817, n26818, n26819, n26820,
         n26821, n26822, n26823, n26824, n26825, n26826, n26827, n26828,
         n26829, n26830, n26831, n26832, n26833, n26834, n26835, n26836,
         n26837, n26838, n26839, n26840, n26841, n26842, n26843, n26844,
         n26845, n26846, n26847, n26848, n26849, n26850, n26851, n26852,
         n26853, n26854, n26855, n26856, n26857, n26858, n26859, n26860,
         n26861, n26862, n26863, n26864, n26865, n26866, n26867, n26868,
         n26869, n26870, n26871, n26872, n26873, n26874, n26875, n26876,
         n26877, n26878, n26879, n26880, n26881, n26882, n26883, n26884,
         n26885, n26886, n26887, n26888, n26889, n26890, n26891, n26892,
         n26893, n26894, n26895, n26896, n26897, n26898, n26899, n26900,
         n26901, n26902, n26903, n26904, n26905, n26906, n26907, n26908,
         n26909, n26910, n26911, n26912, n26913, n26914, n26915, n26916,
         n26917, n26918, n26919, n26920, n26921, n26922, n26923, n26924,
         n26925, n26926, n26927, n26928, n26929, n26930, n26931, n26932,
         n26933, n26934, n26935, n26936, n26937, n26938, n26939, n26940,
         n26941, n26942, n26943, n26944, n26945, n26946, n26947, n26948,
         n26949, n26950, n26951, n26952, n26953, n26954, n26955, n26956,
         n26957, n26958, n26959, n26960, n26961, n26962, n26963, n26964,
         n26965, n26966, n26967, n26968, n26969, n26970, n26971, n26972,
         n26973, n26974, n26975, n26976, n26977, n26978, n26979, n26980,
         n26981, n26982, n26983, n26984, n26985, n26986, n26987, n26988,
         n26989, n26990, n26991, n26992, n26993, n26994, n26995, n26996,
         n26997, n26998, n26999, n27000, n27001, n27002, n27003, n27004,
         n27005, n27006, n27007, n27008, n27009, n27010, n27011, n27012,
         n27013, n27014, n27015, n27016, n27017, n27018, n27019, n27020,
         n27021, n27022, n27023, n27024, n27025, n27026, n27027, n27028,
         n27029, n27030, n27031, n27032, n27033, n27034, n27035, n27036,
         n27037, n27038, n27039, n27040, n27041, n27042, n27043, n27044,
         n27045, n27046, n27047, n27048, n27049, n27050, n27051, n27052,
         n27053, n27054, n27055, n27056, n27057, n27058, n27059, n27060,
         n27061, n27062, n27063, n27064, n27065, n27066, n27067, n27068,
         n27069, n27070, n27071, n27072, n27073, n27074, n27075, n27076,
         n27077, n27078, n27079, n27080, n27081, n27082, n27083, n27084,
         n27085, n27086, n27087, n27088, n27089, n27090, n27091, n27092,
         n27093, n27094, n27095, n27096, n27097, n27098, n27099, n27100,
         n27101, n27102, n27103, n27104, n27105, n27106, n27107, n27108,
         n27109, n27110, n27111, n27112, n27113, n27114, n27115, n27116,
         n27117, n27118, n27119, n27120, n27121, n27122, n27123, n27124,
         n27125, n27126, n27127, n27128, n27129, n27130, n27131, n27132,
         n27133, n27134, n27135, n27136, n27137, n27138, n27139, n27140,
         n27141, n27142, n27143, n27144, n27145, n27146, n27147, n27148,
         n27149, n27150, n27151, n27152, n27153, n27154, n27155, n27156,
         n27157, n27158, n27159, n27160, n27161, n27162, n27163, n27164,
         n27165, n27166, n27167, n27168, n27169, n27170, n27171, n27172,
         n27173, n27174, n27175, n27176, n27177, n27178, n27179, n27180,
         n27181, n27182, n27183, n27184, n27185, n27186, n27187, n27188,
         n27189, n27190, n27191, n27192, n27193, n27194, n27195, n27196,
         n27197, n27198, n27199, n27200, n27201, n27202, n27203, n27204,
         n27205, n27206, n27207, n27208, n27209, n27210, n27211, n27212,
         n27213, n27214, n27215, n27216, n27217, n27218, n27219, n27220,
         n27221, n27222, n27223, n27224, n27225, n27226, n27227, n27228,
         n27229, n27230, n27231, n27232, n27233, n27234, n27235, n27236,
         n27237, n27238, n27239, n27240, n27241, n27242, n27243, n27244,
         n27245, n27246, n27247, n27248, n27249, n27250, n27251, n27252,
         n27253, n27254, n27255, n27256, n27257, n27258, n27259, n27260,
         n27261, n27262, n27263, n27264, n27265, n27266, n27267, n27268,
         n27269, n27270, n27271, n27272, n27273, n27274, n27275, n27276,
         n27277, n27278, n27279, n27280, n27281, n27282, n27283, n27284,
         n27285, n27286, n27287, n27288, n27289, n27290, n27291, n27292,
         n27293, n27294, n27295, n27296, n27297, n27298, n27299, n27300,
         n27301, n27302, n27303, n27304, n27305, n27306, n27307, n27308,
         n27309, n27310, n27311, n27312, n27313, n27314, n27315, n27316,
         n27317, n27318, n27319, n27320, n27321, n27322, n27323, n27324,
         n27325, n27326, n27327, n27328, n27329, n27330, n27331, n27332,
         n27333, n27334, n27335, n27336, n27337, n27338, n27339, n27340,
         n27341, n27342, n27343, n27344, n27345, n27346, n27347, n27348,
         n27349, n27350, n27351, n27352, n27353, n27354, n27355, n27356,
         n27357, n27358, n27359, n27360, n27361, n27362, n27363, n27364,
         n27365, n27366, n27367, n27368, n27369, n27370, n27371, n27372,
         n27373, n27374, n27375, n27376, n27377, n27378, n27379, n27380,
         n27381, n27382, n27383, n27384, n27385, n27386, n27387, n27388,
         n27389, n27390, n27391, n27392, n27393, n27394, n27395, n27396,
         n27397, n27398, n27399, n27400, n27401, n27402, n27403, n27404,
         n27405, n27406, n27407, n27408, n27409, n27410, n27411, n27412,
         n27413, n27414, n27415, n27416, n27417, n27418, n27419, n27420,
         n27421, n27422, n27423, n27424, n27425, n27426, n27427, n27428,
         n27429, n27430, n27431, n27432, n27433, n27434, n27435, n27436,
         n27437, n27438, n27439, n27440, n27441, n27442, n27443, n27444,
         n27445, n27446, n27447, n27448, n27449, n27450, n27451, n27452,
         n27453, n27454, n27455, n27456, n27457, n27458, n27459, n27460,
         n27461, n27462, n27463, n27464, n27465, n27466, n27467, n27468,
         n27469, n27470, n27471, n27472, n27473, n27474, n27475, n27476,
         n27477, n27478, n27479, n27480, n27481, n27482, n27483, n27484,
         n27485, n27486, n27487, n27488, n27489, n27490, n27491, n27492,
         n27493, n27494, n27495, n27496, n27497, n27498, n27499, n27500,
         n27501, n27502, n27503, n27504, n27505, n27506, n27507, n27508,
         n27509, n27510, n27511, n27512, n27513, n27514, n27515, n27516,
         n27517, n27518, n27519, n27520, n27521, n27522, n27523, n27524,
         n27525, n27526, n27527, n27528, n27529, n27530, n27531, n27532,
         n27533, n27534, n27535, n27536, n27537, n27538, n27539, n27540,
         n27541, n27542, n27543, n27544, n27545, n27546, n27547, n27548,
         n27549, n27550, n27551, n27552, n27553, n27554, n27555, n27556,
         n27557, n27558, n27559, n27560, n27561, n27562, n27563, n27564,
         n27565, n27566, n27567, n27568, n27569, n27570, n27571, n27572,
         n27573, n27574, n27575, n27576, n27577, n27578, n27579, n27580,
         n27581, n27582, n27583, n27584, n27585, n27586, n27587, n27588,
         n27589, n27590, n27591, n27592, n27593, n27594, n27595, n27596,
         n27597, n27598, n27599, n27600, n27601, n27602, n27603, n27604,
         n27605, n27606, n27607, n27608, n27609, n27610, n27611, n27612,
         n27613, n27614, n27615, n27616, n27617, n27618, n27619, n27620,
         n27621, n27622, n27623, n27624, n27625, n27626, n27627, n27628,
         n27629, n27630, n27631, n27632, n27633, n27634, n27635, n27636,
         n27637, n27638, n27639, n27640, n27641, n27642, n27643, n27644,
         n27645, n27646, n27647, n27648, n27649, n27650, n27651, n27652,
         n27653, n27654, n27655, n27656, n27657, n27658, n27659, n27660,
         n27661, n27662, n27663, n27664, n27665, n27666, n27667, n27668,
         n27669, n27670, n27671, n27672, n27673, n27674, n27675, n27676,
         n27677, n27678, n27679, n27680, n27681, n27682, n27683, n27684,
         n27685, n27686, n27687, n27688, n27689, n27690, n27691, n27692,
         n27693, n27694, n27695, n27696, n27697, n27698, n27699, n27700,
         n27701, n27702, n27703, n27704, n27705, n27706, n27707, n27708,
         n27709, n27710, n27711, n27712, n27713, n27714, n27715, n27716,
         n27717, n27718, n27719, n27720, n27721, n27722, n27723, n27724,
         n27725, n27726, n27727, n27728, n27729, n27730, n27731, n27732,
         n27733, n27734, n27735, n27736, n27737, n27738, n27739, n27740,
         n27741, n27742, n27743, n27744, n27745, n27746, n27747, n27748,
         n27749, n27750, n27751, n27752, n27753, n27754, n27755, n27756,
         n27757, n27758, n27759, n27760, n27761, n27762, n27763, n27764,
         n27765, n27766, n27767, n27768, n27769, n27770, n27771, n27772,
         n27773, n27774, n27775, n27776, n27777, n27778, n27779, n27780,
         n27781, n27782, n27783, n27784, n27785, n27786, n27787, n27788,
         n27789, n27790, n27791, n27792, n27793, n27794, n27795, n27796,
         n27797, n27798, n27799, n27800, n27801, n27802, n27803, n27804,
         n27805, n27806, n27807, n27808, n27809, n27810, n27811, n27812,
         n27813, n27814, n27815, n27816, n27817, n27818, n27819, n27820,
         n27821, n27822, n27823, n27824, n27825, n27826, n27827, n27828,
         n27829, n27830, n27831, n27832, n27833, n27834, n27835, n27836,
         n27837, n27838, n27839, n27840, n27841, n27842, n27843, n27844,
         n27845, n27846, n27847, n27848, n27849, n27850, n27851, n27852,
         n27853, n27854, n27855, n27856, n27857, n27858, n27859, n27860,
         n27861, n27862, n27863, n27864, n27865, n27866, n27867, n27868,
         n27869, n27870, n27871, n27872, n27873, n27874, n27875, n27876,
         n27877, n27878, n27879, n27880, n27881, n27882, n27883, n27884,
         n27885, n27886, n27887, n27888, n27889, n27890, n27891, n27892,
         n27893, n27894, n27895, n27896, n27897, n27898, n27899, n27900,
         n27901, n27902, n27903, n27904, n27905, n27906, n27907, n27908,
         n27909, n27910, n27911, n27912, n27913, n27914, n27915, n27916,
         n27917, n27918, n27919, n27920, n27921, n27922, n27923, n27924,
         n27925, n27926, n27927, n27928, n27929, n27930, n27931, n27932,
         n27933, n27934, n27935, n27936, n27937, n27938, n27939, n27940,
         n27941, n27942, n27943, n27944, n27945, n27946, n27947, n27948,
         n27949, n27950, n27951, n27952, n27953, n27954, n27955, n27956,
         n27957, n27958, n27959, n27960, n27961, n27962, n27963, n27964,
         n27965, n27966, n27967, n27968, n27969, n27970, n27971, n27972,
         n27973, n27974, n27975, n27976, n27977, n27978, n27979, n27980,
         n27981, n27982, n27983, n27984, n27985, n27986, n27987, n27988,
         n27989, n27990, n27991, n27992, n27993, n27994, n27995, n27996,
         n27997, n27998, n27999, n28000, n28001, n28002, n28003, n28004,
         n28005, n28006, n28007, n28008, n28009, n28010, n28011, n28012,
         n28013, n28014, n28015, n28016, n28017, n28018, n28019, n28020,
         n28021, n28022, n28023, n28024, n28025, n28026, n28027, n28028,
         n28029, n28030, n28031, n28032, n28033, n28034, n28035, n28036,
         n28037, n28038, n28039, n28040, n28041, n28042, n28043, n28044,
         n28045, n28046, n28047, n28048, n28049, n28050, n28051, n28052,
         n28053, n28054, n28055, n28056, n28057, n28058, n28059, n28060,
         n28061, n28062, n28063, n28064, n28065, n28066, n28067, n28068,
         n28069, n28070, n28071, n28072, n28073, n28074, n28075, n28076,
         n28077, n28078, n28079, n28080, n28081, n28082, n28083, n28084,
         n28085, n28086, n28087, n28088, n28089, n28090, n28091, n28092,
         n28093, n28094, n28095, n28096, n28097, n28098, n28099, n28100,
         n28101, n28102, n28103, n28104, n28105, n28106, n28107, n28108,
         n28109, n28110, n28111, n28112, n28113, n28114, n28115, n28116,
         n28117, n28118, n28119, n28120, n28121, n28122, n28123, n28124,
         n28125, n28126, n28127, n28128, n28129, n28130, n28131, n28132,
         n28133, n28134, n28135, n28136, n28137, n28138, n28139, n28140,
         n28141, n28142, n28143, n28144, n28145, n28146, n28147, n28148,
         n28149, n28150, n28151, n28152, n28153, n28154, n28155, n28156,
         n28157, n28158, n28159, n28160, n28161, n28162, n28163, n28164,
         n28165, n28166, n28167, n28168, n28169, n28170, n28171, n28172,
         n28173, n28174, n28175, n28176, n28177, n28178, n28179, n28180,
         n28181, n28182, n28183, n28184, n28185, n28186, n28187, n28188,
         n28189, n28190, n28191, n28192, n28193, n28194, n28195, n28196,
         n28197, n28198, n28199, n28200, n28201, n28202, n28203, n28204,
         n28205, n28206, n28207, n28208, n28209, n28210, n28211, n28212,
         n28213, n28214, n28215, n28216, n28217, n28218, n28219, n28220,
         n28221, n28222, n28223, n28224, n28225, n28226, n28227, n28228,
         n28229, n28230, n28231, n28232, n28233, n28234, n28235, n28236,
         n28237, n28238, n28239, n28240, n28241, n28242, n28243, n28244,
         n28245, n28246, n28247, n28248, n28249, n28250, n28251, n28252,
         n28253, n28254, n28255, n28256, n28257, n28258, n28259, n28260,
         n28261, n28262, n28263, n28264, n28265, n28266, n28267, n28268,
         n28269, n28270, n28271, n28272, n28273, n28274, n28275, n28276,
         n28277, n28278, n28279, n28280, n28281, n28282, n28283, n28284,
         n28285, n28286, n28287, n28288, n28289, n28290, n28291, n28292,
         n28293, n28294, n28295, n28296, n28297, n28298, n28299, n28300,
         n28301, n28302, n28303, n28304, n28305, n28306, n28307, n28308,
         n28309, n28310, n28311, n28312, n28313, n28314, n28315, n28316,
         n28317, n28318, n28319, n28320, n28321, n28322, n28323, n28324,
         n28325, n28326, n28327, n28328, n28329, n28330, n28331, n28332,
         n28333, n28334, n28335, n28336, n28337, n28338, n28339, n28340,
         n28341, n28342, n28343, n28344, n28345, n28346, n28347, n28348,
         n28349, n28350, n28351, n28352, n28353, n28354, n28355, n28356,
         n28357, n28358, n28359, n28360, n28361, n28362, n28363, n28364,
         n28365, n28366, n28367, n28368, n28369, n28370, n28371, n28372,
         n28373, n28374, n28375, n28376, n28377, n28378, n28379, n28380,
         n28381, n28382, n28383, n28384, n28385, n28386, n28387, n28388,
         n28389, n28390, n28391, n28392, n28393, n28394, n28395, n28396,
         n28397, n28398, n28399, n28400, n28401, n28402, n28403, n28404,
         n28405, n28406, n28407, n28408, n28409, n28410, n28411, n28412,
         n28413, n28414, n28415, n28416, n28417, n28418, n28419, n28420,
         n28421, n28422, n28423, n28424, n28425, n28426, n28427, n28428,
         n28429, n28430, n28431, n28432, n28433, n28434, n28435, n28436,
         n28437, n28438, n28439, n28440, n28441, n28442, n28443, n28444,
         n28445, n28446, n28447, n28448, n28449, n28450, n28451, n28452,
         n28453, n28454, n28455, n28456, n28457, n28458, n28459, n28460,
         n28461, n28462, n28463, n28464, n28465, n28466, n28467, n28468,
         n28469, n28470, n28471, n28472, n28473, n28474, n28475, n28476,
         n28477, n28478, n28479, n28480, n28481, n28482, n28483, n28484,
         n28485, n28486, n28487, n28488, n28489, n28490, n28491, n28492,
         n28493, n28494, n28495, n28496, n28497, n28498, n28499, n28500,
         n28501, n28502, n28503, n28504, n28505, n28506, n28507, n28508,
         n28509, n28510, n28511, n28512, n28513, n28514, n28515, n28516,
         n28517, n28518, n28519, n28520, n28521, n28522, n28523, n28524,
         n28525, n28526, n28527, n28528, n28529, n28530, n28531, n28532,
         n28533, n28534, n28535, n28536, n28537, n28538, n28539, n28540,
         n28541, n28542, n28543, n28544, n28545, n28546, n28547, n28548,
         n28549, n28550, n28551, n28552, n28553, n28554, n28555, n28556,
         n28557, n28558, n28559, n28560, n28561, n28562, n28563, n28564,
         n28565, n28566, n28567, n28568, n28569, n28570, n28571, n28572,
         n28573, n28574, n28575, n28576, n28577, n28578, n28579, n28580,
         n28581, n28582, n28583, n28584, n28585, n28586, n28587, n28588,
         n28589, n28590, n28591, n28592, n28593, n28594, n28595, n28596,
         n28597, n28598, n28599, n28600, n28601, n28602, n28603, n28604,
         n28605, n28606, n28607, n28608, n28609, n28610, n28611, n28612,
         n28613, n28614, n28615, n28616, n28617, n28618, n28619, n28620,
         n28621, n28622, n28623, n28624, n28625, n28626, n28627, n28628,
         n28629, n28630, n28631, n28632, n28633, n28634, n28635, n28636,
         n28637, n28638, n28639, n28640, n28641, n28642, n28643, n28644,
         n28645, n28646, n28647, n28648, n28649, n28650, n28651, n28652,
         n28653, n28654, n28655, n28656, n28657, n28658, n28659, n28660,
         n28661, n28662, n28663, n28664, n28665, n28666, n28667, n28668,
         n28669, n28670, n28671, n28672, n28673, n28674, n28675, n28676,
         n28677, n28678, n28679, n28680, n28681, n28682, n28683, n28684,
         n28685, n28686, n28687, n28688, n28689, n28690, n28691, n28692,
         n28693, n28694, n28695, n28696, n28697, n28698, n28699, n28700,
         n28701, n28702, n28703, n28704, n28705, n28706, n28707, n28708,
         n28709, n28710, n28711, n28712, n28713, n28714, n28715, n28716,
         n28717, n28718, n28719, n28720, n28721, n28722, n28723, n28724,
         n28725, n28726, n28727, n28728, n28729, n28730, n28731, n28732,
         n28733, n28734, n28735, n28736, n28737, n28738, n28739, n28740,
         n28741, n28742, n28743, n28744, n28745, n28746, n28747, n28748,
         n28749, n28750, n28751, n28752, n28753, n28754, n28755, n28756,
         n28757, n28758, n28759, n28760, n28761, n28762, n28763, n28764,
         n28765, n28766, n28767, n28768, n28769, n28770, n28771, n28772,
         n28773, n28774, n28775, n28776, n28777, n28778, n28779, n28780,
         n28781, n28782, n28783, n28784, n28785, n28786, n28787, n28788,
         n28789, n28790, n28791, n28792, n28793, n28794, n28795, n28796,
         n28797, n28798, n28799, n28800, n28801, n28802, n28803, n28804,
         n28805, n28806, n28807, n28808, n28809, n28810, n28811, n28812,
         n28813, n28814, n28815, n28816, n28817, n28818, n28819, n28820,
         n28821, n28822, n28823, n28824, n28825, n28826, n28827, n28828,
         n28829, n28830, n28831, n28832, n28833, n28834, n28835, n28836,
         n28837, n28838, n28839, n28840, n28841, n28842, n28843, n28844,
         n28845, n28846, n28847, n28848, n28849, n28850, n28851, n28852,
         n28853, n28854, n28855, n28856, n28857, n28858, n28859, n28860,
         n28861, n28862, n28863, n28864, n28865, n28866, n28867, n28868,
         n28869, n28870, n28871, n28872, n28873, n28874, n28875, n28876,
         n28877, n28878, n28879, n28880, n28881, n28882, n28883, n28884,
         n28885, n28886, n28887, n28888, n28889, n28890, n28891, n28892,
         n28893, n28894, n28895, n28896, n28897, n28898, n28899, n28900,
         n28901, n28902, n28903, n28904, n28905, n28906, n28907, n28908,
         n28909, n28910, n28911, n28912, n28913, n28914, n28915, n28916,
         n28917, n28918, n28919, n28920, n28921, n28922, n28923, n28924,
         n28925, n28926, n28927, n28928, n28929, n28930, n28931, n28932,
         n28933, n28934, n28935, n28936, n28937, n28938, n28939, n28940,
         n28941, n28942, n28943, n28944, n28945, n28946, n28947, n28948,
         n28949, n28950, n28951, n28952, n28953, n28954, n28955, n28956,
         n28957, n28958, n28959, n28960, n28961, n28962, n28963, n28964,
         n28965, n28966, n28967, n28968, n28969, n28970, n28971, n28972,
         n28973, n28974, n28975, n28976, n28977, n28978, n28979, n28980,
         n28981, n28982, n28983, n28984, n28985, n28986, n28987, n28988,
         n28989, n28990, n28991, n28992, n28993, n28994, n28995, n28996,
         n28997, n28998, n28999, n29000, n29001, n29002, n29003, n29004,
         n29005, n29006, n29007, n29008, n29009, n29010, n29011, n29012,
         n29013, n29014, n29015, n29016, n29017, n29018, n29019, n29020,
         n29021, n29022, n29023, n29024, n29025, n29026, n29027, n29028,
         n29029, n29030, n29031, n29032, n29033, n29034, n29035, n29036,
         n29037, n29038, n29039, n29040, n29041, n29042, n29043, n29044,
         n29045, n29046, n29047, n29048, n29049, n29050, n29051, n29052;
  wire   [16:1] ao1;
  wire   [16:1] go1;
  wire   [16:1] bo1;
  wire   [1:15] poh1;
  wire   [1:15] pov1;
  wire   [16:1] ao2;
  wire   [16:1] go2;
  wire   [16:1] bo2;
  wire   [1:15] poh2;
  wire   [16:1] ao3;
  wire   [16:1] go3;
  wire   [16:1] bo3;
  wire   [1:15] poh3;
  wire   [1:15] pov3;
  wire   [16:1] ao4;
  wire   [16:1] go4;
  wire   [16:1] bo4;
  wire   [1:15] poh4;
  wire   [1:15] pov4;
  wire   [16:1] ao5;
  wire   [16:1] go5;
  wire   [16:1] bo5;
  wire   [1:15] poh5;
  wire   [1:15] pov5;
  wire   [16:1] ao6;
  wire   [16:1] go6;
  wire   [16:1] bo6;
  wire   [1:15] poh6;
  wire   [1:15] pov6;
  wire   [16:1] ao7;
  wire   [16:1] go7;
  wire   [16:1] bo7;
  wire   [1:15] poh7;
  wire   [16:1] ao8;
  wire   [16:1] go8;
  wire   [16:1] bo8;
  wire   [1:15] poh8;
  wire   [1:15] pov8;
  wire   [16:1] ao9;
  wire   [16:1] go9;
  wire   [16:1] bo9;
  wire   [1:15] poh9;
  wire   [1:15] pov9;
  wire   [16:1] ao10;
  wire   [16:1] go10;
  wire   [16:1] bo10;
  wire   [1:15] poh10;
  wire   [1:15] pov10;
  wire   [16:1] bo11;
  wire   [1:15] poh11;
  wire   [1:15] \pe1/poht ;
  wire   [16:1] \pe1/got ;
  wire   [16:1] \pe1/aot ;
  wire   [1:15] \pe1/ti_7t ;
  wire   [1:15] \pe2/poht ;
  wire   [16:1] \pe2/got ;
  wire   [16:1] \pe2/aot ;
  wire   [1:15] \pe2/ti_7t ;
  wire   [1:15] \pe2/phq ;
  wire   [1:15] \pe2/pvq ;
  wire   [1:15] \pe3/poht ;
  wire   [16:1] \pe3/got ;
  wire   [16:1] \pe3/aot ;
  wire   [1:15] \pe3/ti_7t ;
  wire   [1:15] \pe3/phq ;
  wire   [1:15] \pe3/pvq ;
  wire   [1:15] \pe4/poht ;
  wire   [16:1] \pe4/got ;
  wire   [16:1] \pe4/aot ;
  wire   [1:15] \pe4/ti_7t ;
  wire   [1:15] \pe4/phq ;
  wire   [1:15] \pe4/pvq ;
  wire   [1:15] \pe5/poht ;
  wire   [16:1] \pe5/got ;
  wire   [16:1] \pe5/aot ;
  wire   [1:15] \pe5/ti_7t ;
  wire   [1:15] \pe5/phq ;
  wire   [1:15] \pe5/pvq ;
  wire   [1:15] \pe6/poht ;
  wire   [16:1] \pe6/got ;
  wire   [16:1] \pe6/aot ;
  wire   [1:15] \pe6/ti_7t ;
  wire   [1:15] \pe6/phq ;
  wire   [1:15] \pe6/pvq ;
  wire   [1:15] \pe7/poht ;
  wire   [16:1] \pe7/got ;
  wire   [16:1] \pe7/aot ;
  wire   [1:15] \pe7/ti_7t ;
  wire   [1:15] \pe7/phq ;
  wire   [1:15] \pe7/pvq ;
  wire   [1:15] \pe8/poht ;
  wire   [16:1] \pe8/got ;
  wire   [16:1] \pe8/aot ;
  wire   [1:15] \pe8/ti_7t ;
  wire   [1:15] \pe8/phq ;
  wire   [1:15] \pe8/pvq ;
  wire   [1:15] \pe9/poht ;
  wire   [16:1] \pe9/got ;
  wire   [16:1] \pe9/aot ;
  wire   [1:15] \pe9/ti_7t ;
  wire   [1:15] \pe9/phq ;
  wire   [1:15] \pe9/pvq ;
  wire   [1:15] \pe10/poht ;
  wire   [16:1] \pe10/got ;
  wire   [16:1] \pe10/aot ;
  wire   [1:15] \pe10/ti_7t ;
  wire   [1:15] \pe10/phq ;
  wire   [1:15] \pe10/pvq ;
  wire   [1:15] \pe11/poht ;
  wire   [16:1] \pe11/got ;
  wire   [16:1] \pe11/aot ;
  wire   [1:15] \pe11/ti_7t ;
  wire   [1:15] \pe11/phq ;
  wire   [1:15] \pe11/pvq ;

  DRNQHSV4 \pe1/pe1/q_reg[16]  ( .D(ai[1]), .CK(clk), .RDN(n28503), .Q(
        \pe1/aot [1]) );
  DRNQHSV4 \pe1/pe1/q_reg[15]  ( .D(ai[2]), .CK(clk), .RDN(n28536), .Q(
        \pe1/aot [2]) );
  DRNQHSV4 \pe1/pe1/q_reg[14]  ( .D(ai[3]), .CK(clk), .RDN(rst), .Q(
        \pe1/aot [3]) );
  DRNQHSV4 \pe1/pe1/q_reg[12]  ( .D(ai[5]), .CK(clk), .RDN(n28490), .Q(
        \pe1/aot [5]) );
  DRNQHSV4 \pe1/pe1/q_reg[10]  ( .D(ai[7]), .CK(clk), .RDN(n28492), .Q(
        \pe1/aot [7]) );
  DRNQHSV4 \pe1/pe1/q_reg[5]  ( .D(ai[12]), .CK(clk), .RDN(rst), .Q(
        \pe1/aot [12]) );
  DRNQHSV4 \pe1/pe1/q_reg[4]  ( .D(ai[13]), .CK(clk), .RDN(n28512), .Q(
        \pe1/aot [13]) );
  DRNQHSV4 \pe1/pe1/q_reg[3]  ( .D(ai[14]), .CK(clk), .RDN(rst), .Q(
        \pe1/aot [14]) );
  DRNQHSV4 \pe1/pe1/q_reg[2]  ( .D(ai[15]), .CK(clk), .RDN(rst), .Q(
        \pe1/aot [15]) );
  DRNQHSV4 \pe1/pe1/q_reg[1]  ( .D(ai[16]), .CK(clk), .RDN(rst), .Q(
        \pe1/aot [16]) );
  DRNQHSV4 \pe1/pe2/q_reg[10]  ( .D(gi[7]), .CK(clk), .RDN(n28498), .Q(
        \pe1/got [7]) );
  DRNQHSV4 \pe1/pe2/q_reg[8]  ( .D(gi[9]), .CK(clk), .RDN(rst), .Q(
        \pe1/got [9]) );
  DRNQHSV4 \pe1/pe2/q_reg[2]  ( .D(gi[15]), .CK(clk), .RDN(n28538), .Q(
        \pe1/got [15]) );
  DRNQHSV4 \pe1/pe2/q_reg[1]  ( .D(gi[16]), .CK(clk), .RDN(rst), .Q(
        \pe1/got [16]) );
  DRNQHSV4 \pe1/pe12/q_reg[16]  ( .D(n28738), .CK(clk), .RDN(n28553), .Q(
        \pe1/bq[1] ) );
  DRNQHSV4 \pe1/pe12/q_reg[15]  ( .D(n28745), .CK(clk), .RDN(n28558), .Q(
        \pe1/bq[2] ) );
  DRNQHSV4 \pe1/pe12/q_reg[14]  ( .D(n28821), .CK(clk), .RDN(n28571), .Q(
        \pe1/bq[3] ) );
  DRNQHSV4 \pe1/pe12/q_reg[13]  ( .D(n28820), .CK(clk), .RDN(n28491), .Q(
        \pe1/bq[4] ) );
  DRNQHSV4 \pe1/pe12/q_reg[12]  ( .D(n28737), .CK(clk), .RDN(n28606), .Q(
        \pe1/bq[5] ) );
  DRNQHSV4 \pe1/pe12/q_reg[11]  ( .D(n28744), .CK(clk), .RDN(n28563), .Q(
        \pe1/bq[6] ) );
  DRNQHSV4 \pe1/pe12/q_reg[10]  ( .D(n28743), .CK(clk), .RDN(n28552), .Q(
        \pe1/bq[7] ) );
  DRNQHSV4 \pe1/pe12/q_reg[9]  ( .D(n28736), .CK(clk), .RDN(n28596), .Q(
        \pe1/bq[8] ) );
  DRNQHSV4 \pe1/pe12/q_reg[8]  ( .D(n28819), .CK(clk), .RDN(n28522), .Q(
        \pe1/bq[9] ) );
  DRNQHSV4 \pe1/pe12/q_reg[7]  ( .D(n28735), .CK(clk), .RDN(n28505), .Q(
        \pe1/bq[10] ) );
  DRNQHSV4 \pe1/pe12/q_reg[6]  ( .D(n28818), .CK(clk), .RDN(n28532), .Q(
        \pe1/bq[11] ) );
  DRNQHSV4 \pe1/pe12/q_reg[5]  ( .D(n28742), .CK(clk), .RDN(n28543), .Q(
        \pe1/bq[12] ) );
  DRNQHSV4 \pe1/pe12/q_reg[4]  ( .D(n28741), .CK(clk), .RDN(n28605), .Q(
        \pe1/bq[13] ) );
  DRNQHSV4 \pe1/pe12/q_reg[3]  ( .D(n28734), .CK(clk), .RDN(n28440), .Q(
        \pe1/bq[14] ) );
  DRNQHSV4 \pe1/pe12/q_reg[2]  ( .D(n28817), .CK(clk), .RDN(n28505), .Q(
        \pe1/bq[15] ) );
  DRNQHSV4 \pe1/pe12/q_reg[1]  ( .D(n28740), .CK(clk), .RDN(n28482), .Q(
        \pe1/bq[16] ) );
  DRNQHSV4 \pe2/pe1/q_reg[16]  ( .D(ao1[1]), .CK(clk), .RDN(n28488), .Q(
        \pe2/aot [1]) );
  DRNQHSV4 \pe2/pe1/q_reg[15]  ( .D(ao1[2]), .CK(clk), .RDN(n28489), .Q(
        \pe2/aot [2]) );
  DRNQHSV4 \pe2/pe1/q_reg[14]  ( .D(ao1[3]), .CK(clk), .RDN(n28574), .Q(
        \pe2/aot [3]) );
  DRNQHSV4 \pe2/pe1/q_reg[13]  ( .D(ao1[4]), .CK(clk), .RDN(n28559), .Q(
        \pe2/aot [4]) );
  DRNQHSV4 \pe2/pe1/q_reg[12]  ( .D(ao1[5]), .CK(clk), .RDN(n28531), .Q(
        \pe2/aot [5]) );
  DRNQHSV4 \pe2/pe1/q_reg[11]  ( .D(ao1[6]), .CK(clk), .RDN(n28507), .Q(
        \pe2/aot [6]) );
  DRNQHSV4 \pe2/pe1/q_reg[10]  ( .D(ao1[7]), .CK(clk), .RDN(n28503), .Q(
        \pe2/aot [7]) );
  DRNQHSV4 \pe2/pe1/q_reg[9]  ( .D(ao1[8]), .CK(clk), .RDN(n28451), .Q(
        \pe2/aot [8]) );
  DRNQHSV4 \pe2/pe1/q_reg[8]  ( .D(ao1[9]), .CK(clk), .RDN(n28525), .Q(
        \pe2/aot [9]) );
  DRNQHSV4 \pe2/pe1/q_reg[7]  ( .D(ao1[10]), .CK(clk), .RDN(n28443), .Q(
        \pe2/aot [10]) );
  DRNQHSV4 \pe2/pe1/q_reg[6]  ( .D(ao1[11]), .CK(clk), .RDN(n28446), .Q(
        \pe2/aot [11]) );
  DRNQHSV4 \pe2/pe1/q_reg[5]  ( .D(ao1[12]), .CK(clk), .RDN(n28477), .Q(
        \pe2/aot [12]) );
  DRNQHSV4 \pe2/pe1/q_reg[4]  ( .D(ao1[13]), .CK(clk), .RDN(n28505), .Q(
        \pe2/aot [13]) );
  DRNQHSV4 \pe2/pe1/q_reg[3]  ( .D(ao1[14]), .CK(clk), .RDN(n28503), .Q(
        \pe2/aot [14]) );
  DRNQHSV4 \pe2/pe1/q_reg[2]  ( .D(ao1[15]), .CK(clk), .RDN(n28522), .Q(
        \pe2/aot [15]) );
  DRNQHSV4 \pe2/pe1/q_reg[1]  ( .D(ao1[16]), .CK(clk), .RDN(n28512), .Q(
        \pe2/aot [16]) );
  DRNQHSV4 \pe2/pe2/q_reg[16]  ( .D(go1[1]), .CK(clk), .RDN(n28497), .Q(
        \pe2/got [1]) );
  DRNQHSV4 \pe2/pe2/q_reg[15]  ( .D(go1[2]), .CK(clk), .RDN(n28494), .Q(
        \pe2/got [2]) );
  DRNQHSV4 \pe2/pe2/q_reg[14]  ( .D(go1[3]), .CK(clk), .RDN(n28515), .Q(
        \pe2/got [3]) );
  DRNQHSV4 \pe2/pe2/q_reg[13]  ( .D(go1[4]), .CK(clk), .RDN(n28477), .Q(
        \pe2/got [4]) );
  DRNQHSV4 \pe2/pe2/q_reg[12]  ( .D(go1[5]), .CK(clk), .RDN(n28448), .Q(
        \pe2/got [5]) );
  DRNQHSV4 \pe2/pe2/q_reg[11]  ( .D(go1[6]), .CK(clk), .RDN(rst), .Q(
        \pe2/got [6]) );
  DRNQHSV4 \pe2/pe2/q_reg[10]  ( .D(go1[7]), .CK(clk), .RDN(n28562), .Q(
        \pe2/got [7]) );
  DRNQHSV4 \pe2/pe2/q_reg[9]  ( .D(go1[8]), .CK(clk), .RDN(n28446), .Q(
        \pe2/got [8]) );
  DRNQHSV4 \pe2/pe2/q_reg[8]  ( .D(go1[9]), .CK(clk), .RDN(n28548), .Q(
        \pe2/got [9]) );
  DRNQHSV4 \pe2/pe2/q_reg[7]  ( .D(go1[10]), .CK(clk), .RDN(n28549), .Q(
        \pe2/got [10]) );
  DRNQHSV4 \pe2/pe2/q_reg[6]  ( .D(go1[11]), .CK(clk), .RDN(n28491), .Q(
        \pe2/got [11]) );
  DRNQHSV4 \pe2/pe2/q_reg[5]  ( .D(go1[12]), .CK(clk), .RDN(n28501), .Q(
        \pe2/got [12]) );
  DRNQHSV4 \pe2/pe2/q_reg[4]  ( .D(go1[13]), .CK(clk), .RDN(n28554), .Q(
        \pe2/got [13]) );
  DRNQHSV4 \pe2/pe2/q_reg[3]  ( .D(go1[14]), .CK(clk), .RDN(n28494), .Q(
        \pe2/got [14]) );
  DRNQHSV4 \pe2/pe2/q_reg[2]  ( .D(go1[15]), .CK(clk), .RDN(n28498), .Q(
        \pe2/got [15]) );
  DRNQHSV4 \pe2/pe2/q_reg[1]  ( .D(go1[16]), .CK(clk), .RDN(n28442), .Q(
        \pe2/got [16]) );
  DRNQHSV4 \pe2/pe5/q_reg[12]  ( .D(pov1[12]), .CK(clk), .RDN(n28504), .Q(
        \pe2/pvq [12]) );
  DRNQHSV4 \pe2/pe5/q_reg[11]  ( .D(n28976), .CK(clk), .RDN(n28606), .Q(
        \pe2/pvq [11]) );
  DRNQHSV4 \pe2/pe5/q_reg[9]  ( .D(n29047), .CK(clk), .RDN(n28539), .Q(
        \pe2/pvq [9]) );
  DRNQHSV4 \pe2/pe5/q_reg[8]  ( .D(n29048), .CK(clk), .RDN(n28482), .Q(
        \pe2/pvq [8]) );
  DRNQHSV4 \pe2/pe5/q_reg[6]  ( .D(pov1[6]), .CK(clk), .RDN(n28574), .Q(
        \pe2/pvq [6]) );
  DRNQHSV4 \pe2/pe5/q_reg[4]  ( .D(n29049), .CK(clk), .RDN(n28482), .Q(
        \pe2/pvq [4]) );
  DRNQHSV4 \pe2/pe5/q_reg[2]  ( .D(n29051), .CK(clk), .RDN(n28531), .Q(
        \pe2/pvq [2]) );
  DRNQHSV4 \pe2/pe6/q_reg[15]  ( .D(poh1[15]), .CK(clk), .RDN(n28516), .Q(
        \pe2/phq [15]) );
  DRNQHSV4 \pe2/pe6/q_reg[14]  ( .D(poh1[14]), .CK(clk), .RDN(n28602), .Q(
        \pe2/phq [14]) );
  DRNQHSV4 \pe2/pe6/q_reg[13]  ( .D(poh1[13]), .CK(clk), .RDN(n28489), .Q(
        \pe2/phq [13]) );
  DRNQHSV4 \pe2/pe6/q_reg[12]  ( .D(poh1[12]), .CK(clk), .RDN(n28572), .Q(
        \pe2/phq [12]) );
  DRNQHSV4 \pe2/pe6/q_reg[11]  ( .D(poh1[11]), .CK(clk), .RDN(n28576), .Q(
        \pe2/phq [11]) );
  DRNQHSV4 \pe2/pe6/q_reg[10]  ( .D(poh1[10]), .CK(clk), .RDN(n28525), .Q(
        \pe2/phq [10]) );
  DRNQHSV4 \pe2/pe6/q_reg[9]  ( .D(poh1[9]), .CK(clk), .RDN(n28488), .Q(
        \pe2/phq [9]) );
  DRNQHSV4 \pe2/pe6/q_reg[8]  ( .D(poh1[8]), .CK(clk), .RDN(n28491), .Q(
        \pe2/phq [8]) );
  DRNQHSV4 \pe2/pe6/q_reg[7]  ( .D(poh1[7]), .CK(clk), .RDN(n28453), .Q(
        \pe2/phq [7]) );
  DRNQHSV4 \pe2/pe6/q_reg[6]  ( .D(poh1[6]), .CK(clk), .RDN(n28513), .Q(
        \pe2/phq [6]) );
  DRNQHSV4 \pe2/pe6/q_reg[5]  ( .D(poh1[5]), .CK(clk), .RDN(n28510), .Q(
        \pe2/phq [5]) );
  DRNQHSV4 \pe2/pe6/q_reg[4]  ( .D(poh1[4]), .CK(clk), .RDN(n28508), .Q(
        \pe2/phq [4]) );
  DRNQHSV4 \pe2/pe6/q_reg[3]  ( .D(poh1[3]), .CK(clk), .RDN(n28453), .Q(
        \pe2/phq [3]) );
  DRNQHSV4 \pe2/pe6/q_reg[2]  ( .D(poh1[2]), .CK(clk), .RDN(n28547), .Q(
        \pe2/phq [2]) );
  DRNQHSV4 \pe2/pe6/q_reg[1]  ( .D(poh1[1]), .CK(clk), .RDN(n28563), .Q(
        \pe2/phq [1]) );
  DRNQHSV4 \pe2/pe7/q_reg  ( .D(n28802), .CK(clk), .RDN(n28571), .Q(\pe2/ctrq ) );
  DRNQHSV4 \pe2/pe12/q_reg[16]  ( .D(n28836), .CK(clk), .RDN(n28510), .Q(
        \pe2/bq[1] ) );
  DRNQHSV4 \pe2/pe12/q_reg[15]  ( .D(n28834), .CK(clk), .RDN(n28577), .Q(
        \pe2/bq[2] ) );
  DRNQHSV4 \pe2/pe12/q_reg[14]  ( .D(n28837), .CK(clk), .RDN(n28451), .Q(
        \pe2/bq[3] ) );
  DRNQHSV4 \pe2/pe12/q_reg[13]  ( .D(n28731), .CK(clk), .RDN(n28563), .Q(
        \pe2/bq[4] ) );
  DRNQHSV4 \pe2/pe12/q_reg[12]  ( .D(n28832), .CK(clk), .RDN(n28573), .Q(
        \pe2/bq[5] ) );
  DRNQHSV4 \pe2/pe12/q_reg[11]  ( .D(n28833), .CK(clk), .RDN(n28529), .Q(
        \pe2/bq[6] ) );
  DRNQHSV4 \pe2/pe12/q_reg[10]  ( .D(n28830), .CK(clk), .RDN(n28556), .Q(
        \pe2/bq[7] ) );
  DRNQHSV4 \pe2/pe12/q_reg[9]  ( .D(n28831), .CK(clk), .RDN(n28534), .Q(
        \pe2/bq[8] ) );
  DRNQHSV4 \pe2/pe12/q_reg[8]  ( .D(n28827), .CK(clk), .RDN(n28515), .Q(
        \pe2/bq[9] ) );
  DRNQHSV4 \pe2/pe12/q_reg[7]  ( .D(n28826), .CK(clk), .RDN(n28560), .Q(
        \pe2/bq[10] ) );
  DRNQHSV4 \pe2/pe12/q_reg[6]  ( .D(n28828), .CK(clk), .RDN(n28493), .Q(
        \pe2/bq[11] ) );
  DRNQHSV4 \pe2/pe12/q_reg[5]  ( .D(n28829), .CK(clk), .RDN(n28525), .Q(
        \pe2/bq[12] ) );
  DRNQHSV4 \pe2/pe12/q_reg[4]  ( .D(n28825), .CK(clk), .RDN(n28541), .Q(
        \pe2/bq[13] ) );
  DRNQHSV4 \pe2/pe12/q_reg[3]  ( .D(n28824), .CK(clk), .RDN(n28563), .Q(
        \pe2/bq[14] ) );
  DRNQHSV4 \pe2/pe12/q_reg[2]  ( .D(n28823), .CK(clk), .RDN(n28534), .Q(
        \pe2/bq[15] ) );
  DRNQHSV4 \pe2/pe12/q_reg[1]  ( .D(n28822), .CK(clk), .RDN(n28555), .Q(
        \pe2/bq[16] ) );
  DRNQHSV4 \pe2/pe13/q_reg  ( .D(\pe2/ti_1t ), .CK(clk), .RDN(n28495), .Q(
        \pe2/ti_1 ) );
  DRNQHSV4 \pe2/pe14/q_reg[2]  ( .D(n28953), .CK(clk), .RDN(n28576), .Q(
        \pe2/ti_7t [2]) );
  DRNQHSV4 \pe3/pe1/q_reg[16]  ( .D(ao2[1]), .CK(clk), .RDN(n28529), .Q(
        \pe3/aot [1]) );
  DRNQHSV4 \pe3/pe1/q_reg[15]  ( .D(ao2[2]), .CK(clk), .RDN(n28452), .Q(
        \pe3/aot [2]) );
  DRNQHSV4 \pe3/pe1/q_reg[14]  ( .D(ao2[3]), .CK(clk), .RDN(n28487), .Q(
        \pe3/aot [3]) );
  DRNQHSV4 \pe3/pe1/q_reg[13]  ( .D(ao2[4]), .CK(clk), .RDN(n28496), .Q(
        \pe3/aot [4]) );
  DRNQHSV4 \pe3/pe1/q_reg[12]  ( .D(ao2[5]), .CK(clk), .RDN(n28439), .Q(
        \pe3/aot [5]) );
  DRNQHSV4 \pe3/pe1/q_reg[11]  ( .D(ao2[6]), .CK(clk), .RDN(n28441), .Q(
        \pe3/aot [6]) );
  DRNQHSV4 \pe3/pe1/q_reg[10]  ( .D(ao2[7]), .CK(clk), .RDN(n28452), .Q(
        \pe3/aot [7]) );
  DRNQHSV4 \pe3/pe1/q_reg[9]  ( .D(ao2[8]), .CK(clk), .RDN(n28596), .Q(
        \pe3/aot [8]) );
  DRNQHSV4 \pe3/pe1/q_reg[8]  ( .D(ao2[9]), .CK(clk), .RDN(n28538), .Q(
        \pe3/aot [9]) );
  DRNQHSV4 \pe3/pe1/q_reg[7]  ( .D(ao2[10]), .CK(clk), .RDN(n28551), .Q(
        \pe3/aot [10]) );
  DRNQHSV4 \pe3/pe1/q_reg[6]  ( .D(ao2[11]), .CK(clk), .RDN(n28442), .Q(
        \pe3/aot [11]) );
  DRNQHSV4 \pe3/pe1/q_reg[5]  ( .D(ao2[12]), .CK(clk), .RDN(n28510), .Q(
        \pe3/aot [12]) );
  DRNQHSV4 \pe3/pe1/q_reg[4]  ( .D(ao2[13]), .CK(clk), .RDN(n28452), .Q(
        \pe3/aot [13]) );
  DRNQHSV4 \pe3/pe1/q_reg[3]  ( .D(ao2[14]), .CK(clk), .RDN(n28554), .Q(
        \pe3/aot [14]) );
  DRNQHSV4 \pe3/pe1/q_reg[2]  ( .D(ao2[15]), .CK(clk), .RDN(n28550), .Q(
        \pe3/aot [15]) );
  DRNQHSV4 \pe3/pe1/q_reg[1]  ( .D(ao2[16]), .CK(clk), .RDN(n28551), .Q(
        \pe3/aot [16]) );
  DRNQHSV4 \pe3/pe2/q_reg[16]  ( .D(go2[1]), .CK(clk), .RDN(n28506), .Q(
        \pe3/got [1]) );
  DRNQHSV4 \pe3/pe2/q_reg[15]  ( .D(go2[2]), .CK(clk), .RDN(n28555), .Q(
        \pe3/got [2]) );
  DRNQHSV4 \pe3/pe2/q_reg[14]  ( .D(go2[3]), .CK(clk), .RDN(n28486), .Q(
        \pe3/got [3]) );
  DRNQHSV4 \pe3/pe2/q_reg[13]  ( .D(go2[4]), .CK(clk), .RDN(n28602), .Q(
        \pe3/got [4]) );
  DRNQHSV4 \pe3/pe2/q_reg[12]  ( .D(go2[5]), .CK(clk), .RDN(n28550), .Q(
        \pe3/got [5]) );
  DRNQHSV4 \pe3/pe2/q_reg[11]  ( .D(go2[6]), .CK(clk), .RDN(n28521), .Q(
        \pe3/got [6]) );
  DRNQHSV4 \pe3/pe2/q_reg[10]  ( .D(go2[7]), .CK(clk), .RDN(n28504), .Q(
        \pe3/got [7]) );
  DRNQHSV4 \pe3/pe2/q_reg[9]  ( .D(go2[8]), .CK(clk), .RDN(n28518), .Q(
        \pe3/got [8]) );
  DRNQHSV4 \pe3/pe2/q_reg[8]  ( .D(go2[9]), .CK(clk), .RDN(n28546), .Q(
        \pe3/got [9]) );
  DRNQHSV4 \pe3/pe2/q_reg[7]  ( .D(go2[10]), .CK(clk), .RDN(n28532), .Q(
        \pe3/got [10]) );
  DRNQHSV4 \pe3/pe2/q_reg[6]  ( .D(go2[11]), .CK(clk), .RDN(n28497), .Q(
        \pe3/got [11]) );
  DRNQHSV4 \pe3/pe2/q_reg[5]  ( .D(go2[12]), .CK(clk), .RDN(n28439), .Q(
        \pe3/got [12]) );
  DRNQHSV4 \pe3/pe2/q_reg[4]  ( .D(go2[13]), .CK(clk), .RDN(n28442), .Q(
        \pe3/got [13]) );
  DRNQHSV4 \pe3/pe2/q_reg[3]  ( .D(go2[14]), .CK(clk), .RDN(n28440), .Q(
        \pe3/got [14]) );
  DRNQHSV4 \pe3/pe2/q_reg[2]  ( .D(go2[15]), .CK(clk), .RDN(n28553), .Q(
        \pe3/got [15]) );
  DRNQHSV4 \pe3/pe2/q_reg[1]  ( .D(go2[16]), .CK(clk), .RDN(n28506), .Q(
        \pe3/got [16]) );
  DRNQHSV4 \pe3/pe5/q_reg[10]  ( .D(\pov2[10] ), .CK(clk), .RDN(n28576), .Q(
        \pe3/pvq [10]) );
  DRNQHSV4 \pe3/pe5/q_reg[7]  ( .D(n29040), .CK(clk), .RDN(n28510), .Q(
        \pe3/pvq [7]) );
  DRNQHSV4 \pe3/pe5/q_reg[5]  ( .D(n29042), .CK(clk), .RDN(n28577), .Q(
        \pe3/pvq [5]) );
  DRNQHSV4 \pe3/pe5/q_reg[2]  ( .D(n29045), .CK(clk), .RDN(n28544), .Q(
        \pe3/pvq [2]) );
  DRNQHSV4 \pe3/pe6/q_reg[15]  ( .D(poh2[15]), .CK(clk), .RDN(n28546), .Q(
        \pe3/phq [15]) );
  DRNQHSV4 \pe3/pe6/q_reg[14]  ( .D(poh2[14]), .CK(clk), .RDN(n28476), .Q(
        \pe3/phq [14]) );
  DRNQHSV4 \pe3/pe6/q_reg[13]  ( .D(poh2[13]), .CK(clk), .RDN(n28560), .Q(
        \pe3/phq [13]) );
  DRNQHSV4 \pe3/pe6/q_reg[12]  ( .D(poh2[12]), .CK(clk), .RDN(n28546), .Q(
        \pe3/phq [12]) );
  DRNQHSV4 \pe3/pe6/q_reg[11]  ( .D(poh2[11]), .CK(clk), .RDN(n28514), .Q(
        \pe3/phq [11]) );
  DRNQHSV4 \pe3/pe6/q_reg[10]  ( .D(poh2[10]), .CK(clk), .RDN(n28502), .Q(
        \pe3/phq [10]) );
  DRNQHSV4 \pe3/pe6/q_reg[9]  ( .D(poh2[9]), .CK(clk), .RDN(n28605), .Q(
        \pe3/phq [9]) );
  DRNQHSV4 \pe3/pe6/q_reg[8]  ( .D(poh2[8]), .CK(clk), .RDN(n28501), .Q(
        \pe3/phq [8]) );
  DRNQHSV4 \pe3/pe6/q_reg[7]  ( .D(poh2[7]), .CK(clk), .RDN(n28484), .Q(
        \pe3/phq [7]) );
  DRNQHSV4 \pe3/pe6/q_reg[6]  ( .D(poh2[6]), .CK(clk), .RDN(n28500), .Q(
        \pe3/phq [6]) );
  DRNQHSV4 \pe3/pe6/q_reg[5]  ( .D(poh2[5]), .CK(clk), .RDN(n28492), .Q(
        \pe3/phq [5]) );
  DRNQHSV4 \pe3/pe6/q_reg[4]  ( .D(poh2[4]), .CK(clk), .RDN(n28527), .Q(
        \pe3/phq [4]) );
  DRNQHSV4 \pe3/pe6/q_reg[3]  ( .D(poh2[3]), .CK(clk), .RDN(n28605), .Q(
        \pe3/phq [3]) );
  DRNQHSV4 \pe3/pe6/q_reg[2]  ( .D(poh2[2]), .CK(clk), .RDN(n28458), .Q(
        \pe3/phq [2]) );
  DRNQHSV4 \pe3/pe6/q_reg[1]  ( .D(poh2[1]), .CK(clk), .RDN(n28534), .Q(
        \pe3/phq [1]) );
  DRNQHSV4 \pe3/pe7/q_reg  ( .D(n28932), .CK(clk), .RDN(n28573), .Q(\pe3/ctrq ) );
  DRNQHSV4 \pe3/pe12/q_reg[16]  ( .D(n28853), .CK(clk), .RDN(n28573), .Q(
        \pe3/bq[1] ) );
  DRNQHSV4 \pe3/pe12/q_reg[15]  ( .D(n28852), .CK(clk), .RDN(n28458), .Q(
        \pe3/bq[2] ) );
  DRNQHSV4 \pe3/pe12/q_reg[14]  ( .D(n28850), .CK(clk), .RDN(n28534), .Q(
        \pe3/bq[3] ) );
  DRNQHSV4 \pe3/pe12/q_reg[13]  ( .D(n28851), .CK(clk), .RDN(n14023), .Q(
        \pe3/bq[4] ) );
  DRNQHSV4 \pe3/pe12/q_reg[12]  ( .D(n28849), .CK(clk), .RDN(n28453), .Q(
        \pe3/bq[5] ) );
  DRNQHSV4 \pe3/pe12/q_reg[11]  ( .D(n28848), .CK(clk), .RDN(n28560), .Q(
        \pe3/bq[6] ) );
  DRNQHSV4 \pe3/pe12/q_reg[10]  ( .D(n28847), .CK(clk), .RDN(n28537), .Q(
        \pe3/bq[7] ) );
  DRNQHSV4 \pe3/pe12/q_reg[9]  ( .D(n28846), .CK(clk), .RDN(n28569), .Q(
        \pe3/bq[8] ) );
  DRNQHSV4 \pe3/pe12/q_reg[8]  ( .D(n28843), .CK(clk), .RDN(rst), .Q(
        \pe3/bq[9] ) );
  DRNQHSV4 \pe3/pe12/q_reg[7]  ( .D(n28844), .CK(clk), .RDN(n14021), .Q(
        \pe3/bq[10] ) );
  DRNQHSV4 \pe3/pe12/q_reg[6]  ( .D(n28845), .CK(clk), .RDN(n28501), .Q(
        \pe3/bq[11] ) );
  DRNQHSV4 \pe3/pe12/q_reg[5]  ( .D(n28840), .CK(clk), .RDN(n28568), .Q(
        \pe3/bq[12] ) );
  DRNQHSV4 \pe3/pe12/q_reg[4]  ( .D(n28839), .CK(clk), .RDN(n28450), .Q(
        \pe3/bq[13] ) );
  DRNQHSV4 \pe3/pe12/q_reg[3]  ( .D(n28841), .CK(clk), .RDN(n28565), .Q(
        \pe3/bq[14] ) );
  DRNQHSV4 \pe3/pe12/q_reg[2]  ( .D(n28842), .CK(clk), .RDN(n28565), .Q(
        \pe3/bq[15] ) );
  DRNQHSV4 \pe3/pe12/q_reg[1]  ( .D(n28838), .CK(clk), .RDN(n28573), .Q(
        \pe3/bq[16] ) );
  DRNQHSV4 \pe3/pe13/q_reg  ( .D(\pe3/ti_1t ), .CK(clk), .RDN(n28516), .Q(
        \pe3/ti_1 ) );
  DRNQHSV4 \pe4/pe1/q_reg[16]  ( .D(ao3[1]), .CK(clk), .RDN(n28494), .Q(
        \pe4/aot [1]) );
  DRNQHSV4 \pe4/pe1/q_reg[15]  ( .D(ao3[2]), .CK(clk), .RDN(n28519), .Q(
        \pe4/aot [2]) );
  DRNQHSV4 \pe4/pe1/q_reg[14]  ( .D(ao3[3]), .CK(clk), .RDN(n28488), .Q(
        \pe4/aot [3]) );
  DRNQHSV4 \pe4/pe1/q_reg[13]  ( .D(ao3[4]), .CK(clk), .RDN(n28501), .Q(
        \pe4/aot [4]) );
  DRNQHSV4 \pe4/pe1/q_reg[12]  ( .D(ao3[5]), .CK(clk), .RDN(n28442), .Q(
        \pe4/aot [5]) );
  DRNQHSV4 \pe4/pe1/q_reg[11]  ( .D(ao3[6]), .CK(clk), .RDN(n28446), .Q(
        \pe4/aot [6]) );
  DRNQHSV4 \pe4/pe1/q_reg[10]  ( .D(ao3[7]), .CK(clk), .RDN(n28577), .Q(
        \pe4/aot [7]) );
  DRNQHSV4 \pe4/pe1/q_reg[9]  ( .D(ao3[8]), .CK(clk), .RDN(n28529), .Q(
        \pe4/aot [8]) );
  DRNQHSV4 \pe4/pe1/q_reg[8]  ( .D(ao3[9]), .CK(clk), .RDN(n28495), .Q(
        \pe4/aot [9]) );
  DRNQHSV4 \pe4/pe1/q_reg[7]  ( .D(ao3[10]), .CK(clk), .RDN(n28538), .Q(
        \pe4/aot [10]) );
  DRNQHSV4 \pe4/pe1/q_reg[6]  ( .D(ao3[11]), .CK(clk), .RDN(n28511), .Q(
        \pe4/aot [11]) );
  DRNQHSV4 \pe4/pe1/q_reg[5]  ( .D(ao3[12]), .CK(clk), .RDN(n28529), .Q(
        \pe4/aot [12]) );
  DRNQHSV4 \pe4/pe1/q_reg[4]  ( .D(ao3[13]), .CK(clk), .RDN(n28517), .Q(
        \pe4/aot [13]) );
  DRNQHSV4 \pe4/pe1/q_reg[3]  ( .D(ao3[14]), .CK(clk), .RDN(n28448), .Q(
        \pe4/aot [14]) );
  DRNQHSV4 \pe4/pe1/q_reg[2]  ( .D(ao3[15]), .CK(clk), .RDN(n28606), .Q(
        \pe4/aot [15]) );
  DRNQHSV4 \pe4/pe1/q_reg[1]  ( .D(ao3[16]), .CK(clk), .RDN(n28515), .Q(
        \pe4/aot [16]) );
  DRNQHSV4 \pe4/pe2/q_reg[16]  ( .D(go3[1]), .CK(clk), .RDN(n28561), .Q(
        \pe4/got [1]) );
  DRNQHSV4 \pe4/pe2/q_reg[15]  ( .D(go3[2]), .CK(clk), .RDN(n28443), .Q(
        \pe4/got [2]) );
  DRNQHSV4 \pe4/pe2/q_reg[14]  ( .D(go3[3]), .CK(clk), .RDN(n28538), .Q(
        \pe4/got [3]) );
  DRNQHSV4 \pe4/pe2/q_reg[13]  ( .D(go3[4]), .CK(clk), .RDN(n28441), .Q(
        \pe4/got [4]) );
  DRNQHSV4 \pe4/pe2/q_reg[12]  ( .D(go3[5]), .CK(clk), .RDN(n28489), .Q(
        \pe4/got [5]) );
  DRNQHSV4 \pe4/pe2/q_reg[11]  ( .D(go3[6]), .CK(clk), .RDN(n28522), .Q(
        \pe4/got [6]) );
  DRNQHSV4 \pe4/pe2/q_reg[10]  ( .D(go3[7]), .CK(clk), .RDN(n28489), .Q(
        \pe4/got [7]) );
  DRNQHSV4 \pe4/pe2/q_reg[9]  ( .D(go3[8]), .CK(clk), .RDN(n28488), .Q(
        \pe4/got [8]) );
  DRNQHSV4 \pe4/pe2/q_reg[8]  ( .D(go3[9]), .CK(clk), .RDN(n28539), .Q(
        \pe4/got [9]) );
  DRNQHSV4 \pe4/pe2/q_reg[7]  ( .D(go3[10]), .CK(clk), .RDN(n28561), .Q(
        \pe4/got [10]) );
  DRNQHSV4 \pe4/pe2/q_reg[6]  ( .D(go3[11]), .CK(clk), .RDN(n28444), .Q(
        \pe4/got [11]) );
  DRNQHSV4 \pe4/pe2/q_reg[5]  ( .D(go3[12]), .CK(clk), .RDN(n28573), .Q(
        \pe4/got [12]) );
  DRNQHSV4 \pe4/pe2/q_reg[4]  ( .D(go3[13]), .CK(clk), .RDN(n28507), .Q(
        \pe4/got [13]) );
  DRNQHSV4 \pe4/pe2/q_reg[3]  ( .D(go3[14]), .CK(clk), .RDN(n28447), .Q(
        \pe4/got [14]) );
  DRNQHSV4 \pe4/pe2/q_reg[2]  ( .D(go3[15]), .CK(clk), .RDN(n28509), .Q(
        \pe4/got [15]) );
  DRNQHSV4 \pe4/pe2/q_reg[1]  ( .D(go3[16]), .CK(clk), .RDN(n28487), .Q(
        \pe4/got [16]) );
  DRNQHSV4 \pe4/pe5/q_reg[11]  ( .D(pov3[11]), .CK(clk), .RDN(n28484), .Q(
        \pe4/pvq [11]) );
  DRNQHSV4 \pe4/pe5/q_reg[6]  ( .D(pov3[6]), .CK(clk), .RDN(n28453), .Q(
        \pe4/pvq [6]) );
  DRNQHSV4 \pe4/pe5/q_reg[3]  ( .D(n28981), .CK(clk), .RDN(n28483), .Q(
        \pe4/pvq [3]) );
  DRNQHSV4 \pe4/pe5/q_reg[2]  ( .D(n29038), .CK(clk), .RDN(n28509), .Q(
        \pe4/pvq [2]) );
  DRNQHSV4 \pe4/pe6/q_reg[15]  ( .D(poh3[15]), .CK(clk), .RDN(n28602), .Q(
        \pe4/phq [15]) );
  DRNQHSV4 \pe4/pe6/q_reg[14]  ( .D(poh3[14]), .CK(clk), .RDN(n28486), .Q(
        \pe4/phq [14]) );
  DRNQHSV4 \pe4/pe6/q_reg[12]  ( .D(poh3[12]), .CK(clk), .RDN(n28482), .Q(
        \pe4/phq [12]) );
  DRNQHSV4 \pe4/pe6/q_reg[11]  ( .D(poh3[11]), .CK(clk), .RDN(n28538), .Q(
        \pe4/phq [11]) );
  DRNQHSV4 \pe4/pe6/q_reg[10]  ( .D(poh3[10]), .CK(clk), .RDN(n28519), .Q(
        \pe4/phq [10]) );
  DRNQHSV4 \pe4/pe6/q_reg[9]  ( .D(poh3[9]), .CK(clk), .RDN(n28482), .Q(
        \pe4/phq [9]) );
  DRNQHSV4 \pe4/pe6/q_reg[8]  ( .D(poh3[8]), .CK(clk), .RDN(n28441), .Q(
        \pe4/phq [8]) );
  DRNQHSV4 \pe4/pe6/q_reg[7]  ( .D(poh3[7]), .CK(clk), .RDN(n28544), .Q(
        \pe4/phq [7]) );
  DRNQHSV4 \pe4/pe6/q_reg[6]  ( .D(poh3[6]), .CK(clk), .RDN(n28529), .Q(
        \pe4/phq [6]) );
  DRNQHSV4 \pe4/pe6/q_reg[5]  ( .D(poh3[5]), .CK(clk), .RDN(n28556), .Q(
        \pe4/phq [5]) );
  DRNQHSV4 \pe4/pe6/q_reg[4]  ( .D(poh3[4]), .CK(clk), .RDN(n28459), .Q(
        \pe4/phq [4]) );
  DRNQHSV4 \pe4/pe6/q_reg[3]  ( .D(poh3[3]), .CK(clk), .RDN(n28439), .Q(
        \pe4/phq [3]) );
  DRNQHSV4 \pe4/pe6/q_reg[2]  ( .D(poh3[2]), .CK(clk), .RDN(n28539), .Q(
        \pe4/phq [2]) );
  DRNQHSV4 \pe4/pe6/q_reg[1]  ( .D(poh3[1]), .CK(clk), .RDN(n28441), .Q(
        \pe4/phq [1]) );
  DRNQHSV4 \pe4/pe7/q_reg  ( .D(n28931), .CK(clk), .RDN(n28528), .Q(\pe4/ctrq ) );
  DRNQHSV4 \pe4/pe8/q_reg  ( .D(n28924), .CK(clk), .RDN(n28451), .Q(ctro4) );
  DRNQHSV4 \pe4/pe12/q_reg[16]  ( .D(n28751), .CK(clk), .RDN(n28539), .Q(
        \pe4/bq[1] ) );
  DRNQHSV4 \pe4/pe12/q_reg[15]  ( .D(n28763), .CK(clk), .RDN(n28534), .Q(
        \pe4/bq[2] ) );
  DRNQHSV4 \pe4/pe12/q_reg[14]  ( .D(n28739), .CK(clk), .RDN(n28545), .Q(
        \pe4/bq[3] ) );
  DRNQHSV4 \pe4/pe12/q_reg[13]  ( .D(n28770), .CK(clk), .RDN(n28441), .Q(
        \pe4/bq[4] ) );
  DRNQHSV4 \pe4/pe12/q_reg[12]  ( .D(n28858), .CK(clk), .RDN(n28575), .Q(
        \pe4/bq[5] ) );
  DRNQHSV4 \pe4/pe12/q_reg[11]  ( .D(n28786), .CK(clk), .RDN(n28530), .Q(
        \pe4/bq[6] ) );
  DRNQHSV4 \pe4/pe12/q_reg[10]  ( .D(n28762), .CK(clk), .RDN(n28577), .Q(
        \pe4/bq[7] ) );
  DRNQHSV4 \pe4/pe12/q_reg[9]  ( .D(n28777), .CK(clk), .RDN(n28442), .Q(
        \pe4/bq[8] ) );
  DRNQHSV4 \pe4/pe12/q_reg[8]  ( .D(n28857), .CK(clk), .RDN(n28450), .Q(
        \pe4/bq[9] ) );
  DRNQHSV4 \pe4/pe12/q_reg[7]  ( .D(n28761), .CK(clk), .RDN(n28576), .Q(
        \pe4/bq[10] ) );
  DRNQHSV4 \pe4/pe12/q_reg[6]  ( .D(n28774), .CK(clk), .RDN(n28544), .Q(
        \pe4/bq[11] ) );
  DRNQHSV4 \pe4/pe12/q_reg[5]  ( .D(n28760), .CK(clk), .RDN(n28445), .Q(
        \pe4/bq[12] ) );
  DRNQHSV4 \pe4/pe12/q_reg[4]  ( .D(n28856), .CK(clk), .RDN(n28497), .Q(
        \pe4/bq[13] ) );
  DRNQHSV4 \pe4/pe12/q_reg[3]  ( .D(n28733), .CK(clk), .RDN(n28518), .Q(
        \pe4/bq[14] ) );
  DRNQHSV4 \pe4/pe12/q_reg[2]  ( .D(n28855), .CK(clk), .RDN(n28516), .Q(
        \pe4/bq[15] ) );
  DRNQHSV4 \pe4/pe12/q_reg[1]  ( .D(n28854), .CK(clk), .RDN(n28517), .Q(
        \pe4/bq[16] ) );
  DRNQHSV4 \pe4/pe13/q_reg  ( .D(\pe4/ti_1t ), .CK(clk), .RDN(n28519), .Q(
        \pe4/ti_1 ) );
  DRNQHSV4 \pe5/pe1/q_reg[16]  ( .D(ao4[1]), .CK(clk), .RDN(n28566), .Q(
        \pe5/aot [1]) );
  DRNQHSV4 \pe5/pe1/q_reg[15]  ( .D(ao4[2]), .CK(clk), .RDN(n28565), .Q(
        \pe5/aot [2]) );
  DRNQHSV4 \pe5/pe1/q_reg[14]  ( .D(ao4[3]), .CK(clk), .RDN(n14021), .Q(
        \pe5/aot [3]) );
  DRNQHSV4 \pe5/pe1/q_reg[13]  ( .D(ao4[4]), .CK(clk), .RDN(n28536), .Q(
        \pe5/aot [4]) );
  DRNQHSV4 \pe5/pe1/q_reg[12]  ( .D(ao4[5]), .CK(clk), .RDN(n28500), .Q(
        \pe5/aot [5]) );
  DRNQHSV4 \pe5/pe1/q_reg[11]  ( .D(ao4[6]), .CK(clk), .RDN(n28565), .Q(
        \pe5/aot [6]) );
  DRNQHSV4 \pe5/pe1/q_reg[10]  ( .D(ao4[7]), .CK(clk), .RDN(n28452), .Q(
        \pe5/aot [7]) );
  DRNQHSV4 \pe5/pe1/q_reg[9]  ( .D(ao4[8]), .CK(clk), .RDN(n28499), .Q(
        \pe5/aot [8]) );
  DRNQHSV4 \pe5/pe1/q_reg[8]  ( .D(ao4[9]), .CK(clk), .RDN(n28524), .Q(
        \pe5/aot [9]) );
  DRNQHSV4 \pe5/pe1/q_reg[7]  ( .D(ao4[10]), .CK(clk), .RDN(n28542), .Q(
        \pe5/aot [10]) );
  DRNQHSV4 \pe5/pe1/q_reg[6]  ( .D(ao4[11]), .CK(clk), .RDN(n28553), .Q(
        \pe5/aot [11]) );
  DRNQHSV4 \pe5/pe1/q_reg[5]  ( .D(ao4[12]), .CK(clk), .RDN(n28494), .Q(
        \pe5/aot [12]) );
  DRNQHSV4 \pe5/pe1/q_reg[4]  ( .D(ao4[13]), .CK(clk), .RDN(n28549), .Q(
        \pe5/aot [13]) );
  DRNQHSV4 \pe5/pe1/q_reg[3]  ( .D(ao4[14]), .CK(clk), .RDN(n28549), .Q(
        \pe5/aot [14]) );
  DRNQHSV4 \pe5/pe1/q_reg[2]  ( .D(ao4[15]), .CK(clk), .RDN(n28553), .Q(
        \pe5/aot [15]) );
  DRNQHSV4 \pe5/pe1/q_reg[1]  ( .D(ao4[16]), .CK(clk), .RDN(n28440), .Q(
        \pe5/aot [16]) );
  DRNQHSV4 \pe5/pe2/q_reg[16]  ( .D(go4[1]), .CK(clk), .RDN(n28458), .Q(
        \pe5/got [1]) );
  DRNQHSV4 \pe5/pe2/q_reg[15]  ( .D(go4[2]), .CK(clk), .RDN(n28569), .Q(
        \pe5/got [2]) );
  DRNQHSV4 \pe5/pe2/q_reg[14]  ( .D(go4[3]), .CK(clk), .RDN(n28533), .Q(
        \pe5/got [3]) );
  DRNQHSV4 \pe5/pe2/q_reg[13]  ( .D(go4[4]), .CK(clk), .RDN(n28537), .Q(
        \pe5/got [4]) );
  DRNQHSV4 \pe5/pe2/q_reg[12]  ( .D(go4[5]), .CK(clk), .RDN(n28521), .Q(
        \pe5/got [5]) );
  DRNQHSV4 \pe5/pe2/q_reg[11]  ( .D(go4[6]), .CK(clk), .RDN(n28502), .Q(
        \pe5/got [6]) );
  DRNQHSV4 \pe5/pe2/q_reg[10]  ( .D(go4[7]), .CK(clk), .RDN(n28553), .Q(
        \pe5/got [7]) );
  DRNQHSV4 \pe5/pe2/q_reg[9]  ( .D(go4[8]), .CK(clk), .RDN(n28494), .Q(
        \pe5/got [8]) );
  DRNQHSV4 \pe5/pe2/q_reg[8]  ( .D(go4[9]), .CK(clk), .RDN(n28528), .Q(
        \pe5/got [9]) );
  DRNQHSV4 \pe5/pe2/q_reg[7]  ( .D(go4[10]), .CK(clk), .RDN(n28483), .Q(
        \pe5/got [10]) );
  DRNQHSV4 \pe5/pe2/q_reg[6]  ( .D(go4[11]), .CK(clk), .RDN(n28525), .Q(
        \pe5/got [11]) );
  DRNQHSV4 \pe5/pe2/q_reg[5]  ( .D(go4[12]), .CK(clk), .RDN(n28542), .Q(
        \pe5/got [12]) );
  DRNQHSV4 \pe5/pe2/q_reg[4]  ( .D(go4[13]), .CK(clk), .RDN(n28442), .Q(
        \pe5/got [13]) );
  DRNQHSV4 \pe5/pe2/q_reg[3]  ( .D(go4[14]), .CK(clk), .RDN(n28605), .Q(
        \pe5/got [14]) );
  DRNQHSV4 \pe5/pe2/q_reg[2]  ( .D(go4[15]), .CK(clk), .RDN(n28525), .Q(
        \pe5/got [15]) );
  DRNQHSV4 \pe5/pe2/q_reg[1]  ( .D(go4[16]), .CK(clk), .RDN(n28490), .Q(
        \pe5/got [16]) );
  DRNQHSV4 \pe5/pe5/q_reg[11]  ( .D(n29029), .CK(clk), .RDN(n14021), .Q(
        \pe5/pvq [11]) );
  DRNQHSV4 \pe5/pe5/q_reg[10]  ( .D(pov4[10]), .CK(clk), .RDN(n28551), .Q(
        \pe5/pvq [10]) );
  DRNQHSV4 \pe5/pe5/q_reg[9]  ( .D(n29030), .CK(clk), .RDN(n28448), .Q(
        \pe5/pvq [9]) );
  DRNQHSV4 \pe5/pe5/q_reg[5]  ( .D(n29032), .CK(clk), .RDN(n28529), .Q(
        \pe5/pvq [5]) );
  DRNQHSV4 \pe5/pe5/q_reg[2]  ( .D(n29034), .CK(clk), .RDN(n28571), .Q(
        \pe5/pvq [2]) );
  DRNQHSV4 \pe5/pe6/q_reg[15]  ( .D(poh4[15]), .CK(clk), .RDN(n28483), .Q(
        \pe5/phq [15]) );
  DRNQHSV4 \pe5/pe6/q_reg[14]  ( .D(poh4[14]), .CK(clk), .RDN(n28533), .Q(
        \pe5/phq [14]) );
  DRNQHSV4 \pe5/pe6/q_reg[13]  ( .D(poh4[13]), .CK(clk), .RDN(n28497), .Q(
        \pe5/phq [13]) );
  DRNQHSV4 \pe5/pe6/q_reg[12]  ( .D(poh4[12]), .CK(clk), .RDN(n28476), .Q(
        \pe5/phq [12]) );
  DRNQHSV4 \pe5/pe6/q_reg[11]  ( .D(poh4[11]), .CK(clk), .RDN(n28446), .Q(
        \pe5/phq [11]) );
  DRNQHSV4 \pe5/pe6/q_reg[10]  ( .D(poh4[10]), .CK(clk), .RDN(n28440), .Q(
        \pe5/phq [10]) );
  DRNQHSV4 \pe5/pe6/q_reg[9]  ( .D(poh4[9]), .CK(clk), .RDN(n28555), .Q(
        \pe5/phq [9]) );
  DRNQHSV4 \pe5/pe6/q_reg[8]  ( .D(poh4[8]), .CK(clk), .RDN(n28494), .Q(
        \pe5/phq [8]) );
  DRNQHSV4 \pe5/pe6/q_reg[7]  ( .D(poh4[7]), .CK(clk), .RDN(n28527), .Q(
        \pe5/phq [7]) );
  DRNQHSV4 \pe5/pe6/q_reg[6]  ( .D(poh4[6]), .CK(clk), .RDN(n28516), .Q(
        \pe5/phq [6]) );
  DRNQHSV4 \pe5/pe6/q_reg[5]  ( .D(poh4[5]), .CK(clk), .RDN(n28505), .Q(
        \pe5/phq [5]) );
  DRNQHSV4 \pe5/pe6/q_reg[4]  ( .D(poh4[4]), .CK(clk), .RDN(n28504), .Q(
        \pe5/phq [4]) );
  DRNQHSV4 \pe5/pe6/q_reg[3]  ( .D(poh4[3]), .CK(clk), .RDN(n14021), .Q(
        \pe5/phq [3]) );
  DRNQHSV4 \pe5/pe6/q_reg[2]  ( .D(poh4[2]), .CK(clk), .RDN(n28483), .Q(
        \pe5/phq [2]) );
  DRNQHSV4 \pe5/pe6/q_reg[1]  ( .D(poh4[1]), .CK(clk), .RDN(n28443), .Q(
        \pe5/phq [1]) );
  DRNQHSV4 \pe5/pe7/q_reg  ( .D(n28812), .CK(clk), .RDN(n28447), .Q(\pe5/ctrq ) );
  DRNQHSV4 \pe5/pe12/q_reg[16]  ( .D(n28866), .CK(clk), .RDN(n28555), .Q(
        \pe5/bq[1] ) );
  DRNQHSV4 \pe5/pe12/q_reg[15]  ( .D(n28716), .CK(clk), .RDN(n28542), .Q(
        \pe5/bq[2] ) );
  DRNQHSV4 \pe5/pe12/q_reg[14]  ( .D(n28715), .CK(clk), .RDN(n28533), .Q(
        \pe5/bq[3] ) );
  DRNQHSV4 \pe5/pe12/q_reg[13]  ( .D(n28865), .CK(clk), .RDN(n28476), .Q(
        \pe5/bq[4] ) );
  DRNQHSV4 \pe5/pe12/q_reg[12]  ( .D(n28864), .CK(clk), .RDN(n28541), .Q(
        \pe5/bq[5] ) );
  DRNQHSV4 \pe5/pe12/q_reg[11]  ( .D(n28714), .CK(clk), .RDN(n28542), .Q(
        \pe5/bq[6] ) );
  DRNQHSV4 \pe5/pe12/q_reg[10]  ( .D(n28863), .CK(clk), .RDN(n28527), .Q(
        \pe5/bq[7] ) );
  DRNQHSV4 \pe5/pe12/q_reg[9]  ( .D(n28862), .CK(clk), .RDN(n28504), .Q(
        \pe5/bq[8] ) );
  DRNQHSV4 \pe5/pe12/q_reg[8]  ( .D(n28713), .CK(clk), .RDN(n28563), .Q(
        \pe5/bq[9] ) );
  DRNQHSV4 \pe5/pe12/q_reg[7]  ( .D(n28712), .CK(clk), .RDN(n28499), .Q(
        \pe5/bq[10] ) );
  DRNQHSV4 \pe5/pe12/q_reg[6]  ( .D(n28711), .CK(clk), .RDN(n28607), .Q(
        \pe5/bq[11] ) );
  DRNQHSV4 \pe5/pe12/q_reg[5]  ( .D(n28861), .CK(clk), .RDN(n28527), .Q(
        \pe5/bq[12] ) );
  DRNQHSV4 \pe5/pe12/q_reg[4]  ( .D(n28710), .CK(clk), .RDN(n28498), .Q(
        \pe5/bq[13] ) );
  DRNQHSV4 \pe5/pe12/q_reg[3]  ( .D(n28859), .CK(clk), .RDN(n28520), .Q(
        \pe5/bq[14] ) );
  DRNQHSV4 \pe5/pe12/q_reg[2]  ( .D(n28860), .CK(clk), .RDN(n28441), .Q(
        \pe5/bq[15] ) );
  DRNQHSV4 \pe5/pe12/q_reg[1]  ( .D(n28709), .CK(clk), .RDN(n28444), .Q(
        \pe5/bq[16] ) );
  DRNQHSV4 \pe5/pe13/q_reg  ( .D(\pe5/ti_1t ), .CK(clk), .RDN(n28499), .Q(
        \pe5/ti_1 ) );
  DRNQHSV4 \pe5/pe14/q_reg[5]  ( .D(n28955), .CK(clk), .RDN(n28569), .Q(
        \pe5/ti_7t [5]) );
  DRNQHSV4 \pe6/pe1/q_reg[16]  ( .D(ao5[1]), .CK(clk), .RDN(n28595), .Q(
        \pe6/aot [1]) );
  DRNQHSV4 \pe6/pe1/q_reg[15]  ( .D(ao5[2]), .CK(clk), .RDN(n28453), .Q(
        \pe6/aot [2]) );
  DRNQHSV4 \pe6/pe1/q_reg[14]  ( .D(ao5[3]), .CK(clk), .RDN(n28570), .Q(
        \pe6/aot [3]) );
  DRNQHSV4 \pe6/pe1/q_reg[13]  ( .D(ao5[4]), .CK(clk), .RDN(n28550), .Q(
        \pe6/aot [4]) );
  DRNQHSV4 \pe6/pe1/q_reg[12]  ( .D(ao5[5]), .CK(clk), .RDN(n28506), .Q(
        \pe6/aot [5]) );
  DRNQHSV4 \pe6/pe1/q_reg[11]  ( .D(ao5[6]), .CK(clk), .RDN(n28513), .Q(
        \pe6/aot [6]) );
  DRNQHSV4 \pe6/pe1/q_reg[10]  ( .D(ao5[7]), .CK(clk), .RDN(n28531), .Q(
        \pe6/aot [7]) );
  DRNQHSV4 \pe6/pe1/q_reg[9]  ( .D(ao5[8]), .CK(clk), .RDN(n28535), .Q(
        \pe6/aot [8]) );
  DRNQHSV4 \pe6/pe1/q_reg[8]  ( .D(ao5[9]), .CK(clk), .RDN(n28564), .Q(
        \pe6/aot [9]) );
  DRNQHSV4 \pe6/pe1/q_reg[7]  ( .D(ao5[10]), .CK(clk), .RDN(n28450), .Q(
        \pe6/aot [10]) );
  DRNQHSV4 \pe6/pe1/q_reg[6]  ( .D(ao5[11]), .CK(clk), .RDN(n28606), .Q(
        \pe6/aot [11]) );
  DRNQHSV4 \pe6/pe1/q_reg[5]  ( .D(ao5[12]), .CK(clk), .RDN(n28571), .Q(
        \pe6/aot [12]) );
  DRNQHSV4 \pe6/pe1/q_reg[4]  ( .D(ao5[13]), .CK(clk), .RDN(n28450), .Q(
        \pe6/aot [13]) );
  DRNQHSV4 \pe6/pe1/q_reg[3]  ( .D(ao5[14]), .CK(clk), .RDN(n28566), .Q(
        \pe6/aot [14]) );
  DRNQHSV4 \pe6/pe1/q_reg[2]  ( .D(ao5[15]), .CK(clk), .RDN(n28529), .Q(
        \pe6/aot [15]) );
  DRNQHSV4 \pe6/pe1/q_reg[1]  ( .D(ao5[16]), .CK(clk), .RDN(n28517), .Q(
        \pe6/aot [16]) );
  DRNQHSV4 \pe6/pe2/q_reg[16]  ( .D(go5[1]), .CK(clk), .RDN(n28595), .Q(
        \pe6/got [1]) );
  DRNQHSV4 \pe6/pe2/q_reg[15]  ( .D(go5[2]), .CK(clk), .RDN(n28501), .Q(
        \pe6/got [2]) );
  DRNQHSV4 \pe6/pe2/q_reg[14]  ( .D(go5[3]), .CK(clk), .RDN(n28444), .Q(
        \pe6/got [3]) );
  DRNQHSV4 \pe6/pe2/q_reg[13]  ( .D(go5[4]), .CK(clk), .RDN(n28496), .Q(
        \pe6/got [4]) );
  DRNQHSV4 \pe6/pe2/q_reg[12]  ( .D(go5[5]), .CK(clk), .RDN(n28508), .Q(
        \pe6/got [5]) );
  DRNQHSV4 \pe6/pe2/q_reg[11]  ( .D(go5[6]), .CK(clk), .RDN(n28596), .Q(
        \pe6/got [6]) );
  DRNQHSV4 \pe6/pe2/q_reg[10]  ( .D(go5[7]), .CK(clk), .RDN(n28496), .Q(
        \pe6/got [7]) );
  DRNQHSV4 \pe6/pe2/q_reg[9]  ( .D(go5[8]), .CK(clk), .RDN(n28440), .Q(
        \pe6/got [8]) );
  DRNQHSV4 \pe6/pe2/q_reg[8]  ( .D(go5[9]), .CK(clk), .RDN(n28565), .Q(
        \pe6/got [9]) );
  DRNQHSV4 \pe6/pe2/q_reg[7]  ( .D(go5[10]), .CK(clk), .RDN(n28569), .Q(
        \pe6/got [10]) );
  DRNQHSV4 \pe6/pe2/q_reg[6]  ( .D(go5[11]), .CK(clk), .RDN(n28499), .Q(
        \pe6/got [11]) );
  DRNQHSV4 \pe6/pe2/q_reg[5]  ( .D(go5[12]), .CK(clk), .RDN(n28550), .Q(
        \pe6/got [12]) );
  DRNQHSV4 \pe6/pe2/q_reg[4]  ( .D(go5[13]), .CK(clk), .RDN(n28562), .Q(
        \pe6/got [13]) );
  DRNQHSV4 \pe6/pe2/q_reg[3]  ( .D(go5[14]), .CK(clk), .RDN(n28531), .Q(
        \pe6/got [14]) );
  DRNQHSV4 \pe6/pe2/q_reg[2]  ( .D(go5[15]), .CK(clk), .RDN(n28506), .Q(
        \pe6/got [15]) );
  DRNQHSV4 \pe6/pe2/q_reg[1]  ( .D(go5[16]), .CK(clk), .RDN(n28492), .Q(
        \pe6/got [16]) );
  DRNQHSV4 \pe6/pe5/q_reg[7]  ( .D(n29025), .CK(clk), .RDN(n28607), .Q(
        \pe6/pvq [7]) );
  DRNQHSV4 \pe6/pe5/q_reg[4]  ( .D(n28992), .CK(clk), .RDN(n28558), .Q(
        \pe6/pvq [4]) );
  DRNQHSV4 \pe6/pe5/q_reg[3]  ( .D(n29026), .CK(clk), .RDN(n28540), .Q(
        \pe6/pvq [3]) );
  DRNQHSV4 \pe6/pe5/q_reg[2]  ( .D(n29027), .CK(clk), .RDN(n28564), .Q(
        \pe6/pvq [2]) );
  DRNQHSV4 \pe6/pe6/q_reg[15]  ( .D(poh5[15]), .CK(clk), .RDN(n28537), .Q(
        \pe6/phq [15]) );
  DRNQHSV4 \pe6/pe6/q_reg[14]  ( .D(poh5[14]), .CK(clk), .RDN(n28505), .Q(
        \pe6/phq [14]) );
  DRNQHSV4 \pe6/pe6/q_reg[13]  ( .D(poh5[13]), .CK(clk), .RDN(n28520), .Q(
        \pe6/phq [13]) );
  DRNQHSV4 \pe6/pe6/q_reg[12]  ( .D(poh5[12]), .CK(clk), .RDN(n28519), .Q(
        \pe6/phq [12]) );
  DRNQHSV4 \pe6/pe6/q_reg[11]  ( .D(poh5[11]), .CK(clk), .RDN(n28553), .Q(
        \pe6/phq [11]) );
  DRNQHSV4 \pe6/pe6/q_reg[10]  ( .D(poh5[10]), .CK(clk), .RDN(n28495), .Q(
        \pe6/phq [10]) );
  DRNQHSV4 \pe6/pe6/q_reg[9]  ( .D(poh5[9]), .CK(clk), .RDN(n28558), .Q(
        \pe6/phq [9]) );
  DRNQHSV4 \pe6/pe6/q_reg[8]  ( .D(poh5[8]), .CK(clk), .RDN(n28524), .Q(
        \pe6/phq [8]) );
  DRNQHSV4 \pe6/pe6/q_reg[7]  ( .D(poh5[7]), .CK(clk), .RDN(n28509), .Q(
        \pe6/phq [7]) );
  DRNQHSV4 \pe6/pe6/q_reg[6]  ( .D(poh5[6]), .CK(clk), .RDN(n28494), .Q(
        \pe6/phq [6]) );
  DRNQHSV4 \pe6/pe6/q_reg[5]  ( .D(poh5[5]), .CK(clk), .RDN(n28496), .Q(
        \pe6/phq [5]) );
  DRNQHSV4 \pe6/pe6/q_reg[4]  ( .D(poh5[4]), .CK(clk), .RDN(n28566), .Q(
        \pe6/phq [4]) );
  DRNQHSV4 \pe6/pe6/q_reg[3]  ( .D(poh5[3]), .CK(clk), .RDN(n28484), .Q(
        \pe6/phq [3]) );
  DRNQHSV4 \pe6/pe6/q_reg[2]  ( .D(poh5[2]), .CK(clk), .RDN(n28444), .Q(
        \pe6/phq [2]) );
  DRNQHSV4 \pe6/pe6/q_reg[1]  ( .D(poh5[1]), .CK(clk), .RDN(n28522), .Q(
        \pe6/phq [1]) );
  DRNQHSV4 \pe6/pe7/q_reg  ( .D(n21345), .CK(clk), .RDN(n28569), .Q(\pe6/ctrq ) );
  DRNQHSV4 \pe6/pe8/q_reg  ( .D(n28867), .CK(clk), .RDN(n28476), .Q(ctro6) );
  DRNQHSV4 \pe6/pe12/q_reg[16]  ( .D(n28773), .CK(clk), .RDN(n28545), .Q(
        \pe6/bq[1] ) );
  DRNQHSV4 \pe6/pe12/q_reg[15]  ( .D(n28783), .CK(clk), .RDN(n28476), .Q(
        \pe6/bq[2] ) );
  DRNQHSV4 \pe6/pe12/q_reg[14]  ( .D(n28750), .CK(clk), .RDN(n28447), .Q(
        \pe6/bq[3] ) );
  DRNQHSV4 \pe6/pe12/q_reg[13]  ( .D(n28875), .CK(clk), .RDN(n28477), .Q(
        \pe6/bq[4] ) );
  DRNQHSV4 \pe6/pe12/q_reg[12]  ( .D(n28747), .CK(clk), .RDN(n14021), .Q(
        \pe6/bq[5] ) );
  DRNQHSV4 \pe6/pe12/q_reg[11]  ( .D(n28749), .CK(clk), .RDN(n28490), .Q(
        \pe6/bq[6] ) );
  DRNQHSV4 \pe6/pe12/q_reg[10]  ( .D(n28746), .CK(clk), .RDN(n28491), .Q(
        \pe6/bq[7] ) );
  DRNQHSV4 \pe6/pe12/q_reg[9]  ( .D(n28748), .CK(clk), .RDN(n28447), .Q(
        \pe6/bq[8] ) );
  DRNQHSV4 \pe6/pe12/q_reg[8]  ( .D(n28874), .CK(clk), .RDN(n28519), .Q(
        \pe6/bq[9] ) );
  DRNQHSV4 \pe6/pe12/q_reg[7]  ( .D(n28873), .CK(clk), .RDN(n28548), .Q(
        \pe6/bq[10] ) );
  DRNQHSV4 \pe6/pe12/q_reg[6]  ( .D(n28872), .CK(clk), .RDN(n28491), .Q(
        \pe6/bq[11] ) );
  DRNQHSV4 \pe6/pe12/q_reg[5]  ( .D(n28871), .CK(clk), .RDN(n28556), .Q(
        \pe6/bq[12] ) );
  DRNQHSV4 \pe6/pe12/q_reg[4]  ( .D(n28870), .CK(clk), .RDN(n28557), .Q(
        \pe6/bq[13] ) );
  DRNQHSV4 \pe6/pe12/q_reg[3]  ( .D(n28869), .CK(clk), .RDN(n28565), .Q(
        \pe6/bq[14] ) );
  DRNQHSV4 \pe6/pe12/q_reg[2]  ( .D(n28868), .CK(clk), .RDN(n28540), .Q(
        \pe6/bq[15] ) );
  DRNQHSV4 \pe6/pe12/q_reg[1]  ( .D(n28732), .CK(clk), .RDN(n28513), .Q(
        \pe6/bq[16] ) );
  DRNQHSV4 \pe6/pe13/q_reg  ( .D(\pe6/ti_1t ), .CK(clk), .RDN(n28563), .Q(
        \pe6/ti_1 ) );
  DRNQHSV4 \pe6/pe14/q_reg[5]  ( .D(n26034), .CK(clk), .RDN(n28490), .Q(
        \pe6/ti_7t [5]) );
  DRNQHSV4 \pe7/pe1/q_reg[16]  ( .D(ao6[1]), .CK(clk), .RDN(n28554), .Q(
        \pe7/aot [1]) );
  DRNQHSV4 \pe7/pe1/q_reg[15]  ( .D(ao6[2]), .CK(clk), .RDN(n28559), .Q(
        \pe7/aot [2]) );
  DRNQHSV4 \pe7/pe1/q_reg[14]  ( .D(ao6[3]), .CK(clk), .RDN(n28557), .Q(
        \pe7/aot [3]) );
  DRNQHSV4 \pe7/pe1/q_reg[13]  ( .D(ao6[4]), .CK(clk), .RDN(n28450), .Q(
        \pe7/aot [4]) );
  DRNQHSV4 \pe7/pe1/q_reg[12]  ( .D(ao6[5]), .CK(clk), .RDN(n28495), .Q(
        \pe7/aot [5]) );
  DRNQHSV4 \pe7/pe1/q_reg[11]  ( .D(ao6[6]), .CK(clk), .RDN(n28556), .Q(
        \pe7/aot [6]) );
  DRNQHSV4 \pe7/pe1/q_reg[10]  ( .D(ao6[7]), .CK(clk), .RDN(n28555), .Q(
        \pe7/aot [7]) );
  DRNQHSV4 \pe7/pe1/q_reg[9]  ( .D(ao6[8]), .CK(clk), .RDN(n28559), .Q(
        \pe7/aot [8]) );
  DRNQHSV4 \pe7/pe1/q_reg[8]  ( .D(ao6[9]), .CK(clk), .RDN(n28605), .Q(
        \pe7/aot [9]) );
  DRNQHSV4 \pe7/pe1/q_reg[7]  ( .D(ao6[10]), .CK(clk), .RDN(n28482), .Q(
        \pe7/aot [10]) );
  DRNQHSV4 \pe7/pe1/q_reg[6]  ( .D(ao6[11]), .CK(clk), .RDN(n28597), .Q(
        \pe7/aot [11]) );
  DRNQHSV4 \pe7/pe1/q_reg[5]  ( .D(ao6[12]), .CK(clk), .RDN(n28557), .Q(
        \pe7/aot [12]) );
  DRNQHSV4 \pe7/pe1/q_reg[4]  ( .D(ao6[13]), .CK(clk), .RDN(n28554), .Q(
        \pe7/aot [13]) );
  DRNQHSV4 \pe7/pe1/q_reg[3]  ( .D(ao6[14]), .CK(clk), .RDN(n28556), .Q(
        \pe7/aot [14]) );
  DRNQHSV4 \pe7/pe1/q_reg[2]  ( .D(ao6[15]), .CK(clk), .RDN(n28448), .Q(
        \pe7/aot [15]) );
  DRNQHSV4 \pe7/pe1/q_reg[1]  ( .D(ao6[16]), .CK(clk), .RDN(n28447), .Q(
        \pe7/aot [16]) );
  DRNQHSV4 \pe7/pe2/q_reg[16]  ( .D(go6[1]), .CK(clk), .RDN(n28560), .Q(
        \pe7/got [1]) );
  DRNQHSV4 \pe7/pe2/q_reg[15]  ( .D(go6[2]), .CK(clk), .RDN(n28530), .Q(
        \pe7/got [2]) );
  DRNQHSV4 \pe7/pe2/q_reg[14]  ( .D(go6[3]), .CK(clk), .RDN(n28605), .Q(
        \pe7/got [3]) );
  DRNQHSV4 \pe7/pe2/q_reg[13]  ( .D(go6[4]), .CK(clk), .RDN(n28577), .Q(
        \pe7/got [4]) );
  DRNQHSV4 \pe7/pe2/q_reg[12]  ( .D(go6[5]), .CK(clk), .RDN(n28606), .Q(
        \pe7/got [5]) );
  DRNQHSV4 \pe7/pe2/q_reg[11]  ( .D(go6[6]), .CK(clk), .RDN(n28532), .Q(
        \pe7/got [6]) );
  DRNQHSV4 \pe7/pe2/q_reg[10]  ( .D(go6[7]), .CK(clk), .RDN(n28570), .Q(
        \pe7/got [7]) );
  DRNQHSV4 \pe7/pe2/q_reg[9]  ( .D(go6[8]), .CK(clk), .RDN(n28530), .Q(
        \pe7/got [8]) );
  DRNQHSV4 \pe7/pe2/q_reg[8]  ( .D(go6[9]), .CK(clk), .RDN(n28552), .Q(
        \pe7/got [9]) );
  DRNQHSV4 \pe7/pe2/q_reg[7]  ( .D(go6[10]), .CK(clk), .RDN(n28543), .Q(
        \pe7/got [10]) );
  DRNQHSV4 \pe7/pe2/q_reg[6]  ( .D(go6[11]), .CK(clk), .RDN(n28595), .Q(
        \pe7/got [11]) );
  DRNQHSV4 \pe7/pe2/q_reg[5]  ( .D(go6[12]), .CK(clk), .RDN(n28512), .Q(
        \pe7/got [12]) );
  DRNQHSV4 \pe7/pe2/q_reg[4]  ( .D(go6[13]), .CK(clk), .RDN(n28551), .Q(
        \pe7/got [13]) );
  DRNQHSV4 \pe7/pe2/q_reg[3]  ( .D(go6[14]), .CK(clk), .RDN(n28542), .Q(
        \pe7/got [14]) );
  DRNQHSV4 \pe7/pe2/q_reg[2]  ( .D(go6[15]), .CK(clk), .RDN(n28448), .Q(
        \pe7/got [15]) );
  DRNQHSV4 \pe7/pe2/q_reg[1]  ( .D(go6[16]), .CK(clk), .RDN(n28537), .Q(
        \pe7/got [16]) );
  DRNQHSV4 \pe7/pe5/q_reg[9]  ( .D(n29022), .CK(clk), .RDN(n28448), .Q(
        \pe7/pvq [9]) );
  DRNQHSV4 \pe7/pe5/q_reg[4]  ( .D(n28991), .CK(clk), .RDN(n28541), .Q(
        \pe7/pvq [4]) );
  DRNQHSV4 \pe7/pe5/q_reg[3]  ( .D(n28993), .CK(clk), .RDN(n28561), .Q(
        \pe7/pvq [3]) );
  DRNQHSV4 \pe7/pe5/q_reg[2]  ( .D(n29024), .CK(clk), .RDN(n28528), .Q(
        \pe7/pvq [2]) );
  DRNQHSV4 \pe7/pe6/q_reg[15]  ( .D(poh6[15]), .CK(clk), .RDN(n28452), .Q(
        \pe7/phq [15]) );
  DRNQHSV4 \pe7/pe6/q_reg[14]  ( .D(poh6[14]), .CK(clk), .RDN(n28576), .Q(
        \pe7/phq [14]) );
  DRNQHSV4 \pe7/pe6/q_reg[13]  ( .D(poh6[13]), .CK(clk), .RDN(n28530), .Q(
        \pe7/phq [13]) );
  DRNQHSV4 \pe7/pe6/q_reg[12]  ( .D(poh6[12]), .CK(clk), .RDN(n28507), .Q(
        \pe7/phq [12]) );
  DRNQHSV4 \pe7/pe6/q_reg[11]  ( .D(poh6[11]), .CK(clk), .RDN(n28602), .Q(
        \pe7/phq [11]) );
  DRNQHSV4 \pe7/pe6/q_reg[10]  ( .D(poh6[10]), .CK(clk), .RDN(n28490), .Q(
        \pe7/phq [10]) );
  DRNQHSV4 \pe7/pe6/q_reg[9]  ( .D(poh6[9]), .CK(clk), .RDN(n28538), .Q(
        \pe7/phq [9]) );
  DRNQHSV4 \pe7/pe6/q_reg[8]  ( .D(poh6[8]), .CK(clk), .RDN(n28451), .Q(
        \pe7/phq [8]) );
  DRNQHSV4 \pe7/pe6/q_reg[7]  ( .D(poh6[7]), .CK(clk), .RDN(n28508), .Q(
        \pe7/phq [7]) );
  DRNQHSV4 \pe7/pe6/q_reg[6]  ( .D(poh6[6]), .CK(clk), .RDN(n28533), .Q(
        \pe7/phq [6]) );
  DRNQHSV4 \pe7/pe6/q_reg[5]  ( .D(poh6[5]), .CK(clk), .RDN(n28561), .Q(
        \pe7/phq [5]) );
  DRNQHSV4 \pe7/pe6/q_reg[4]  ( .D(poh6[4]), .CK(clk), .RDN(n28443), .Q(
        \pe7/phq [4]) );
  DRNQHSV4 \pe7/pe6/q_reg[3]  ( .D(poh6[3]), .CK(clk), .RDN(n28537), .Q(
        \pe7/phq [3]) );
  DRNQHSV4 \pe7/pe6/q_reg[2]  ( .D(poh6[2]), .CK(clk), .RDN(n28552), .Q(
        \pe7/phq [2]) );
  DRNQHSV4 \pe7/pe6/q_reg[1]  ( .D(poh6[1]), .CK(clk), .RDN(n28540), .Q(
        \pe7/phq [1]) );
  DRNQHSV4 \pe7/pe7/q_reg  ( .D(n19068), .CK(clk), .RDN(n28532), .Q(\pe7/ctrq ) );
  DRNQHSV4 \pe7/pe12/q_reg[16]  ( .D(n28772), .CK(clk), .RDN(n28506), .Q(
        \pe7/bq[1] ) );
  DRNQHSV4 \pe7/pe12/q_reg[15]  ( .D(n28759), .CK(clk), .RDN(n28445), .Q(
        \pe7/bq[2] ) );
  DRNQHSV4 \pe7/pe12/q_reg[14]  ( .D(n28776), .CK(clk), .RDN(n28605), .Q(
        \pe7/bq[3] ) );
  DRNQHSV4 \pe7/pe12/q_reg[13]  ( .D(n28785), .CK(clk), .RDN(n14023), .Q(
        \pe7/bq[4] ) );
  DRNQHSV4 \pe7/pe12/q_reg[12]  ( .D(n28775), .CK(clk), .RDN(n28498), .Q(
        \pe7/bq[5] ) );
  DRNQHSV4 \pe7/pe12/q_reg[11]  ( .D(n28880), .CK(clk), .RDN(n28540), .Q(
        \pe7/bq[6] ) );
  DRNQHSV4 \pe7/pe12/q_reg[10]  ( .D(n28758), .CK(clk), .RDN(n28486), .Q(
        \pe7/bq[7] ) );
  DRNQHSV4 \pe7/pe12/q_reg[9]  ( .D(n28878), .CK(clk), .RDN(n28530), .Q(
        \pe7/bq[8] ) );
  DRNQHSV4 \pe7/pe12/q_reg[8]  ( .D(n28879), .CK(clk), .RDN(n28528), .Q(
        \pe7/bq[9] ) );
  DRNQHSV4 \pe7/pe12/q_reg[7]  ( .D(n28769), .CK(clk), .RDN(n28561), .Q(
        \pe7/bq[10] ) );
  DRNQHSV4 \pe7/pe12/q_reg[6]  ( .D(n28757), .CK(clk), .RDN(n28538), .Q(
        \pe7/bq[11] ) );
  DRNQHSV4 \pe7/pe12/q_reg[5]  ( .D(n28877), .CK(clk), .RDN(n28604), .Q(
        \pe7/bq[12] ) );
  DRNQHSV4 \pe7/pe12/q_reg[4]  ( .D(n28784), .CK(clk), .RDN(n28489), .Q(
        \pe7/bq[13] ) );
  DRNQHSV4 \pe7/pe12/q_reg[3]  ( .D(n28782), .CK(clk), .RDN(n28567), .Q(
        \pe7/bq[14] ) );
  DRNQHSV4 \pe7/pe12/q_reg[2]  ( .D(n28756), .CK(clk), .RDN(n28545), .Q(
        \pe7/bq[15] ) );
  DRNQHSV4 \pe7/pe12/q_reg[1]  ( .D(n28768), .CK(clk), .RDN(n28604), .Q(
        \pe7/bq[16] ) );
  DRNQHSV4 \pe7/pe13/q_reg  ( .D(\pe7/ti_1t ), .CK(clk), .RDN(n28453), .Q(
        \pe7/ti_1 ) );
  DRNQHSV4 \pe8/pe1/q_reg[16]  ( .D(ao7[1]), .CK(clk), .RDN(n28451), .Q(
        \pe8/aot [1]) );
  DRNQHSV4 \pe8/pe1/q_reg[15]  ( .D(ao7[2]), .CK(clk), .RDN(n28604), .Q(
        \pe8/aot [2]) );
  DRNQHSV4 \pe8/pe1/q_reg[14]  ( .D(ao7[3]), .CK(clk), .RDN(n28522), .Q(
        \pe8/aot [3]) );
  DRNQHSV4 \pe8/pe1/q_reg[13]  ( .D(ao7[4]), .CK(clk), .RDN(n28531), .Q(
        \pe8/aot [4]) );
  DRNQHSV4 \pe8/pe1/q_reg[12]  ( .D(ao7[5]), .CK(clk), .RDN(n28596), .Q(
        \pe8/aot [5]) );
  DRNQHSV4 \pe8/pe1/q_reg[11]  ( .D(ao7[6]), .CK(clk), .RDN(n28567), .Q(
        \pe8/aot [6]) );
  DRNQHSV4 \pe8/pe1/q_reg[10]  ( .D(ao7[7]), .CK(clk), .RDN(n28501), .Q(
        \pe8/aot [7]) );
  DRNQHSV4 \pe8/pe1/q_reg[9]  ( .D(ao7[8]), .CK(clk), .RDN(n28595), .Q(
        \pe8/aot [8]) );
  DRNQHSV4 \pe8/pe1/q_reg[8]  ( .D(ao7[9]), .CK(clk), .RDN(n28498), .Q(
        \pe8/aot [9]) );
  DRNQHSV4 \pe8/pe1/q_reg[7]  ( .D(ao7[10]), .CK(clk), .RDN(n28514), .Q(
        \pe8/aot [10]) );
  DRNQHSV4 \pe8/pe1/q_reg[6]  ( .D(ao7[11]), .CK(clk), .RDN(n28549), .Q(
        \pe8/aot [11]) );
  DRNQHSV4 \pe8/pe1/q_reg[5]  ( .D(ao7[12]), .CK(clk), .RDN(n28566), .Q(
        \pe8/aot [12]) );
  DRNQHSV4 \pe8/pe1/q_reg[4]  ( .D(ao7[13]), .CK(clk), .RDN(n28573), .Q(
        \pe8/aot [13]) );
  DRNQHSV4 \pe8/pe1/q_reg[3]  ( .D(ao7[14]), .CK(clk), .RDN(n28596), .Q(
        \pe8/aot [14]) );
  DRNQHSV4 \pe8/pe1/q_reg[2]  ( .D(ao7[15]), .CK(clk), .RDN(n28452), .Q(
        \pe8/aot [15]) );
  DRNQHSV4 \pe8/pe1/q_reg[1]  ( .D(ao7[16]), .CK(clk), .RDN(n28514), .Q(
        \pe8/aot [16]) );
  DRNQHSV4 \pe8/pe2/q_reg[16]  ( .D(go7[1]), .CK(clk), .RDN(n28514), .Q(
        \pe8/got [1]) );
  DRNQHSV4 \pe8/pe2/q_reg[15]  ( .D(go7[2]), .CK(clk), .RDN(n28449), .Q(
        \pe8/got [2]) );
  DRNQHSV4 \pe8/pe2/q_reg[14]  ( .D(go7[3]), .CK(clk), .RDN(n28496), .Q(
        \pe8/got [3]) );
  DRNQHSV4 \pe8/pe2/q_reg[13]  ( .D(go7[4]), .CK(clk), .RDN(n28496), .Q(
        \pe8/got [4]) );
  DRNQHSV4 \pe8/pe2/q_reg[12]  ( .D(go7[5]), .CK(clk), .RDN(n28522), .Q(
        \pe8/got [5]) );
  DRNQHSV4 \pe8/pe2/q_reg[11]  ( .D(go7[6]), .CK(clk), .RDN(n28566), .Q(
        \pe8/got [6]) );
  DRNQHSV4 \pe8/pe2/q_reg[10]  ( .D(go7[7]), .CK(clk), .RDN(n28439), .Q(
        \pe8/got [7]) );
  DRNQHSV4 \pe8/pe2/q_reg[9]  ( .D(go7[8]), .CK(clk), .RDN(n28512), .Q(
        \pe8/got [8]) );
  DRNQHSV4 \pe8/pe2/q_reg[8]  ( .D(go7[9]), .CK(clk), .RDN(n28514), .Q(
        \pe8/got [9]) );
  DRNQHSV4 \pe8/pe2/q_reg[7]  ( .D(go7[10]), .CK(clk), .RDN(n28529), .Q(
        \pe8/got [10]) );
  DRNQHSV4 \pe8/pe2/q_reg[6]  ( .D(go7[11]), .CK(clk), .RDN(n28512), .Q(
        \pe8/got [11]) );
  DRNQHSV4 \pe8/pe2/q_reg[5]  ( .D(go7[12]), .CK(clk), .RDN(n28450), .Q(
        \pe8/got [12]) );
  DRNQHSV4 \pe8/pe2/q_reg[4]  ( .D(go7[13]), .CK(clk), .RDN(n28491), .Q(
        \pe8/got [13]) );
  DRNQHSV4 \pe8/pe2/q_reg[3]  ( .D(go7[14]), .CK(clk), .RDN(n28554), .Q(
        \pe8/got [14]) );
  DRNQHSV4 \pe8/pe5/q_reg[12]  ( .D(n28975), .CK(clk), .RDN(n28576), .Q(
        \pe8/pvq [12]) );
  DRNQHSV4 \pe8/pe5/q_reg[11]  ( .D(n28977), .CK(clk), .RDN(n28446), .Q(
        \pe8/pvq [11]) );
  DRNQHSV4 \pe8/pe5/q_reg[10]  ( .D(\pov7[10] ), .CK(clk), .RDN(n28498), .Q(
        \pe8/pvq [10]) );
  DRNQHSV4 \pe8/pe5/q_reg[9]  ( .D(n28983), .CK(clk), .RDN(n28513), .Q(
        \pe8/pvq [9]) );
  DRNQHSV4 \pe8/pe5/q_reg[8]  ( .D(n29014), .CK(clk), .RDN(n28494), .Q(
        \pe8/pvq [8]) );
  DRNQHSV4 \pe8/pe5/q_reg[6]  ( .D(n29015), .CK(clk), .RDN(n14023), .Q(
        \pe8/pvq [6]) );
  DRNQHSV4 \pe8/pe5/q_reg[5]  ( .D(n28987), .CK(clk), .RDN(n28448), .Q(
        \pe8/pvq [5]) );
  DRNQHSV4 \pe8/pe5/q_reg[4]  ( .D(n28960), .CK(clk), .RDN(n28449), .Q(
        \pe8/pvq [4]) );
  DRNQHSV4 \pe8/pe5/q_reg[3]  ( .D(n29016), .CK(clk), .RDN(n28452), .Q(
        \pe8/pvq [3]) );
  DRNQHSV4 \pe8/pe5/q_reg[2]  ( .D(n29017), .CK(clk), .RDN(n28512), .Q(
        \pe8/pvq [2]) );
  DRNQHSV4 \pe8/pe6/q_reg[15]  ( .D(poh7[15]), .CK(clk), .RDN(n28568), .Q(
        \pe8/phq [15]) );
  DRNQHSV4 \pe8/pe6/q_reg[14]  ( .D(poh7[14]), .CK(clk), .RDN(n28446), .Q(
        \pe8/phq [14]) );
  DRNQHSV4 \pe8/pe6/q_reg[13]  ( .D(poh7[13]), .CK(clk), .RDN(n28511), .Q(
        \pe8/phq [13]) );
  DRNQHSV4 \pe8/pe6/q_reg[12]  ( .D(poh7[12]), .CK(clk), .RDN(n28499), .Q(
        \pe8/phq [12]) );
  DRNQHSV4 \pe8/pe6/q_reg[11]  ( .D(poh7[11]), .CK(clk), .RDN(n28570), .Q(
        \pe8/phq [11]) );
  DRNQHSV4 \pe8/pe6/q_reg[8]  ( .D(poh7[8]), .CK(clk), .RDN(n28477), .Q(
        \pe8/phq [8]) );
  DRNQHSV4 \pe8/pe6/q_reg[7]  ( .D(poh7[7]), .CK(clk), .RDN(n28567), .Q(
        \pe8/phq [7]) );
  DRNQHSV4 \pe8/pe6/q_reg[6]  ( .D(poh7[6]), .CK(clk), .RDN(n28551), .Q(
        \pe8/phq [6]) );
  DRNQHSV4 \pe8/pe6/q_reg[5]  ( .D(poh7[5]), .CK(clk), .RDN(n28556), .Q(
        \pe8/phq [5]) );
  DRNQHSV4 \pe8/pe6/q_reg[4]  ( .D(poh7[4]), .CK(clk), .RDN(n28493), .Q(
        \pe8/phq [4]) );
  DRNQHSV4 \pe8/pe6/q_reg[3]  ( .D(poh7[3]), .CK(clk), .RDN(n28556), .Q(
        \pe8/phq [3]) );
  DRNQHSV4 \pe8/pe6/q_reg[2]  ( .D(poh7[2]), .CK(clk), .RDN(n28595), .Q(
        \pe8/phq [2]) );
  DRNQHSV4 \pe8/pe6/q_reg[1]  ( .D(poh7[1]), .CK(clk), .RDN(n28559), .Q(
        \pe8/phq [1]) );
  DRNQHSV4 \pe8/pe8/q_reg  ( .D(n25625), .CK(clk), .RDN(n28557), .Q(ctro8) );
  DRNQHSV4 \pe8/pe12/q_reg[16]  ( .D(n28895), .CK(clk), .RDN(n28442), .Q(
        \pe8/bq[1] ) );
  DRNQHSV4 \pe8/pe12/q_reg[15]  ( .D(n28896), .CK(clk), .RDN(n28539), .Q(
        \pe8/bq[2] ) );
  DRNQHSV4 \pe8/pe12/q_reg[14]  ( .D(n28891), .CK(clk), .RDN(n28602), .Q(
        \pe8/bq[3] ) );
  DRNQHSV4 \pe8/pe12/q_reg[13]  ( .D(n28893), .CK(clk), .RDN(n28555), .Q(
        \pe8/bq[4] ) );
  DRNQHSV4 \pe8/pe12/q_reg[12]  ( .D(n28892), .CK(clk), .RDN(n28604), .Q(
        \pe8/bq[5] ) );
  DRNQHSV4 \pe8/pe12/q_reg[11]  ( .D(n28894), .CK(clk), .RDN(n28573), .Q(
        \pe8/bq[6] ) );
  DRNQHSV4 \pe8/pe12/q_reg[10]  ( .D(n28890), .CK(clk), .RDN(n28541), .Q(
        \pe8/bq[7] ) );
  DRNQHSV4 \pe8/pe12/q_reg[9]  ( .D(n28889), .CK(clk), .RDN(n28535), .Q(
        \pe8/bq[8] ) );
  DRNQHSV4 \pe8/pe12/q_reg[8]  ( .D(n28888), .CK(clk), .RDN(n28556), .Q(
        \pe8/bq[9] ) );
  DRNQHSV4 \pe8/pe12/q_reg[7]  ( .D(n28887), .CK(clk), .RDN(n28554), .Q(
        \pe8/bq[10] ) );
  DRNQHSV4 \pe8/pe12/q_reg[6]  ( .D(n28883), .CK(clk), .RDN(n28486), .Q(
        \pe8/bq[11] ) );
  DRNQHSV4 \pe8/pe12/q_reg[5]  ( .D(n28885), .CK(clk), .RDN(n28530), .Q(
        \pe8/bq[12] ) );
  DRNQHSV4 \pe8/pe12/q_reg[4]  ( .D(n28886), .CK(clk), .RDN(n28459), .Q(
        \pe8/bq[13] ) );
  DRNQHSV4 \pe8/pe12/q_reg[3]  ( .D(n28882), .CK(clk), .RDN(n28607), .Q(
        \pe8/bq[14] ) );
  DRNQHSV4 \pe8/pe12/q_reg[2]  ( .D(n28881), .CK(clk), .RDN(n28446), .Q(
        \pe8/bq[15] ) );
  DRNQHSV4 \pe8/pe13/q_reg  ( .D(\pe8/ti_1t ), .CK(clk), .RDN(n28559), .Q(
        \pe8/ti_1 ) );
  DRNQHSV4 \pe8/pe14/q_reg[4]  ( .D(n16445), .CK(clk), .RDN(n28459), .Q(
        \pe8/ti_7t [4]) );
  DRNQHSV4 \pe8/pe14/q_reg[7]  ( .D(n28947), .CK(clk), .RDN(n28540), .Q(
        \pe8/ti_7t [7]) );
  DRNQHSV4 \pe9/pe1/q_reg[16]  ( .D(ao8[1]), .CK(clk), .RDN(n28498), .Q(
        \pe9/aot [1]) );
  DRNQHSV4 \pe9/pe1/q_reg[15]  ( .D(ao8[2]), .CK(clk), .RDN(n28515), .Q(
        \pe9/aot [2]) );
  DRNQHSV4 \pe9/pe1/q_reg[14]  ( .D(ao8[3]), .CK(clk), .RDN(n28453), .Q(
        \pe9/aot [3]) );
  DRNQHSV4 \pe9/pe1/q_reg[13]  ( .D(ao8[4]), .CK(clk), .RDN(n28439), .Q(
        \pe9/aot [4]) );
  DRNQHSV4 \pe9/pe1/q_reg[12]  ( .D(ao8[5]), .CK(clk), .RDN(n28449), .Q(
        \pe9/aot [5]) );
  DRNQHSV4 \pe9/pe1/q_reg[11]  ( .D(ao8[6]), .CK(clk), .RDN(n28544), .Q(
        \pe9/aot [6]) );
  DRNQHSV4 \pe9/pe1/q_reg[10]  ( .D(ao8[7]), .CK(clk), .RDN(n28545), .Q(
        \pe9/aot [7]) );
  DRNQHSV4 \pe9/pe1/q_reg[9]  ( .D(ao8[8]), .CK(clk), .RDN(n28562), .Q(
        \pe9/aot [8]) );
  DRNQHSV4 \pe9/pe1/q_reg[8]  ( .D(ao8[9]), .CK(clk), .RDN(n28493), .Q(
        \pe9/aot [9]) );
  DRNQHSV4 \pe9/pe1/q_reg[7]  ( .D(ao8[10]), .CK(clk), .RDN(n28560), .Q(
        \pe9/aot [10]) );
  DRNQHSV4 \pe9/pe1/q_reg[6]  ( .D(ao8[11]), .CK(clk), .RDN(n28502), .Q(
        \pe9/aot [11]) );
  DRNQHSV4 \pe9/pe1/q_reg[5]  ( .D(ao8[12]), .CK(clk), .RDN(n28502), .Q(
        \pe9/aot [12]) );
  DRNQHSV4 \pe9/pe1/q_reg[4]  ( .D(ao8[13]), .CK(clk), .RDN(n28524), .Q(
        \pe9/aot [13]) );
  DRNQHSV4 \pe9/pe1/q_reg[3]  ( .D(ao8[14]), .CK(clk), .RDN(n28483), .Q(
        \pe9/aot [14]) );
  DRNQHSV4 \pe9/pe1/q_reg[2]  ( .D(ao8[15]), .CK(clk), .RDN(n28555), .Q(
        \pe9/aot [15]) );
  DRNQHSV4 \pe9/pe1/q_reg[1]  ( .D(ao8[16]), .CK(clk), .RDN(n28496), .Q(
        \pe9/aot [16]) );
  DRNQHSV4 \pe9/pe2/q_reg[16]  ( .D(go8[1]), .CK(clk), .RDN(n28531), .Q(
        \pe9/got [1]) );
  DRNQHSV4 \pe9/pe2/q_reg[15]  ( .D(go8[2]), .CK(clk), .RDN(n28446), .Q(
        \pe9/got [2]) );
  DRNQHSV4 \pe9/pe2/q_reg[14]  ( .D(go8[3]), .CK(clk), .RDN(n28483), .Q(
        \pe9/got [3]) );
  DRNQHSV4 \pe9/pe2/q_reg[13]  ( .D(go8[4]), .CK(clk), .RDN(n28554), .Q(
        \pe9/got [4]) );
  DRNQHSV4 \pe9/pe2/q_reg[12]  ( .D(go8[5]), .CK(clk), .RDN(n28532), .Q(
        \pe9/got [5]) );
  DRNQHSV4 \pe9/pe2/q_reg[11]  ( .D(go8[6]), .CK(clk), .RDN(n28532), .Q(
        \pe9/got [6]) );
  DRNQHSV4 \pe9/pe2/q_reg[10]  ( .D(go8[7]), .CK(clk), .RDN(n28440), .Q(
        \pe9/got [7]) );
  DRNQHSV4 \pe9/pe2/q_reg[9]  ( .D(go8[8]), .CK(clk), .RDN(n28573), .Q(
        \pe9/got [8]) );
  DRNQHSV4 \pe9/pe2/q_reg[8]  ( .D(go8[9]), .CK(clk), .RDN(n28533), .Q(
        \pe9/got [9]) );
  DRNQHSV4 \pe9/pe2/q_reg[7]  ( .D(go8[10]), .CK(clk), .RDN(n28547), .Q(
        \pe9/got [10]) );
  DRNQHSV4 \pe9/pe2/q_reg[6]  ( .D(go8[11]), .CK(clk), .RDN(n28558), .Q(
        \pe9/got [11]) );
  DRNQHSV4 \pe9/pe2/q_reg[5]  ( .D(go8[12]), .CK(clk), .RDN(n28506), .Q(
        \pe9/got [12]) );
  DRNQHSV4 \pe9/pe2/q_reg[4]  ( .D(go8[13]), .CK(clk), .RDN(n28499), .Q(
        \pe9/got [13]) );
  DRNQHSV4 \pe9/pe2/q_reg[3]  ( .D(go8[14]), .CK(clk), .RDN(n28574), .Q(
        \pe9/got [14]) );
  DRNQHSV4 \pe9/pe2/q_reg[2]  ( .D(go8[15]), .CK(clk), .RDN(n28539), .Q(
        \pe9/got [15]) );
  DRNQHSV4 \pe9/pe2/q_reg[1]  ( .D(go8[16]), .CK(clk), .RDN(n28567), .Q(
        \pe9/got [16]) );
  DRNQHSV4 \pe9/pe5/q_reg[11]  ( .D(n29005), .CK(clk), .RDN(n28595), .Q(
        \pe9/pvq [11]) );
  DRNQHSV4 \pe9/pe5/q_reg[6]  ( .D(n29008), .CK(clk), .RDN(n28496), .Q(
        \pe9/pvq [6]) );
  DRNQHSV4 \pe9/pe5/q_reg[4]  ( .D(n29009), .CK(clk), .RDN(n28507), .Q(
        \pe9/pvq [4]) );
  DRNQHSV4 \pe9/pe5/q_reg[3]  ( .D(n29010), .CK(clk), .RDN(n28445), .Q(
        \pe9/pvq [3]) );
  DRNQHSV4 \pe9/pe5/q_reg[2]  ( .D(n29011), .CK(clk), .RDN(n28549), .Q(
        \pe9/pvq [2]) );
  DRNQHSV4 \pe9/pe6/q_reg[15]  ( .D(poh8[15]), .CK(clk), .RDN(n28508), .Q(
        \pe9/phq [15]) );
  DRNQHSV4 \pe9/pe6/q_reg[14]  ( .D(poh8[14]), .CK(clk), .RDN(n28569), .Q(
        \pe9/phq [14]) );
  DRNQHSV4 \pe9/pe6/q_reg[13]  ( .D(poh8[13]), .CK(clk), .RDN(n28569), .Q(
        \pe9/phq [13]) );
  DRNQHSV4 \pe9/pe6/q_reg[12]  ( .D(poh8[12]), .CK(clk), .RDN(n28533), .Q(
        \pe9/phq [12]) );
  DRNQHSV4 \pe9/pe6/q_reg[11]  ( .D(poh8[11]), .CK(clk), .RDN(n28547), .Q(
        \pe9/phq [11]) );
  DRNQHSV4 \pe9/pe6/q_reg[10]  ( .D(poh8[10]), .CK(clk), .RDN(n28508), .Q(
        \pe9/phq [10]) );
  DRNQHSV4 \pe9/pe6/q_reg[9]  ( .D(poh8[9]), .CK(clk), .RDN(n28567), .Q(
        \pe9/phq [9]) );
  DRNQHSV4 \pe9/pe6/q_reg[8]  ( .D(poh8[8]), .CK(clk), .RDN(n28519), .Q(
        \pe9/phq [8]) );
  DRNQHSV4 \pe9/pe6/q_reg[7]  ( .D(poh8[7]), .CK(clk), .RDN(n28509), .Q(
        \pe9/phq [7]) );
  DRNQHSV4 \pe9/pe6/q_reg[6]  ( .D(poh8[6]), .CK(clk), .RDN(n28459), .Q(
        \pe9/phq [6]) );
  DRNQHSV4 \pe9/pe6/q_reg[5]  ( .D(poh8[5]), .CK(clk), .RDN(n28509), .Q(
        \pe9/phq [5]) );
  DRNQHSV4 \pe9/pe6/q_reg[4]  ( .D(poh8[4]), .CK(clk), .RDN(n28521), .Q(
        \pe9/phq [4]) );
  DRNQHSV4 \pe9/pe6/q_reg[3]  ( .D(poh8[3]), .CK(clk), .RDN(n28458), .Q(
        \pe9/phq [3]) );
  DRNQHSV4 \pe9/pe6/q_reg[2]  ( .D(poh8[2]), .CK(clk), .RDN(n28567), .Q(
        \pe9/phq [2]) );
  DRNQHSV4 \pe9/pe6/q_reg[1]  ( .D(poh8[1]), .CK(clk), .RDN(n28535), .Q(
        \pe9/phq [1]) );
  DRNQHSV4 \pe9/pe7/q_reg  ( .D(n22138), .CK(clk), .RDN(n28528), .Q(\pe9/ctrq ) );
  DRNQHSV4 \pe9/pe8/q_reg  ( .D(n23530), .CK(clk), .RDN(n28483), .Q(ctro9) );
  DRNQHSV4 \pe9/pe12/q_reg[16]  ( .D(n28755), .CK(clk), .RDN(n28574), .Q(
        \pe9/bq[1] ) );
  DRNQHSV4 \pe9/pe12/q_reg[15]  ( .D(n28779), .CK(clk), .RDN(n28503), .Q(
        \pe9/bq[2] ) );
  DRNQHSV4 \pe9/pe12/q_reg[14]  ( .D(n28767), .CK(clk), .RDN(n28512), .Q(
        \pe9/bq[3] ) );
  DRNQHSV4 \pe9/pe12/q_reg[13]  ( .D(n28766), .CK(clk), .RDN(n28525), .Q(
        \pe9/bq[4] ) );
  DRNQHSV4 \pe9/pe12/q_reg[12]  ( .D(n28752), .CK(clk), .RDN(n28484), .Q(
        \pe9/bq[5] ) );
  DRNQHSV4 \pe9/pe12/q_reg[11]  ( .D(n28898), .CK(clk), .RDN(n28504), .Q(
        \pe9/bq[6] ) );
  DRNQHSV4 \pe9/pe12/q_reg[10]  ( .D(n28781), .CK(clk), .RDN(n28520), .Q(
        \pe9/bq[7] ) );
  DRNQHSV4 \pe9/pe12/q_reg[9]  ( .D(n28765), .CK(clk), .RDN(n28449), .Q(
        \pe9/bq[8] ) );
  DRNQHSV4 \pe9/pe12/q_reg[8]  ( .D(n28771), .CK(clk), .RDN(n28530), .Q(
        \pe9/bq[9] ) );
  DRNQHSV4 \pe9/pe12/q_reg[7]  ( .D(n28764), .CK(clk), .RDN(n28570), .Q(
        \pe9/bq[10] ) );
  DRNQHSV4 \pe9/pe12/q_reg[6]  ( .D(n28897), .CK(clk), .RDN(n28568), .Q(
        \pe9/bq[11] ) );
  DRNQHSV4 \pe9/pe12/q_reg[5]  ( .D(n28778), .CK(clk), .RDN(n28489), .Q(
        \pe9/bq[12] ) );
  DRNQHSV4 \pe9/pe12/q_reg[4]  ( .D(n28754), .CK(clk), .RDN(n28488), .Q(
        \pe9/bq[13] ) );
  DRNQHSV4 \pe9/pe12/q_reg[3]  ( .D(n28780), .CK(clk), .RDN(n28495), .Q(
        \pe9/bq[14] ) );
  DRNQHSV4 \pe9/pe12/q_reg[2]  ( .D(n28730), .CK(clk), .RDN(n28543), .Q(
        \pe9/bq[15] ) );
  DRNQHSV4 \pe9/pe12/q_reg[1]  ( .D(n28753), .CK(clk), .RDN(n28440), .Q(
        \pe9/bq[16] ) );
  DRNQHSV4 \pe9/pe13/q_reg  ( .D(\pe9/ti_1t ), .CK(clk), .RDN(n28531), .Q(
        \pe9/ti_1 ) );
  DRNQHSV4 \pe10/pe1/q_reg[16]  ( .D(ao9[1]), .CK(clk), .RDN(n28449), .Q(
        \pe10/aot [1]) );
  DRNQHSV4 \pe10/pe1/q_reg[15]  ( .D(ao9[2]), .CK(clk), .RDN(n28513), .Q(
        \pe10/aot [2]) );
  DRNQHSV4 \pe10/pe1/q_reg[14]  ( .D(ao9[3]), .CK(clk), .RDN(n28513), .Q(
        \pe10/aot [3]) );
  DRNQHSV4 \pe10/pe1/q_reg[13]  ( .D(ao9[4]), .CK(clk), .RDN(n28572), .Q(
        \pe10/aot [4]) );
  DRNQHSV4 \pe10/pe1/q_reg[12]  ( .D(ao9[5]), .CK(clk), .RDN(n14023), .Q(
        \pe10/aot [5]) );
  DRNQHSV4 \pe10/pe1/q_reg[11]  ( .D(ao9[6]), .CK(clk), .RDN(n28477), .Q(
        \pe10/aot [6]) );
  DRNQHSV4 \pe10/pe1/q_reg[10]  ( .D(ao9[7]), .CK(clk), .RDN(n28535), .Q(
        \pe10/aot [7]) );
  DRNQHSV4 \pe10/pe1/q_reg[9]  ( .D(ao9[8]), .CK(clk), .RDN(n28560), .Q(
        \pe10/aot [8]) );
  DRNQHSV4 \pe10/pe1/q_reg[8]  ( .D(ao9[9]), .CK(clk), .RDN(n28439), .Q(
        \pe10/aot [9]) );
  DRNQHSV4 \pe10/pe1/q_reg[7]  ( .D(ao9[10]), .CK(clk), .RDN(n28574), .Q(
        \pe10/aot [10]) );
  DRNQHSV4 \pe10/pe1/q_reg[6]  ( .D(ao9[11]), .CK(clk), .RDN(n28488), .Q(
        \pe10/aot [11]) );
  DRNQHSV4 \pe10/pe1/q_reg[5]  ( .D(ao9[12]), .CK(clk), .RDN(n28567), .Q(
        \pe10/aot [12]) );
  DRNQHSV4 \pe10/pe1/q_reg[4]  ( .D(ao9[13]), .CK(clk), .RDN(n28449), .Q(
        \pe10/aot [13]) );
  DRNQHSV4 \pe10/pe1/q_reg[3]  ( .D(ao9[14]), .CK(clk), .RDN(n28495), .Q(
        \pe10/aot [14]) );
  DRNQHSV4 \pe10/pe1/q_reg[2]  ( .D(ao9[15]), .CK(clk), .RDN(n28477), .Q(
        \pe10/aot [15]) );
  DRNQHSV4 \pe10/pe1/q_reg[1]  ( .D(ao9[16]), .CK(clk), .RDN(n28494), .Q(
        \pe10/aot [16]) );
  DRNQHSV4 \pe10/pe2/q_reg[16]  ( .D(go9[1]), .CK(clk), .RDN(n28510), .Q(
        \pe10/got [1]) );
  DRNQHSV4 \pe10/pe2/q_reg[15]  ( .D(go9[2]), .CK(clk), .RDN(n28596), .Q(
        \pe10/got [2]) );
  DRNQHSV4 \pe10/pe2/q_reg[14]  ( .D(go9[3]), .CK(clk), .RDN(n28524), .Q(
        \pe10/got [3]) );
  DRNQHSV4 \pe10/pe2/q_reg[13]  ( .D(go9[4]), .CK(clk), .RDN(n28556), .Q(
        \pe10/got [4]) );
  DRNQHSV4 \pe10/pe2/q_reg[12]  ( .D(go9[5]), .CK(clk), .RDN(n28560), .Q(
        \pe10/got [5]) );
  DRNQHSV4 \pe10/pe2/q_reg[11]  ( .D(go9[6]), .CK(clk), .RDN(n28543), .Q(
        \pe10/got [6]) );
  DRNQHSV4 \pe10/pe2/q_reg[10]  ( .D(go9[7]), .CK(clk), .RDN(n28493), .Q(
        \pe10/got [7]) );
  DRNQHSV4 \pe10/pe2/q_reg[9]  ( .D(go9[8]), .CK(clk), .RDN(n28490), .Q(
        \pe10/got [8]) );
  DRNQHSV4 \pe10/pe2/q_reg[8]  ( .D(go9[9]), .CK(clk), .RDN(n28507), .Q(
        \pe10/got [9]) );
  DRNQHSV4 \pe10/pe2/q_reg[7]  ( .D(go9[10]), .CK(clk), .RDN(n28487), .Q(
        \pe10/got [10]) );
  DRNQHSV4 \pe10/pe2/q_reg[6]  ( .D(go9[11]), .CK(clk), .RDN(n28521), .Q(
        \pe10/got [11]) );
  DRNQHSV4 \pe10/pe2/q_reg[5]  ( .D(go9[12]), .CK(clk), .RDN(n28510), .Q(
        \pe10/got [12]) );
  DRNQHSV4 \pe10/pe2/q_reg[4]  ( .D(go9[13]), .CK(clk), .RDN(n28449), .Q(
        \pe10/got [13]) );
  DRNQHSV4 \pe10/pe2/q_reg[3]  ( .D(go9[14]), .CK(clk), .RDN(n28577), .Q(
        \pe10/got [14]) );
  DRNQHSV4 \pe10/pe2/q_reg[2]  ( .D(go9[15]), .CK(clk), .RDN(n28559), .Q(
        \pe10/got [15]) );
  DRNQHSV4 \pe10/pe2/q_reg[1]  ( .D(go9[16]), .CK(clk), .RDN(n28537), .Q(
        \pe10/got [16]) );
  DRNQHSV4 \pe10/pe5/q_reg[11]  ( .D(pov9[11]), .CK(clk), .RDN(n28484), .Q(
        \pe10/pvq [11]) );
  DRNQHSV4 \pe10/pe5/q_reg[8]  ( .D(n28999), .CK(clk), .RDN(n28449), .Q(
        \pe10/pvq [8]) );
  DRNQHSV4 \pe10/pe5/q_reg[6]  ( .D(n28962), .CK(clk), .RDN(n28441), .Q(
        \pe10/pvq [6]) );
  DRNQHSV4 \pe10/pe5/q_reg[3]  ( .D(n29002), .CK(clk), .RDN(n28500), .Q(
        \pe10/pvq [3]) );
  DRNQHSV4 \pe10/pe5/q_reg[2]  ( .D(n29003), .CK(clk), .RDN(n28548), .Q(
        \pe10/pvq [2]) );
  DRNQHSV4 \pe10/pe5/q_reg[1]  ( .D(n28691), .CK(clk), .RDN(n28542), .Q(
        \pe10/pvq [1]) );
  DRNQHSV4 \pe10/pe6/q_reg[15]  ( .D(poh9[15]), .CK(clk), .RDN(n28564), .Q(
        \pe10/phq [15]) );
  DRNQHSV4 \pe10/pe6/q_reg[14]  ( .D(poh9[14]), .CK(clk), .RDN(n28551), .Q(
        \pe10/phq [14]) );
  DRNQHSV4 \pe10/pe6/q_reg[13]  ( .D(poh9[13]), .CK(clk), .RDN(n28513), .Q(
        \pe10/phq [13]) );
  DRNQHSV4 \pe10/pe6/q_reg[12]  ( .D(poh9[12]), .CK(clk), .RDN(n28503), .Q(
        \pe10/phq [12]) );
  DRNQHSV4 \pe10/pe6/q_reg[11]  ( .D(poh9[11]), .CK(clk), .RDN(n28447), .Q(
        \pe10/phq [11]) );
  DRNQHSV4 \pe10/pe6/q_reg[10]  ( .D(poh9[10]), .CK(clk), .RDN(n28571), .Q(
        \pe10/phq [10]) );
  DRNQHSV4 \pe10/pe6/q_reg[9]  ( .D(poh9[9]), .CK(clk), .RDN(n28536), .Q(
        \pe10/phq [9]) );
  DRNQHSV4 \pe10/pe6/q_reg[8]  ( .D(poh9[8]), .CK(clk), .RDN(n28567), .Q(
        \pe10/phq [8]) );
  DRNQHSV4 \pe10/pe6/q_reg[7]  ( .D(poh9[7]), .CK(clk), .RDN(n28554), .Q(
        \pe10/phq [7]) );
  DRNQHSV4 \pe10/pe6/q_reg[6]  ( .D(poh9[6]), .CK(clk), .RDN(n28546), .Q(
        \pe10/phq [6]) );
  DRNQHSV4 \pe10/pe6/q_reg[5]  ( .D(poh9[5]), .CK(clk), .RDN(n28568), .Q(
        \pe10/phq [5]) );
  DRNQHSV4 \pe10/pe6/q_reg[4]  ( .D(poh9[4]), .CK(clk), .RDN(n28515), .Q(
        \pe10/phq [4]) );
  DRNQHSV4 \pe10/pe6/q_reg[3]  ( .D(poh9[3]), .CK(clk), .RDN(n28554), .Q(
        \pe10/phq [3]) );
  DRNQHSV4 \pe10/pe6/q_reg[2]  ( .D(poh9[2]), .CK(clk), .RDN(n28558), .Q(
        \pe10/phq [2]) );
  DRNQHSV4 \pe10/pe6/q_reg[1]  ( .D(poh9[1]), .CK(clk), .RDN(n28490), .Q(
        \pe10/phq [1]) );
  DRNQHSV4 \pe10/pe7/q_reg  ( .D(n18641), .CK(clk), .RDN(n28531), .Q(
        \pe10/ctrq ) );
  DRNQHSV4 \pe10/pe12/q_reg[16]  ( .D(n28912), .CK(clk), .RDN(n28483), .Q(
        \pe10/bq[1] ) );
  DRNQHSV4 \pe10/pe12/q_reg[15]  ( .D(n28913), .CK(clk), .RDN(n28534), .Q(
        \pe10/bq[2] ) );
  DRNQHSV4 \pe10/pe12/q_reg[14]  ( .D(n28914), .CK(clk), .RDN(n28450), .Q(
        \pe10/bq[3] ) );
  DRNQHSV4 \pe10/pe12/q_reg[13]  ( .D(n28911), .CK(clk), .RDN(n28597), .Q(
        \pe10/bq[4] ) );
  DRNQHSV4 \pe10/pe12/q_reg[12]  ( .D(n28910), .CK(clk), .RDN(n28557), .Q(
        \pe10/bq[5] ) );
  DRNQHSV4 \pe10/pe12/q_reg[11]  ( .D(n28909), .CK(clk), .RDN(n28574), .Q(
        \pe10/bq[6] ) );
  DRNQHSV4 \pe10/pe12/q_reg[10]  ( .D(n28908), .CK(clk), .RDN(n28574), .Q(
        \pe10/bq[7] ) );
  DRNQHSV4 \pe10/pe12/q_reg[9]  ( .D(n28907), .CK(clk), .RDN(n28566), .Q(
        \pe10/bq[8] ) );
  DRNQHSV4 \pe10/pe12/q_reg[8]  ( .D(n28906), .CK(clk), .RDN(n28443), .Q(
        \pe10/bq[9] ) );
  DRNQHSV4 \pe10/pe12/q_reg[7]  ( .D(n28905), .CK(clk), .RDN(n28487), .Q(
        \pe10/bq[10] ) );
  DRNQHSV4 \pe10/pe12/q_reg[6]  ( .D(n28904), .CK(clk), .RDN(n28597), .Q(
        \pe10/bq[11] ) );
  DRNQHSV4 \pe10/pe12/q_reg[5]  ( .D(n28903), .CK(clk), .RDN(n28562), .Q(
        \pe10/bq[12] ) );
  DRNQHSV4 \pe10/pe12/q_reg[4]  ( .D(n28902), .CK(clk), .RDN(n28476), .Q(
        \pe10/bq[13] ) );
  DRNQHSV4 \pe10/pe12/q_reg[3]  ( .D(n28900), .CK(clk), .RDN(n28562), .Q(
        \pe10/bq[14] ) );
  DRNQHSV4 \pe10/pe12/q_reg[2]  ( .D(n28899), .CK(clk), .RDN(n28601), .Q(
        \pe10/bq[15] ) );
  DRNQHSV4 \pe10/pe12/q_reg[1]  ( .D(n28901), .CK(clk), .RDN(n28518), .Q(
        \pe10/bq[16] ) );
  DRNQHSV4 \pe11/pe1/q_reg[16]  ( .D(ao10[1]), .CK(clk), .RDN(n28546), .Q(
        \pe11/aot [1]) );
  DRNQHSV4 \pe11/pe1/q_reg[15]  ( .D(ao10[2]), .CK(clk), .RDN(n28458), .Q(
        \pe11/aot [2]) );
  DRNQHSV4 \pe11/pe1/q_reg[14]  ( .D(ao10[3]), .CK(clk), .RDN(n28544), .Q(
        \pe11/aot [3]) );
  DRNQHSV4 \pe11/pe1/q_reg[13]  ( .D(ao10[4]), .CK(clk), .RDN(n28446), .Q(
        \pe11/aot [4]) );
  DRNQHSV4 \pe11/pe1/q_reg[12]  ( .D(ao10[5]), .CK(clk), .RDN(n28541), .Q(
        \pe11/aot [5]) );
  DRNQHSV4 \pe11/pe1/q_reg[11]  ( .D(ao10[6]), .CK(clk), .RDN(n28486), .Q(
        \pe11/aot [6]) );
  DRNQHSV4 \pe11/pe1/q_reg[10]  ( .D(ao10[7]), .CK(clk), .RDN(n28488), .Q(
        \pe11/aot [7]) );
  DRNQHSV4 \pe11/pe1/q_reg[9]  ( .D(ao10[8]), .CK(clk), .RDN(n28521), .Q(
        \pe11/aot [8]) );
  DRNQHSV4 \pe11/pe1/q_reg[8]  ( .D(ao10[9]), .CK(clk), .RDN(n28492), .Q(
        \pe11/aot [9]) );
  DRNQHSV4 \pe11/pe1/q_reg[7]  ( .D(ao10[10]), .CK(clk), .RDN(n28496), .Q(
        \pe11/aot [10]) );
  DRNQHSV4 \pe11/pe1/q_reg[6]  ( .D(ao10[11]), .CK(clk), .RDN(n28546), .Q(
        \pe11/aot [11]) );
  DRNQHSV4 \pe11/pe1/q_reg[5]  ( .D(ao10[12]), .CK(clk), .RDN(n28451), .Q(
        \pe11/aot [12]) );
  DRNQHSV4 \pe11/pe1/q_reg[4]  ( .D(ao10[13]), .CK(clk), .RDN(n28510), .Q(
        \pe11/aot [13]) );
  DRNQHSV4 \pe11/pe1/q_reg[3]  ( .D(ao10[14]), .CK(clk), .RDN(n28446), .Q(
        \pe11/aot [14]) );
  DRNQHSV4 \pe11/pe1/q_reg[2]  ( .D(ao10[15]), .CK(clk), .RDN(n28504), .Q(
        \pe11/aot [15]) );
  DRNQHSV4 \pe11/pe1/q_reg[1]  ( .D(ao10[16]), .CK(clk), .RDN(n28552), .Q(
        \pe11/aot [16]) );
  DRNQHSV4 \pe11/pe2/q_reg[16]  ( .D(go10[1]), .CK(clk), .RDN(n28605), .Q(
        \pe11/got [1]) );
  DRNQHSV4 \pe11/pe2/q_reg[15]  ( .D(go10[2]), .CK(clk), .RDN(n28571), .Q(
        \pe11/got [2]) );
  DRNQHSV4 \pe11/pe2/q_reg[14]  ( .D(go10[3]), .CK(clk), .RDN(n28553), .Q(
        \pe11/got [3]) );
  DRNQHSV4 \pe11/pe2/q_reg[13]  ( .D(go10[4]), .CK(clk), .RDN(n28490), .Q(
        \pe11/got [4]) );
  DRNQHSV4 \pe11/pe2/q_reg[12]  ( .D(go10[5]), .CK(clk), .RDN(n28575), .Q(
        \pe11/got [5]) );
  DRNQHSV4 \pe11/pe2/q_reg[11]  ( .D(go10[6]), .CK(clk), .RDN(n28491), .Q(
        \pe11/got [6]) );
  DRNQHSV4 \pe11/pe2/q_reg[10]  ( .D(go10[7]), .CK(clk), .RDN(n28607), .Q(
        \pe11/got [7]) );
  DRNQHSV4 \pe11/pe2/q_reg[9]  ( .D(go10[8]), .CK(clk), .RDN(n28477), .Q(
        \pe11/got [8]) );
  DRNQHSV4 \pe11/pe2/q_reg[8]  ( .D(go10[9]), .CK(clk), .RDN(n28517), .Q(
        \pe11/got [9]) );
  DRNQHSV4 \pe11/pe2/q_reg[7]  ( .D(go10[10]), .CK(clk), .RDN(n28443), .Q(
        \pe11/got [10]) );
  DRNQHSV4 \pe11/pe2/q_reg[6]  ( .D(go10[11]), .CK(clk), .RDN(n28443), .Q(
        \pe11/got [11]) );
  DRNQHSV4 \pe11/pe2/q_reg[5]  ( .D(go10[12]), .CK(clk), .RDN(n28439), .Q(
        \pe11/got [12]) );
  DRNQHSV4 \pe11/pe2/q_reg[4]  ( .D(go10[13]), .CK(clk), .RDN(n28515), .Q(
        \pe11/got [13]) );
  DRNQHSV4 \pe11/pe2/q_reg[3]  ( .D(go10[14]), .CK(clk), .RDN(n28534), .Q(
        \pe11/got [14]) );
  DRNQHSV4 \pe11/pe2/q_reg[2]  ( .D(go10[15]), .CK(clk), .RDN(n28535), .Q(
        \pe11/got [15]) );
  DRNQHSV4 \pe11/pe2/q_reg[1]  ( .D(go10[16]), .CK(clk), .RDN(n28495), .Q(
        \pe11/got [16]) );
  DRNQHSV4 \pe11/pe5/q_reg[12]  ( .D(n28995), .CK(clk), .RDN(n28557), .Q(
        \pe11/pvq [12]) );
  DRNQHSV4 \pe11/pe5/q_reg[10]  ( .D(pov10[10]), .CK(clk), .RDN(n28521), .Q(
        \pe11/pvq [10]) );
  DRNQHSV4 \pe11/pe5/q_reg[5]  ( .D(n28982), .CK(clk), .RDN(n28514), .Q(
        \pe11/pvq [5]) );
  DRNQHSV4 \pe11/pe5/q_reg[3]  ( .D(n28944), .CK(clk), .RDN(n28544), .Q(
        \pe11/pvq [3]) );
  DRNQHSV4 \pe11/pe5/q_reg[2]  ( .D(n28998), .CK(clk), .RDN(n28568), .Q(
        \pe11/pvq [2]) );
  DRNQHSV4 \pe11/pe6/q_reg[15]  ( .D(poh10[15]), .CK(clk), .RDN(n28597), .Q(
        \pe11/phq [15]) );
  DRNQHSV4 \pe11/pe6/q_reg[14]  ( .D(poh10[14]), .CK(clk), .RDN(n28547), .Q(
        \pe11/phq [14]) );
  DRNQHSV4 \pe11/pe6/q_reg[13]  ( .D(poh10[13]), .CK(clk), .RDN(n28570), .Q(
        \pe11/phq [13]) );
  DRNQHSV4 \pe11/pe6/q_reg[12]  ( .D(poh10[12]), .CK(clk), .RDN(n28519), .Q(
        \pe11/phq [12]) );
  DRNQHSV4 \pe11/pe6/q_reg[11]  ( .D(poh10[11]), .CK(clk), .RDN(n28572), .Q(
        \pe11/phq [11]) );
  DRNQHSV4 \pe11/pe6/q_reg[10]  ( .D(poh10[10]), .CK(clk), .RDN(n28552), .Q(
        \pe11/phq [10]) );
  DRNQHSV4 \pe11/pe6/q_reg[9]  ( .D(poh10[9]), .CK(clk), .RDN(n28541), .Q(
        \pe11/phq [9]) );
  DRNQHSV4 \pe11/pe6/q_reg[8]  ( .D(poh10[8]), .CK(clk), .RDN(n28505), .Q(
        \pe11/phq [8]) );
  DRNQHSV4 \pe11/pe6/q_reg[7]  ( .D(poh10[7]), .CK(clk), .RDN(n28595), .Q(
        \pe11/phq [7]) );
  DRNQHSV4 \pe11/pe6/q_reg[6]  ( .D(poh10[6]), .CK(clk), .RDN(n28520), .Q(
        \pe11/phq [6]) );
  DRNQHSV4 \pe11/pe6/q_reg[5]  ( .D(poh10[5]), .CK(clk), .RDN(n28569), .Q(
        \pe11/phq [5]) );
  DRNQHSV4 \pe11/pe6/q_reg[4]  ( .D(poh10[4]), .CK(clk), .RDN(n28571), .Q(
        \pe11/phq [4]) );
  DRNQHSV4 \pe11/pe6/q_reg[3]  ( .D(poh10[3]), .CK(clk), .RDN(n28528), .Q(
        \pe11/phq [3]) );
  DRNQHSV4 \pe11/pe6/q_reg[2]  ( .D(poh10[2]), .CK(clk), .RDN(n28518), .Q(
        \pe11/phq [2]) );
  DRNQHSV4 \pe11/pe6/q_reg[1]  ( .D(poh10[1]), .CK(clk), .RDN(n28528), .Q(
        \pe11/phq [1]) );
  DRNQHSV4 \pe11/pe7/q_reg  ( .D(n20148), .CK(clk), .RDN(n28506), .Q(
        \pe11/ctrq ) );
  DRNQHSV4 \pe11/pe12/q_reg[16]  ( .D(n28727), .CK(clk), .RDN(n28532), .Q(
        \pe11/bq[1] ) );
  DRNQHSV4 \pe11/pe12/q_reg[15]  ( .D(n28721), .CK(clk), .RDN(n28564), .Q(
        \pe11/bq[2] ) );
  DRNQHSV4 \pe11/pe12/q_reg[14]  ( .D(n28720), .CK(clk), .RDN(n28571), .Q(
        \pe11/bq[3] ) );
  DRNQHSV4 \pe11/pe12/q_reg[13]  ( .D(n28723), .CK(clk), .RDN(n28601), .Q(
        \pe11/bq[4] ) );
  DRNQHSV4 \pe11/pe12/q_reg[12]  ( .D(n28722), .CK(clk), .RDN(n28506), .Q(
        \pe11/bq[5] ) );
  DRNQHSV4 \pe11/pe12/q_reg[11]  ( .D(n28724), .CK(clk), .RDN(n28509), .Q(
        \pe11/bq[6] ) );
  DRNQHSV4 \pe11/pe12/q_reg[10]  ( .D(n28719), .CK(clk), .RDN(n28448), .Q(
        \pe11/bq[7] ) );
  DRNQHSV4 \pe11/pe12/q_reg[9]  ( .D(n28718), .CK(clk), .RDN(n28444), .Q(
        \pe11/bq[8] ) );
  DRNQHSV4 \pe11/pe12/q_reg[8]  ( .D(n28917), .CK(clk), .RDN(n28566), .Q(
        \pe11/bq[9] ) );
  DRNQHSV4 \pe11/pe12/q_reg[7]  ( .D(n28916), .CK(clk), .RDN(n28595), .Q(
        \pe11/bq[10] ) );
  DRNQHSV4 \pe11/pe12/q_reg[6]  ( .D(n28728), .CK(clk), .RDN(n28518), .Q(
        \pe11/bq[11] ) );
  DRNQHSV4 \pe11/pe12/q_reg[5]  ( .D(n28915), .CK(clk), .RDN(n28524), .Q(
        \pe11/bq[12] ) );
  DRNQHSV4 \pe11/pe12/q_reg[4]  ( .D(n28726), .CK(clk), .RDN(n28486), .Q(
        \pe11/bq[13] ) );
  DRNQHSV4 \pe11/pe12/q_reg[3]  ( .D(n28717), .CK(clk), .RDN(n28570), .Q(
        \pe11/bq[14] ) );
  DRNQHSV4 \pe11/pe12/q_reg[2]  ( .D(n28725), .CK(clk), .RDN(n28507), .Q(
        \pe11/bq[15] ) );
  DRNQHSV4 \pe11/pe12/q_reg[1]  ( .D(n28729), .CK(clk), .RDN(n14021), .Q(
        \pe11/bq[16] ) );
  DRNQHSV4 \pe11/pe13/q_reg  ( .D(\pe11/ti_1t ), .CK(clk), .RDN(n28577), .Q(
        \pe11/ti_1 ) );
  DRNQHSV1 \pe7/pe14/q_reg[8]  ( .D(n28587), .CK(clk), .RDN(n28517), .Q(
        \pe7/ti_7t [8]) );
  DRNQHSV1 \pe6/pe5/q_reg[13]  ( .D(n28969), .CK(clk), .RDN(n28574), .Q(
        \pe6/pvq [13]) );
  DRNQHSV2 \pe4/pe14/q_reg[2]  ( .D(n28671), .CK(clk), .RDN(n28512), .Q(
        \pe4/ti_7t [2]) );
  DRNQHSV1 \pe6/pe5/q_reg[6]  ( .D(pov5[6]), .CK(clk), .RDN(n28458), .Q(
        \pe6/pvq [6]) );
  DRNQHSV2 \pe8/pe5/q_reg[7]  ( .D(n28985), .CK(clk), .RDN(n28552), .Q(
        \pe8/pvq [7]) );
  DRNQHSV1 \pe8/pe14/q_reg[2]  ( .D(n28788), .CK(clk), .RDN(n28493), .Q(
        \pe8/ti_7t [2]) );
  DRNQHSV2 \pe7/pe14/q_reg[9]  ( .D(n28430), .CK(clk), .RDN(n28503), .Q(
        \pe7/ti_7t [9]) );
  DRNQHSV1 \pe7/pe14/q_reg[14]  ( .D(n28703), .CK(clk), .RDN(n28500), .Q(
        \pe7/ti_7t [14]) );
  DRNQHSV2 \pe8/pe6/q_reg[10]  ( .D(poh7[10]), .CK(clk), .RDN(n28502), .Q(
        \pe8/phq [10]) );
  DRNQHSV1 \pe10/pe5/q_reg[12]  ( .D(n28705), .CK(clk), .RDN(n14023), .Q(
        \pe10/pvq [12]) );
  DRNQHSV1 \pe10/pe5/q_reg[10]  ( .D(n28964), .CK(clk), .RDN(n28447), .Q(
        \pe10/pvq [10]) );
  DRNQHSV1 \pe4/pe14/q_reg[4]  ( .D(n28923), .CK(clk), .RDN(n28575), .Q(
        \pe4/ti_7t [4]) );
  DRNQHSV1 \pe7/pe5/q_reg[6]  ( .D(n28966), .CK(clk), .RDN(n28527), .Q(
        \pe7/pvq [6]) );
  DRNQHSV1 \pe6/pe14/q_reg[15]  ( .D(n25784), .CK(clk), .RDN(n28607), .Q(
        \pe6/ti_7t [15]) );
  DRNQHSV4 \pe1/pe8/q_reg  ( .D(n28598), .CK(clk), .RDN(n28575), .Q(ctro1) );
  DRNQHSV1 \pe2/pe17/q_reg[3]  ( .D(\pe2/poht [3]), .CK(clk), .RDN(n28491), 
        .Q(poh2[3]) );
  DRNQHSV2 \pe4/pe14/q_reg[10]  ( .D(n28583), .CK(clk), .RDN(n28548), .Q(
        \pe4/ti_7t [10]) );
  DRNQHSV2 \pe11/pe3/q_reg[16]  ( .D(bo10[1]), .CK(clk), .RDN(n28486), .Q(
        bo11[1]) );
  DRNQHSV2 \pe11/pe3/q_reg[15]  ( .D(bo10[2]), .CK(clk), .RDN(n14021), .Q(
        bo11[2]) );
  DRNQHSV2 \pe11/pe3/q_reg[14]  ( .D(bo10[3]), .CK(clk), .RDN(n28524), .Q(
        bo11[3]) );
  DRNQHSV2 \pe11/pe3/q_reg[13]  ( .D(bo10[4]), .CK(clk), .RDN(n28539), .Q(
        bo11[4]) );
  DRNQHSV2 \pe11/pe3/q_reg[12]  ( .D(bo10[5]), .CK(clk), .RDN(n28511), .Q(
        bo11[5]) );
  DRNQHSV2 \pe11/pe3/q_reg[11]  ( .D(bo10[6]), .CK(clk), .RDN(n28458), .Q(
        bo11[6]) );
  DRNQHSV2 \pe11/pe3/q_reg[10]  ( .D(bo10[7]), .CK(clk), .RDN(n28574), .Q(
        bo11[7]) );
  DRNQHSV2 \pe11/pe3/q_reg[9]  ( .D(bo10[8]), .CK(clk), .RDN(n28532), .Q(
        bo11[8]) );
  DRNQHSV2 \pe11/pe3/q_reg[6]  ( .D(bo10[11]), .CK(clk), .RDN(n28529), .Q(
        bo11[11]) );
  DRNQHSV2 \pe11/pe3/q_reg[4]  ( .D(bo10[13]), .CK(clk), .RDN(n28498), .Q(
        bo11[13]) );
  DRNQHSV2 \pe11/pe3/q_reg[3]  ( .D(bo10[14]), .CK(clk), .RDN(n28533), .Q(
        bo11[14]) );
  DRNQHSV2 \pe11/pe3/q_reg[2]  ( .D(bo10[15]), .CK(clk), .RDN(n28543), .Q(
        bo11[15]) );
  DRNQHSV2 \pe11/pe3/q_reg[1]  ( .D(bo10[16]), .CK(clk), .RDN(n28494), .Q(
        bo11[16]) );
  DRNQHSV1 \pe1/pe14/q_reg[13]  ( .D(n28700), .CK(clk), .RDN(n28512), .Q(
        \pe1/ti_7t [13]) );
  DRNQHSV1 \pe3/pe14/q_reg[13]  ( .D(n28652), .CK(clk), .RDN(n28575), .Q(
        \pe3/ti_7t [13]) );
  DRNQHSV1 \pe7/pe14/q_reg[15]  ( .D(n28659), .CK(clk), .RDN(n28493), .Q(
        \pe7/ti_7t [15]) );
  DRNQHSV1 \pe8/pe14/q_reg[15]  ( .D(n28420), .CK(clk), .RDN(n28447), .Q(
        \pe8/ti_7t [15]) );
  DRNQHSV1 \pe1/pe15/q_reg[16]  ( .D(\pe1/aot [1]), .CK(clk), .RDN(n28497), 
        .Q(ao1[1]) );
  DRNQHSV1 \pe1/pe15/q_reg[15]  ( .D(\pe1/aot [2]), .CK(clk), .RDN(n28451), 
        .Q(ao1[2]) );
  DRNQHSV1 \pe1/pe15/q_reg[14]  ( .D(\pe1/aot [3]), .CK(clk), .RDN(n28484), 
        .Q(ao1[3]) );
  DRNQHSV1 \pe1/pe15/q_reg[13]  ( .D(\pe1/aot [4]), .CK(clk), .RDN(n28458), 
        .Q(ao1[4]) );
  DRNQHSV1 \pe1/pe15/q_reg[12]  ( .D(\pe1/aot [5]), .CK(clk), .RDN(n28441), 
        .Q(ao1[5]) );
  DRNQHSV1 \pe1/pe15/q_reg[11]  ( .D(\pe1/aot [6]), .CK(clk), .RDN(n28563), 
        .Q(ao1[6]) );
  DRNQHSV1 \pe1/pe15/q_reg[10]  ( .D(\pe1/aot [7]), .CK(clk), .RDN(n28558), 
        .Q(ao1[7]) );
  DRNQHSV1 \pe1/pe15/q_reg[9]  ( .D(\pe1/aot [8]), .CK(clk), .RDN(n28557), .Q(
        ao1[8]) );
  DRNQHSV1 \pe1/pe15/q_reg[8]  ( .D(\pe1/aot [9]), .CK(clk), .RDN(n28442), .Q(
        ao1[9]) );
  DRNQHSV1 \pe1/pe15/q_reg[7]  ( .D(\pe1/aot [10]), .CK(clk), .RDN(n28552), 
        .Q(ao1[10]) );
  DRNQHSV1 \pe1/pe15/q_reg[6]  ( .D(\pe1/aot [11]), .CK(clk), .RDN(n28520), 
        .Q(ao1[11]) );
  DRNQHSV1 \pe1/pe15/q_reg[5]  ( .D(\pe1/aot [12]), .CK(clk), .RDN(n28533), 
        .Q(ao1[12]) );
  DRNQHSV1 \pe1/pe15/q_reg[4]  ( .D(\pe1/aot [13]), .CK(clk), .RDN(n28517), 
        .Q(ao1[13]) );
  DRNQHSV1 \pe1/pe15/q_reg[3]  ( .D(\pe1/aot [14]), .CK(clk), .RDN(n28601), 
        .Q(ao1[14]) );
  DRNQHSV1 \pe1/pe15/q_reg[2]  ( .D(n28468), .CK(clk), .RDN(n28521), .Q(
        ao1[15]) );
  DRNQHSV1 \pe1/pe15/q_reg[1]  ( .D(n28485), .CK(clk), .RDN(n28577), .Q(
        ao1[16]) );
  DRNQHSV1 \pe1/pe16/q_reg[16]  ( .D(\pe1/got [1]), .CK(clk), .RDN(n28558), 
        .Q(go1[1]) );
  DRNQHSV1 \pe1/pe16/q_reg[15]  ( .D(\pe1/got [2]), .CK(clk), .RDN(n28494), 
        .Q(go1[2]) );
  DRNQHSV1 \pe1/pe16/q_reg[14]  ( .D(\pe1/got [3]), .CK(clk), .RDN(n28459), 
        .Q(go1[3]) );
  DRNQHSV1 \pe1/pe16/q_reg[13]  ( .D(n28435), .CK(clk), .RDN(n28597), .Q(
        go1[4]) );
  DRNQHSV1 \pe1/pe16/q_reg[12]  ( .D(\pe1/got [5]), .CK(clk), .RDN(n28572), 
        .Q(go1[5]) );
  DRNQHSV1 \pe1/pe16/q_reg[11]  ( .D(n28434), .CK(clk), .RDN(n28597), .Q(
        go1[6]) );
  DRNQHSV1 \pe1/pe16/q_reg[10]  ( .D(\pe1/got [7]), .CK(clk), .RDN(n28542), 
        .Q(go1[7]) );
  DRNQHSV1 \pe1/pe16/q_reg[9]  ( .D(\pe1/got [8]), .CK(clk), .RDN(n28525), .Q(
        go1[8]) );
  DRNQHSV1 \pe1/pe16/q_reg[8]  ( .D(\pe1/got [9]), .CK(clk), .RDN(n28522), .Q(
        go1[9]) );
  DRNQHSV1 \pe1/pe16/q_reg[7]  ( .D(n28615), .CK(clk), .RDN(n28512), .Q(
        go1[10]) );
  DRNQHSV1 \pe1/pe16/q_reg[6]  ( .D(\pe1/got [11]), .CK(clk), .RDN(n28562), 
        .Q(go1[11]) );
  DRNQHSV1 \pe1/pe16/q_reg[5]  ( .D(n28425), .CK(clk), .RDN(n28498), .Q(
        go1[12]) );
  DRNQHSV1 \pe1/pe16/q_reg[4]  ( .D(\pe1/got [13]), .CK(clk), .RDN(n28545), 
        .Q(go1[13]) );
  DRNQHSV1 \pe1/pe16/q_reg[3]  ( .D(\pe1/got [14]), .CK(clk), .RDN(n28511), 
        .Q(go1[14]) );
  DRNQHSV1 \pe1/pe16/q_reg[2]  ( .D(\pe1/got [15]), .CK(clk), .RDN(n28539), 
        .Q(go1[15]) );
  DRNQHSV1 \pe1/pe16/q_reg[1]  ( .D(n28422), .CK(clk), .RDN(n28561), .Q(
        go1[16]) );
  DRNQHSV2 \pe1/pe17/q_reg[15]  ( .D(\pe1/poht [15]), .CK(clk), .RDN(n28544), 
        .Q(poh1[15]) );
  DRNQHSV2 \pe1/pe17/q_reg[13]  ( .D(\pe1/poht [13]), .CK(clk), .RDN(n28545), 
        .Q(poh1[13]) );
  DRNQHSV2 \pe1/pe17/q_reg[11]  ( .D(\pe1/poht [11]), .CK(clk), .RDN(n28511), 
        .Q(poh1[11]) );
  DRNQHSV2 \pe1/pe17/q_reg[8]  ( .D(\pe1/poht [8]), .CK(clk), .RDN(n28544), 
        .Q(poh1[8]) );
  DRNQHSV2 \pe1/pe17/q_reg[6]  ( .D(\pe1/poht [6]), .CK(clk), .RDN(n28508), 
        .Q(poh1[6]) );
  DRNQHSV2 \pe1/pe17/q_reg[3]  ( .D(\pe1/poht [3]), .CK(clk), .RDN(n28503), 
        .Q(poh1[3]) );
  DRNQHSV1 \pe2/pe15/q_reg[16]  ( .D(\pe2/aot [1]), .CK(clk), .RDN(n28568), 
        .Q(ao2[1]) );
  DRNQHSV1 \pe2/pe15/q_reg[15]  ( .D(\pe2/aot [2]), .CK(clk), .RDN(n28440), 
        .Q(ao2[2]) );
  DRNQHSV1 \pe2/pe15/q_reg[14]  ( .D(\pe2/aot [3]), .CK(clk), .RDN(n28487), 
        .Q(ao2[3]) );
  DRNQHSV1 \pe2/pe15/q_reg[13]  ( .D(\pe2/aot [4]), .CK(clk), .RDN(n28451), 
        .Q(ao2[4]) );
  DRNQHSV1 \pe2/pe15/q_reg[12]  ( .D(\pe2/aot [5]), .CK(clk), .RDN(n28515), 
        .Q(ao2[5]) );
  DRNQHSV1 \pe2/pe15/q_reg[11]  ( .D(\pe2/aot [6]), .CK(clk), .RDN(n28548), 
        .Q(ao2[6]) );
  DRNQHSV1 \pe2/pe15/q_reg[10]  ( .D(\pe2/aot [7]), .CK(clk), .RDN(n28537), 
        .Q(ao2[7]) );
  DRNQHSV1 \pe2/pe15/q_reg[9]  ( .D(\pe2/aot [8]), .CK(clk), .RDN(n28452), .Q(
        ao2[8]) );
  DRNQHSV1 \pe2/pe15/q_reg[8]  ( .D(\pe2/aot [9]), .CK(clk), .RDN(n28575), .Q(
        ao2[9]) );
  DRNQHSV1 \pe2/pe15/q_reg[7]  ( .D(\pe2/aot [10]), .CK(clk), .RDN(n28568), 
        .Q(ao2[10]) );
  DRNQHSV1 \pe2/pe15/q_reg[6]  ( .D(\pe2/aot [11]), .CK(clk), .RDN(n28540), 
        .Q(ao2[11]) );
  DRNQHSV1 \pe2/pe15/q_reg[5]  ( .D(\pe2/aot [12]), .CK(clk), .RDN(n28604), 
        .Q(ao2[12]) );
  DRNQHSV1 \pe2/pe15/q_reg[4]  ( .D(\pe2/aot [13]), .CK(clk), .RDN(n28606), 
        .Q(ao2[13]) );
  DRNQHSV1 \pe2/pe15/q_reg[3]  ( .D(n14020), .CK(clk), .RDN(n28516), .Q(
        ao2[14]) );
  DRNQHSV1 \pe2/pe15/q_reg[2]  ( .D(\pe2/aot [15]), .CK(clk), .RDN(n28553), 
        .Q(ao2[15]) );
  DRNQHSV1 \pe2/pe15/q_reg[1]  ( .D(n11953), .CK(clk), .RDN(n28568), .Q(
        ao2[16]) );
  DRNQHSV1 \pe2/pe16/q_reg[16]  ( .D(\pe2/got [1]), .CK(clk), .RDN(n28459), 
        .Q(go2[1]) );
  DRNQHSV1 \pe2/pe16/q_reg[15]  ( .D(\pe2/got [2]), .CK(clk), .RDN(n28560), 
        .Q(go2[2]) );
  DRNQHSV1 \pe2/pe16/q_reg[14]  ( .D(n14062), .CK(clk), .RDN(n28540), .Q(
        go2[3]) );
  DRNQHSV1 \pe2/pe16/q_reg[13]  ( .D(n28634), .CK(clk), .RDN(n28572), .Q(
        go2[4]) );
  DRNQHSV1 \pe2/pe16/q_reg[12]  ( .D(\pe2/got [5]), .CK(clk), .RDN(n28544), 
        .Q(go2[5]) );
  DRNQHSV1 \pe2/pe16/q_reg[11]  ( .D(n14006), .CK(clk), .RDN(n28543), .Q(
        go2[6]) );
  DRNQHSV1 \pe2/pe16/q_reg[10]  ( .D(\pe2/got [7]), .CK(clk), .RDN(n28450), 
        .Q(go2[7]) );
  DRNQHSV1 \pe2/pe16/q_reg[9]  ( .D(\pe2/got [8]), .CK(clk), .RDN(n28540), .Q(
        go2[8]) );
  DRNQHSV1 \pe2/pe16/q_reg[8]  ( .D(n28636), .CK(clk), .RDN(n14023), .Q(go2[9]) );
  DRNQHSV1 \pe2/pe16/q_reg[7]  ( .D(\pe2/got [10]), .CK(clk), .RDN(n28495), 
        .Q(go2[10]) );
  DRNQHSV1 \pe2/pe16/q_reg[6]  ( .D(\pe2/got [11]), .CK(clk), .RDN(n28522), 
        .Q(go2[11]) );
  DRNQHSV1 \pe2/pe16/q_reg[5]  ( .D(\pe2/got [12]), .CK(clk), .RDN(n28536), 
        .Q(go2[12]) );
  DRNQHSV1 \pe2/pe16/q_reg[4]  ( .D(n28429), .CK(clk), .RDN(n28536), .Q(
        go2[13]) );
  DRNQHSV1 \pe2/pe16/q_reg[3]  ( .D(\pe2/got [14]), .CK(clk), .RDN(n28497), 
        .Q(go2[14]) );
  DRNQHSV1 \pe2/pe16/q_reg[2]  ( .D(n28421), .CK(clk), .RDN(n28606), .Q(
        go2[15]) );
  DRNQHSV1 \pe2/pe16/q_reg[1]  ( .D(n28693), .CK(clk), .RDN(n28536), .Q(
        go2[16]) );
  DRNQHSV2 \pe2/pe17/q_reg[15]  ( .D(\pe2/poht [15]), .CK(clk), .RDN(n28484), 
        .Q(poh2[15]) );
  DRNQHSV1 \pe2/pe17/q_reg[9]  ( .D(\pe2/poht [9]), .CK(clk), .RDN(n14023), 
        .Q(poh2[9]) );
  DRNQHSV1 \pe2/pe17/q_reg[4]  ( .D(\pe2/poht [4]), .CK(clk), .RDN(n28527), 
        .Q(poh2[4]) );
  DRNQHSV1 \pe2/pe17/q_reg[2]  ( .D(\pe2/poht [2]), .CK(clk), .RDN(n28520), 
        .Q(poh2[2]) );
  DRNQHSV1 \pe2/pe17/q_reg[1]  ( .D(\pe2/poht [1]), .CK(clk), .RDN(n28451), 
        .Q(poh2[1]) );
  DRNQHSV1 \pe3/pe15/q_reg[16]  ( .D(\pe3/aot [1]), .CK(clk), .RDN(n28450), 
        .Q(ao3[1]) );
  DRNQHSV1 \pe3/pe15/q_reg[15]  ( .D(\pe3/aot [2]), .CK(clk), .RDN(n28536), 
        .Q(ao3[2]) );
  DRNQHSV1 \pe3/pe15/q_reg[14]  ( .D(\pe3/aot [3]), .CK(clk), .RDN(n28529), 
        .Q(ao3[3]) );
  DRNQHSV1 \pe3/pe15/q_reg[13]  ( .D(\pe3/aot [4]), .CK(clk), .RDN(n28484), 
        .Q(ao3[4]) );
  DRNQHSV1 \pe3/pe15/q_reg[12]  ( .D(\pe3/aot [5]), .CK(clk), .RDN(n28497), 
        .Q(ao3[5]) );
  DRNQHSV1 \pe3/pe15/q_reg[11]  ( .D(\pe3/aot [6]), .CK(clk), .RDN(n28451), 
        .Q(ao3[6]) );
  DRNQHSV1 \pe3/pe15/q_reg[10]  ( .D(\pe3/aot [7]), .CK(clk), .RDN(n28565), 
        .Q(ao3[7]) );
  DRNQHSV1 \pe3/pe15/q_reg[9]  ( .D(\pe3/aot [8]), .CK(clk), .RDN(n28535), .Q(
        ao3[8]) );
  DRNQHSV1 \pe3/pe15/q_reg[8]  ( .D(\pe3/aot [9]), .CK(clk), .RDN(n28518), .Q(
        ao3[9]) );
  DRNQHSV1 \pe3/pe15/q_reg[7]  ( .D(\pe3/aot [10]), .CK(clk), .RDN(n28508), 
        .Q(ao3[10]) );
  DRNQHSV1 \pe3/pe15/q_reg[6]  ( .D(\pe3/aot [11]), .CK(clk), .RDN(n28538), 
        .Q(ao3[11]) );
  DRNQHSV1 \pe3/pe15/q_reg[5]  ( .D(\pe3/aot [12]), .CK(clk), .RDN(n28448), 
        .Q(ao3[12]) );
  DRNQHSV1 \pe3/pe15/q_reg[4]  ( .D(n11932), .CK(clk), .RDN(n28476), .Q(
        ao3[13]) );
  DRNQHSV1 \pe3/pe15/q_reg[3]  ( .D(\pe3/aot [14]), .CK(clk), .RDN(n28564), 
        .Q(ao3[14]) );
  DRNQHSV1 \pe3/pe15/q_reg[2]  ( .D(\pe3/aot [15]), .CK(clk), .RDN(n28511), 
        .Q(ao3[15]) );
  DRNQHSV1 \pe3/pe15/q_reg[1]  ( .D(n14040), .CK(clk), .RDN(n28459), .Q(
        ao3[16]) );
  DRNQHSV1 \pe3/pe16/q_reg[16]  ( .D(\pe3/got [1]), .CK(clk), .RDN(n28553), 
        .Q(go3[1]) );
  DRNQHSV1 \pe3/pe16/q_reg[15]  ( .D(\pe3/got [2]), .CK(clk), .RDN(n28499), 
        .Q(go3[2]) );
  DRNQHSV1 \pe3/pe16/q_reg[14]  ( .D(\pe3/got [3]), .CK(clk), .RDN(n28504), 
        .Q(go3[3]) );
  DRNQHSV1 \pe3/pe16/q_reg[13]  ( .D(\pe3/got [4]), .CK(clk), .RDN(n28447), 
        .Q(go3[4]) );
  DRNQHSV1 \pe3/pe16/q_reg[12]  ( .D(\pe3/got [5]), .CK(clk), .RDN(n28451), 
        .Q(go3[5]) );
  DRNQHSV1 \pe3/pe16/q_reg[11]  ( .D(\pe3/got [6]), .CK(clk), .RDN(n28602), 
        .Q(go3[6]) );
  DRNQHSV1 \pe3/pe16/q_reg[10]  ( .D(\pe3/got [7]), .CK(clk), .RDN(n28556), 
        .Q(go3[7]) );
  DRNQHSV1 \pe3/pe16/q_reg[9]  ( .D(n14074), .CK(clk), .RDN(n28601), .Q(go3[8]) );
  DRNQHSV1 \pe3/pe16/q_reg[8]  ( .D(\pe3/got [9]), .CK(clk), .RDN(n28550), .Q(
        go3[9]) );
  DRNQHSV1 \pe3/pe16/q_reg[7]  ( .D(\pe3/got [10]), .CK(clk), .RDN(n28539), 
        .Q(go3[10]) );
  DRNQHSV1 \pe3/pe16/q_reg[6]  ( .D(\pe3/got [11]), .CK(clk), .RDN(n28562), 
        .Q(go3[11]) );
  DRNQHSV1 \pe3/pe16/q_reg[5]  ( .D(n11891), .CK(clk), .RDN(n28534), .Q(
        go3[12]) );
  DRNQHSV1 \pe3/pe16/q_reg[4]  ( .D(n28628), .CK(clk), .RDN(n28547), .Q(
        go3[13]) );
  DRNQHSV1 \pe3/pe16/q_reg[3]  ( .D(n15086), .CK(clk), .RDN(n28500), .Q(
        go3[14]) );
  DRNQHSV2 \pe3/pe17/q_reg[15]  ( .D(\pe3/poht [15]), .CK(clk), .RDN(n28525), 
        .Q(poh3[15]) );
  DRNQHSV2 \pe3/pe17/q_reg[14]  ( .D(\pe3/poht [14]), .CK(clk), .RDN(n28521), 
        .Q(poh3[14]) );
  DRNQHSV2 \pe3/pe17/q_reg[13]  ( .D(\pe3/poht [13]), .CK(clk), .RDN(n28537), 
        .Q(poh3[13]) );
  DRNQHSV2 \pe3/pe17/q_reg[6]  ( .D(\pe3/poht [6]), .CK(clk), .RDN(n28519), 
        .Q(poh3[6]) );
  DRNQHSV1 \pe4/pe15/q_reg[16]  ( .D(\pe4/aot [1]), .CK(clk), .RDN(n28488), 
        .Q(ao4[1]) );
  DRNQHSV1 \pe4/pe15/q_reg[15]  ( .D(\pe4/aot [2]), .CK(clk), .RDN(n28476), 
        .Q(ao4[2]) );
  DRNQHSV1 \pe4/pe15/q_reg[14]  ( .D(\pe4/aot [3]), .CK(clk), .RDN(n28507), 
        .Q(ao4[3]) );
  DRNQHSV1 \pe4/pe15/q_reg[13]  ( .D(\pe4/aot [4]), .CK(clk), .RDN(n28565), 
        .Q(ao4[4]) );
  DRNQHSV1 \pe4/pe15/q_reg[12]  ( .D(\pe4/aot [5]), .CK(clk), .RDN(n28538), 
        .Q(ao4[5]) );
  DRNQHSV1 \pe4/pe15/q_reg[11]  ( .D(\pe4/aot [6]), .CK(clk), .RDN(n28534), 
        .Q(ao4[6]) );
  DRNQHSV1 \pe4/pe15/q_reg[10]  ( .D(\pe4/aot [7]), .CK(clk), .RDN(n28528), 
        .Q(ao4[7]) );
  DRNQHSV1 \pe4/pe15/q_reg[9]  ( .D(\pe4/aot [8]), .CK(clk), .RDN(n28606), .Q(
        ao4[8]) );
  DRNQHSV1 \pe4/pe15/q_reg[8]  ( .D(\pe4/aot [9]), .CK(clk), .RDN(n28445), .Q(
        ao4[9]) );
  DRNQHSV1 \pe4/pe15/q_reg[7]  ( .D(\pe4/aot [10]), .CK(clk), .RDN(n28541), 
        .Q(ao4[10]) );
  DRNQHSV1 \pe4/pe15/q_reg[6]  ( .D(\pe4/aot [11]), .CK(clk), .RDN(n28486), 
        .Q(ao4[11]) );
  DRNQHSV1 \pe4/pe15/q_reg[5]  ( .D(\pe4/aot [12]), .CK(clk), .RDN(n28539), 
        .Q(ao4[12]) );
  DRNQHSV1 \pe4/pe15/q_reg[4]  ( .D(\pe4/aot [13]), .CK(clk), .RDN(n28459), 
        .Q(ao4[13]) );
  DRNQHSV1 \pe4/pe15/q_reg[2]  ( .D(n28433), .CK(clk), .RDN(n28490), .Q(
        ao4[15]) );
  DRNQHSV1 \pe4/pe16/q_reg[16]  ( .D(n28624), .CK(clk), .RDN(n28501), .Q(
        go4[1]) );
  DRNQHSV1 \pe4/pe16/q_reg[15]  ( .D(n28591), .CK(clk), .RDN(n28504), .Q(
        go4[2]) );
  DRNQHSV1 \pe4/pe16/q_reg[13]  ( .D(\pe4/got [4]), .CK(clk), .RDN(n28541), 
        .Q(go4[4]) );
  DRNQHSV1 \pe4/pe16/q_reg[12]  ( .D(\pe4/got [5]), .CK(clk), .RDN(n28604), 
        .Q(go4[5]) );
  DRNQHSV1 \pe4/pe16/q_reg[11]  ( .D(\pe4/got [6]), .CK(clk), .RDN(n28533), 
        .Q(go4[6]) );
  DRNQHSV1 \pe4/pe16/q_reg[10]  ( .D(n14000), .CK(clk), .RDN(n28500), .Q(
        go4[7]) );
  DRNQHSV1 \pe4/pe16/q_reg[9]  ( .D(\pe4/got [8]), .CK(clk), .RDN(n28519), .Q(
        go4[8]) );
  DRNQHSV1 \pe4/pe16/q_reg[8]  ( .D(\pe4/got [9]), .CK(clk), .RDN(n28524), .Q(
        go4[9]) );
  DRNQHSV1 \pe4/pe16/q_reg[7]  ( .D(\pe4/got [10]), .CK(clk), .RDN(n28545), 
        .Q(go4[10]) );
  DRNQHSV1 \pe4/pe16/q_reg[6]  ( .D(\pe4/got [11]), .CK(clk), .RDN(n28517), 
        .Q(go4[11]) );
  DRNQHSV1 \pe4/pe16/q_reg[5]  ( .D(n28428), .CK(clk), .RDN(n14021), .Q(
        go4[12]) );
  DRNQHSV1 \pe4/pe16/q_reg[4]  ( .D(n28463), .CK(clk), .RDN(n28528), .Q(
        go4[13]) );
  DRNQHSV1 \pe4/pe16/q_reg[3]  ( .D(n28612), .CK(clk), .RDN(n28575), .Q(
        go4[14]) );
  DRNQHSV1 \pe4/pe16/q_reg[2]  ( .D(n28592), .CK(clk), .RDN(n28505), .Q(
        go4[15]) );
  DRNQHSV1 \pe4/pe16/q_reg[1]  ( .D(\pe4/got [16]), .CK(clk), .RDN(n28539), 
        .Q(go4[16]) );
  DRNQHSV2 \pe4/pe17/q_reg[14]  ( .D(\pe4/poht [14]), .CK(clk), .RDN(n28545), 
        .Q(poh4[14]) );
  DRNQHSV1 \pe4/pe17/q_reg[13]  ( .D(\pe4/poht [13]), .CK(clk), .RDN(n28506), 
        .Q(poh4[13]) );
  DRNQHSV1 \pe4/pe17/q_reg[10]  ( .D(\pe4/poht [10]), .CK(clk), .RDN(n28546), 
        .Q(poh4[10]) );
  DRNQHSV1 \pe4/pe17/q_reg[9]  ( .D(\pe4/poht [9]), .CK(clk), .RDN(n28491), 
        .Q(poh4[9]) );
  DRNQHSV2 \pe4/pe17/q_reg[8]  ( .D(\pe4/poht [8]), .CK(clk), .RDN(n28550), 
        .Q(poh4[8]) );
  DRNQHSV1 \pe4/pe17/q_reg[6]  ( .D(\pe4/poht [6]), .CK(clk), .RDN(n28453), 
        .Q(poh4[6]) );
  DRNQHSV1 \pe4/pe17/q_reg[5]  ( .D(\pe4/poht [5]), .CK(clk), .RDN(n28576), 
        .Q(poh4[5]) );
  DRNQHSV1 \pe4/pe17/q_reg[4]  ( .D(\pe4/poht [4]), .CK(clk), .RDN(n28549), 
        .Q(poh4[4]) );
  DRNQHSV1 \pe4/pe17/q_reg[3]  ( .D(\pe4/poht [3]), .CK(clk), .RDN(n28550), 
        .Q(poh4[3]) );
  DRNQHSV1 \pe4/pe17/q_reg[1]  ( .D(\pe4/poht [1]), .CK(clk), .RDN(n28499), 
        .Q(poh4[1]) );
  DRNQHSV1 \pe5/pe15/q_reg[16]  ( .D(\pe5/aot [1]), .CK(clk), .RDN(n28577), 
        .Q(ao5[1]) );
  DRNQHSV1 \pe5/pe15/q_reg[15]  ( .D(\pe5/aot [2]), .CK(clk), .RDN(n28604), 
        .Q(ao5[2]) );
  DRNQHSV1 \pe5/pe15/q_reg[14]  ( .D(\pe5/aot [3]), .CK(clk), .RDN(n28505), 
        .Q(ao5[3]) );
  DRNQHSV1 \pe5/pe15/q_reg[13]  ( .D(\pe5/aot [4]), .CK(clk), .RDN(n28491), 
        .Q(ao5[4]) );
  DRNQHSV1 \pe5/pe15/q_reg[12]  ( .D(\pe5/aot [5]), .CK(clk), .RDN(n28551), 
        .Q(ao5[5]) );
  DRNQHSV1 \pe5/pe15/q_reg[11]  ( .D(\pe5/aot [6]), .CK(clk), .RDN(n28575), 
        .Q(ao5[6]) );
  DRNQHSV1 \pe5/pe15/q_reg[10]  ( .D(\pe5/aot [7]), .CK(clk), .RDN(n28535), 
        .Q(ao5[7]) );
  DRNQHSV1 \pe5/pe15/q_reg[9]  ( .D(\pe5/aot [8]), .CK(clk), .RDN(n28513), .Q(
        ao5[8]) );
  DRNQHSV1 \pe5/pe15/q_reg[8]  ( .D(\pe5/aot [9]), .CK(clk), .RDN(n28544), .Q(
        ao5[9]) );
  DRNQHSV1 \pe5/pe15/q_reg[7]  ( .D(\pe5/aot [10]), .CK(clk), .RDN(n28507), 
        .Q(ao5[10]) );
  DRNQHSV1 \pe5/pe15/q_reg[6]  ( .D(\pe5/aot [11]), .CK(clk), .RDN(n28525), 
        .Q(ao5[11]) );
  DRNQHSV1 \pe5/pe15/q_reg[5]  ( .D(\pe5/aot [12]), .CK(clk), .RDN(n28539), 
        .Q(ao5[12]) );
  DRNQHSV1 \pe5/pe15/q_reg[4]  ( .D(n14019), .CK(clk), .RDN(n28501), .Q(
        ao5[13]) );
  DRNQHSV1 \pe5/pe15/q_reg[3]  ( .D(\pe5/aot [14]), .CK(clk), .RDN(n28497), 
        .Q(ao5[14]) );
  DRNQHSV1 \pe5/pe15/q_reg[2]  ( .D(n14031), .CK(clk), .RDN(n28575), .Q(
        ao5[15]) );
  DRNQHSV1 \pe5/pe15/q_reg[1]  ( .D(n21488), .CK(clk), .RDN(n28549), .Q(
        ao5[16]) );
  DRNQHSV1 \pe5/pe16/q_reg[16]  ( .D(n28640), .CK(clk), .RDN(n28448), .Q(
        go5[1]) );
  DRNQHSV1 \pe5/pe16/q_reg[15]  ( .D(\pe5/got [2]), .CK(clk), .RDN(n28504), 
        .Q(go5[2]) );
  DRNQHSV1 \pe5/pe16/q_reg[14]  ( .D(\pe5/got [3]), .CK(clk), .RDN(n28550), 
        .Q(go5[3]) );
  DRNQHSV1 \pe5/pe16/q_reg[13]  ( .D(n13999), .CK(clk), .RDN(n28458), .Q(
        go5[4]) );
  DRNQHSV1 \pe5/pe16/q_reg[12]  ( .D(n14072), .CK(clk), .RDN(n28560), .Q(
        go5[5]) );
  DRNQHSV1 \pe5/pe16/q_reg[11]  ( .D(n28647), .CK(clk), .RDN(n28484), .Q(
        go5[6]) );
  DRNQHSV1 \pe5/pe16/q_reg[10]  ( .D(n28645), .CK(clk), .RDN(n28488), .Q(
        go5[7]) );
  DRNQHSV1 \pe5/pe16/q_reg[9]  ( .D(n28632), .CK(clk), .RDN(n28567), .Q(go5[8]) );
  DRNQHSV1 \pe5/pe16/q_reg[8]  ( .D(n14071), .CK(clk), .RDN(n28569), .Q(go5[9]) );
  DRNQHSV1 \pe5/pe16/q_reg[7]  ( .D(\pe5/got [10]), .CK(clk), .RDN(n28604), 
        .Q(go5[10]) );
  DRNQHSV1 \pe5/pe16/q_reg[6]  ( .D(\pe5/got [11]), .CK(clk), .RDN(n28477), 
        .Q(go5[11]) );
  DRNQHSV1 \pe5/pe16/q_reg[5]  ( .D(\pe5/got [12]), .CK(clk), .RDN(n28605), 
        .Q(go5[12]) );
  DRNQHSV1 \pe5/pe16/q_reg[4]  ( .D(n14852), .CK(clk), .RDN(n28476), .Q(
        go5[13]) );
  DRNQHSV1 \pe5/pe16/q_reg[3]  ( .D(\pe5/got [14]), .CK(clk), .RDN(n28549), 
        .Q(go5[14]) );
  DRNQHSV1 \pe5/pe16/q_reg[2]  ( .D(\pe5/got [15]), .CK(clk), .RDN(n28543), 
        .Q(go5[15]) );
  DRNQHSV1 \pe5/pe16/q_reg[1]  ( .D(\pe5/got [16]), .CK(clk), .RDN(n28493), 
        .Q(go5[16]) );
  DRNQHSV2 \pe5/pe17/q_reg[11]  ( .D(\pe5/poht [11]), .CK(clk), .RDN(n28534), 
        .Q(poh5[11]) );
  DRNQHSV2 \pe5/pe17/q_reg[10]  ( .D(\pe5/poht [10]), .CK(clk), .RDN(n28558), 
        .Q(poh5[10]) );
  DRNQHSV2 \pe5/pe17/q_reg[5]  ( .D(\pe5/poht [5]), .CK(clk), .RDN(n28559), 
        .Q(poh5[5]) );
  DRNQHSV2 \pe5/pe17/q_reg[3]  ( .D(\pe5/poht [3]), .CK(clk), .RDN(n28445), 
        .Q(poh5[3]) );
  DRNQHSV1 \pe6/pe15/q_reg[16]  ( .D(\pe6/aot [1]), .CK(clk), .RDN(n28562), 
        .Q(ao6[1]) );
  DRNQHSV1 \pe6/pe15/q_reg[15]  ( .D(\pe6/aot [2]), .CK(clk), .RDN(n28477), 
        .Q(ao6[2]) );
  DRNQHSV1 \pe6/pe15/q_reg[14]  ( .D(\pe6/aot [3]), .CK(clk), .RDN(n28520), 
        .Q(ao6[3]) );
  DRNQHSV1 \pe6/pe15/q_reg[13]  ( .D(\pe6/aot [4]), .CK(clk), .RDN(n14021), 
        .Q(ao6[4]) );
  DRNQHSV1 \pe6/pe15/q_reg[12]  ( .D(\pe6/aot [5]), .CK(clk), .RDN(n28535), 
        .Q(ao6[5]) );
  DRNQHSV1 \pe6/pe15/q_reg[11]  ( .D(\pe6/aot [6]), .CK(clk), .RDN(n28444), 
        .Q(ao6[6]) );
  DRNQHSV1 \pe6/pe15/q_reg[10]  ( .D(\pe6/aot [7]), .CK(clk), .RDN(n14023), 
        .Q(ao6[7]) );
  DRNQHSV1 \pe6/pe15/q_reg[9]  ( .D(\pe6/aot [8]), .CK(clk), .RDN(n28596), .Q(
        ao6[8]) );
  DRNQHSV1 \pe6/pe15/q_reg[8]  ( .D(\pe6/aot [9]), .CK(clk), .RDN(n28476), .Q(
        ao6[9]) );
  DRNQHSV1 \pe6/pe15/q_reg[7]  ( .D(\pe6/aot [10]), .CK(clk), .RDN(n28562), 
        .Q(ao6[10]) );
  DRNQHSV1 \pe6/pe15/q_reg[6]  ( .D(\pe6/aot [11]), .CK(clk), .RDN(n28497), 
        .Q(ao6[11]) );
  DRNQHSV1 \pe6/pe15/q_reg[5]  ( .D(\pe6/aot [12]), .CK(clk), .RDN(n28440), 
        .Q(ao6[12]) );
  DRNQHSV1 \pe6/pe15/q_reg[4]  ( .D(\pe6/aot [13]), .CK(clk), .RDN(n28559), 
        .Q(ao6[13]) );
  DRNQHSV1 \pe6/pe15/q_reg[3]  ( .D(\pe6/aot [14]), .CK(clk), .RDN(n28562), 
        .Q(ao6[14]) );
  DRNQHSV1 \pe6/pe15/q_reg[2]  ( .D(n28680), .CK(clk), .RDN(n28452), .Q(
        ao6[15]) );
  DRNQHSV1 \pe6/pe15/q_reg[1]  ( .D(n28681), .CK(clk), .RDN(n28607), .Q(
        ao6[16]) );
  DRNQHSV1 \pe6/pe16/q_reg[16]  ( .D(n28608), .CK(clk), .RDN(n28503), .Q(
        go6[1]) );
  DRNQHSV1 \pe6/pe16/q_reg[15]  ( .D(\pe6/got [2]), .CK(clk), .RDN(n28601), 
        .Q(go6[2]) );
  DRNQHSV1 \pe6/pe16/q_reg[14]  ( .D(\pe6/got [3]), .CK(clk), .RDN(n28547), 
        .Q(go6[3]) );
  DRNQHSV1 \pe6/pe16/q_reg[13]  ( .D(\pe6/got [4]), .CK(clk), .RDN(n28564), 
        .Q(go6[4]) );
  DRNQHSV1 \pe6/pe16/q_reg[12]  ( .D(\pe6/got [5]), .CK(clk), .RDN(n28484), 
        .Q(go6[5]) );
  DRNQHSV1 \pe6/pe16/q_reg[11]  ( .D(\pe6/got [6]), .CK(clk), .RDN(n28527), 
        .Q(go6[6]) );
  DRNQHSV1 \pe6/pe16/q_reg[10]  ( .D(\pe6/got [7]), .CK(clk), .RDN(n28555), 
        .Q(go6[7]) );
  DRNQHSV1 \pe6/pe16/q_reg[9]  ( .D(\pe6/got [8]), .CK(clk), .RDN(n28555), .Q(
        go6[8]) );
  DRNQHSV1 \pe6/pe16/q_reg[8]  ( .D(\pe6/got [9]), .CK(clk), .RDN(n28509), .Q(
        go6[9]) );
  DRNQHSV1 \pe6/pe16/q_reg[7]  ( .D(\pe6/got [10]), .CK(clk), .RDN(n28483), 
        .Q(go6[10]) );
  DRNQHSV1 \pe6/pe16/q_reg[6]  ( .D(n28586), .CK(clk), .RDN(n28487), .Q(
        go6[11]) );
  DRNQHSV1 \pe6/pe16/q_reg[5]  ( .D(n28593), .CK(clk), .RDN(n28542), .Q(
        go6[12]) );
  DRNQHSV1 \pe6/pe16/q_reg[4]  ( .D(n14236), .CK(clk), .RDN(n28552), .Q(
        go6[13]) );
  DRNQHSV1 \pe6/pe16/q_reg[3]  ( .D(n28686), .CK(clk), .RDN(n28520), .Q(
        go6[14]) );
  DRNQHSV1 \pe6/pe16/q_reg[1]  ( .D(n28472), .CK(clk), .RDN(n28499), .Q(
        go6[16]) );
  DRNQHSV2 \pe6/pe17/q_reg[11]  ( .D(\pe6/poht [11]), .CK(clk), .RDN(n28602), 
        .Q(poh6[11]) );
  DRNQHSV2 \pe6/pe17/q_reg[9]  ( .D(\pe6/poht [9]), .CK(clk), .RDN(n28510), 
        .Q(poh6[9]) );
  DRNQHSV1 \pe6/pe17/q_reg[6]  ( .D(\pe6/poht [6]), .CK(clk), .RDN(n28506), 
        .Q(poh6[6]) );
  DRNQHSV2 \pe6/pe17/q_reg[4]  ( .D(\pe6/poht [4]), .CK(clk), .RDN(n28507), 
        .Q(poh6[4]) );
  DRNQHSV2 \pe6/pe17/q_reg[3]  ( .D(\pe6/poht [3]), .CK(clk), .RDN(n28509), 
        .Q(poh6[3]) );
  DRNQHSV1 \pe6/pe17/q_reg[2]  ( .D(\pe6/poht [2]), .CK(clk), .RDN(n28444), 
        .Q(poh6[2]) );
  DRNQHSV1 \pe7/pe15/q_reg[16]  ( .D(\pe7/aot [1]), .CK(clk), .RDN(n28546), 
        .Q(ao7[1]) );
  DRNQHSV1 \pe7/pe15/q_reg[15]  ( .D(\pe7/aot [2]), .CK(clk), .RDN(n28537), 
        .Q(ao7[2]) );
  DRNQHSV1 \pe7/pe15/q_reg[14]  ( .D(\pe7/aot [3]), .CK(clk), .RDN(n28509), 
        .Q(ao7[3]) );
  DRNQHSV1 \pe7/pe15/q_reg[13]  ( .D(\pe7/aot [4]), .CK(clk), .RDN(n28504), 
        .Q(ao7[4]) );
  DRNQHSV1 \pe7/pe15/q_reg[12]  ( .D(\pe7/aot [5]), .CK(clk), .RDN(n28534), 
        .Q(ao7[5]) );
  DRNQHSV1 \pe7/pe15/q_reg[11]  ( .D(\pe7/aot [6]), .CK(clk), .RDN(n28495), 
        .Q(ao7[6]) );
  DRNQHSV1 \pe7/pe15/q_reg[10]  ( .D(\pe7/aot [7]), .CK(clk), .RDN(n28547), 
        .Q(ao7[7]) );
  DRNQHSV1 \pe7/pe15/q_reg[9]  ( .D(\pe7/aot [8]), .CK(clk), .RDN(n28551), .Q(
        ao7[8]) );
  DRNQHSV1 \pe7/pe15/q_reg[8]  ( .D(\pe7/aot [9]), .CK(clk), .RDN(n28507), .Q(
        ao7[9]) );
  DRNQHSV1 \pe7/pe15/q_reg[7]  ( .D(\pe7/aot [10]), .CK(clk), .RDN(n28558), 
        .Q(ao7[10]) );
  DRNQHSV1 \pe7/pe15/q_reg[6]  ( .D(\pe7/aot [11]), .CK(clk), .RDN(n28546), 
        .Q(ao7[11]) );
  DRNQHSV1 \pe7/pe15/q_reg[5]  ( .D(\pe7/aot [12]), .CK(clk), .RDN(n28487), 
        .Q(ao7[12]) );
  DRNQHSV1 \pe7/pe15/q_reg[4]  ( .D(n14050), .CK(clk), .RDN(n28486), .Q(
        ao7[13]) );
  DRNQHSV1 \pe7/pe15/q_reg[3]  ( .D(\pe7/aot [14]), .CK(clk), .RDN(n14023), 
        .Q(ao7[14]) );
  DRNQHSV1 \pe7/pe15/q_reg[2]  ( .D(\pe7/aot [15]), .CK(clk), .RDN(n28575), 
        .Q(ao7[15]) );
  DRNQHSV1 \pe7/pe15/q_reg[1]  ( .D(n14078), .CK(clk), .RDN(n28575), .Q(
        ao7[16]) );
  DRNQHSV1 \pe7/pe16/q_reg[16]  ( .D(\pe7/got [1]), .CK(clk), .RDN(n28548), 
        .Q(go7[1]) );
  DRNQHSV1 \pe7/pe16/q_reg[15]  ( .D(\pe7/got [2]), .CK(clk), .RDN(n28551), 
        .Q(go7[2]) );
  DRNQHSV1 \pe7/pe16/q_reg[14]  ( .D(\pe7/got [3]), .CK(clk), .RDN(n28512), 
        .Q(go7[3]) );
  DRNQHSV1 \pe7/pe16/q_reg[13]  ( .D(\pe7/got [4]), .CK(clk), .RDN(n28506), 
        .Q(go7[4]) );
  DRNQHSV1 \pe7/pe16/q_reg[12]  ( .D(\pe7/got [5]), .CK(clk), .RDN(n28548), 
        .Q(go7[5]) );
  DRNQHSV1 \pe7/pe16/q_reg[11]  ( .D(\pe7/got [6]), .CK(clk), .RDN(n28511), 
        .Q(go7[6]) );
  DRNQHSV1 \pe7/pe16/q_reg[10]  ( .D(\pe7/got [7]), .CK(clk), .RDN(n28439), 
        .Q(go7[7]) );
  DRNQHSV1 \pe7/pe16/q_reg[9]  ( .D(\pe7/got [8]), .CK(clk), .RDN(n28573), .Q(
        go7[8]) );
  DRNQHSV1 \pe7/pe16/q_reg[8]  ( .D(\pe7/got [9]), .CK(clk), .RDN(n28548), .Q(
        go7[9]) );
  DRNQHSV1 \pe7/pe16/q_reg[7]  ( .D(n24214), .CK(clk), .RDN(n28532), .Q(
        go7[10]) );
  DRNQHSV1 \pe7/pe16/q_reg[6]  ( .D(n14022), .CK(clk), .RDN(n28499), .Q(
        go7[11]) );
  DRNQHSV1 \pe7/pe16/q_reg[5]  ( .D(\pe7/got [12]), .CK(clk), .RDN(n28511), 
        .Q(go7[12]) );
  DRNQHSV1 \pe7/pe16/q_reg[4]  ( .D(\pe7/got [13]), .CK(clk), .RDN(n28548), 
        .Q(go7[13]) );
  DRNQHSV1 \pe7/pe16/q_reg[3]  ( .D(n24271), .CK(clk), .RDN(n28560), .Q(
        go7[14]) );
  DRNQHSV1 \pe7/pe16/q_reg[2]  ( .D(n28816), .CK(clk), .RDN(n14023), .Q(
        go7[15]) );
  DRNQHSV1 \pe7/pe16/q_reg[1]  ( .D(n28610), .CK(clk), .RDN(n28554), .Q(
        go7[16]) );
  DRNQHSV1 \pe7/pe17/q_reg[15]  ( .D(\pe7/poht [15]), .CK(clk), .RDN(n28452), 
        .Q(poh7[15]) );
  DRNQHSV2 \pe7/pe17/q_reg[11]  ( .D(\pe7/poht [11]), .CK(clk), .RDN(n28515), 
        .Q(poh7[11]) );
  DRNQHSV2 \pe7/pe17/q_reg[9]  ( .D(\pe7/poht [9]), .CK(clk), .RDN(n28596), 
        .Q(poh7[9]) );
  DRNQHSV2 \pe7/pe17/q_reg[8]  ( .D(\pe7/poht [8]), .CK(clk), .RDN(n28534), 
        .Q(poh7[8]) );
  DRNQHSV2 \pe7/pe17/q_reg[7]  ( .D(\pe7/poht [7]), .CK(clk), .RDN(n28477), 
        .Q(poh7[7]) );
  DRNQHSV2 \pe7/pe17/q_reg[6]  ( .D(\pe7/poht [6]), .CK(clk), .RDN(n28448), 
        .Q(poh7[6]) );
  DRNQHSV2 \pe7/pe17/q_reg[5]  ( .D(\pe7/poht [5]), .CK(clk), .RDN(n28517), 
        .Q(poh7[5]) );
  DRNQHSV2 \pe7/pe17/q_reg[4]  ( .D(\pe7/poht [4]), .CK(clk), .RDN(n28556), 
        .Q(poh7[4]) );
  DRNQHSV2 \pe7/pe17/q_reg[3]  ( .D(\pe7/poht [3]), .CK(clk), .RDN(n28490), 
        .Q(poh7[3]) );
  DRNQHSV2 \pe7/pe17/q_reg[2]  ( .D(\pe7/poht [2]), .CK(clk), .RDN(n28571), 
        .Q(poh7[2]) );
  DRNQHSV2 \pe7/pe17/q_reg[1]  ( .D(\pe7/poht [1]), .CK(clk), .RDN(n28532), 
        .Q(poh7[1]) );
  DRNQHSV1 \pe8/pe15/q_reg[16]  ( .D(\pe8/aot [1]), .CK(clk), .RDN(n28487), 
        .Q(ao8[1]) );
  DRNQHSV1 \pe8/pe15/q_reg[15]  ( .D(\pe8/aot [2]), .CK(clk), .RDN(n28517), 
        .Q(ao8[2]) );
  DRNQHSV1 \pe8/pe15/q_reg[14]  ( .D(\pe8/aot [3]), .CK(clk), .RDN(n28502), 
        .Q(ao8[3]) );
  DRNQHSV1 \pe8/pe15/q_reg[13]  ( .D(\pe8/aot [4]), .CK(clk), .RDN(n28576), 
        .Q(ao8[4]) );
  DRNQHSV1 \pe8/pe15/q_reg[12]  ( .D(\pe8/aot [5]), .CK(clk), .RDN(n28482), 
        .Q(ao8[5]) );
  DRNQHSV1 \pe8/pe15/q_reg[11]  ( .D(\pe8/aot [6]), .CK(clk), .RDN(n28536), 
        .Q(ao8[6]) );
  DRNQHSV1 \pe8/pe15/q_reg[10]  ( .D(\pe8/aot [7]), .CK(clk), .RDN(n28545), 
        .Q(ao8[7]) );
  DRNQHSV1 \pe8/pe15/q_reg[9]  ( .D(\pe8/aot [8]), .CK(clk), .RDN(n28512), .Q(
        ao8[8]) );
  DRNQHSV1 \pe8/pe15/q_reg[8]  ( .D(\pe8/aot [9]), .CK(clk), .RDN(n28500), .Q(
        ao8[9]) );
  DRNQHSV1 \pe8/pe15/q_reg[7]  ( .D(\pe8/aot [10]), .CK(clk), .RDN(n28530), 
        .Q(ao8[10]) );
  DRNQHSV1 \pe8/pe15/q_reg[6]  ( .D(\pe8/aot [11]), .CK(clk), .RDN(n28450), 
        .Q(ao8[11]) );
  DRNQHSV1 \pe8/pe15/q_reg[5]  ( .D(\pe8/aot [12]), .CK(clk), .RDN(n28607), 
        .Q(ao8[12]) );
  DRNQHSV1 \pe8/pe15/q_reg[4]  ( .D(\pe8/aot [13]), .CK(clk), .RDN(n28527), 
        .Q(ao8[13]) );
  DRNQHSV1 \pe8/pe15/q_reg[3]  ( .D(\pe8/aot [14]), .CK(clk), .RDN(n28459), 
        .Q(ao8[14]) );
  DRNQHSV1 \pe8/pe15/q_reg[2]  ( .D(\pe8/aot [15]), .CK(clk), .RDN(n28515), 
        .Q(ao8[15]) );
  DRNQHSV1 \pe8/pe15/q_reg[1]  ( .D(n28627), .CK(clk), .RDN(n28451), .Q(
        ao8[16]) );
  DRNQHSV1 \pe8/pe16/q_reg[16]  ( .D(\pe8/got [1]), .CK(clk), .RDN(n28447), 
        .Q(go8[1]) );
  DRNQHSV1 \pe8/pe16/q_reg[15]  ( .D(\pe8/got [2]), .CK(clk), .RDN(n28565), 
        .Q(go8[2]) );
  DRNQHSV1 \pe8/pe16/q_reg[14]  ( .D(\pe8/got [3]), .CK(clk), .RDN(n28548), 
        .Q(go8[3]) );
  DRNQHSV1 \pe8/pe16/q_reg[13]  ( .D(n25577), .CK(clk), .RDN(n28542), .Q(
        go8[4]) );
  DRNQHSV1 \pe8/pe16/q_reg[12]  ( .D(\pe8/got [5]), .CK(clk), .RDN(n28566), 
        .Q(go8[5]) );
  DRNQHSV1 \pe8/pe16/q_reg[11]  ( .D(\pe8/got [6]), .CK(clk), .RDN(n28569), 
        .Q(go8[6]) );
  DRNQHSV1 \pe8/pe16/q_reg[10]  ( .D(n14068), .CK(clk), .RDN(n28550), .Q(
        go8[7]) );
  DRNQHSV1 \pe8/pe16/q_reg[8]  ( .D(\pe8/got [9]), .CK(clk), .RDN(n28514), .Q(
        go8[9]) );
  DRNQHSV1 \pe8/pe16/q_reg[7]  ( .D(\pe8/got [10]), .CK(clk), .RDN(n28569), 
        .Q(go8[10]) );
  DRNQHSV1 \pe8/pe16/q_reg[6]  ( .D(n28618), .CK(clk), .RDN(n28505), .Q(
        go8[11]) );
  DRNQHSV1 \pe8/pe16/q_reg[5]  ( .D(\pe8/got [12]), .CK(clk), .RDN(n28595), 
        .Q(go8[12]) );
  DRNQHSV1 \pe8/pe16/q_reg[4]  ( .D(\pe8/got [13]), .CK(clk), .RDN(n28562), 
        .Q(go8[13]) );
  DRNQHSV1 \pe8/pe16/q_reg[3]  ( .D(n28599), .CK(clk), .RDN(n28558), .Q(
        go8[14]) );
  DRNQHSV1 \pe8/pe16/q_reg[2]  ( .D(n28625), .CK(clk), .RDN(n28459), .Q(
        go8[15]) );
  DRNQHSV2 \pe8/pe17/q_reg[3]  ( .D(\pe8/poht [3]), .CK(clk), .RDN(n28577), 
        .Q(poh8[3]) );
  DRNQHSV1 \pe9/pe15/q_reg[16]  ( .D(\pe9/aot [1]), .CK(clk), .RDN(n28502), 
        .Q(ao9[1]) );
  DRNQHSV1 \pe9/pe15/q_reg[15]  ( .D(\pe9/aot [2]), .CK(clk), .RDN(n28496), 
        .Q(ao9[2]) );
  DRNQHSV1 \pe9/pe15/q_reg[14]  ( .D(\pe9/aot [3]), .CK(clk), .RDN(n28442), 
        .Q(ao9[3]) );
  DRNQHSV1 \pe9/pe15/q_reg[13]  ( .D(\pe9/aot [4]), .CK(clk), .RDN(n28596), 
        .Q(ao9[4]) );
  DRNQHSV1 \pe9/pe15/q_reg[12]  ( .D(\pe9/aot [5]), .CK(clk), .RDN(n28524), 
        .Q(ao9[5]) );
  DRNQHSV1 \pe9/pe15/q_reg[11]  ( .D(\pe9/aot [6]), .CK(clk), .RDN(n28540), 
        .Q(ao9[6]) );
  DRNQHSV1 \pe9/pe15/q_reg[10]  ( .D(\pe9/aot [7]), .CK(clk), .RDN(n28604), 
        .Q(ao9[7]) );
  DRNQHSV1 \pe9/pe15/q_reg[9]  ( .D(\pe9/aot [8]), .CK(clk), .RDN(n28574), .Q(
        ao9[8]) );
  DRNQHSV1 \pe9/pe15/q_reg[8]  ( .D(\pe9/aot [9]), .CK(clk), .RDN(n28518), .Q(
        ao9[9]) );
  DRNQHSV1 \pe9/pe15/q_reg[7]  ( .D(\pe9/aot [10]), .CK(clk), .RDN(n28566), 
        .Q(ao9[10]) );
  DRNQHSV1 \pe9/pe15/q_reg[6]  ( .D(\pe9/aot [11]), .CK(clk), .RDN(n28532), 
        .Q(ao9[11]) );
  DRNQHSV1 \pe9/pe15/q_reg[5]  ( .D(\pe9/aot [12]), .CK(clk), .RDN(n28442), 
        .Q(ao9[12]) );
  DRNQHSV1 \pe9/pe15/q_reg[4]  ( .D(\pe9/aot [13]), .CK(clk), .RDN(n28441), 
        .Q(ao9[13]) );
  DRNQHSV1 \pe9/pe15/q_reg[3]  ( .D(\pe9/aot [14]), .CK(clk), .RDN(n28519), 
        .Q(ao9[14]) );
  DRNQHSV1 \pe9/pe15/q_reg[2]  ( .D(n14079), .CK(clk), .RDN(n28451), .Q(
        ao9[15]) );
  DRNQHSV1 \pe9/pe15/q_reg[1]  ( .D(n12618), .CK(clk), .RDN(n28566), .Q(
        ao9[16]) );
  DRNQHSV1 \pe9/pe16/q_reg[16]  ( .D(n28658), .CK(clk), .RDN(n28453), .Q(
        go9[1]) );
  DRNQHSV1 \pe9/pe16/q_reg[15]  ( .D(n28654), .CK(clk), .RDN(n28517), .Q(
        go9[2]) );
  DRNQHSV1 \pe9/pe16/q_reg[14]  ( .D(n28405), .CK(clk), .RDN(n28595), .Q(
        go9[3]) );
  DRNQHSV1 \pe9/pe16/q_reg[13]  ( .D(\pe9/got [4]), .CK(clk), .RDN(n28444), 
        .Q(go9[4]) );
  DRNQHSV1 \pe9/pe16/q_reg[12]  ( .D(n28643), .CK(clk), .RDN(n28570), .Q(
        go9[5]) );
  DRNQHSV1 \pe9/pe16/q_reg[11]  ( .D(\pe9/got [6]), .CK(clk), .RDN(n28561), 
        .Q(go9[6]) );
  DRNQHSV1 \pe9/pe16/q_reg[10]  ( .D(\pe9/got [7]), .CK(clk), .RDN(n28516), 
        .Q(go9[7]) );
  DRNQHSV1 \pe9/pe16/q_reg[9]  ( .D(\pe9/got [8]), .CK(clk), .RDN(n28489), .Q(
        go9[8]) );
  DRNQHSV1 \pe9/pe16/q_reg[8]  ( .D(\pe9/got [9]), .CK(clk), .RDN(n28443), .Q(
        go9[9]) );
  DRNQHSV1 \pe9/pe16/q_reg[7]  ( .D(\pe9/got [10]), .CK(clk), .RDN(n28535), 
        .Q(go9[10]) );
  DRNQHSV1 \pe9/pe16/q_reg[5]  ( .D(\pe9/got [12]), .CK(clk), .RDN(n28449), 
        .Q(go9[12]) );
  DRNQHSV1 \pe9/pe16/q_reg[4]  ( .D(n18029), .CK(clk), .RDN(n28492), .Q(
        go9[13]) );
  DRNQHSV1 \pe9/pe16/q_reg[2]  ( .D(\pe9/got [15]), .CK(clk), .RDN(n28596), 
        .Q(go9[15]) );
  DRNQHSV1 \pe10/pe15/q_reg[16]  ( .D(\pe10/aot [1]), .CK(clk), .RDN(n28518), 
        .Q(ao10[1]) );
  DRNQHSV1 \pe10/pe15/q_reg[15]  ( .D(\pe10/aot [2]), .CK(clk), .RDN(n28449), 
        .Q(ao10[2]) );
  DRNQHSV1 \pe10/pe15/q_reg[14]  ( .D(\pe10/aot [3]), .CK(clk), .RDN(n28452), 
        .Q(ao10[3]) );
  DRNQHSV1 \pe10/pe15/q_reg[13]  ( .D(\pe10/aot [4]), .CK(clk), .RDN(n28553), 
        .Q(ao10[4]) );
  DRNQHSV1 \pe10/pe15/q_reg[12]  ( .D(\pe10/aot [5]), .CK(clk), .RDN(n28535), 
        .Q(ao10[5]) );
  DRNQHSV1 \pe10/pe15/q_reg[11]  ( .D(\pe10/aot [6]), .CK(clk), .RDN(n28516), 
        .Q(ao10[6]) );
  DRNQHSV1 \pe10/pe15/q_reg[10]  ( .D(\pe10/aot [7]), .CK(clk), .RDN(n28547), 
        .Q(ao10[7]) );
  DRNQHSV1 \pe10/pe15/q_reg[9]  ( .D(\pe10/aot [8]), .CK(clk), .RDN(n28513), 
        .Q(ao10[8]) );
  DRNQHSV1 \pe10/pe15/q_reg[8]  ( .D(\pe10/aot [9]), .CK(clk), .RDN(n28521), 
        .Q(ao10[9]) );
  DRNQHSV1 \pe10/pe15/q_reg[7]  ( .D(\pe10/aot [10]), .CK(clk), .RDN(n28524), 
        .Q(ao10[10]) );
  DRNQHSV1 \pe10/pe15/q_reg[6]  ( .D(\pe10/aot [11]), .CK(clk), .RDN(n28491), 
        .Q(ao10[11]) );
  DRNQHSV1 \pe10/pe15/q_reg[5]  ( .D(\pe10/aot [12]), .CK(clk), .RDN(n28549), 
        .Q(ao10[12]) );
  DRNQHSV1 \pe10/pe15/q_reg[4]  ( .D(\pe10/aot [13]), .CK(clk), .RDN(n28509), 
        .Q(ao10[13]) );
  DRNQHSV1 \pe10/pe15/q_reg[3]  ( .D(\pe10/aot [14]), .CK(clk), .RDN(n28557), 
        .Q(ao10[14]) );
  DRNQHSV1 \pe10/pe15/q_reg[2]  ( .D(n16973), .CK(clk), .RDN(n28532), .Q(
        ao10[15]) );
  DRNQHSV1 \pe10/pe15/q_reg[1]  ( .D(n28424), .CK(clk), .RDN(n28459), .Q(
        ao10[16]) );
  DRNQHSV1 \pe10/pe16/q_reg[16]  ( .D(n28633), .CK(clk), .RDN(n28540), .Q(
        go10[1]) );
  DRNQHSV1 \pe10/pe16/q_reg[15]  ( .D(n28637), .CK(clk), .RDN(n28504), .Q(
        go10[2]) );
  DRNQHSV1 \pe10/pe16/q_reg[14]  ( .D(\pe10/got [3]), .CK(clk), .RDN(n28597), 
        .Q(go10[3]) );
  DRNQHSV1 \pe10/pe16/q_reg[13]  ( .D(\pe10/got [4]), .CK(clk), .RDN(n28547), 
        .Q(go10[4]) );
  DRNQHSV1 \pe10/pe16/q_reg[12]  ( .D(\pe10/got [5]), .CK(clk), .RDN(n28486), 
        .Q(go10[5]) );
  DRNQHSV1 \pe10/pe16/q_reg[11]  ( .D(\pe10/got [6]), .CK(clk), .RDN(n28597), 
        .Q(go10[6]) );
  DRNQHSV1 \pe10/pe16/q_reg[10]  ( .D(\pe10/got [7]), .CK(clk), .RDN(n28498), 
        .Q(go10[7]) );
  DRNQHSV1 \pe10/pe16/q_reg[9]  ( .D(n28642), .CK(clk), .RDN(n28542), .Q(
        go10[8]) );
  DRNQHSV1 \pe10/pe16/q_reg[8]  ( .D(\pe10/got [9]), .CK(clk), .RDN(n28537), 
        .Q(go10[9]) );
  DRNQHSV1 \pe10/pe16/q_reg[7]  ( .D(n28644), .CK(clk), .RDN(n28449), .Q(
        go10[10]) );
  DRNQHSV1 \pe10/pe16/q_reg[6]  ( .D(\pe10/got [11]), .CK(clk), .RDN(n28531), 
        .Q(go10[11]) );
  DRNQHSV1 \pe10/pe16/q_reg[5]  ( .D(n16876), .CK(clk), .RDN(n14023), .Q(
        go10[12]) );
  DRNQHSV1 \pe10/pe16/q_reg[4]  ( .D(n28479), .CK(clk), .RDN(n28533), .Q(
        go10[13]) );
  DRNQHSV1 \pe10/pe16/q_reg[3]  ( .D(\pe10/got [14]), .CK(clk), .RDN(n28560), 
        .Q(go10[14]) );
  DRNQHSV1 \pe10/pe16/q_reg[2]  ( .D(\pe10/got [15]), .CK(clk), .RDN(n28565), 
        .Q(go10[15]) );
  DRNQHSV1 \pe10/pe16/q_reg[1]  ( .D(n28810), .CK(clk), .RDN(n28570), .Q(
        go10[16]) );
  DRNQHSV2 \pe10/pe17/q_reg[11]  ( .D(\pe10/poht [11]), .CK(clk), .RDN(n28597), 
        .Q(poh10[11]) );
  DRNQHSV2 \pe10/pe17/q_reg[9]  ( .D(\pe10/poht [9]), .CK(clk), .RDN(n28533), 
        .Q(poh10[9]) );
  DRNQHSV2 \pe10/pe17/q_reg[8]  ( .D(\pe10/poht [8]), .CK(clk), .RDN(n28570), 
        .Q(poh10[8]) );
  DRNQHSV2 \pe10/pe17/q_reg[6]  ( .D(\pe10/poht [6]), .CK(clk), .RDN(n28551), 
        .Q(poh10[6]) );
  DRNQHSV2 \pe10/pe17/q_reg[5]  ( .D(\pe10/poht [5]), .CK(clk), .RDN(n28561), 
        .Q(poh10[5]) );
  DRNQHSV2 \pe10/pe17/q_reg[3]  ( .D(\pe10/poht [3]), .CK(clk), .RDN(n28540), 
        .Q(poh10[3]) );
  DRNQHSV2 \pe10/pe17/q_reg[1]  ( .D(\pe10/poht [1]), .CK(clk), .RDN(n28540), 
        .Q(poh10[1]) );
  DRNQHSV2 \pe11/pe3/q_reg[8]  ( .D(bo10[9]), .CK(clk), .RDN(n28514), .Q(
        bo11[9]) );
  DRNQHSV2 \pe11/pe3/q_reg[7]  ( .D(bo10[10]), .CK(clk), .RDN(n28449), .Q(
        bo11[10]) );
  DRNQHSV2 \pe11/pe3/q_reg[5]  ( .D(bo10[12]), .CK(clk), .RDN(n28513), .Q(
        bo11[12]) );
  DRNQHSV2 \pe11/pe17/q_reg[15]  ( .D(\pe11/poht [15]), .CK(clk), .RDN(n28525), 
        .Q(poh11[15]) );
  DRNQHSV2 \pe11/pe17/q_reg[13]  ( .D(\pe11/poht [13]), .CK(clk), .RDN(n28488), 
        .Q(poh11[13]) );
  DRNQHSV2 \pe11/pe17/q_reg[6]  ( .D(\pe11/poht [6]), .CK(clk), .RDN(n28489), 
        .Q(poh11[6]) );
  DRNQHSV2 \pe11/pe17/q_reg[4]  ( .D(\pe11/poht [4]), .CK(clk), .RDN(n28520), 
        .Q(poh11[4]) );
  DRNQHSV2 \pe11/pe17/q_reg[3]  ( .D(\pe11/poht [3]), .CK(clk), .RDN(n28550), 
        .Q(poh11[3]) );
  DRNQHSV2 \pe11/pe17/q_reg[2]  ( .D(\pe11/poht [2]), .CK(clk), .RDN(n28517), 
        .Q(poh11[2]) );
  DRNQHSV2 \pe11/pe17/q_reg[1]  ( .D(\pe11/poht [1]), .CK(clk), .RDN(n28489), 
        .Q(poh11[1]) );
  DRNQHSV1 \pe1/pe14/q_reg[14]  ( .D(n26909), .CK(clk), .RDN(n28522), .Q(
        \pe1/ti_7t [14]) );
  DRNQHSV1 \pe3/pe14/q_reg[14]  ( .D(n28801), .CK(clk), .RDN(n28534), .Q(
        \pe3/ti_7t [14]) );
  DRNQHSV1 \pe4/pe14/q_reg[15]  ( .D(n28461), .CK(clk), .RDN(n28514), .Q(
        \pe4/ti_7t [15]) );
  DRNQHSV1 \pe5/pe14/q_reg[13]  ( .D(n12517), .CK(clk), .RDN(n28572), .Q(
        \pe5/ti_7t [13]) );
  DRNQHSV1 \pe5/pe14/q_reg[15]  ( .D(n28436), .CK(clk), .RDN(n28493), .Q(
        \pe5/ti_7t [15]) );
  DRNQHSV2 \pe9/pe14/q_reg[14]  ( .D(\pe9/ti_7[14] ), .CK(clk), .RDN(n28535), 
        .Q(\pe9/ti_7t [14]) );
  DRNQHSV1 \pe10/pe14/q_reg[13]  ( .D(n22718), .CK(clk), .RDN(n28547), .Q(
        \pe10/ti_7t [13]) );
  DRNQHSV1 \pe11/pe14/q_reg[14]  ( .D(n28936), .CK(clk), .RDN(n28536), .Q(
        \pe11/ti_7t [14]) );
  DRNQHSV1 \pe11/pe14/q_reg[15]  ( .D(n28927), .CK(clk), .RDN(n28530), .Q(
        \pe11/ti_7t [15]) );
  DRNQHSV2 \pe3/pe3/q_reg[2]  ( .D(bo2[15]), .CK(clk), .RDN(n28525), .Q(
        bo3[15]) );
  DRNQHSV2 \pe4/pe3/q_reg[2]  ( .D(bo3[15]), .CK(clk), .RDN(n28482), .Q(
        bo4[15]) );
  DRNQHSV2 \pe6/pe3/q_reg[13]  ( .D(bo5[4]), .CK(clk), .RDN(n28502), .Q(bo6[4]) );
  DRNQHSV2 \pe7/pe3/q_reg[5]  ( .D(bo6[12]), .CK(clk), .RDN(n28531), .Q(
        bo7[12]) );
  DRNQHSV2 \pe11/pe17/q_reg[11]  ( .D(\pe11/poht [11]), .CK(clk), .RDN(n28551), 
        .Q(poh11[11]) );
  DRNQHSV2 \pe11/pe17/q_reg[9]  ( .D(\pe11/poht [9]), .CK(clk), .RDN(n28561), 
        .Q(poh11[9]) );
  DRNQHSV2 \pe1/pe3/q_reg[16]  ( .D(bi[1]), .CK(clk), .RDN(n28536), .Q(bo1[1])
         );
  DRNQHSV2 \pe1/pe3/q_reg[15]  ( .D(bi[2]), .CK(clk), .RDN(rst), .Q(bo1[2]) );
  DRNQHSV2 \pe1/pe3/q_reg[12]  ( .D(bi[5]), .CK(clk), .RDN(n28535), .Q(bo1[5])
         );
  DRNQHSV2 \pe1/pe3/q_reg[11]  ( .D(bi[6]), .CK(clk), .RDN(rst), .Q(bo1[6]) );
  DRNQHSV2 \pe1/pe3/q_reg[7]  ( .D(bi[10]), .CK(clk), .RDN(n28576), .Q(bo1[10]) );
  DRNQHSV2 \pe1/pe3/q_reg[5]  ( .D(bi[12]), .CK(clk), .RDN(n28442), .Q(bo1[12]) );
  DRNQHSV2 \pe1/pe3/q_reg[4]  ( .D(bi[13]), .CK(clk), .RDN(n28571), .Q(bo1[13]) );
  DRNQHSV2 \pe1/pe3/q_reg[3]  ( .D(bi[14]), .CK(clk), .RDN(n28507), .Q(bo1[14]) );
  DRNQHSV2 \pe2/pe3/q_reg[13]  ( .D(bo1[4]), .CK(clk), .RDN(n28490), .Q(bo2[4]) );
  DRNQHSV2 \pe4/pe3/q_reg[16]  ( .D(bo3[1]), .CK(clk), .RDN(n28500), .Q(bo4[1]) );
  DRNQHSV2 \pe4/pe3/q_reg[15]  ( .D(bo3[2]), .CK(clk), .RDN(n28576), .Q(bo4[2]) );
  DRNQHSV2 \pe4/pe3/q_reg[14]  ( .D(bo3[3]), .CK(clk), .RDN(n28539), .Q(bo4[3]) );
  DRNQHSV2 \pe4/pe3/q_reg[13]  ( .D(bo3[4]), .CK(clk), .RDN(n28488), .Q(bo4[4]) );
  DRNQHSV2 \pe4/pe3/q_reg[11]  ( .D(bo3[6]), .CK(clk), .RDN(n14021), .Q(bo4[6]) );
  DRNQHSV2 \pe4/pe3/q_reg[10]  ( .D(bo3[7]), .CK(clk), .RDN(n28530), .Q(bo4[7]) );
  DRNQHSV2 \pe4/pe3/q_reg[9]  ( .D(bo3[8]), .CK(clk), .RDN(n28492), .Q(bo4[8])
         );
  DRNQHSV2 \pe4/pe3/q_reg[7]  ( .D(bo3[10]), .CK(clk), .RDN(n28440), .Q(
        bo4[10]) );
  DRNQHSV2 \pe4/pe3/q_reg[6]  ( .D(bo3[11]), .CK(clk), .RDN(n28604), .Q(
        bo4[11]) );
  DRNQHSV2 \pe4/pe3/q_reg[5]  ( .D(bo3[12]), .CK(clk), .RDN(n28570), .Q(
        bo4[12]) );
  DRNQHSV2 \pe4/pe3/q_reg[3]  ( .D(bo3[14]), .CK(clk), .RDN(n28550), .Q(
        bo4[14]) );
  DRNQHSV2 \pe6/pe3/q_reg[16]  ( .D(bo5[1]), .CK(clk), .RDN(n28514), .Q(bo6[1]) );
  DRNQHSV2 \pe6/pe3/q_reg[15]  ( .D(bo5[2]), .CK(clk), .RDN(n28489), .Q(bo6[2]) );
  DRNQHSV2 \pe6/pe3/q_reg[12]  ( .D(bo5[5]), .CK(clk), .RDN(n28555), .Q(bo6[5]) );
  DRNQHSV2 \pe6/pe3/q_reg[11]  ( .D(bo5[6]), .CK(clk), .RDN(n28607), .Q(bo6[6]) );
  DRNQHSV2 \pe6/pe3/q_reg[10]  ( .D(bo5[7]), .CK(clk), .RDN(n28545), .Q(bo6[7]) );
  DRNQHSV2 \pe6/pe3/q_reg[9]  ( .D(bo5[8]), .CK(clk), .RDN(n28602), .Q(bo6[8])
         );
  DRNQHSV2 \pe6/pe3/q_reg[1]  ( .D(bo5[16]), .CK(clk), .RDN(n28513), .Q(
        bo6[16]) );
  DRNQHSV2 \pe7/pe3/q_reg[16]  ( .D(bo6[1]), .CK(clk), .RDN(n28568), .Q(bo7[1]) );
  DRNQHSV2 \pe7/pe3/q_reg[15]  ( .D(bo6[2]), .CK(clk), .RDN(n28537), .Q(bo7[2]) );
  DRNQHSV2 \pe7/pe3/q_reg[14]  ( .D(bo6[3]), .CK(clk), .RDN(n28558), .Q(bo7[3]) );
  DRNQHSV2 \pe7/pe3/q_reg[13]  ( .D(bo6[4]), .CK(clk), .RDN(n28541), .Q(bo7[4]) );
  DRNQHSV2 \pe7/pe3/q_reg[12]  ( .D(bo6[5]), .CK(clk), .RDN(n28452), .Q(bo7[5]) );
  DRNQHSV2 \pe7/pe3/q_reg[10]  ( .D(bo6[7]), .CK(clk), .RDN(n28558), .Q(bo7[7]) );
  DRNQHSV2 \pe7/pe3/q_reg[7]  ( .D(bo6[10]), .CK(clk), .RDN(n28521), .Q(
        bo7[10]) );
  DRNQHSV2 \pe7/pe3/q_reg[6]  ( .D(bo6[11]), .CK(clk), .RDN(n28542), .Q(
        bo7[11]) );
  DRNQHSV2 \pe7/pe3/q_reg[4]  ( .D(bo6[13]), .CK(clk), .RDN(n28507), .Q(
        bo7[13]) );
  DRNQHSV2 \pe7/pe3/q_reg[3]  ( .D(bo6[14]), .CK(clk), .RDN(n28552), .Q(
        bo7[14]) );
  DRNQHSV2 \pe7/pe3/q_reg[2]  ( .D(bo6[15]), .CK(clk), .RDN(n28574), .Q(
        bo7[15]) );
  DRNQHSV2 \pe7/pe3/q_reg[1]  ( .D(bo6[16]), .CK(clk), .RDN(n28522), .Q(
        bo7[16]) );
  DRNQHSV2 \pe9/pe3/q_reg[16]  ( .D(bo8[1]), .CK(clk), .RDN(n28516), .Q(bo9[1]) );
  DRNQHSV2 \pe9/pe3/q_reg[15]  ( .D(bo8[2]), .CK(clk), .RDN(n28459), .Q(bo9[2]) );
  DRNQHSV2 \pe9/pe3/q_reg[14]  ( .D(bo8[3]), .CK(clk), .RDN(n28482), .Q(bo9[3]) );
  DRNQHSV2 \pe9/pe3/q_reg[13]  ( .D(bo8[4]), .CK(clk), .RDN(n28508), .Q(bo9[4]) );
  DRNQHSV2 \pe9/pe3/q_reg[10]  ( .D(bo8[7]), .CK(clk), .RDN(n28543), .Q(bo9[7]) );
  DRNQHSV2 \pe9/pe3/q_reg[9]  ( .D(bo8[8]), .CK(clk), .RDN(n28567), .Q(bo9[8])
         );
  DRNQHSV2 \pe9/pe3/q_reg[8]  ( .D(bo8[9]), .CK(clk), .RDN(n28601), .Q(bo9[9])
         );
  DRNQHSV2 \pe9/pe3/q_reg[7]  ( .D(bo8[10]), .CK(clk), .RDN(n28500), .Q(
        bo9[10]) );
  DRNQHSV2 \pe9/pe3/q_reg[5]  ( .D(bo8[12]), .CK(clk), .RDN(n28521), .Q(
        bo9[12]) );
  DRNQHSV2 \pe9/pe3/q_reg[4]  ( .D(bo8[13]), .CK(clk), .RDN(n28504), .Q(
        bo9[13]) );
  DRNQHSV2 \pe9/pe3/q_reg[3]  ( .D(bo8[14]), .CK(clk), .RDN(n28504), .Q(
        bo9[14]) );
  DRNQHSV2 \pe9/pe3/q_reg[2]  ( .D(bo8[15]), .CK(clk), .RDN(n28446), .Q(
        bo9[15]) );
  DRNQHSV2 \pe9/pe3/q_reg[1]  ( .D(bo8[16]), .CK(clk), .RDN(n28575), .Q(
        bo9[16]) );
  DRNQHSV2 \pe5/pe3/q_reg[15]  ( .D(bo4[2]), .CK(clk), .RDN(n28552), .Q(bo5[2]) );
  DRNQHSV2 \pe5/pe3/q_reg[14]  ( .D(bo4[3]), .CK(clk), .RDN(n28491), .Q(bo5[3]) );
  DRNQHSV2 \pe5/pe3/q_reg[11]  ( .D(bo4[6]), .CK(clk), .RDN(n28492), .Q(bo5[6]) );
  DRNQHSV2 \pe5/pe3/q_reg[8]  ( .D(bo4[9]), .CK(clk), .RDN(n28602), .Q(bo5[9])
         );
  DRNQHSV2 \pe5/pe3/q_reg[7]  ( .D(bo4[10]), .CK(clk), .RDN(n28511), .Q(
        bo5[10]) );
  DRNQHSV2 \pe5/pe3/q_reg[6]  ( .D(bo4[11]), .CK(clk), .RDN(n28604), .Q(
        bo5[11]) );
  DRNQHSV2 \pe5/pe3/q_reg[4]  ( .D(bo4[13]), .CK(clk), .RDN(n28533), .Q(
        bo5[13]) );
  DRNQHSV2 \pe6/pe3/q_reg[14]  ( .D(bo5[3]), .CK(clk), .RDN(n28561), .Q(bo6[3]) );
  DRNQHSV2 \pe9/pe3/q_reg[12]  ( .D(bo8[5]), .CK(clk), .RDN(n28491), .Q(bo9[5]) );
  DRNQHSV2 \pe1/pe3/q_reg[14]  ( .D(bi[3]), .CK(clk), .RDN(rst), .Q(bo1[3]) );
  DRNQHSV2 \pe1/pe3/q_reg[13]  ( .D(bi[4]), .CK(clk), .RDN(n28498), .Q(bo1[4])
         );
  DRNQHSV2 \pe1/pe3/q_reg[6]  ( .D(bi[11]), .CK(clk), .RDN(n28445), .Q(bo1[11]) );
  DRNQHSV2 \pe2/pe3/q_reg[16]  ( .D(bo1[1]), .CK(clk), .RDN(n28573), .Q(bo2[1]) );
  DRNQHSV2 \pe2/pe3/q_reg[15]  ( .D(bo1[2]), .CK(clk), .RDN(n28441), .Q(bo2[2]) );
  DRNQHSV2 \pe2/pe3/q_reg[14]  ( .D(bo1[3]), .CK(clk), .RDN(n28549), .Q(bo2[3]) );
  DRNQHSV2 \pe2/pe3/q_reg[12]  ( .D(bo1[5]), .CK(clk), .RDN(n28530), .Q(bo2[5]) );
  DRNQHSV2 \pe2/pe3/q_reg[11]  ( .D(bo1[6]), .CK(clk), .RDN(n28503), .Q(bo2[6]) );
  DRNQHSV2 \pe2/pe3/q_reg[10]  ( .D(bo1[7]), .CK(clk), .RDN(n28500), .Q(bo2[7]) );
  DRNQHSV2 \pe2/pe3/q_reg[9]  ( .D(bo1[8]), .CK(clk), .RDN(n28527), .Q(bo2[8])
         );
  DRNQHSV2 \pe2/pe3/q_reg[8]  ( .D(bo1[9]), .CK(clk), .RDN(n28532), .Q(bo2[9])
         );
  DRNQHSV2 \pe2/pe3/q_reg[7]  ( .D(bo1[10]), .CK(clk), .RDN(n28484), .Q(
        bo2[10]) );
  DRNQHSV2 \pe2/pe3/q_reg[6]  ( .D(bo1[11]), .CK(clk), .RDN(n28575), .Q(
        bo2[11]) );
  DRNQHSV2 \pe2/pe3/q_reg[5]  ( .D(bo1[12]), .CK(clk), .RDN(n28573), .Q(
        bo2[12]) );
  DRNQHSV2 \pe2/pe3/q_reg[4]  ( .D(bo1[13]), .CK(clk), .RDN(n28574), .Q(
        bo2[13]) );
  DRNQHSV2 \pe2/pe3/q_reg[3]  ( .D(bo1[14]), .CK(clk), .RDN(n28498), .Q(
        bo2[14]) );
  DRNQHSV2 \pe2/pe3/q_reg[2]  ( .D(bo1[15]), .CK(clk), .RDN(n28534), .Q(
        bo2[15]) );
  DRNQHSV2 \pe2/pe3/q_reg[1]  ( .D(bo1[16]), .CK(clk), .RDN(n28528), .Q(
        bo2[16]) );
  DRNQHSV2 \pe3/pe3/q_reg[16]  ( .D(bo2[1]), .CK(clk), .RDN(n28549), .Q(bo3[1]) );
  DRNQHSV2 \pe3/pe3/q_reg[15]  ( .D(bo2[2]), .CK(clk), .RDN(n28440), .Q(bo3[2]) );
  DRNQHSV2 \pe3/pe3/q_reg[14]  ( .D(bo2[3]), .CK(clk), .RDN(n28503), .Q(bo3[3]) );
  DRNQHSV1 \pe3/pe3/q_reg[13]  ( .D(bo2[4]), .CK(clk), .RDN(n28536), .Q(bo3[4]) );
  DRNQHSV2 \pe3/pe3/q_reg[12]  ( .D(bo2[5]), .CK(clk), .RDN(n28511), .Q(bo3[5]) );
  DRNQHSV2 \pe3/pe3/q_reg[10]  ( .D(bo2[7]), .CK(clk), .RDN(n28490), .Q(bo3[7]) );
  DRNQHSV2 \pe3/pe3/q_reg[9]  ( .D(bo2[8]), .CK(clk), .RDN(n28566), .Q(bo3[8])
         );
  DRNQHSV2 \pe3/pe3/q_reg[8]  ( .D(bo2[9]), .CK(clk), .RDN(n28524), .Q(bo3[9])
         );
  DRNQHSV2 \pe3/pe3/q_reg[7]  ( .D(bo2[10]), .CK(clk), .RDN(n28508), .Q(
        bo3[10]) );
  DRNQHSV2 \pe3/pe3/q_reg[6]  ( .D(bo2[11]), .CK(clk), .RDN(n28536), .Q(
        bo3[11]) );
  DRNQHSV2 \pe3/pe3/q_reg[5]  ( .D(bo2[12]), .CK(clk), .RDN(n28607), .Q(
        bo3[12]) );
  DRNQHSV2 \pe3/pe3/q_reg[4]  ( .D(bo2[13]), .CK(clk), .RDN(n28528), .Q(
        bo3[13]) );
  DRNQHSV2 \pe3/pe3/q_reg[3]  ( .D(bo2[14]), .CK(clk), .RDN(n28573), .Q(
        bo3[14]) );
  DRNQHSV2 \pe3/pe3/q_reg[1]  ( .D(bo2[16]), .CK(clk), .RDN(n28538), .Q(
        bo3[16]) );
  DRNQHSV2 \pe4/pe3/q_reg[12]  ( .D(bo3[5]), .CK(clk), .RDN(n28520), .Q(bo4[5]) );
  DRNQHSV2 \pe4/pe3/q_reg[8]  ( .D(bo3[9]), .CK(clk), .RDN(n28496), .Q(bo4[9])
         );
  DRNQHSV2 \pe4/pe3/q_reg[4]  ( .D(bo3[13]), .CK(clk), .RDN(n14021), .Q(
        bo4[13]) );
  DRNQHSV2 \pe4/pe3/q_reg[1]  ( .D(bo3[16]), .CK(clk), .RDN(n28539), .Q(
        bo4[16]) );
  DRNQHSV2 \pe6/pe3/q_reg[8]  ( .D(bo5[9]), .CK(clk), .RDN(n28492), .Q(bo6[9])
         );
  DRNQHSV2 \pe6/pe3/q_reg[7]  ( .D(bo5[10]), .CK(clk), .RDN(n28517), .Q(
        bo6[10]) );
  DRNQHSV2 \pe6/pe3/q_reg[6]  ( .D(bo5[11]), .CK(clk), .RDN(n28541), .Q(
        bo6[11]) );
  DRNQHSV2 \pe6/pe3/q_reg[5]  ( .D(bo5[12]), .CK(clk), .RDN(n28495), .Q(
        bo6[12]) );
  DRNQHSV2 \pe6/pe3/q_reg[4]  ( .D(bo5[13]), .CK(clk), .RDN(n28453), .Q(
        bo6[13]) );
  DRNQHSV2 \pe6/pe3/q_reg[3]  ( .D(bo5[14]), .CK(clk), .RDN(n28543), .Q(
        bo6[14]) );
  DRNQHSV2 \pe6/pe3/q_reg[2]  ( .D(bo5[15]), .CK(clk), .RDN(n28511), .Q(
        bo6[15]) );
  DRNQHSV2 \pe7/pe3/q_reg[11]  ( .D(bo6[6]), .CK(clk), .RDN(n28516), .Q(bo7[6]) );
  DRNQHSV2 \pe7/pe3/q_reg[9]  ( .D(bo6[8]), .CK(clk), .RDN(n28575), .Q(bo7[8])
         );
  DRNQHSV2 \pe7/pe3/q_reg[8]  ( .D(bo6[9]), .CK(clk), .RDN(n28601), .Q(bo7[9])
         );
  DRNQHSV1 \pe8/pe3/q_reg[16]  ( .D(bo7[1]), .CK(clk), .RDN(n28493), .Q(bo8[1]) );
  DRNQHSV2 \pe8/pe3/q_reg[15]  ( .D(bo7[2]), .CK(clk), .RDN(n28493), .Q(bo8[2]) );
  DRNQHSV1 \pe8/pe3/q_reg[14]  ( .D(bo7[3]), .CK(clk), .RDN(n28548), .Q(bo8[3]) );
  DRNQHSV2 \pe8/pe3/q_reg[13]  ( .D(bo7[4]), .CK(clk), .RDN(n28575), .Q(bo8[4]) );
  DRNQHSV2 \pe8/pe3/q_reg[12]  ( .D(bo7[5]), .CK(clk), .RDN(n28530), .Q(bo8[5]) );
  DRNQHSV2 \pe8/pe3/q_reg[11]  ( .D(bo7[6]), .CK(clk), .RDN(n28558), .Q(bo8[6]) );
  DRNQHSV2 \pe8/pe3/q_reg[10]  ( .D(bo7[7]), .CK(clk), .RDN(n28562), .Q(bo8[7]) );
  DRNQHSV2 \pe8/pe3/q_reg[9]  ( .D(bo7[8]), .CK(clk), .RDN(n28537), .Q(bo8[8])
         );
  DRNQHSV2 \pe8/pe3/q_reg[8]  ( .D(bo7[9]), .CK(clk), .RDN(n28576), .Q(bo8[9])
         );
  DRNQHSV2 \pe8/pe3/q_reg[7]  ( .D(bo7[10]), .CK(clk), .RDN(n28527), .Q(
        bo8[10]) );
  DRNQHSV2 \pe8/pe3/q_reg[6]  ( .D(bo7[11]), .CK(clk), .RDN(n28566), .Q(
        bo8[11]) );
  DRNQHSV2 \pe8/pe3/q_reg[5]  ( .D(bo7[12]), .CK(clk), .RDN(n28459), .Q(
        bo8[12]) );
  DRNQHSV2 \pe8/pe3/q_reg[4]  ( .D(bo7[13]), .CK(clk), .RDN(n28527), .Q(
        bo8[13]) );
  DRNQHSV1 \pe8/pe3/q_reg[3]  ( .D(bo7[14]), .CK(clk), .RDN(n28576), .Q(
        bo8[14]) );
  DRNQHSV1 \pe8/pe3/q_reg[2]  ( .D(bo7[15]), .CK(clk), .RDN(n28527), .Q(
        bo8[15]) );
  DRNQHSV1 \pe8/pe3/q_reg[1]  ( .D(bo7[16]), .CK(clk), .RDN(n28550), .Q(
        bo8[16]) );
  DRNQHSV2 \pe9/pe3/q_reg[11]  ( .D(bo8[6]), .CK(clk), .RDN(n28516), .Q(bo9[6]) );
  DRNQHSV2 \pe9/pe3/q_reg[6]  ( .D(bo8[11]), .CK(clk), .RDN(n28572), .Q(
        bo9[11]) );
  DRNQHSV2 \pe10/pe3/q_reg[16]  ( .D(bo9[1]), .CK(clk), .RDN(n28540), .Q(
        bo10[1]) );
  DRNQHSV1 \pe10/pe3/q_reg[15]  ( .D(bo9[2]), .CK(clk), .RDN(n28511), .Q(
        bo10[2]) );
  DRNQHSV2 \pe10/pe3/q_reg[14]  ( .D(bo9[3]), .CK(clk), .RDN(n28601), .Q(
        bo10[3]) );
  DRNQHSV2 \pe10/pe3/q_reg[13]  ( .D(bo9[4]), .CK(clk), .RDN(n28450), .Q(
        bo10[4]) );
  DRNQHSV2 \pe10/pe3/q_reg[12]  ( .D(bo9[5]), .CK(clk), .RDN(n28448), .Q(
        bo10[5]) );
  DRNQHSV2 \pe10/pe3/q_reg[11]  ( .D(bo9[6]), .CK(clk), .RDN(n28549), .Q(
        bo10[6]) );
  DRNQHSV2 \pe10/pe3/q_reg[10]  ( .D(bo9[7]), .CK(clk), .RDN(n28511), .Q(
        bo10[7]) );
  DRNQHSV2 \pe10/pe3/q_reg[9]  ( .D(bo9[8]), .CK(clk), .RDN(n28601), .Q(
        bo10[8]) );
  DRNQHSV2 \pe10/pe3/q_reg[8]  ( .D(bo9[9]), .CK(clk), .RDN(n28476), .Q(
        bo10[9]) );
  DRNQHSV2 \pe10/pe3/q_reg[7]  ( .D(bo9[10]), .CK(clk), .RDN(n28513), .Q(
        bo10[10]) );
  DRNQHSV2 \pe10/pe3/q_reg[6]  ( .D(bo9[11]), .CK(clk), .RDN(n28483), .Q(
        bo10[11]) );
  DRNQHSV2 \pe10/pe3/q_reg[5]  ( .D(bo9[12]), .CK(clk), .RDN(n28543), .Q(
        bo10[12]) );
  DRNQHSV2 \pe10/pe3/q_reg[4]  ( .D(bo9[13]), .CK(clk), .RDN(n28566), .Q(
        bo10[13]) );
  DRNQHSV2 \pe10/pe3/q_reg[3]  ( .D(bo9[14]), .CK(clk), .RDN(n28498), .Q(
        bo10[14]) );
  DRNQHSV1 \pe10/pe3/q_reg[2]  ( .D(bo9[15]), .CK(clk), .RDN(n28520), .Q(
        bo10[15]) );
  DRNQHSV1 \pe10/pe3/q_reg[1]  ( .D(bo9[16]), .CK(clk), .RDN(n28543), .Q(
        bo10[16]) );
  DRNQHSV2 \pe5/pe3/q_reg[16]  ( .D(bo4[1]), .CK(clk), .RDN(n28571), .Q(bo5[1]) );
  DRNQHSV2 \pe5/pe3/q_reg[13]  ( .D(bo4[4]), .CK(clk), .RDN(n28541), .Q(bo5[4]) );
  DRNQHSV2 \pe5/pe3/q_reg[12]  ( .D(bo4[5]), .CK(clk), .RDN(n28544), .Q(bo5[5]) );
  DRNQHSV2 \pe5/pe3/q_reg[10]  ( .D(bo4[7]), .CK(clk), .RDN(n28602), .Q(bo5[7]) );
  DRNQHSV2 \pe5/pe3/q_reg[9]  ( .D(bo4[8]), .CK(clk), .RDN(n28515), .Q(bo5[8])
         );
  DRNQHSV2 \pe5/pe3/q_reg[5]  ( .D(bo4[12]), .CK(clk), .RDN(n28525), .Q(
        bo5[12]) );
  DRNQHSV2 \pe5/pe3/q_reg[3]  ( .D(bo4[14]), .CK(clk), .RDN(n28503), .Q(
        bo5[14]) );
  DRNQHSV1 \pe5/pe3/q_reg[2]  ( .D(bo4[15]), .CK(clk), .RDN(n28442), .Q(
        bo5[15]) );
  DRNQHSV1 \pe2/pe14/q_reg[15]  ( .D(n28456), .CK(clk), .RDN(n28548), .Q(
        \pe2/ti_7t [15]) );
  DRNQHSV1 \pe10/pe14/q_reg[14]  ( .D(n25060), .CK(clk), .RDN(n28500), .Q(
        \pe10/ti_7t [14]) );
  DRNQHSV1 \pe6/pe14/q_reg[13]  ( .D(n28699), .CK(clk), .RDN(n28562), .Q(
        \pe6/ti_7t [13]) );
  DRNQHSV1 \pe9/pe14/q_reg[13]  ( .D(n28475), .CK(clk), .RDN(n28491), .Q(
        \pe9/ti_7t [13]) );
  DRNQHSV1 \pe5/pe14/q_reg[14]  ( .D(n28946), .CK(clk), .RDN(n28505), .Q(
        \pe5/ti_7t [14]) );
  DRNQHSV1 \pe6/pe14/q_reg[14]  ( .D(n28787), .CK(clk), .RDN(n28576), .Q(
        \pe6/ti_7t [14]) );
  DRNQHSV2 \pe7/pe14/q_reg[13]  ( .D(n28934), .CK(clk), .RDN(n28546), .Q(
        \pe7/ti_7t [13]) );
  DRNQHSV2 \pe4/pe14/q_reg[14]  ( .D(n28941), .CK(clk), .RDN(n28577), .Q(
        \pe4/ti_7t [14]) );
  DRNQHSV1 \pe8/pe14/q_reg[13]  ( .D(n28426), .CK(clk), .RDN(n28452), .Q(
        \pe8/ti_7t [13]) );
  DRNQHSV1 \pe5/pe14/q_reg[12]  ( .D(n28473), .CK(clk), .RDN(n28448), .Q(
        \pe5/ti_7t [12]) );
  DRNQHSV1 \pe4/pe14/q_reg[13]  ( .D(n28480), .CK(clk), .RDN(n28524), .Q(
        \pe4/ti_7t [13]) );
  DRNQHSV1 \pe2/pe14/q_reg[14]  ( .D(n28701), .CK(clk), .RDN(n28525), .Q(
        \pe2/ti_7t [14]) );
  DRNQHSV1 \pe3/pe14/q_reg[8]  ( .D(n23327), .CK(clk), .RDN(n28441), .Q(
        \pe3/ti_7t [8]) );
  DRNQHSV2 \pe5/pe14/q_reg[9]  ( .D(n21554), .CK(clk), .RDN(n28497), .Q(
        \pe5/ti_7t [9]) );
  DRNQHSV1 \pe5/pe14/q_reg[11]  ( .D(n28803), .CK(clk), .RDN(n28441), .Q(
        \pe5/ti_7t [11]) );
  DRNQHSV1 \pe6/pe14/q_reg[8]  ( .D(n23041), .CK(clk), .RDN(n28548), .Q(
        \pe6/ti_7t [8]) );
  DRNQHSV1 \pe6/pe14/q_reg[12]  ( .D(n28467), .CK(clk), .RDN(n28451), .Q(
        \pe6/ti_7t [12]) );
  DRNQHSV1 \pe7/pe14/q_reg[11]  ( .D(n28665), .CK(clk), .RDN(n28602), .Q(
        \pe7/ti_7t [11]) );
  DRNQHSV1 \pe8/pe14/q_reg[10]  ( .D(n14059), .CK(clk), .RDN(n28572), .Q(
        \pe8/ti_7t [10]) );
  DRNQHSV1 \pe9/pe14/q_reg[8]  ( .D(n28790), .CK(clk), .RDN(n28452), .Q(
        \pe9/ti_7t [8]) );
  DRNQHSV1 \pe11/pe14/q_reg[11]  ( .D(n25137), .CK(clk), .RDN(n28520), .Q(
        \pe11/ti_7t [11]) );
  DRNQHSV1 \pe1/pe14/q_reg[9]  ( .D(n26854), .CK(clk), .RDN(n28552), .Q(
        \pe1/ti_7t [9]) );
  DRNQHSV1 \pe1/pe14/q_reg[12]  ( .D(n28460), .CK(clk), .RDN(n28551), .Q(
        \pe1/ti_7t [12]) );
  DRNQHSV1 \pe2/pe14/q_reg[10]  ( .D(n28474), .CK(clk), .RDN(n28515), .Q(
        \pe2/ti_7t [10]) );
  DRNQHSV1 \pe2/pe14/q_reg[11]  ( .D(n27657), .CK(clk), .RDN(n28559), .Q(
        \pe2/ti_7t [11]) );
  DRNQHSV1 \pe2/pe14/q_reg[12]  ( .D(n28702), .CK(clk), .RDN(n28559), .Q(
        \pe2/ti_7t [12]) );
  DRNQHSV1 \pe3/pe14/q_reg[10]  ( .D(n28945), .CK(clk), .RDN(n28535), .Q(
        \pe3/ti_7t [10]) );
  DRNQHSV1 \pe4/pe14/q_reg[11]  ( .D(n14038), .CK(clk), .RDN(n28568), .Q(
        \pe4/ti_7t [11]) );
  DRNQHSV1 \pe7/pe14/q_reg[10]  ( .D(n28656), .CK(clk), .RDN(n28531), .Q(
        \pe7/ti_7t [10]) );
  DRNQHSV1 \pe8/pe14/q_reg[11]  ( .D(n28706), .CK(clk), .RDN(n28489), .Q(
        \pe8/ti_7t [11]) );
  DRNQHSV1 \pe9/pe14/q_reg[10]  ( .D(n28317), .CK(clk), .RDN(n28515), .Q(
        \pe9/ti_7t [10]) );
  DRNQHSV1 \pe10/pe14/q_reg[12]  ( .D(n28469), .CK(clk), .RDN(n28495), .Q(
        \pe10/ti_7t [12]) );
  DRNQHSV1 \pe11/pe14/q_reg[10]  ( .D(n14064), .CK(clk), .RDN(n28501), .Q(
        \pe11/ti_7t [10]) );
  DRNQHSV1 \pe6/pe14/q_reg[9]  ( .D(n26068), .CK(clk), .RDN(n28495), .Q(
        \pe6/ti_7t [9]) );
  DRNQHSV1 \pe8/pe14/q_reg[8]  ( .D(n28616), .CK(clk), .RDN(n28557), .Q(
        \pe8/ti_7t [8]) );
  DRNQHSV1 \pe1/pe14/q_reg[8]  ( .D(n28589), .CK(clk), .RDN(n28561), .Q(
        \pe1/ti_7t [8]) );
  DRNQHSV2 \pe3/pe14/q_reg[12]  ( .D(n28939), .CK(clk), .RDN(n28447), .Q(
        \pe3/ti_7t [12]) );
  DRNQHSV1 \pe11/pe14/q_reg[12]  ( .D(n28919), .CK(clk), .RDN(n28570), .Q(
        \pe11/ti_7t [12]) );
  DRNQHSV1 \pe5/pe14/q_reg[8]  ( .D(n28800), .CK(clk), .RDN(n28499), .Q(
        \pe5/ti_7t [8]) );
  DRNQHSV1 \pe4/pe14/q_reg[8]  ( .D(n28578), .CK(clk), .RDN(n28576), .Q(
        \pe4/ti_7t [8]) );
  DRNQHSV2 \pe10/pe14/q_reg[11]  ( .D(n26215), .CK(clk), .RDN(n28521), .Q(
        \pe10/ti_7t [11]) );
  DRNQHSV1 \pe1/pe14/q_reg[11]  ( .D(n26416), .CK(clk), .RDN(n28597), .Q(
        \pe1/ti_7t [11]) );
  DRNQHSV1 \pe9/pe14/q_reg[11]  ( .D(n28419), .CK(clk), .RDN(n28557), .Q(
        \pe9/ti_7t [11]) );
  DRNQHSV1 \pe3/pe14/q_reg[9]  ( .D(n28438), .CK(clk), .RDN(n14023), .Q(
        \pe3/ti_7t [9]) );
  DRNQHSV1 \pe5/pe14/q_reg[10]  ( .D(\pe5/ti_7[10] ), .CK(clk), .RDN(n28557), 
        .Q(\pe5/ti_7t [10]) );
  DRNQHSV1 \pe1/pe14/q_reg[10]  ( .D(n26418), .CK(clk), .RDN(n28597), .Q(
        \pe1/ti_7t [10]) );
  DRNQHSV1 \pe6/pe14/q_reg[11]  ( .D(n28937), .CK(clk), .RDN(n28505), .Q(
        \pe6/ti_7t [11]) );
  DRNQHSV1 \pe4/pe14/q_reg[12]  ( .D(n25079), .CK(clk), .RDN(n28577), .Q(
        \pe4/ti_7t [12]) );
  DRNQHSV1 \pe2/pe14/q_reg[9]  ( .D(n28805), .CK(clk), .RDN(n28500), .Q(
        \pe2/ti_7t [9]) );
  DRNQHSV1 \pe10/pe14/q_reg[8]  ( .D(n28620), .CK(clk), .RDN(n28541), .Q(
        \pe10/ti_7t [8]) );
  DRNQHSV1 \pe7/pe14/q_reg[3]  ( .D(n28621), .CK(clk), .RDN(n28554), .Q(
        \pe7/ti_7t [3]) );
  DRNQHSV1 \pe9/pe14/q_reg[5]  ( .D(n28638), .CK(clk), .RDN(n28542), .Q(
        \pe9/ti_7t [5]) );
  DRNQHSV1 \pe9/pe14/q_reg[6]  ( .D(n28689), .CK(clk), .RDN(n28535), .Q(
        \pe9/ti_7t [6]) );
  DRNQHSV1 \pe5/pe14/q_reg[4]  ( .D(n28664), .CK(clk), .RDN(n28443), .Q(
        \pe5/ti_7t [4]) );
  DRNQHSV1 \pe2/pe14/q_reg[5]  ( .D(n28809), .CK(clk), .RDN(n28595), .Q(
        \pe2/ti_7t [5]) );
  DRNQHSV1 \pe1/pe14/q_reg[6]  ( .D(n28418), .CK(clk), .RDN(n28501), .Q(
        \pe1/ti_7t [6]) );
  DRNQHSV2 \pe2/pe5/q_reg[15]  ( .D(n29046), .CK(clk), .RDN(n28493), .Q(
        \pe2/pvq [15]) );
  DRNQHSV1 \pe2/pe5/q_reg[14]  ( .D(n13962), .CK(clk), .RDN(n28493), .Q(
        \pe2/pvq [14]) );
  DRNQHSV1 \pe2/pe5/q_reg[13]  ( .D(n28958), .CK(clk), .RDN(n28483), .Q(
        \pe2/pvq [13]) );
  DRNQHSV1 \pe2/pe14/q_reg[4]  ( .D(n28427), .CK(clk), .RDN(n28444), .Q(
        \pe2/ti_7t [4]) );
  DRNQHSV1 \pe2/pe14/q_reg[7]  ( .D(n28617), .CK(clk), .RDN(n28525), .Q(
        \pe2/ti_7t [7]) );
  DRNQHSV2 \pe3/pe5/q_reg[15]  ( .D(n28970), .CK(clk), .RDN(n28536), .Q(
        \pe3/pvq [15]) );
  DRNQHSV2 \pe3/pe5/q_reg[13]  ( .D(n28986), .CK(clk), .RDN(n28563), .Q(
        \pe3/pvq [13]) );
  DRNQHSV1 \pe3/pe5/q_reg[12]  ( .D(n28972), .CK(clk), .RDN(n28565), .Q(
        \pe3/pvq [12]) );
  DRNQHSV1 \pe3/pe5/q_reg[11]  ( .D(n28950), .CK(clk), .RDN(n28529), .Q(
        \pe3/pvq [11]) );
  DRNQHSV1 \pe3/pe5/q_reg[9]  ( .D(n28956), .CK(clk), .RDN(n28520), .Q(
        \pe3/pvq [9]) );
  DRNQHSV2 \pe4/pe5/q_reg[15]  ( .D(n28979), .CK(clk), .RDN(n28509), .Q(
        \pe4/pvq [15]) );
  DRNQHSV1 \pe4/pe5/q_reg[14]  ( .D(n29035), .CK(clk), .RDN(n28549), .Q(
        \pe4/pvq [14]) );
  DRNQHSV1 \pe4/pe5/q_reg[13]  ( .D(n28963), .CK(clk), .RDN(n28458), .Q(
        \pe4/pvq [13]) );
  DRNQHSV1 \pe4/pe5/q_reg[12]  ( .D(n21312), .CK(clk), .RDN(n28528), .Q(
        \pe4/pvq [12]) );
  DRNQHSV2 \pe5/pe5/q_reg[15]  ( .D(pov4[15]), .CK(clk), .RDN(n28595), .Q(
        \pe5/pvq [15]) );
  DRNQHSV1 \pe5/pe5/q_reg[14]  ( .D(pov4[14]), .CK(clk), .RDN(n28538), .Q(
        \pe5/pvq [14]) );
  DRNQHSV1 \pe5/pe5/q_reg[13]  ( .D(pov4[13]), .CK(clk), .RDN(n28492), .Q(
        \pe5/pvq [13]) );
  DRNQHSV1 \pe5/pe5/q_reg[12]  ( .D(n29028), .CK(clk), .RDN(n28601), .Q(
        \pe5/pvq [12]) );
  DRNQHSV1 \pe6/pe5/q_reg[15]  ( .D(pov5[15]), .CK(clk), .RDN(n28508), .Q(
        \pe6/pvq [15]) );
  DRNQHSV1 \pe6/pe5/q_reg[14]  ( .D(n28965), .CK(clk), .RDN(n28445), .Q(
        \pe6/pvq [14]) );
  DRNQHSV1 \pe6/pe5/q_reg[12]  ( .D(n28973), .CK(clk), .RDN(n28458), .Q(
        \pe6/pvq [12]) );
  DRNQHSV1 \pe6/pe5/q_reg[11]  ( .D(n28971), .CK(clk), .RDN(n28602), .Q(
        \pe6/pvq [11]) );
  DRNQHSV1 \pe6/pe14/q_reg[3]  ( .D(n28793), .CK(clk), .RDN(n28486), .Q(
        \pe6/ti_7t [3]) );
  DRNQHSV1 \pe6/pe14/q_reg[4]  ( .D(n28792), .CK(clk), .RDN(n28547), .Q(
        \pe6/ti_7t [4]) );
  DRNQHSV1 \pe6/pe14/q_reg[6]  ( .D(n28526), .CK(clk), .RDN(n28548), .Q(
        \pe6/ti_7t [6]) );
  DRNQHSV1 \pe7/pe5/q_reg[15]  ( .D(pov6[15]), .CK(clk), .RDN(n28518), .Q(
        \pe7/pvq [15]) );
  DRNQHSV2 \pe7/pe5/q_reg[14]  ( .D(n29018), .CK(clk), .RDN(n28495), .Q(
        \pe7/pvq [14]) );
  DRNQHSV1 \pe7/pe5/q_reg[13]  ( .D(n29019), .CK(clk), .RDN(n28572), .Q(
        \pe7/pvq [13]) );
  DRNQHSV1 \pe7/pe5/q_reg[12]  ( .D(n29020), .CK(clk), .RDN(n28551), .Q(
        \pe7/pvq [12]) );
  DRNQHSV1 \pe7/pe5/q_reg[11]  ( .D(pov6[11]), .CK(clk), .RDN(n28563), .Q(
        \pe7/pvq [11]) );
  DRNQHSV1 \pe7/pe5/q_reg[10]  ( .D(n29021), .CK(clk), .RDN(n28568), .Q(
        \pe7/pvq [10]) );
  DRNQHSV1 \pe7/pe14/q_reg[4]  ( .D(n11936), .CK(clk), .RDN(n28560), .Q(
        \pe7/ti_7t [4]) );
  DRNQHSV1 \pe8/pe5/q_reg[15]  ( .D(n28978), .CK(clk), .RDN(n28520), .Q(
        \pe8/pvq [15]) );
  DRNQHSV2 \pe8/pe5/q_reg[14]  ( .D(n29013), .CK(clk), .RDN(n28502), .Q(
        \pe8/pvq [14]) );
  DRNQHSV1 \pe8/pe5/q_reg[13]  ( .D(n28948), .CK(clk), .RDN(n28565), .Q(
        \pe8/pvq [13]) );
  DRNQHSV1 \pe8/pe14/q_reg[6]  ( .D(n14042), .CK(clk), .RDN(n28447), .Q(
        \pe8/ti_7t [6]) );
  DRNQHSV1 \pe9/pe5/q_reg[15]  ( .D(n29004), .CK(clk), .RDN(n28516), .Q(
        \pe9/pvq [15]) );
  DRNQHSV1 \pe9/pe5/q_reg[12]  ( .D(pov8[12]), .CK(clk), .RDN(n28538), .Q(
        \pe9/pvq [12]) );
  DRNQHSV2 \pe10/pe5/q_reg[15]  ( .D(pov9[15]), .CK(clk), .RDN(n28543), .Q(
        \pe10/pvq [15]) );
  DRNQHSV1 \pe10/pe5/q_reg[14]  ( .D(pov9[14]), .CK(clk), .RDN(n28607), .Q(
        \pe10/pvq [14]) );
  DRNQHSV2 \pe10/pe5/q_reg[13]  ( .D(pov9[13]), .CK(clk), .RDN(n28497), .Q(
        \pe10/pvq [13]) );
  DRNQHSV1 \pe10/pe14/q_reg[3]  ( .D(n28679), .CK(clk), .RDN(n28447), .Q(
        \pe10/ti_7t [3]) );
  DRNQHSV1 \pe10/pe14/q_reg[5]  ( .D(n26131), .CK(clk), .RDN(n28524), .Q(
        \pe10/ti_7t [5]) );
  DRNQHSV2 \pe11/pe5/q_reg[15]  ( .D(n28980), .CK(clk), .RDN(n28596), .Q(
        \pe11/pvq [15]) );
  DRNQHSV2 \pe11/pe5/q_reg[14]  ( .D(pov10[14]), .CK(clk), .RDN(n28522), .Q(
        \pe11/pvq [14]) );
  DRNQHSV1 \pe11/pe5/q_reg[13]  ( .D(n12263), .CK(clk), .RDN(n28518), .Q(
        \pe11/pvq [13]) );
  DRNQHSV1 \pe11/pe5/q_reg[11]  ( .D(n28996), .CK(clk), .RDN(n28564), .Q(
        \pe11/pvq [11]) );
  DRNQHSV1 \pe11/pe14/q_reg[3]  ( .D(n28807), .CK(clk), .RDN(n28476), .Q(
        \pe11/ti_7t [3]) );
  DRNQHSV1 \pe11/pe14/q_reg[4]  ( .D(n20467), .CK(clk), .RDN(n28516), .Q(
        \pe11/ti_7t [4]) );
  DRNQHSV1 \pe11/pe14/q_reg[7]  ( .D(n28791), .CK(clk), .RDN(n28501), .Q(
        \pe11/ti_7t [7]) );
  DRNQHSV1 \pe7/pe14/q_reg[5]  ( .D(n28657), .CK(clk), .RDN(n28541), .Q(
        \pe7/ti_7t [5]) );
  DRNQHSV1 \pe8/pe14/q_reg[3]  ( .D(n28799), .CK(clk), .RDN(n28606), .Q(
        \pe8/ti_7t [3]) );
  DRNQHSV1 \pe5/pe14/q_reg[7]  ( .D(n28806), .CK(clk), .RDN(n28499), .Q(
        \pe5/ti_7t [7]) );
  DRNQHSV1 \pe4/pe14/q_reg[6]  ( .D(n28933), .CK(clk), .RDN(n28484), .Q(
        \pe4/ti_7t [6]) );
  DRNQHSV1 \pe2/pe14/q_reg[6]  ( .D(n27271), .CK(clk), .RDN(n28459), .Q(
        \pe2/ti_7t [6]) );
  DRNQHSV2 \pe5/pe4/q_reg  ( .D(po4), .CK(clk), .RDN(n28486), .Q(\pe5/pq ) );
  DRNQHSV2 \pe6/pe4/q_reg  ( .D(po5), .CK(clk), .RDN(n28549), .Q(\pe6/pq ) );
  DRNQHSV2 \pe9/pe4/q_reg  ( .D(po8), .CK(clk), .RDN(n28564), .Q(\pe9/pq ) );
  DRNQHSV1 \pe3/pe14/q_reg[5]  ( .D(n28432), .CK(clk), .RDN(n28497), .Q(
        \pe3/ti_7t [5]) );
  DRNQHSV1 \pe4/pe14/q_reg[7]  ( .D(\pe4/ti_7[7] ), .CK(clk), .RDN(n28545), 
        .Q(\pe4/ti_7t [7]) );
  DRNQHSV1 \pe1/pe14/q_reg[5]  ( .D(n28649), .CK(clk), .RDN(n28542), .Q(
        \pe1/ti_7t [5]) );
  DRNQHSV1 \pe9/pe14/q_reg[7]  ( .D(n28952), .CK(clk), .RDN(n28492), .Q(
        \pe9/ti_7t [7]) );
  DRNQHSV1 \pe1/pe14/q_reg[7]  ( .D(n28609), .CK(clk), .RDN(n28574), .Q(
        \pe1/ti_7t [7]) );
  DRNQHSV1 \pe4/pe14/q_reg[5]  ( .D(n28696), .CK(clk), .RDN(n28602), .Q(
        \pe4/ti_7t [5]) );
  DRNQHSV1 \pe8/pe14/q_reg[5]  ( .D(n28462), .CK(clk), .RDN(n28439), .Q(
        \pe8/ti_7t [5]) );
  DRNQHSV1 \pe10/pe14/q_reg[4]  ( .D(n28794), .CK(clk), .RDN(n28561), .Q(
        \pe10/ti_7t [4]) );
  DRNQHSV1 \pe11/pe14/q_reg[6]  ( .D(n28471), .CK(clk), .RDN(n28482), .Q(
        \pe11/ti_7t [6]) );
  DRNQHSV1 \pe5/pe14/q_reg[6]  ( .D(n28478), .CK(clk), .RDN(n28488), .Q(
        \pe5/ti_7t [6]) );
  DRNQHSV1 \pe3/pe14/q_reg[7]  ( .D(n28588), .CK(clk), .RDN(n28506), .Q(
        \pe3/ti_7t [7]) );
  DRNQHSV1 \pe3/pe14/q_reg[3]  ( .D(n28920), .CK(clk), .RDN(n28554), .Q(
        \pe3/ti_7t [3]) );
  DRNQHSV1 \pe2/pe14/q_reg[3]  ( .D(n28954), .CK(clk), .RDN(n28500), .Q(
        \pe2/ti_7t [3]) );
  DRNQHSV1 \pe9/pe14/q_reg[3]  ( .D(n28804), .CK(clk), .RDN(n28496), .Q(
        \pe9/ti_7t [3]) );
  DRNQHSV1 \pe4/pe14/q_reg[3]  ( .D(n28951), .CK(clk), .RDN(n28519), .Q(
        \pe4/ti_7t [3]) );
  DRNQHSV1 \pe9/pe14/q_reg[4]  ( .D(n28949), .CK(clk), .RDN(n28488), .Q(
        \pe9/ti_7t [4]) );
  DRNQHSV2 \pe1/pe2/q_reg[16]  ( .D(gi[1]), .CK(clk), .RDN(n28604), .Q(
        \pe1/got [1]) );
  DRNQHSV2 \pe1/pe2/q_reg[14]  ( .D(gi[3]), .CK(clk), .RDN(n28604), .Q(
        \pe1/got [3]) );
  DRNQHSV2 \pe1/pe2/q_reg[12]  ( .D(gi[5]), .CK(clk), .RDN(n28601), .Q(
        \pe1/got [5]) );
  DRNQHSV1 \pe2/pe14/q_reg[1]  ( .D(n28697), .CK(clk), .RDN(n28494), .Q(
        \pe2/ti_7t [1]) );
  DRNQHSV1 \pe3/pe14/q_reg[2]  ( .D(n15979), .CK(clk), .RDN(n28497), .Q(
        \pe3/ti_7t [2]) );
  DRNQHSV1 \pe10/pe14/q_reg[2]  ( .D(n28630), .CK(clk), .RDN(n28555), .Q(
        \pe10/ti_7t [2]) );
  DRNQHSV1 \pe1/pe14/q_reg[2]  ( .D(n28814), .CK(clk), .RDN(n28597), .Q(
        \pe1/ti_7t [2]) );
  DRNQHSV1 \pe11/pe14/q_reg[2]  ( .D(n20505), .CK(clk), .RDN(n28544), .Q(
        \pe11/ti_7t [2]) );
  DRNQHSV1 \pe2/pe5/q_reg[7]  ( .D(pov1[7]), .CK(clk), .RDN(n14021), .Q(
        \pe2/pvq [7]) );
  DRNQHSV1 \pe2/pe5/q_reg[5]  ( .D(pov1[5]), .CK(clk), .RDN(n28606), .Q(
        \pe2/pvq [5]) );
  DRNQHSV1 \pe3/pe5/q_reg[8]  ( .D(n14033), .CK(clk), .RDN(n28606), .Q(
        \pe3/pvq [8]) );
  DRNQHSV1 \pe3/pe5/q_reg[6]  ( .D(n29041), .CK(clk), .RDN(n28517), .Q(
        \pe3/pvq [6]) );
  DRNQHSV1 \pe3/pe5/q_reg[3]  ( .D(n29044), .CK(clk), .RDN(n28563), .Q(
        \pe3/pvq [3]) );
  DRNQHSV1 \pe4/pe5/q_reg[10]  ( .D(n28708), .CK(clk), .RDN(n28511), .Q(
        \pe4/pvq [10]) );
  DRNQHSV1 \pe4/pe5/q_reg[9]  ( .D(n14054), .CK(clk), .RDN(n28486), .Q(
        \pe4/pvq [9]) );
  DRNQHSV1 \pe4/pe5/q_reg[8]  ( .D(n28611), .CK(clk), .RDN(n28538), .Q(
        \pe4/pvq [8]) );
  DRNQHSV1 \pe4/pe5/q_reg[7]  ( .D(n28613), .CK(clk), .RDN(n28512), .Q(
        \pe4/pvq [7]) );
  DRNQHSV1 \pe4/pe5/q_reg[5]  ( .D(n29036), .CK(clk), .RDN(n28483), .Q(
        \pe4/pvq [5]) );
  DRNQHSV1 \pe4/pe5/q_reg[4]  ( .D(n14041), .CK(clk), .RDN(n28482), .Q(
        \pe4/pvq [4]) );
  DRNQHSV2 \pe5/pe5/q_reg[7]  ( .D(n28957), .CK(clk), .RDN(n28492), .Q(
        \pe5/pvq [7]) );
  DRNQHSV1 \pe5/pe5/q_reg[6]  ( .D(n28581), .CK(clk), .RDN(n28559), .Q(
        \pe5/pvq [6]) );
  DRNQHSV1 \pe5/pe5/q_reg[4]  ( .D(n28974), .CK(clk), .RDN(n28492), .Q(
        \pe5/pvq [4]) );
  DRNQHSV1 \pe5/pe14/q_reg[2]  ( .D(n28594), .CK(clk), .RDN(n28574), .Q(
        \pe5/ti_7t [2]) );
  DRNQHSV1 \pe6/pe5/q_reg[10]  ( .D(pov5[10]), .CK(clk), .RDN(n28503), .Q(
        \pe6/pvq [10]) );
  DRNQHSV1 \pe6/pe5/q_reg[9]  ( .D(pov5[9]), .CK(clk), .RDN(n28505), .Q(
        \pe6/pvq [9]) );
  DRNQHSV1 \pe6/pe5/q_reg[5]  ( .D(n28990), .CK(clk), .RDN(n28547), .Q(
        \pe6/pvq [5]) );
  DRNQHSV1 \pe6/pe14/q_reg[2]  ( .D(n28798), .CK(clk), .RDN(n28607), .Q(
        \pe6/ti_7t [2]) );
  DRNQHSV1 \pe7/pe5/q_reg[8]  ( .D(n28676), .CK(clk), .RDN(n28556), .Q(
        \pe7/pvq [8]) );
  DRNQHSV1 \pe7/pe5/q_reg[7]  ( .D(n29023), .CK(clk), .RDN(n28572), .Q(
        \pe7/pvq [7]) );
  DRNQHSV1 \pe9/pe5/q_reg[9]  ( .D(n29006), .CK(clk), .RDN(n28572), .Q(
        \pe9/pvq [9]) );
  DRNQHSV1 \pe9/pe5/q_reg[7]  ( .D(n29007), .CK(clk), .RDN(n28516), .Q(
        \pe9/pvq [7]) );
  DRNQHSV1 \pe9/pe5/q_reg[5]  ( .D(n28984), .CK(clk), .RDN(n14023), .Q(
        \pe9/pvq [5]) );
  DRNQHSV1 \pe9/pe14/q_reg[1]  ( .D(n28688), .CK(clk), .RDN(n28533), .Q(
        \pe9/ti_7t [1]) );
  DRNQHSV1 \pe10/pe5/q_reg[9]  ( .D(pov9[9]), .CK(clk), .RDN(n28563), .Q(
        \pe10/pvq [9]) );
  DRNQHSV1 \pe10/pe5/q_reg[7]  ( .D(n29000), .CK(clk), .RDN(n28477), .Q(
        \pe10/pvq [7]) );
  DRNQHSV1 \pe10/pe5/q_reg[5]  ( .D(n29001), .CK(clk), .RDN(n28442), .Q(
        \pe10/pvq [5]) );
  DRNQHSV1 \pe10/pe5/q_reg[4]  ( .D(n28961), .CK(clk), .RDN(n28459), .Q(
        \pe10/pvq [4]) );
  DRNQHSV1 \pe11/pe5/q_reg[6]  ( .D(n28997), .CK(clk), .RDN(n28439), .Q(
        \pe11/pvq [6]) );
  DRNQHSV1 \pe11/pe5/q_reg[4]  ( .D(n28959), .CK(clk), .RDN(n28564), .Q(
        \pe11/pvq [4]) );
  DRNQHSV1 \pe9/pe5/q_reg[1]  ( .D(n29012), .CK(clk), .RDN(n28504), .Q(
        \pe9/pvq [1]) );
  DRNQHSV1 \pe5/pe14/q_reg[3]  ( .D(n14848), .CK(clk), .RDN(n28596), .Q(
        \pe5/ti_7t [3]) );
  DRNQHSV1 \pe7/pe14/q_reg[2]  ( .D(n28808), .CK(clk), .RDN(n28439), .Q(
        \pe7/ti_7t [2]) );
  DRNQHSV1 \pe5/pe14/q_reg[1]  ( .D(n14474), .CK(clk), .RDN(n28514), .Q(
        \pe5/ti_7t [1]) );
  DRNQHSV1 \pe3/pe8/q_reg  ( .D(\pe3/ctrq ), .CK(clk), .RDN(n28563), .Q(ctro3)
         );
  DRNQHSV1 \pe8/pe14/q_reg[1]  ( .D(n28796), .CK(clk), .RDN(n28508), .Q(
        \pe8/ti_7t [1]) );
  DRNQHSV1 \pe3/pe5/q_reg[4]  ( .D(n29043), .CK(clk), .RDN(n28453), .Q(
        \pe3/pvq [4]) );
  DRNQHSV1 \pe3/pe14/q_reg[1]  ( .D(n26255), .CK(clk), .RDN(n28500), .Q(
        \pe3/ti_7t [1]) );
  DRNQHSV1 \pe6/pe14/q_reg[1]  ( .D(\pe6/ti_7[1] ), .CK(clk), .RDN(n28519), 
        .Q(\pe6/ti_7t [1]) );
  DRNQHSV1 \pe7/pe14/q_reg[1]  ( .D(n11858), .CK(clk), .RDN(n28553), .Q(
        \pe7/ti_7t [1]) );
  DRNQHSV2 \pe6/pe5/q_reg[8]  ( .D(n28989), .CK(clk), .RDN(n28493), .Q(
        \pe6/pvq [8]) );
  DRNQHSV1 \pe8/pe17/q_reg[8]  ( .D(\pe8/poht [8]), .CK(clk), .RDN(n28552), 
        .Q(poh8[8]) );
  DRNQHSV4 \pe6/pe5/q_reg[1]  ( .D(n28455), .CK(clk), .RDN(n28508), .Q(
        \pe6/pvq [1]) );
  DRNQHSV1 \pe8/pe17/q_reg[9]  ( .D(\pe8/poht [9]), .CK(clk), .RDN(n28568), 
        .Q(poh8[9]) );
  DRNQHSV2 \pe2/pe5/q_reg[1]  ( .D(n12023), .CK(clk), .RDN(n28477), .Q(
        \pe2/pvq [1]) );
  DRNQHSV4 \pe11/pe17/q_reg[14]  ( .D(\pe11/poht [14]), .CK(clk), .RDN(n28572), 
        .Q(poh11[14]) );
  DRNQHSV4 \pe9/pe5/q_reg[14]  ( .D(pov8[14]), .CK(clk), .RDN(n28445), .Q(
        \pe9/pvq [14]) );
  DRNQHSV4 \pe9/pe5/q_reg[13]  ( .D(n28994), .CK(clk), .RDN(n28489), .Q(
        \pe9/pvq [13]) );
  DRNQHSV2 \pe8/pe17/q_reg[6]  ( .D(\pe8/poht [6]), .CK(clk), .RDN(n28510), 
        .Q(poh8[6]) );
  DRNQHSV2 \pe8/pe17/q_reg[7]  ( .D(\pe8/poht [7]), .CK(clk), .RDN(n28439), 
        .Q(poh8[7]) );
  DRNQHSV1 \pe3/pe17/q_reg[9]  ( .D(\pe3/poht [9]), .CK(clk), .RDN(n28522), 
        .Q(poh3[9]) );
  DRNQHSV1 \pe3/pe17/q_reg[8]  ( .D(\pe3/poht [8]), .CK(clk), .RDN(n28557), 
        .Q(poh3[8]) );
  DRNQHSV1 \pe3/pe17/q_reg[3]  ( .D(\pe3/poht [3]), .CK(clk), .RDN(n28550), 
        .Q(poh3[3]) );
  DRNQHSV1 \pe3/pe17/q_reg[4]  ( .D(\pe3/poht [4]), .CK(clk), .RDN(n28487), 
        .Q(poh3[4]) );
  DRNQHSV1 \pe3/pe17/q_reg[7]  ( .D(\pe3/poht [7]), .CK(clk), .RDN(n28557), 
        .Q(poh3[7]) );
  DRNQHSV4 \pe7/pe8/q_reg  ( .D(n28876), .CK(clk), .RDN(n28558), .Q(ctro7) );
  DRNQHSV4 \pe10/pe8/q_reg  ( .D(n28811), .CK(clk), .RDN(n28568), .Q(ctro10)
         );
  DRNQHSV4 \pe11/pe17/q_reg[7]  ( .D(\pe11/poht [7]), .CK(clk), .RDN(n28482), 
        .Q(poh11[7]) );
  DRNQHSV4 \pe11/pe17/q_reg[5]  ( .D(\pe11/poht [5]), .CK(clk), .RDN(n28564), 
        .Q(poh11[5]) );
  DRNQHSV1 \pe2/pe17/q_reg[14]  ( .D(\pe2/poht [14]), .CK(clk), .RDN(n28450), 
        .Q(poh2[14]) );
  DRNQHSV1 \pe2/pe17/q_reg[12]  ( .D(\pe2/poht [12]), .CK(clk), .RDN(n28517), 
        .Q(poh2[12]) );
  DRNQHSV4 \pe1/pe1/q_reg[6]  ( .D(ai[11]), .CK(clk), .RDN(rst), .Q(
        \pe1/aot [11]) );
  DRNQHSV2 \pe5/pe5/q_reg[3]  ( .D(n29033), .CK(clk), .RDN(n28561), .Q(
        \pe5/pvq [3]) );
  DRNQHSV1 \pe1/pe17/q_reg[2]  ( .D(\pe1/poht [2]), .CK(clk), .RDN(n28544), 
        .Q(poh1[2]) );
  DRNQHSV4 \pe11/pe17/q_reg[8]  ( .D(\pe11/poht [8]), .CK(clk), .RDN(n28540), 
        .Q(poh11[8]) );
  DRNQHSV4 \pe11/pe17/q_reg[10]  ( .D(\pe11/poht [10]), .CK(clk), .RDN(n28564), 
        .Q(poh11[10]) );
  DRNQHSV4 \pe11/pe17/q_reg[12]  ( .D(\pe11/poht [12]), .CK(clk), .RDN(n28502), 
        .Q(poh11[12]) );
  DRNQHSV1 \pe3/pe17/q_reg[5]  ( .D(\pe3/poht [5]), .CK(clk), .RDN(n28519), 
        .Q(poh3[5]) );
  DRNQHSV4 \pe8/pe4/q_reg  ( .D(po7), .CK(clk), .RDN(n28502), .Q(\pe8/pq ) );
  DRNQHSV1 \pe4/pe4/q_reg  ( .D(po3), .CK(clk), .RDN(n28487), .Q(\pe4/pq ) );
  DRNQHSV4 \pe2/pe8/q_reg  ( .D(n28835), .CK(clk), .RDN(n28568), .Q(ctro2) );
  DRNQHSV2 \pe8/pe17/q_reg[10]  ( .D(\pe8/poht [10]), .CK(clk), .RDN(n28607), 
        .Q(poh8[10]) );
  DRNQHSV4 \pe10/pe13/q_reg  ( .D(\pe10/ti_1t ), .CK(clk), .RDN(n28514), .Q(
        \pe10/ti_1 ) );
  DRNQHSV2 \pe8/pe17/q_reg[15]  ( .D(\pe8/poht [15]), .CK(clk), .RDN(n28572), 
        .Q(poh8[15]) );
  DRNQHSV4 \pe7/pe5/q_reg[1]  ( .D(n28579), .CK(clk), .RDN(n28445), .Q(
        \pe7/pvq [1]) );
  DRNQHSV1 \pe8/pe17/q_reg[1]  ( .D(\pe8/poht [1]), .CK(clk), .RDN(n28487), 
        .Q(poh8[1]) );
  DRNQHSV1 \pe8/pe17/q_reg[13]  ( .D(\pe8/poht [13]), .CK(clk), .RDN(n28510), 
        .Q(poh8[13]) );
  DRNQHSV2 \pe8/pe17/q_reg[11]  ( .D(\pe8/poht [11]), .CK(clk), .RDN(n28453), 
        .Q(poh8[11]) );
  DSNHSV4 \pe8/pe7/q_reg  ( .D(n28789), .CK(clk), .SDN(n28444), .Q(n28623), 
        .QN(\pe8/ctrq ) );
  DSNHSV4 \pe8/pe2/q_reg[1]  ( .D(n28670), .CK(clk), .SDN(n28483), .Q(n28667), 
        .QN(\pe8/got [16]) );
  DRNQHSV4 \pe10/pe14/q_reg[1]  ( .D(n28666), .CK(clk), .RDN(n28527), .Q(
        \pe10/ti_7t [1]) );
  DRNQHSV2 \pe9/pe14/q_reg[12]  ( .D(n28580), .CK(clk), .RDN(n28562), .Q(
        \pe9/ti_7t [12]) );
  DRNQHSV4 \pe1/pe14/q_reg[3]  ( .D(n28481), .CK(clk), .RDN(n28542), .Q(
        \pe1/ti_7t [3]) );
  DRNQHSV4 \pe1/pe3/q_reg[1]  ( .D(bi[16]), .CK(clk), .RDN(n28492), .Q(bo1[16]) );
  DRNQHSV4 \pe1/pe3/q_reg[2]  ( .D(bi[15]), .CK(clk), .RDN(n28482), .Q(bo1[15]) );
  DRNQHSV4 \pe1/pe3/q_reg[10]  ( .D(bi[7]), .CK(clk), .RDN(n28507), .Q(bo1[7])
         );
  DRNQHSV4 \pe1/pe3/q_reg[8]  ( .D(bi[9]), .CK(clk), .RDN(n28503), .Q(bo1[9])
         );
  DRNQHSV4 \pe1/pe3/q_reg[9]  ( .D(bi[8]), .CK(clk), .RDN(rst), .Q(bo1[8]) );
  DRNQHSV4 \pe1/pe2/q_reg[9]  ( .D(gi[8]), .CK(clk), .RDN(rst), .Q(
        \pe1/got [8]) );
  DRNQHSV1 \pe1/pe17/q_reg[5]  ( .D(\pe1/poht [5]), .CK(clk), .RDN(n28516), 
        .Q(poh1[5]) );
  DRNQHSV4 \pe1/pe7/q_reg  ( .D(ctr), .CK(clk), .RDN(n28499), .Q(\pe1/ctrq )
         );
  DRNQHSV4 \pe1/pe1/q_reg[7]  ( .D(ai[10]), .CK(clk), .RDN(n28443), .Q(
        \pe1/aot [10]) );
  DRNQHSV4 \pe1/pe1/q_reg[9]  ( .D(ai[8]), .CK(clk), .RDN(n28606), .Q(
        \pe1/aot [8]) );
  DRNQHSV1 \pe9/pe17/q_reg[2]  ( .D(\pe9/poht [2]), .CK(clk), .RDN(n28551), 
        .Q(poh9[2]) );
  DRNQHSV1 \pe9/pe17/q_reg[3]  ( .D(\pe9/poht [3]), .CK(clk), .RDN(n28560), 
        .Q(poh9[3]) );
  DRNQHSV4 \pe1/pe1/q_reg[13]  ( .D(ai[4]), .CK(clk), .RDN(rst), .Q(
        \pe1/aot [4]) );
  DRNQHSV4 \pe1/pe1/q_reg[11]  ( .D(ai[6]), .CK(clk), .RDN(rst), .Q(
        \pe1/aot [6]) );
  DRNQHSV4 \pe4/pe14/q_reg[1]  ( .D(n28653), .CK(clk), .RDN(n28446), .Q(
        \pe4/ti_7t [1]) );
  DRNQHSV4 \pe1/pe2/q_reg[5]  ( .D(gi[12]), .CK(clk), .RDN(n28607), .Q(
        \pe1/got [12]) );
  DRNQHSV4 \pe1/pe2/q_reg[7]  ( .D(gi[10]), .CK(clk), .RDN(rst), .Q(
        \pe1/got [10]) );
  DRNQHSV4 \pe1/pe2/q_reg[6]  ( .D(gi[11]), .CK(clk), .RDN(n28606), .Q(
        \pe1/got [11]) );
  DRNQHSV4 \pe1/pe2/q_reg[13]  ( .D(gi[4]), .CK(clk), .RDN(n28601), .Q(
        \pe1/got [4]) );
  DRNQHSV4 \pe1/pe2/q_reg[11]  ( .D(gi[6]), .CK(clk), .RDN(n28601), .Q(
        \pe1/got [6]) );
  DRNQHSV4 \pe1/pe1/q_reg[8]  ( .D(ai[9]), .CK(clk), .RDN(n28440), .Q(
        \pe1/aot [9]) );
  DRNQHSV1 \pe9/pe17/q_reg[7]  ( .D(\pe9/poht [7]), .CK(clk), .RDN(n28567), 
        .Q(poh9[7]) );
  DRNQHSV1 \pe9/pe17/q_reg[4]  ( .D(\pe9/poht [4]), .CK(clk), .RDN(n28555), 
        .Q(poh9[4]) );
  DRNQHSV1 \pe9/pe17/q_reg[1]  ( .D(\pe9/poht [1]), .CK(clk), .RDN(n28531), 
        .Q(poh9[1]) );
  DRNQHSV2 \pe11/pe14/q_reg[9]  ( .D(n28464), .CK(clk), .RDN(n28489), .Q(
        \pe11/ti_7t [9]) );
  DRNQHSV1 \pe9/pe17/q_reg[12]  ( .D(\pe9/poht [12]), .CK(clk), .RDN(n28494), 
        .Q(poh9[12]) );
  DRNQHSV4 \pe11/pe8/q_reg  ( .D(n28639), .CK(clk), .RDN(n28501), .Q(ctro11)
         );
  DRNQHSV4 \pe3/pe14/q_reg[4]  ( .D(n16112), .CK(clk), .RDN(n28439), .Q(
        \pe3/ti_7t [4]) );
  DRNQHSV4 \pe1/pe14/q_reg[1]  ( .D(n28622), .CK(clk), .RDN(n28546), .Q(
        \pe1/ti_7t [1]) );
  DRNQHSV4 \pe4/pe5/q_reg[1]  ( .D(n28619), .CK(clk), .RDN(n28546), .Q(
        \pe4/pvq [1]) );
  DRNQHSV4 \pe1/pe2/q_reg[3]  ( .D(gi[14]), .CK(clk), .RDN(n28607), .Q(
        \pe1/got [14]) );
  DRNQHSV4 \pe6/pe14/q_reg[10]  ( .D(n28662), .CK(clk), .RDN(n28493), .Q(
        \pe6/ti_7t [10]) );
  DRNQHSV4 \pe1/pe2/q_reg[4]  ( .D(gi[13]), .CK(clk), .RDN(n28441), .Q(
        \pe1/got [13]) );
  DRNQHSV2 \pe11/pe14/q_reg[13]  ( .D(n28922), .CK(clk), .RDN(n28501), .Q(
        \pe11/ti_7t [13]) );
  DRNQHSV2 \pe3/pe14/q_reg[15]  ( .D(n28661), .CK(clk), .RDN(n28565), .Q(
        \pe3/ti_7t [15]) );
  DRNQHSV2 \pe1/pe14/q_reg[4]  ( .D(n28635), .CK(clk), .RDN(n28444), .Q(
        \pe1/ti_7t [4]) );
  DRNQHSV2 \pe9/pe14/q_reg[2]  ( .D(n11863), .CK(clk), .RDN(n28543), .Q(
        \pe9/ti_7t [2]) );
  DRNQHSV4 \pe3/pe14/q_reg[11]  ( .D(n28584), .CK(clk), .RDN(n28509), .Q(
        \pe3/ti_7t [11]) );
  DRNQHSV2 \pe9/pe16/q_reg[1]  ( .D(n28669), .CK(clk), .RDN(n28486), .Q(
        go9[16]) );
  DRNQHSV1 \pe11/pe14/q_reg[8]  ( .D(n28935), .CK(clk), .RDN(n28572), .Q(
        \pe11/ti_7t [8]) );
  DRNQHSV2 \pe3/pe17/q_reg[11]  ( .D(\pe3/poht [11]), .CK(clk), .RDN(n28502), 
        .Q(poh3[11]) );
  DRNQHSV4 \pe5/pe3/q_reg[1]  ( .D(bo4[16]), .CK(clk), .RDN(n28563), .Q(
        bo5[16]) );
  DRNQHSV2 \pe4/pe15/q_reg[1]  ( .D(n28683), .CK(clk), .RDN(n28524), .Q(
        ao4[16]) );
  DRNQHSV1 \pe7/pe17/q_reg[12]  ( .D(\pe7/poht [12]), .CK(clk), .RDN(n28559), 
        .Q(poh7[12]) );
  DRNQHSV2 \pe8/pe6/q_reg[9]  ( .D(poh7[9]), .CK(clk), .RDN(n28511), .Q(
        \pe8/phq [9]) );
  DRNQHSV1 \pe9/pe17/q_reg[13]  ( .D(\pe9/poht [13]), .CK(clk), .RDN(n28492), 
        .Q(poh9[13]) );
  DRNQHSV1 \pe9/pe17/q_reg[14]  ( .D(\pe9/poht [14]), .CK(clk), .RDN(n28527), 
        .Q(poh9[14]) );
  DRNQHSV1 \pe9/pe17/q_reg[5]  ( .D(\pe9/poht [5]), .CK(clk), .RDN(n28449), 
        .Q(poh9[5]) );
  DRNQHSV1 \pe9/pe17/q_reg[8]  ( .D(\pe9/poht [8]), .CK(clk), .RDN(n28602), 
        .Q(poh9[8]) );
  DRNQHSV1 \pe10/pe4/q_reg  ( .D(po9), .CK(clk), .RDN(n28543), .Q(\pe10/pq )
         );
  DRNQHSV1 \pe9/pe17/q_reg[6]  ( .D(\pe9/poht [6]), .CK(clk), .RDN(n28565), 
        .Q(poh9[6]) );
  DRNQHSV1 \pe5/pe5/q_reg[8]  ( .D(n29031), .CK(clk), .RDN(n28567), .Q(
        \pe5/pvq [8]) );
  DSNHSV1 \pe8/pe14/q_reg[14]  ( .D(n28692), .CK(clk), .SDN(n28530), .Q(n28685) );
  DRNQHSV2 \pe10/pe17/q_reg[13]  ( .D(\pe10/poht [13]), .CK(clk), .RDN(n28514), 
        .Q(poh10[13]) );
  DRNQHSV1 \pe10/pe14/q_reg[9]  ( .D(n28585), .CK(clk), .RDN(n28548), .Q(
        \pe10/ti_7t [9]) );
  DRNQHSV4 \pe1/pe2/q_reg[15]  ( .D(gi[2]), .CK(clk), .RDN(n28604), .Q(
        \pe1/got [2]) );
  DRNQHSV1 \pe6/pe17/q_reg[1]  ( .D(\pe6/poht [1]), .CK(clk), .RDN(n28555), 
        .Q(poh6[1]) );
  DRNQHSV1 \pe7/pe4/q_reg  ( .D(po6), .CK(clk), .RDN(n28458), .Q(\pe7/pq ) );
  DRNQHSV1 \pe6/pe17/q_reg[13]  ( .D(\pe6/poht [13]), .CK(clk), .RDN(n28476), 
        .Q(poh6[13]) );
  DRNQHSV1 \pe3/pe5/q_reg[14]  ( .D(n28967), .CK(clk), .RDN(n28508), .Q(
        \pe3/pvq [14]) );
  DRNQHSV4 \pe9/pe14/q_reg[9]  ( .D(n28437), .CK(clk), .RDN(n28596), .Q(
        \pe9/ti_7t [9]) );
  DRNQHSV1 \pe3/pe14/q_reg[6]  ( .D(n28707), .CK(clk), .RDN(n28547), .Q(
        \pe3/ti_7t [6]) );
  DRNQHSV1 \pe11/pe14/q_reg[5]  ( .D(n14043), .CK(clk), .RDN(n28509), .Q(
        \pe11/ti_7t [5]) );
  DRNQHSV4 \pe8/pe14/q_reg[12]  ( .D(n28698), .CK(clk), .RDN(n28552), .Q(
        \pe8/ti_7t [12]) );
  DRNQHSV1 \pe5/pe17/q_reg[15]  ( .D(\pe5/poht [15]), .CK(clk), .RDN(n28541), 
        .Q(poh5[15]) );
  DRNQHSV1 \pe9/pe17/q_reg[10]  ( .D(\pe9/poht [10]), .CK(clk), .RDN(n28605), 
        .Q(poh9[10]) );
  DRNQHSV1 \pe9/pe17/q_reg[15]  ( .D(\pe9/poht [15]), .CK(clk), .RDN(n28443), 
        .Q(poh9[15]) );
  DRNQHSV2 \pe4/pe6/q_reg[13]  ( .D(poh3[13]), .CK(clk), .RDN(n28545), .Q(
        \pe4/phq [13]) );
  DRNQHSV2 \pe3/pe5/q_reg[1]  ( .D(n28454), .CK(clk), .RDN(n28510), .Q(
        \pe3/pvq [1]) );
  DRNQHSV2 \pe10/pe17/q_reg[4]  ( .D(\pe10/poht [4]), .CK(clk), .RDN(n28444), 
        .Q(poh10[4]) );
  DSNHSV1 \pe9/pe5/q_reg[8]  ( .D(n28815), .CK(clk), .SDN(n28444), .QN(
        \pe9/pvq [8]) );
  DSNHSV1 \pe9/pe5/q_reg[10]  ( .D(n28690), .CK(clk), .SDN(n28445), .QN(
        \pe9/pvq [10]) );
  DSNHSV2 \pe11/pe5/q_reg[9]  ( .D(n28694), .CK(clk), .SDN(n28444), .QN(
        \pe11/pvq [9]) );
  DRNQHSV1 \pe6/pe14/q_reg[7]  ( .D(\pe6/ti_7[7] ), .CK(clk), .RDN(n28553), 
        .Q(\pe6/ti_7t [7]) );
  DRNQHSV1 \pe4/pe17/q_reg[11]  ( .D(\pe4/poht [11]), .CK(clk), .RDN(n28487), 
        .Q(poh4[11]) );
  DRNQHSV1 \pe7/pe14/q_reg[12]  ( .D(n14030), .CK(clk), .RDN(n28500), .Q(
        \pe7/ti_7t [12]) );
  DRNQHSV1 \pe4/pe17/q_reg[7]  ( .D(\pe4/poht [7]), .CK(clk), .RDN(n28550), 
        .Q(poh4[7]) );
  DRNQHSV1 \pe2/pe17/q_reg[11]  ( .D(\pe2/poht [11]), .CK(clk), .RDN(n28529), 
        .Q(poh2[11]) );
  DRNQHSV1 \pe2/pe17/q_reg[8]  ( .D(\pe2/poht [8]), .CK(clk), .RDN(n28458), 
        .Q(poh2[8]) );
  DRNQHSV1 \pe7/pe14/q_reg[7]  ( .D(n14067), .CK(clk), .RDN(n28476), .Q(
        \pe7/ti_7t [7]) );
  DRNQHSV1 \pe3/pe17/q_reg[12]  ( .D(\pe3/poht [12]), .CK(clk), .RDN(n28537), 
        .Q(poh3[12]) );
  DRNQHSV1 \pe2/pe17/q_reg[10]  ( .D(\pe2/poht [10]), .CK(clk), .RDN(n28567), 
        .Q(poh2[10]) );
  DRNQHSV1 \pe2/pe17/q_reg[13]  ( .D(\pe2/poht [13]), .CK(clk), .RDN(n28529), 
        .Q(poh2[13]) );
  DRNQHSV1 \pe1/pe14/q_reg[15]  ( .D(n28600), .CK(clk), .RDN(n28559), .Q(
        \pe1/ti_7t [15]) );
  DRNQHSV1 \pe8/pe14/q_reg[9]  ( .D(n28631), .CK(clk), .RDN(n28518), .Q(
        \pe8/ti_7t [9]) );
  DRNQHSV4 \pe3/pe3/q_reg[11]  ( .D(bo2[6]), .CK(clk), .RDN(n28518), .Q(bo3[6]) );
  DRNQHSV1 \pe2/pe17/q_reg[6]  ( .D(\pe2/poht [6]), .CK(clk), .RDN(n28502), 
        .Q(poh2[6]) );
  DRNQHSV1 \pe22/q_reg  ( .D(po11), .CK(clk), .RDN(n28572), .Q(po[1]) );
  DRNQHSV1 \pe6/pe16/q_reg[2]  ( .D(\pe6/got [15]), .CK(clk), .RDN(n28573), 
        .Q(go6[15]) );
  DSNHSV1 \pe8/pe16/q_reg[9]  ( .D(n28655), .CK(clk), .SDN(n28444), .QN(go8[8]) );
  DSNHSV1 \pe3/pe16/q_reg[1]  ( .D(n28929), .CK(clk), .SDN(n28501), .QN(
        go3[16]) );
  DSNHSV4 \pe10/pe14/q_reg[7]  ( .D(n28675), .CK(clk), .SDN(n28597), .QN(
        \pe10/ti_7t [7]) );
  DRNQHSV2 \pe9/pe16/q_reg[6]  ( .D(n28423), .CK(clk), .RDN(n28554), .Q(
        go9[11]) );
  DRNQHSV1 \pe4/pe17/q_reg[12]  ( .D(\pe4/poht [12]), .CK(clk), .RDN(n28510), 
        .Q(poh4[12]) );
  DRNQHSV2 \pe8/pe16/q_reg[1]  ( .D(n25523), .CK(clk), .RDN(n28556), .Q(
        go8[16]) );
  DRNQHSV2 \pe3/pe16/q_reg[2]  ( .D(n26240), .CK(clk), .RDN(n28564), .Q(
        go3[15]) );
  DRNQHSV2 \pe4/pe16/q_reg[14]  ( .D(n28626), .CK(clk), .RDN(n28528), .Q(
        go4[3]) );
  DRNQHSV2 \pe4/pe15/q_reg[3]  ( .D(n28660), .CK(clk), .RDN(n28513), .Q(
        ao4[14]) );
  DRNQHSV1 \pe7/pe5/q_reg[5]  ( .D(n28678), .CK(clk), .RDN(n28520), .Q(
        \pe7/pvq [5]) );
  DSNHSV2 \pe11/pe5/q_reg[7]  ( .D(n28672), .CK(clk), .SDN(n28445), .QN(
        \pe11/pvq [7]) );
  DRNQHSV2 \pe9/pe17/q_reg[9]  ( .D(\pe9/poht [9]), .CK(clk), .RDN(n14023), 
        .Q(poh9[9]) );
  DRNQHSV4 \pe3/pe17/q_reg[10]  ( .D(\pe3/poht [10]), .CK(clk), .RDN(n28547), 
        .Q(poh3[10]) );
  DRNQHSV2 \pe4/pe17/q_reg[2]  ( .D(\pe4/poht [2]), .CK(clk), .RDN(n28545), 
        .Q(poh4[2]) );
  DRNQHSV2 \pe9/pe17/q_reg[11]  ( .D(\pe9/poht [11]), .CK(clk), .RDN(n28577), 
        .Q(poh9[11]) );
  DRNQHSV2 \pe9/pe16/q_reg[3]  ( .D(n28928), .CK(clk), .RDN(n28484), .Q(
        go9[14]) );
  DRNQHSV1 \pe1/pe17/q_reg[12]  ( .D(\pe1/poht [12]), .CK(clk), .RDN(n28544), 
        .Q(poh1[12]) );
  DRNQHSV1 \pe4/pe17/q_reg[15]  ( .D(\pe4/poht [15]), .CK(clk), .RDN(n28510), 
        .Q(poh4[15]) );
  DRNQHSV1 \pe11/pe14/q_reg[1]  ( .D(n28629), .CK(clk), .RDN(n28570), .Q(
        \pe11/ti_7t [1]) );
  DRNHSV2 \pe8/pe2/q_reg[2]  ( .D(go7[15]), .CK(clk), .RDN(n28524), .Q(n28695), 
        .QN(n28646) );
  DRNQHSV1 \pe4/pe14/q_reg[9]  ( .D(n27877), .CK(clk), .RDN(n28505), .Q(
        \pe4/ti_7t [9]) );
  DRNQHSV1 \pe1/pe17/q_reg[4]  ( .D(\pe1/poht [4]), .CK(clk), .RDN(n28505), 
        .Q(poh1[4]) );
  DRNQHSV1 \pe7/pe14/q_reg[6]  ( .D(n28466), .CK(clk), .RDN(n28546), .Q(
        \pe7/ti_7t [6]) );
  DRNQHSV2 \pe10/pe14/q_reg[6]  ( .D(n20074), .CK(clk), .RDN(n28601), .Q(
        \pe10/ti_7t [6]) );
  DRNQHSV4 \pe5/pe8/q_reg  ( .D(n28682), .CK(clk), .RDN(n28443), .Q(ctro5) );
  DRNQHSV2 \pe5/pe17/q_reg[8]  ( .D(\pe5/poht [8]), .CK(clk), .RDN(n28570), 
        .Q(poh5[8]) );
  DSNHSV2 \pe10/pe14/q_reg[10]  ( .D(n28674), .CK(clk), .SDN(n28445), .QN(
        \pe10/ti_7t [10]) );
  DRNQHSV1 \pe2/pe17/q_reg[5]  ( .D(\pe2/poht [5]), .CK(clk), .RDN(n28453), 
        .Q(poh2[5]) );
  DRNQHSV2 \pe11/pe4/q_reg  ( .D(po10), .CK(clk), .RDN(n28569), .Q(\pe11/pq )
         );
  DRNQHSV1 \pe2/pe14/q_reg[8]  ( .D(n21816), .CK(clk), .RDN(n28571), .Q(
        \pe2/ti_7t [8]) );
  DRNQHSV1 \pe3/pe4/q_reg  ( .D(po2), .CK(clk), .RDN(n28533), .Q(\pe3/pq ) );
  DRNQHSV1 \pe2/pe5/q_reg[10]  ( .D(n28968), .CK(clk), .RDN(n28515), .Q(
        \pe2/pvq [10]) );
  DRNQHSV1 \pe10/pe14/q_reg[15]  ( .D(n23219), .CK(clk), .RDN(n28605), .Q(
        \pe10/ti_7t [15]) );
  DRNQHSV1 \pe1/pe17/q_reg[7]  ( .D(\pe1/poht [7]), .CK(clk), .RDN(n28518), 
        .Q(poh1[7]) );
  DSNHSV4 \pe11/pe5/q_reg[8]  ( .D(n28431), .CK(clk), .SDN(n28445), .QN(
        \pe11/pvq [8]) );
  DRNQHSV4 \pe9/pe14/q_reg[15]  ( .D(n28943), .CK(clk), .RDN(n28447), .Q(
        \pe9/ti_7t [15]) );
  DRNQHSV1 \pe2/pe17/q_reg[7]  ( .D(\pe2/poht [7]), .CK(clk), .RDN(n28564), 
        .Q(poh2[7]) );
  DRNQHSV1 \pe8/pe17/q_reg[2]  ( .D(\pe8/poht [2]), .CK(clk), .RDN(n28569), 
        .Q(poh8[2]) );
  DRNQHSV1 \pe7/pe17/q_reg[13]  ( .D(\pe7/poht [13]), .CK(clk), .RDN(n28571), 
        .Q(poh7[13]) );
  DRNQHSV1 \pe1/pe17/q_reg[14]  ( .D(\pe1/poht [14]), .CK(clk), .RDN(n28497), 
        .Q(poh1[14]) );
  DRNQHSV1 \pe1/pe17/q_reg[1]  ( .D(\pe1/poht [1]), .CK(clk), .RDN(n28530), 
        .Q(poh1[1]) );
  DRNQHSV2 \pe11/pe5/q_reg[1]  ( .D(n28704), .CK(clk), .RDN(n28521), .Q(
        \pe11/pvq [1]) );
  DRNQHSV1 \pe1/pe17/q_reg[9]  ( .D(\pe1/poht [9]), .CK(clk), .RDN(n28545), 
        .Q(poh1[9]) );
  DRNQHSV1 \pe7/pe17/q_reg[10]  ( .D(\pe7/poht [10]), .CK(clk), .RDN(n28445), 
        .Q(poh7[10]) );
  DRNQHSV1 \pe2/pe14/q_reg[13]  ( .D(n27731), .CK(clk), .RDN(n28515), .Q(
        \pe2/ti_7t [13]) );
  DRNQHSV4 \pe5/pe5/q_reg[1]  ( .D(n15428), .CK(clk), .RDN(n28519), .Q(
        \pe5/pvq [1]) );
  DRNQHSV2 \pe6/pe17/q_reg[14]  ( .D(\pe6/poht [14]), .CK(clk), .RDN(n28477), 
        .Q(poh6[14]) );
  DRNQHSV2 \pe6/pe17/q_reg[8]  ( .D(\pe6/poht [8]), .CK(clk), .RDN(n28553), 
        .Q(poh6[8]) );
  DRNQHSV2 \pe8/pe17/q_reg[14]  ( .D(\pe8/poht [14]), .CK(clk), .RDN(n14023), 
        .Q(poh8[14]) );
  DRNQHSV4 \pe8/pe5/q_reg[1]  ( .D(n28797), .CK(clk), .RDN(n28518), .Q(
        \pe8/pvq [1]) );
  DRNQHSV2 \pe5/pe17/q_reg[7]  ( .D(\pe5/poht [7]), .CK(clk), .RDN(n28522), 
        .Q(poh5[7]) );
  DRNQHSV2 \pe5/pe17/q_reg[6]  ( .D(\pe5/poht [6]), .CK(clk), .RDN(n28450), 
        .Q(poh5[6]) );
  DRNQHSV2 \pe5/pe17/q_reg[9]  ( .D(\pe5/poht [9]), .CK(clk), .RDN(n28507), 
        .Q(poh5[9]) );
  DRNQHSV2 \pe5/pe17/q_reg[12]  ( .D(\pe5/poht [12]), .CK(clk), .RDN(n28538), 
        .Q(poh5[12]) );
  DRNQHSV2 \pe5/pe17/q_reg[4]  ( .D(\pe5/poht [4]), .CK(clk), .RDN(n28536), 
        .Q(poh5[4]) );
  DRNQHSV2 \pe10/pe17/q_reg[15]  ( .D(\pe10/poht [15]), .CK(clk), .RDN(n28484), 
        .Q(poh10[15]) );
  DRNQHSV2 \pe2/pe5/q_reg[3]  ( .D(n29050), .CK(clk), .RDN(n28536), .Q(
        \pe2/pvq [3]) );
  DRNQHSV2 \pe3/pe17/q_reg[1]  ( .D(\pe3/poht [1]), .CK(clk), .RDN(n28506), 
        .Q(poh3[1]) );
  DRNQHSV2 \pe3/pe17/q_reg[2]  ( .D(\pe3/poht [2]), .CK(clk), .RDN(n28559), 
        .Q(poh3[2]) );
  DRNQHSV2 \pe10/pe17/q_reg[12]  ( .D(\pe10/poht [12]), .CK(clk), .RDN(n28531), 
        .Q(poh10[12]) );
  DRNQHSV2 \pe5/pe17/q_reg[13]  ( .D(\pe5/poht [13]), .CK(clk), .RDN(n28566), 
        .Q(poh5[13]) );
  DRNQHSV1 \pe5/pe17/q_reg[2]  ( .D(\pe5/poht [2]), .CK(clk), .RDN(n28522), 
        .Q(poh5[2]) );
  DRNHSV4 \pe8/pe12/q_reg[1]  ( .D(n28884), .CK(clk), .RDN(n28597), .Q(n28663), 
        .QN(n28813) );
  DRNQHSV2 \pe8/pe17/q_reg[5]  ( .D(\pe8/poht [5]), .CK(clk), .RDN(n28503), 
        .Q(poh8[5]) );
  DRNQHSV2 \pe10/pe17/q_reg[14]  ( .D(\pe10/poht [14]), .CK(clk), .RDN(n28487), 
        .Q(poh10[14]) );
  DRNQHSV2 \pe6/pe17/q_reg[5]  ( .D(\pe6/poht [5]), .CK(clk), .RDN(n28557), 
        .Q(poh6[5]) );
  DRNQHSV2 \pe10/pe17/q_reg[2]  ( .D(\pe10/poht [2]), .CK(clk), .RDN(n28440), 
        .Q(poh10[2]) );
  DRNQHSV4 \pe6/pe17/q_reg[12]  ( .D(\pe6/poht [12]), .CK(clk), .RDN(n28605), 
        .Q(poh6[12]) );
  DRNQHSV2 \pe6/pe17/q_reg[15]  ( .D(\pe6/poht [15]), .CK(clk), .RDN(n28445), 
        .Q(poh6[15]) );
  DRNQHSV4 \pe10/pe17/q_reg[10]  ( .D(\pe10/poht [10]), .CK(clk), .RDN(n28605), 
        .Q(poh10[10]) );
  DRNQHSV2 \pe8/pe17/q_reg[4]  ( .D(\pe8/poht [4]), .CK(clk), .RDN(n28502), 
        .Q(poh8[4]) );
  DRNQHSV2 \pe7/pe17/q_reg[14]  ( .D(\pe7/poht [14]), .CK(clk), .RDN(n28512), 
        .Q(poh7[14]) );
  DRNQHSV4 \pe10/pe17/q_reg[7]  ( .D(\pe10/poht [7]), .CK(clk), .RDN(n28490), 
        .Q(poh10[7]) );
  DRNQHSV2 \pe8/pe17/q_reg[12]  ( .D(\pe8/poht [12]), .CK(clk), .RDN(n28458), 
        .Q(poh8[12]) );
  DRNQHSV4 \pe5/pe17/q_reg[1]  ( .D(\pe5/poht [1]), .CK(clk), .RDN(n14021), 
        .Q(poh5[1]) );
  DRNQHSV1 \pe1/pe17/q_reg[10]  ( .D(\pe1/poht [10]), .CK(clk), .RDN(n28521), 
        .Q(poh1[10]) );
  DRNQHSV1 \pe2/pe4/q_reg  ( .D(po1), .CK(clk), .RDN(n28596), .Q(\pe2/pq ) );
  DRNQHSV4 \pe6/pe17/q_reg[7]  ( .D(\pe6/poht [7]), .CK(clk), .RDN(n28487), 
        .Q(poh6[7]) );
  DRNQHSV2 \pe6/pe17/q_reg[10]  ( .D(\pe6/poht [10]), .CK(clk), .RDN(n28561), 
        .Q(poh6[10]) );
  DRNQHSV2 \pe5/pe17/q_reg[14]  ( .D(\pe5/poht [14]), .CK(clk), .RDN(n28510), 
        .Q(poh5[14]) );
  INHSV4 U12493 ( .I(n12309), .ZN(n20928) );
  INHSV4 U12494 ( .I(n14478), .ZN(n13992) );
  NOR2HSV4 U12495 ( .A1(n12194), .A2(n19947), .ZN(n12193) );
  NAND2HSV4 U12496 ( .A1(n12193), .A2(n19951), .ZN(n19963) );
  CLKNAND2HSV4 U12497 ( .A1(n14458), .A2(n14457), .ZN(n28455) );
  NAND3HSV2 U12498 ( .A1(n14572), .A2(n14488), .A3(n14573), .ZN(n14489) );
  BUFHSV4 U12499 ( .I(\pe5/got [1]), .Z(n28640) );
  CLKNAND2HSV2 U12500 ( .A1(n13061), .A2(n13060), .ZN(n13062) );
  OAI21HSV2 U12501 ( .A1(n13757), .A2(n13758), .B(n13759), .ZN(\pe5/poht [10])
         );
  NAND2HSV4 U12502 ( .A1(n28946), .A2(n24636), .ZN(n23952) );
  NAND2HSV2 U12503 ( .A1(n21464), .A2(n21463), .ZN(n28946) );
  CLKNAND2HSV2 U12504 ( .A1(n28473), .A2(n14072), .ZN(n23270) );
  CLKXOR2HSV2 U12505 ( .A1(n23270), .A2(n23269), .Z(n23271) );
  CLKNAND2HSV2 U12506 ( .A1(n25137), .A2(\pe11/got [9]), .ZN(n24740) );
  XNOR2HSV2 U12507 ( .A1(n24740), .A2(n24739), .ZN(n24742) );
  INHSV4 U12508 ( .I(n16184), .ZN(n16185) );
  INHSV4 U12509 ( .I(n20868), .ZN(n20862) );
  CLKNAND2HSV4 U12510 ( .A1(n21062), .A2(n21063), .ZN(n12127) );
  CLKNAND2HSV8 U12511 ( .A1(n29006), .A2(n22129), .ZN(n18786) );
  CLKNAND2HSV8 U12512 ( .A1(n18786), .A2(n18785), .ZN(n21322) );
  XOR2HSV4 U12513 ( .A1(n21212), .A2(n12012), .Z(n21213) );
  NAND2HSV2 U12514 ( .A1(n17785), .A2(\pe2/bq[11] ), .ZN(n17786) );
  CLKXOR2HSV2 U12515 ( .A1(n17787), .A2(n17786), .Z(n17788) );
  CLKNAND2HSV4 U12516 ( .A1(n12654), .A2(n21424), .ZN(\pe5/ti_7[10] ) );
  OR2HSV8 U12517 ( .A1(n18604), .A2(n28085), .Z(n18605) );
  CLKNAND2HSV4 U12518 ( .A1(n21693), .A2(n21641), .ZN(n22080) );
  CLKNAND2HSV8 U12519 ( .A1(n22080), .A2(n22079), .ZN(n21815) );
  NAND2HSV2 U12520 ( .A1(n27106), .A2(n28647), .ZN(n21569) );
  NAND2HSV0 U12521 ( .A1(n11801), .A2(n11800), .ZN(n21884) );
  INHSV2 U12522 ( .I(n25357), .ZN(n11800) );
  NOR2HSV2 U12523 ( .A1(n28950), .A2(n11802), .ZN(n11801) );
  CLKNAND2HSV4 U12524 ( .A1(n23445), .A2(n17767), .ZN(n11802) );
  CLKNHSV6 U12525 ( .I(\pe6/ti_1 ), .ZN(n18955) );
  CLKNAND2HSV4 U12526 ( .A1(\pe6/bq[15] ), .A2(\pe6/aot [15]), .ZN(n14124) );
  NAND2HSV4 U12527 ( .A1(n19992), .A2(n19940), .ZN(n19941) );
  CLKNAND2HSV2 U12528 ( .A1(n28936), .A2(\pe11/got [9]), .ZN(n12305) );
  CLKNAND2HSV2 U12529 ( .A1(n28473), .A2(n24636), .ZN(n24694) );
  NAND2HSV2 U12530 ( .A1(n18841), .A2(n18842), .ZN(n11911) );
  INHSV4 U12531 ( .I(n11803), .ZN(n18842) );
  NAND2HSV4 U12532 ( .A1(n19992), .A2(n28695), .ZN(n11803) );
  NOR2HSV4 U12533 ( .A1(n21970), .A2(n21969), .ZN(n21972) );
  NAND2HSV4 U12534 ( .A1(n21972), .A2(n21971), .ZN(n26925) );
  INHSV4 U12535 ( .I(n14209), .ZN(n14207) );
  CLKNAND2HSV4 U12536 ( .A1(n14241), .A2(n14240), .ZN(n14243) );
  BUFHSV8 U12537 ( .I(n26634), .Z(n26752) );
  CLKBUFHSV12 U12538 ( .I(n24966), .Z(n11804) );
  CLKNAND2HSV4 U12539 ( .A1(n14119), .A2(n25647), .ZN(n14178) );
  CLKNAND2HSV4 U12540 ( .A1(n14178), .A2(n14285), .ZN(n14147) );
  INHSV2 U12541 ( .I(n21941), .ZN(n20355) );
  CLKNAND2HSV2 U12542 ( .A1(n20356), .A2(n20355), .ZN(n20359) );
  NAND2HSV2 U12543 ( .A1(n13040), .A2(n13038), .ZN(n13041) );
  CLKNAND2HSV4 U12544 ( .A1(n29037), .A2(n23664), .ZN(n15147) );
  CLKNAND2HSV8 U12545 ( .A1(n15147), .A2(n15146), .ZN(n15241) );
  INHSV2 U12546 ( .I(n14643), .ZN(n24637) );
  INHSV8 U12547 ( .I(n21643), .ZN(n17829) );
  CLKXOR2HSV4 U12548 ( .A1(n21568), .A2(n21569), .Z(n12981) );
  CLKNAND2HSV2 U12549 ( .A1(n15853), .A2(n25131), .ZN(n15618) );
  OAI21HSV2 U12550 ( .A1(n13820), .A2(n13821), .B(n13822), .ZN(\pe5/poht [11])
         );
  CLKNAND2HSV2 U12551 ( .A1(n24975), .A2(\pe11/got [9]), .ZN(n20383) );
  NAND2HSV4 U12552 ( .A1(n20455), .A2(n20454), .ZN(n20499) );
  INHSV4 U12553 ( .I(n20499), .ZN(n20502) );
  INHSV4 U12554 ( .I(n27904), .ZN(n27999) );
  OR2HSV2 U12555 ( .A1(n27999), .A2(n28000), .Z(n25077) );
  INHSV4 U12556 ( .I(n12319), .ZN(n18270) );
  XNOR2HSV4 U12557 ( .A1(n11806), .A2(n11805), .ZN(n21639) );
  XNOR2HSV4 U12558 ( .A1(n21216), .A2(n21215), .ZN(n11805) );
  AOI22HSV4 U12559 ( .A1(n21176), .A2(n21177), .B1(n21179), .B2(n21178), .ZN(
        n11806) );
  CLKNHSV6 U12560 ( .I(n19831), .ZN(n19840) );
  NAND2HSV4 U12561 ( .A1(n23320), .A2(n23319), .ZN(n24957) );
  NAND2HSV2 U12562 ( .A1(n24957), .A2(\pe11/got [9]), .ZN(n24958) );
  INHSV8 U12563 ( .I(\pe6/ctrq ), .ZN(n14048) );
  INHSV6 U12564 ( .I(n14048), .ZN(n14220) );
  NOR2HSV8 U12565 ( .A1(n16712), .A2(n16711), .ZN(n16880) );
  INHSV6 U12566 ( .I(n16880), .ZN(n16837) );
  NAND2HSV4 U12567 ( .A1(n28611), .A2(n15333), .ZN(n15906) );
  NAND2HSV4 U12568 ( .A1(n27877), .A2(n11807), .ZN(n15836) );
  CLKNHSV2 U12569 ( .I(n15835), .ZN(n11807) );
  CLKNAND2HSV8 U12570 ( .A1(n12724), .A2(n18463), .ZN(n28133) );
  CLKNAND2HSV4 U12571 ( .A1(n28133), .A2(n18464), .ZN(n18465) );
  CLKNAND2HSV8 U12572 ( .A1(n21003), .A2(\pe5/ti_7t [14]), .ZN(n21463) );
  NAND2HSV1 U12573 ( .A1(n27112), .A2(n13993), .ZN(n13155) );
  NAND2HSV2 U12574 ( .A1(n28473), .A2(n20977), .ZN(n24430) );
  NOR2HSV8 U12575 ( .A1(n23110), .A2(n23109), .ZN(n12663) );
  OAI21HSV4 U12576 ( .A1(n23425), .A2(n12663), .B(n23180), .ZN(n23187) );
  CLKNAND2HSV2 U12577 ( .A1(n11808), .A2(n15403), .ZN(n12570) );
  CLKNHSV2 U12578 ( .I(n11809), .ZN(n11808) );
  CLKNAND2HSV2 U12579 ( .A1(n15404), .A2(n12574), .ZN(n11809) );
  CLKNAND2HSV4 U12580 ( .A1(n17979), .A2(n17978), .ZN(n17980) );
  MUX2NHSV4 U12581 ( .I0(n17600), .I1(n13292), .S(n17599), .ZN(n17616) );
  OAI21HSV4 U12582 ( .A1(n17616), .A2(n28422), .B(n17601), .ZN(n17611) );
  CLKNAND2HSV2 U12583 ( .A1(n13820), .A2(n13821), .ZN(n13822) );
  XNOR2HSV4 U12584 ( .A1(n11810), .A2(n24338), .ZN(n13820) );
  CLKNHSV2 U12585 ( .I(n24339), .ZN(n11810) );
  NAND2HSV2 U12586 ( .A1(n11811), .A2(n16950), .ZN(n16951) );
  NOR2HSV2 U12587 ( .A1(n16946), .A2(n16947), .ZN(n11811) );
  NAND2HSV4 U12588 ( .A1(n21419), .A2(n21420), .ZN(n12215) );
  XNOR2HSV4 U12589 ( .A1(n27111), .A2(n11812), .ZN(\pe5/poht [14]) );
  XNOR2HSV4 U12590 ( .A1(n27110), .A2(n27109), .ZN(n11812) );
  XNOR2HSV4 U12591 ( .A1(n21689), .A2(n21688), .ZN(n21691) );
  NOR2HSV4 U12592 ( .A1(n11813), .A2(n21906), .ZN(n21907) );
  XNOR2HSV4 U12593 ( .A1(n23433), .A2(n11814), .ZN(n11813) );
  CLKNHSV2 U12594 ( .I(n21904), .ZN(n11814) );
  NAND3HSV4 U12595 ( .A1(n18450), .A2(n18451), .A3(n18452), .ZN(n18453) );
  INHSV4 U12596 ( .I(n18453), .ZN(n13481) );
  CLKNAND2HSV4 U12597 ( .A1(n28948), .A2(n28789), .ZN(n23190) );
  NAND2HSV4 U12598 ( .A1(n23118), .A2(n23119), .ZN(n28948) );
  CLKNAND2HSV4 U12599 ( .A1(n20399), .A2(n20398), .ZN(n20445) );
  CLKNHSV0 U12600 ( .I(n13784), .ZN(n13785) );
  AO32HSV4 U12601 ( .A1(n13785), .A2(n28664), .A3(n14852), .B1(n13784), .B2(
        n14671), .Z(n14672) );
  CLKNHSV12 U12602 ( .I(n27190), .ZN(n14045) );
  INAND2HSV4 U12603 ( .A1(n22125), .B1(\pe8/ti_7t [10]), .ZN(n21317) );
  CLKNAND2HSV3 U12604 ( .A1(n12380), .A2(n16991), .ZN(n20068) );
  INHSV2 U12605 ( .I(n20547), .ZN(n20453) );
  NAND2HSV4 U12606 ( .A1(n11815), .A2(n20360), .ZN(n20361) );
  CLKNAND2HSV4 U12607 ( .A1(n20359), .A2(n20358), .ZN(n11815) );
  NAND2HSV4 U12608 ( .A1(n24284), .A2(\pe7/got [2]), .ZN(n24283) );
  CLKNAND2HSV2 U12609 ( .A1(n18762), .A2(n12481), .ZN(n18763) );
  CLKNAND2HSV4 U12610 ( .A1(n18918), .A2(n18853), .ZN(n12488) );
  CLKNAND2HSV4 U12611 ( .A1(n12488), .A2(n18854), .ZN(n11816) );
  CLKNHSV4 U12612 ( .I(n16632), .ZN(n16635) );
  CLKNAND2HSV0 U12613 ( .A1(n27112), .A2(n24636), .ZN(n13061) );
  CLKNHSV6 U12614 ( .I(n15532), .ZN(n15704) );
  CLKNAND2HSV2 U12615 ( .A1(n28787), .A2(n14061), .ZN(n26079) );
  XOR2HSV4 U12616 ( .A1(n17108), .A2(n11838), .Z(n17109) );
  NAND2HSV4 U12617 ( .A1(n20125), .A2(n12379), .ZN(n12380) );
  NAND2HSV4 U12618 ( .A1(n12336), .A2(n12339), .ZN(n15567) );
  CLKNAND2HSV4 U12619 ( .A1(n11816), .A2(n18919), .ZN(n19132) );
  CLKXOR2HSV2 U12620 ( .A1(n22984), .A2(n22983), .Z(n22985) );
  INHSV2 U12621 ( .I(n11817), .ZN(n22914) );
  CLKNAND2HSV2 U12622 ( .A1(n22904), .A2(n22905), .ZN(n11817) );
  CLKNAND2HSV4 U12623 ( .A1(n11818), .A2(n12160), .ZN(n16999) );
  NAND2HSV4 U12624 ( .A1(n12159), .A2(n12158), .ZN(n11818) );
  NAND2HSV2 U12625 ( .A1(n28969), .A2(n21347), .ZN(n21418) );
  NAND2HSV2 U12626 ( .A1(n21418), .A2(n21417), .ZN(n21419) );
  NAND2HSV4 U12627 ( .A1(n16349), .A2(n16348), .ZN(n16350) );
  CLKNAND2HSV2 U12628 ( .A1(\pe4/bq[15] ), .A2(\pe4/aot [16]), .ZN(n13367) );
  MUX2NHSV4 U12629 ( .I0(n13366), .I1(\pe4/phq [2]), .S(n13367), .ZN(n15365)
         );
  NAND2HSV4 U12630 ( .A1(n28436), .A2(n24635), .ZN(n24436) );
  CLKAND2HSV4 U12631 ( .A1(n19234), .A2(n19263), .Z(n19240) );
  CLKNAND2HSV2 U12632 ( .A1(n11819), .A2(\pe4/pvq [2]), .ZN(n15366) );
  CLKNHSV2 U12633 ( .I(n15502), .ZN(n11819) );
  XOR2HSV2 U12634 ( .A1(n11820), .A2(n15521), .Z(n15522) );
  AOI21HSV4 U12635 ( .A1(n15520), .A2(n15519), .B(n15518), .ZN(n11820) );
  CLKNAND2HSV2 U12636 ( .A1(n24284), .A2(\pe7/got [12]), .ZN(n23908) );
  NAND2HSV4 U12637 ( .A1(n20611), .A2(n20690), .ZN(n20691) );
  CLKNHSV6 U12638 ( .I(n24220), .ZN(n28659) );
  NAND2HSV2 U12639 ( .A1(n11821), .A2(n18076), .ZN(n18143) );
  CLKNHSV2 U12640 ( .I(n18027), .ZN(n11821) );
  CLKNAND2HSV2 U12641 ( .A1(n18077), .A2(n17955), .ZN(n18027) );
  CLKNAND2HSV2 U12642 ( .A1(n13293), .A2(n15408), .ZN(n15405) );
  CLKNHSV0 U12643 ( .I(n15405), .ZN(n15483) );
  NOR2HSV4 U12644 ( .A1(n25340), .A2(n25339), .ZN(n25341) );
  CLKNAND2HSV4 U12645 ( .A1(n21875), .A2(n21876), .ZN(n21877) );
  CLKNAND2HSV4 U12646 ( .A1(n29020), .A2(n25420), .ZN(n19133) );
  NAND2HSV2 U12647 ( .A1(n19132), .A2(n19131), .ZN(n29020) );
  NAND3HSV3 U12648 ( .A1(n15822), .A2(n15636), .A3(n15823), .ZN(n15637) );
  CLKNAND2HSV2 U12649 ( .A1(n26213), .A2(n13039), .ZN(n13040) );
  OAI21HSV4 U12650 ( .A1(n13038), .A2(n13040), .B(n13041), .ZN(n13042) );
  XNOR2HSV4 U12651 ( .A1(n11823), .A2(n11822), .ZN(n19257) );
  AOI21HSV4 U12652 ( .A1(n19253), .A2(n25494), .B(n19252), .ZN(n11822) );
  XNOR2HSV4 U12653 ( .A1(n19254), .A2(n11960), .ZN(n11823) );
  MUX2NHSV2 U12654 ( .I0(n15713), .I1(n15708), .S(n15714), .ZN(n15709) );
  CLKNAND2HSV2 U12655 ( .A1(n15853), .A2(n28428), .ZN(n15714) );
  NAND2HSV2 U12656 ( .A1(n27344), .A2(n27231), .ZN(n21690) );
  CLKNAND2HSV4 U12657 ( .A1(n19064), .A2(n19065), .ZN(n12141) );
  NAND2HSV2 U12658 ( .A1(n16447), .A2(n25649), .ZN(n16448) );
  NAND2HSV2 U12659 ( .A1(n17989), .A2(n18326), .ZN(n17990) );
  INAND2HSV2 U12660 ( .A1(n19794), .B1(n18199), .ZN(n18206) );
  CLKNAND2HSV2 U12661 ( .A1(n19226), .A2(n19475), .ZN(n19183) );
  INHSV2 U12662 ( .I(n23373), .ZN(n14053) );
  NAND2HSV2 U12663 ( .A1(n28699), .A2(\pe6/got [2]), .ZN(n23710) );
  CLKNAND2HSV8 U12664 ( .A1(n17417), .A2(n17214), .ZN(n22075) );
  XNOR2HSV4 U12665 ( .A1(n21863), .A2(n21862), .ZN(n21864) );
  CLKNAND2HSV2 U12666 ( .A1(n13718), .A2(n11824), .ZN(n13719) );
  CLKNAND2HSV2 U12667 ( .A1(n11826), .A2(n11825), .ZN(n11824) );
  CLKNHSV2 U12668 ( .I(n13716), .ZN(n11825) );
  CLKNHSV2 U12669 ( .I(n13717), .ZN(n11826) );
  INHSV2 U12670 ( .I(n28988), .ZN(n20144) );
  INHSV4 U12671 ( .I(n19900), .ZN(n25597) );
  CLKNHSV1 U12672 ( .I(n22594), .ZN(n22592) );
  OAI21HSV1 U12673 ( .A1(n13060), .A2(n13061), .B(n13062), .ZN(\pe5/poht [4])
         );
  NAND2HSV2 U12674 ( .A1(n11884), .A2(n11950), .ZN(\pe10/poht [10]) );
  OAI21HSV1 U12675 ( .A1(n13154), .A2(n13155), .B(n13156), .ZN(\pe5/poht [12])
         );
  NAND2HSV4 U12676 ( .A1(n11828), .A2(n11827), .ZN(n16786) );
  INHSV2 U12677 ( .I(n16785), .ZN(n11827) );
  INHSV4 U12678 ( .I(n16784), .ZN(n11828) );
  XOR2HSV2 U12679 ( .A1(n12452), .A2(n11829), .Z(n13750) );
  AOI31HSV2 U12680 ( .A1(n13748), .A2(n12129), .A3(\pe11/got [1]), .B(n13749), 
        .ZN(n11829) );
  INHSV4 U12681 ( .I(n12369), .ZN(n16673) );
  CLKNAND2HSV4 U12682 ( .A1(n16781), .A2(n22508), .ZN(n12369) );
  NAND2HSV4 U12683 ( .A1(n16761), .A2(\pe10/got [12]), .ZN(n16681) );
  CLKNHSV6 U12684 ( .I(n28692), .ZN(n25525) );
  CLKNHSV6 U12685 ( .I(n28692), .ZN(n26231) );
  CLKXOR2HSV4 U12686 ( .A1(n27448), .A2(n27447), .Z(n27451) );
  CLKNAND2HSV4 U12687 ( .A1(n19949), .A2(n18783), .ZN(n21316) );
  CLKNAND2HSV8 U12688 ( .A1(n21316), .A2(n21317), .ZN(n19992) );
  NAND2HSV2 U12689 ( .A1(n24322), .A2(n20977), .ZN(n13681) );
  CLKNAND2HSV2 U12690 ( .A1(n24277), .A2(n25271), .ZN(n23218) );
  XNOR2HSV2 U12691 ( .A1(n23218), .A2(n23217), .ZN(\pe7/poht [9]) );
  NAND2HSV2 U12692 ( .A1(n28603), .A2(\pe10/got [5]), .ZN(n12397) );
  NAND2HSV2 U12693 ( .A1(n15376), .A2(n15375), .ZN(n12572) );
  NAND3HSV4 U12694 ( .A1(n20440), .A2(n20438), .A3(n20373), .ZN(n20393) );
  IOA21HSV4 U12695 ( .A1(n25597), .A2(n19835), .B(n18839), .ZN(n19990) );
  NAND2HSV2 U12696 ( .A1(\pe8/bq[12] ), .A2(\pe8/aot [15]), .ZN(n16372) );
  INHSV4 U12697 ( .I(n20998), .ZN(n21000) );
  NAND3HSV4 U12698 ( .A1(n12910), .A2(n19679), .A3(n19678), .ZN(n19617) );
  CLKNHSV6 U12699 ( .I(n28813), .ZN(n16464) );
  XNOR2HSV4 U12700 ( .A1(n24428), .A2(n24427), .ZN(n24429) );
  CLKXOR2HSV2 U12701 ( .A1(n24430), .A2(n24429), .Z(n24431) );
  CLKXOR2HSV4 U12702 ( .A1(n20269), .A2(n20268), .Z(n20270) );
  NAND2HSV4 U12703 ( .A1(n12075), .A2(n18262), .ZN(n18266) );
  XNOR2HSV4 U12704 ( .A1(n13823), .A2(n13824), .ZN(n13825) );
  NOR2HSV2 U12705 ( .A1(n11831), .A2(n11830), .ZN(n12594) );
  CLKNAND2HSV2 U12706 ( .A1(n28950), .A2(n21697), .ZN(n11830) );
  CLKNHSV2 U12707 ( .I(n25357), .ZN(n11831) );
  CLKXOR2HSV4 U12708 ( .A1(n17179), .A2(n17178), .Z(n17193) );
  XNOR2HSV2 U12709 ( .A1(n17193), .A2(n17192), .ZN(n17194) );
  MUX2NHSV2 U12710 ( .I0(n27209), .I1(n27208), .S(n11832), .ZN(n13796) );
  NOR2HSV4 U12711 ( .A1(n11834), .A2(n11833), .ZN(n11832) );
  CLKNHSV2 U12712 ( .I(\pe10/got [3]), .ZN(n11833) );
  CLKNHSV2 U12713 ( .I(n28603), .ZN(n11834) );
  XNOR2HSV4 U12714 ( .A1(n24699), .A2(n11835), .ZN(\pe5/poht [1]) );
  XNOR2HSV4 U12715 ( .A1(n24698), .A2(n24697), .ZN(n11835) );
  INHSV4 U12716 ( .I(n13290), .ZN(n16883) );
  NAND2HSV4 U12717 ( .A1(n19575), .A2(n27131), .ZN(n12077) );
  NAND2HSV4 U12718 ( .A1(n12489), .A2(n11836), .ZN(n19131) );
  INHSV4 U12719 ( .I(n18919), .ZN(n11836) );
  NAND2HSV4 U12720 ( .A1(n24075), .A2(n23107), .ZN(n23425) );
  CLKNAND2HSV2 U12721 ( .A1(n28801), .A2(n23414), .ZN(n23669) );
  XOR2HSV4 U12722 ( .A1(n23661), .A2(n23660), .Z(n23662) );
  XNOR2HSV2 U12723 ( .A1(n19895), .A2(n19894), .ZN(n19979) );
  XNOR2HSV4 U12724 ( .A1(n27489), .A2(n27488), .ZN(n27491) );
  XNOR2HSV4 U12725 ( .A1(n18309), .A2(n11837), .ZN(n13076) );
  XNOR2HSV4 U12726 ( .A1(n18306), .A2(n18307), .ZN(n11837) );
  INHSV2 U12727 ( .I(n15974), .ZN(n12820) );
  CLKNAND2HSV2 U12728 ( .A1(n20055), .A2(n21004), .ZN(n25606) );
  NAND2HSV4 U12729 ( .A1(n25607), .A2(n25606), .ZN(n12217) );
  NAND2HSV2 U12730 ( .A1(n21244), .A2(n21245), .ZN(n21295) );
  NOR2HSV4 U12731 ( .A1(n19569), .A2(n25628), .ZN(n19571) );
  CLKNHSV0 U12732 ( .I(n19571), .ZN(n27131) );
  CLKNAND2HSV4 U12733 ( .A1(n28949), .A2(n28137), .ZN(n18179) );
  NAND2HSV4 U12734 ( .A1(n14132), .A2(n14131), .ZN(n14134) );
  INHSV4 U12735 ( .I(n14134), .ZN(n14135) );
  NOR2HSV4 U12736 ( .A1(n19831), .A2(n13987), .ZN(n19834) );
  NOR2HSV8 U12737 ( .A1(n17302), .A2(n17374), .ZN(n14975) );
  NAND2HSV2 U12738 ( .A1(n18206), .A2(n18543), .ZN(n18208) );
  INHSV4 U12739 ( .I(n27271), .ZN(n27527) );
  CLKAND2HSV2 U12740 ( .A1(n27271), .A2(\pe2/got [9]), .Z(n21684) );
  CLKNAND2HSV2 U12741 ( .A1(n12370), .A2(n17066), .ZN(n11838) );
  CLKXOR2HSV2 U12742 ( .A1(n23600), .A2(n23599), .Z(n23601) );
  XNOR2HSV4 U12743 ( .A1(n20388), .A2(n20387), .ZN(n20390) );
  CLKNHSV4 U12744 ( .I(n16648), .ZN(n16734) );
  INHSV6 U12745 ( .I(n22230), .ZN(n25577) );
  BUFHSV12 U12746 ( .I(\pe8/got [1]), .Z(n26230) );
  INHSV2 U12747 ( .I(n16700), .ZN(n16698) );
  NAND2HSV2 U12748 ( .A1(n21162), .A2(n21161), .ZN(n12047) );
  INHSV2 U12749 ( .I(n23555), .ZN(n25374) );
  NAND2HSV2 U12750 ( .A1(n26231), .A2(\pe8/got [3]), .ZN(n23786) );
  NOR2HSV2 U12751 ( .A1(n19978), .A2(n11839), .ZN(n19984) );
  INHSV2 U12752 ( .I(n11840), .ZN(n11839) );
  NAND2HSV2 U12753 ( .A1(n19975), .A2(n19979), .ZN(n11840) );
  NAND2HSV4 U12754 ( .A1(n25597), .A2(n19835), .ZN(n18840) );
  INHSV2 U12755 ( .I(n18840), .ZN(n18844) );
  XNOR2HSV4 U12756 ( .A1(n12030), .A2(n16934), .ZN(n25677) );
  NAND2HSV2 U12757 ( .A1(n12031), .A2(n25677), .ZN(n16936) );
  NAND2HSV2 U12758 ( .A1(\pe5/ti_7[10] ), .A2(n14072), .ZN(n24369) );
  XNOR2HSV2 U12759 ( .A1(n24369), .A2(n24368), .ZN(n24371) );
  XOR2HSV4 U12760 ( .A1(n26157), .A2(n16891), .Z(n16842) );
  CLKNAND2HSV4 U12761 ( .A1(n16888), .A2(n16845), .ZN(n26157) );
  INHSV4 U12762 ( .I(n23550), .ZN(n24284) );
  CLKXOR2HSV4 U12763 ( .A1(n24627), .A2(n24626), .Z(n24631) );
  CLKXOR2HSV2 U12764 ( .A1(n16718), .A2(n16717), .Z(n16726) );
  NAND2HSV4 U12765 ( .A1(n16761), .A2(\pe10/got [13]), .ZN(n16649) );
  XNOR2HSV4 U12766 ( .A1(n11841), .A2(n23904), .ZN(n23907) );
  XNOR2HSV4 U12767 ( .A1(n23905), .A2(n23906), .ZN(n11841) );
  NAND2HSV2 U12768 ( .A1(n12517), .A2(n14071), .ZN(n21458) );
  NAND2HSV4 U12769 ( .A1(n28959), .A2(n16755), .ZN(n16756) );
  INHSV4 U12770 ( .I(n16756), .ZN(n16789) );
  NAND3HSV4 U12771 ( .A1(n24074), .A2(n24075), .A3(n24073), .ZN(n28703) );
  NAND2HSV2 U12772 ( .A1(n28703), .A2(\pe7/got [7]), .ZN(n24035) );
  CLKNAND2HSV2 U12773 ( .A1(n29044), .A2(n11842), .ZN(n17800) );
  CLKNHSV2 U12774 ( .I(n17797), .ZN(n11842) );
  XNOR2HSV4 U12775 ( .A1(n17749), .A2(n17748), .ZN(n29044) );
  NAND2HSV2 U12776 ( .A1(n26634), .A2(n11891), .ZN(n23379) );
  XOR2HSV4 U12777 ( .A1(n23379), .A2(n23378), .Z(n23381) );
  XOR2HSV2 U12778 ( .A1(n20434), .A2(n20435), .Z(n20437) );
  CLKNAND2HSV0 U12779 ( .A1(n26221), .A2(n27196), .ZN(n25695) );
  CLKNHSV4 U12780 ( .I(n14266), .ZN(n12065) );
  NAND2HSV4 U12781 ( .A1(n19967), .A2(n22125), .ZN(n22118) );
  INHSV4 U12782 ( .I(n23277), .ZN(n21570) );
  CLKXOR2HSV4 U12783 ( .A1(n21460), .A2(n21459), .Z(n13680) );
  XNOR2HSV4 U12784 ( .A1(n24376), .A2(n11843), .ZN(n13221) );
  CLKXOR2HSV4 U12785 ( .A1(n24375), .A2(n11844), .Z(n11843) );
  INHSV2 U12786 ( .I(n24374), .ZN(n11844) );
  NAND3HSV4 U12787 ( .A1(n14338), .A2(n14337), .A3(n14339), .ZN(n14283) );
  INHSV2 U12788 ( .I(n20401), .ZN(n20364) );
  NAND2HSV4 U12789 ( .A1(n16168), .A2(n24516), .ZN(n23400) );
  XNOR2HSV4 U12790 ( .A1(n14085), .A2(n11845), .ZN(n14090) );
  XOR2HSV2 U12791 ( .A1(n14084), .A2(n14083), .Z(n11845) );
  CLKNAND2HSV2 U12792 ( .A1(n19794), .A2(n18464), .ZN(n18139) );
  NAND2HSV4 U12793 ( .A1(n19573), .A2(n19572), .ZN(n19574) );
  CLKNHSV2 U12794 ( .I(n11846), .ZN(n19985) );
  CLKNAND2HSV2 U12795 ( .A1(n19984), .A2(n19983), .ZN(n11846) );
  INHSV6 U12796 ( .I(n19809), .ZN(n18625) );
  CLKNAND2HSV4 U12797 ( .A1(n28657), .A2(n11896), .ZN(n27213) );
  BUFHSV6 U12798 ( .I(n28706), .Z(n25204) );
  AND2HSV4 U12799 ( .A1(n19516), .A2(n25664), .Z(n19521) );
  XNOR2HSV4 U12800 ( .A1(n27968), .A2(n27967), .ZN(n27972) );
  OR2HSV8 U12801 ( .A1(n25374), .A2(n24128), .Z(n12269) );
  CLKXOR2HSV4 U12802 ( .A1(n17105), .A2(n17104), .Z(n17107) );
  NAND2HSV4 U12803 ( .A1(n12450), .A2(n12451), .ZN(n12447) );
  INAND2HSV4 U12804 ( .A1(n12211), .B1(n12447), .ZN(n12210) );
  OAI21HSV4 U12805 ( .A1(n14628), .A2(\pe5/ti_7t [12]), .B(n14045), .ZN(n20866) );
  CLKNAND2HSV3 U12806 ( .A1(n16794), .A2(n16793), .ZN(n16800) );
  CLKNAND2HSV4 U12807 ( .A1(n16748), .A2(n16747), .ZN(n16752) );
  NOR2HSV8 U12808 ( .A1(n16805), .A2(n25261), .ZN(n16806) );
  NAND2HSV4 U12809 ( .A1(n17063), .A2(n20070), .ZN(n17062) );
  XNOR2HSV4 U12810 ( .A1(n22559), .A2(n22558), .ZN(n22562) );
  XNOR2HSV4 U12811 ( .A1(n24304), .A2(n24303), .ZN(\pe7/poht [11]) );
  CLKNHSV6 U12812 ( .I(n22198), .ZN(n26229) );
  INHSV4 U12813 ( .I(n16837), .ZN(n16746) );
  NAND2HSV4 U12814 ( .A1(n16746), .A2(n16745), .ZN(n16748) );
  NAND2HSV4 U12815 ( .A1(n11938), .A2(n11847), .ZN(n11937) );
  AOI21HSV4 U12816 ( .A1(n17818), .A2(n17736), .B(n21701), .ZN(n11847) );
  OAI21HSV4 U12817 ( .A1(n18767), .A2(n29004), .B(n13799), .ZN(n13808) );
  XNOR2HSV2 U12818 ( .A1(n22276), .A2(n22275), .ZN(n22279) );
  INHSV2 U12819 ( .I(n22279), .ZN(n22277) );
  NAND2HSV4 U12820 ( .A1(n28679), .A2(n16876), .ZN(n16833) );
  NAND2HSV4 U12821 ( .A1(n12440), .A2(n12438), .ZN(n14110) );
  INHSV4 U12822 ( .I(n14110), .ZN(n11959) );
  NOR2HSV8 U12823 ( .A1(n24286), .A2(n19242), .ZN(n24273) );
  XOR3HSV4 U12824 ( .A1(n24274), .A2(n24273), .A3(n24272), .Z(n24275) );
  NAND2HSV2 U12825 ( .A1(\pe6/bq[16] ), .A2(\pe6/aot [12]), .ZN(n14215) );
  INHSV2 U12826 ( .I(n14215), .ZN(n12155) );
  AND2HSV2 U12827 ( .A1(n23555), .A2(\pe7/got [8]), .Z(n24077) );
  CLKXOR2HSV2 U12828 ( .A1(n23659), .A2(n23658), .Z(n23660) );
  XOR2HSV2 U12829 ( .A1(n21582), .A2(n21583), .Z(n13154) );
  NOR2HSV4 U12830 ( .A1(n29031), .A2(n15700), .ZN(n15846) );
  XNOR2HSV4 U12831 ( .A1(n11848), .A2(n15688), .ZN(n29031) );
  CLKNHSV2 U12832 ( .I(n15628), .ZN(n11848) );
  NAND2HSV4 U12833 ( .A1(n24893), .A2(\pe11/got [2]), .ZN(n12615) );
  CLKNAND2HSV4 U12834 ( .A1(n25634), .A2(n17917), .ZN(n18022) );
  CLKNAND2HSV4 U12835 ( .A1(n21815), .A2(n27231), .ZN(n21873) );
  INHSV4 U12836 ( .I(n21873), .ZN(n21876) );
  CLKNAND2HSV4 U12837 ( .A1(n22248), .A2(n22247), .ZN(n28698) );
  OAI22HSV2 U12838 ( .A1(n19235), .A2(n19262), .B1(n25309), .B2(n19189), .ZN(
        n19190) );
  CLKNAND2HSV2 U12839 ( .A1(\pe10/aot [15]), .A2(\pe10/bq[13] ), .ZN(n16687)
         );
  NAND2HSV4 U12840 ( .A1(n16897), .A2(\pe10/aot [13]), .ZN(n16682) );
  XOR2HSV4 U12841 ( .A1(n16682), .A2(n16681), .Z(n16686) );
  NAND2HSV4 U12842 ( .A1(n21452), .A2(n24635), .ZN(n12548) );
  INHSV4 U12843 ( .I(n12548), .ZN(n20994) );
  CLKXOR2HSV4 U12844 ( .A1(n19412), .A2(n19411), .Z(n19413) );
  CLKBUFHSV4 U12845 ( .I(n14506), .Z(n21342) );
  CLKNHSV1 U12846 ( .I(n16458), .ZN(n16456) );
  NAND2HSV2 U12847 ( .A1(n27112), .A2(n28647), .ZN(n13758) );
  INHSV4 U12848 ( .I(n16798), .ZN(n16712) );
  NAND2HSV4 U12849 ( .A1(n12620), .A2(n12619), .ZN(n16798) );
  INHSV4 U12850 ( .I(n14048), .ZN(n12437) );
  INHSV2 U12851 ( .I(n14047), .ZN(n21764) );
  XNOR2HSV4 U12852 ( .A1(n24696), .A2(n24695), .ZN(n24697) );
  BUFHSV4 U12853 ( .I(n22375), .Z(n18399) );
  CLKNHSV6 U12854 ( .I(n18104), .ZN(n18002) );
  NAND2HSV4 U12855 ( .A1(n12404), .A2(n22136), .ZN(n16579) );
  CLKNAND2HSV4 U12856 ( .A1(n21571), .A2(n21570), .ZN(n24322) );
  CLKNAND2HSV2 U12857 ( .A1(n24322), .A2(n14503), .ZN(n23954) );
  CLKAND2HSV4 U12858 ( .A1(n21738), .A2(n22418), .Z(n16996) );
  CLKNAND2HSV2 U12859 ( .A1(n24377), .A2(n24340), .ZN(n21553) );
  NAND2HSV4 U12860 ( .A1(n19140), .A2(n11849), .ZN(n12226) );
  NAND2HSV4 U12861 ( .A1(n12109), .A2(n19150), .ZN(n11849) );
  INHSV2 U12862 ( .I(n14787), .ZN(n14790) );
  CLKNAND2HSV2 U12863 ( .A1(n14790), .A2(n14789), .ZN(n14791) );
  NAND2HSV4 U12864 ( .A1(n18266), .A2(n18265), .ZN(n18269) );
  CLKNAND2HSV4 U12865 ( .A1(n27439), .A2(n27544), .ZN(n21871) );
  NAND2HSV2 U12866 ( .A1(n28134), .A2(n28689), .ZN(n13077) );
  AOI21HSV4 U12867 ( .A1(n17614), .A2(n13962), .B(n11850), .ZN(n25874) );
  CLKNAND2HSV2 U12868 ( .A1(n17612), .A2(n17613), .ZN(n11850) );
  CLKNAND2HSV2 U12869 ( .A1(n28807), .A2(n20707), .ZN(n20351) );
  DELHS1 U12870 ( .I(n20171), .Z(n11851) );
  CLKXOR2HSV4 U12871 ( .A1(n23675), .A2(n23674), .Z(n12925) );
  CLKBUFHSV12 U12872 ( .I(n20601), .Z(n11852) );
  CLKNAND2HSV3 U12873 ( .A1(n20929), .A2(n20928), .ZN(n11908) );
  CLKNHSV6 U12874 ( .I(n21909), .ZN(n24893) );
  OR2HSV4 U12875 ( .A1(n18920), .A2(n18993), .Z(n18921) );
  INHSV6 U12876 ( .I(n22880), .ZN(n25134) );
  CLKXOR2HSV2 U12877 ( .A1(n25947), .A2(n25946), .Z(n25948) );
  CLKNAND2HSV2 U12878 ( .A1(n22431), .A2(n20135), .ZN(n20139) );
  CLKNAND2HSV2 U12879 ( .A1(n20132), .A2(n20142), .ZN(n22431) );
  CLKNHSV6 U12880 ( .I(n11853), .ZN(n21879) );
  INHSV6 U12881 ( .I(n28950), .ZN(n11853) );
  INHSV4 U12882 ( .I(n11854), .ZN(n19670) );
  INHSV2 U12883 ( .I(n19610), .ZN(n11854) );
  INHSV2 U12884 ( .I(n12569), .ZN(n21151) );
  BUFHSV2 U12885 ( .I(n14077), .Z(n11855) );
  NOR2HSV8 U12886 ( .A1(n28674), .A2(n26156), .ZN(n17060) );
  XOR2HSV0 U12887 ( .A1(n23322), .A2(n23321), .Z(\pe11/poht [11]) );
  AND2HSV8 U12888 ( .A1(n15455), .A2(n15452), .Z(n13972) );
  NAND2HSV4 U12889 ( .A1(n13972), .A2(n15640), .ZN(n15499) );
  XNOR2HSV4 U12890 ( .A1(n16278), .A2(n16277), .ZN(n16279) );
  NAND2HSV2 U12891 ( .A1(n24965), .A2(\pe11/got [4]), .ZN(n24874) );
  NOR2HSV4 U12892 ( .A1(n16788), .A2(n12345), .ZN(n16836) );
  NAND2HSV2 U12893 ( .A1(n13199), .A2(n12573), .ZN(n15493) );
  NAND2HSV2 U12894 ( .A1(n15493), .A2(n15484), .ZN(n15485) );
  NAND2HSV2 U12895 ( .A1(n16287), .A2(n16286), .ZN(n17171) );
  NAND2HSV4 U12896 ( .A1(n28430), .A2(\pe7/got [12]), .ZN(n19750) );
  XOR2HSV0 U12897 ( .A1(n25747), .A2(n25748), .Z(\pe6/poht [3]) );
  NAND2HSV2 U12898 ( .A1(\pe11/aot [14]), .A2(\pe11/bq[14] ), .ZN(n20273) );
  INHSV6 U12899 ( .I(\pe11/ti_1 ), .ZN(n20151) );
  CLKNHSV6 U12900 ( .I(n20151), .ZN(n20272) );
  CLKNAND2HSV4 U12901 ( .A1(n11856), .A2(n17806), .ZN(n17805) );
  NAND2HSV2 U12902 ( .A1(n17804), .A2(n28421), .ZN(n11856) );
  NOR2HSV2 U12903 ( .A1(n12570), .A2(n12571), .ZN(n15492) );
  INHSV4 U12904 ( .I(\pe11/pvq [2]), .ZN(n20166) );
  NAND2HSV2 U12905 ( .A1(n22597), .A2(n22596), .ZN(\pe10/poht [8]) );
  CLKNAND2HSV2 U12906 ( .A1(n14646), .A2(\pe5/pvq [7]), .ZN(n14585) );
  NAND2HSV2 U12907 ( .A1(n22635), .A2(n22634), .ZN(\pe10/poht [7]) );
  CLKNAND2HSV2 U12908 ( .A1(n21322), .A2(n22136), .ZN(n19938) );
  CLKNAND2HSV4 U12909 ( .A1(n14619), .A2(n14635), .ZN(n14623) );
  NAND2HSV4 U12910 ( .A1(n14623), .A2(n14622), .ZN(n28990) );
  XOR2HSV4 U12911 ( .A1(n12015), .A2(n25341), .Z(n12014) );
  NAND2HSV2 U12912 ( .A1(n17639), .A2(n11857), .ZN(n17650) );
  NAND4HSV2 U12913 ( .A1(\pe2/pvq [1]), .A2(\pe2/aot [16]), .A3(\pe2/bq[16] ), 
        .A4(\pe2/ctrq ), .ZN(n11857) );
  CLKNAND2HSV2 U12914 ( .A1(n23482), .A2(n25131), .ZN(n15467) );
  CLKNAND2HSV4 U12915 ( .A1(n21817), .A2(n27231), .ZN(n17854) );
  CLKNAND2HSV2 U12916 ( .A1(n17084), .A2(\pe10/aot [13]), .ZN(n16650) );
  NAND2HSV4 U12917 ( .A1(n20774), .A2(n20773), .ZN(n20779) );
  INHSV4 U12918 ( .I(n12110), .ZN(n12109) );
  NOR2HSV2 U12919 ( .A1(n18549), .A2(n18545), .ZN(n18546) );
  INHSV4 U12920 ( .I(\pe7/bq[16] ), .ZN(n19246) );
  NOR2HSV2 U12921 ( .A1(n19247), .A2(n19246), .ZN(n19249) );
  DELHS1 U12922 ( .I(\pe7/ti_7[1] ), .Z(n11858) );
  CLKNAND2HSV2 U12923 ( .A1(n16837), .A2(n17112), .ZN(n12021) );
  XNOR2HSV4 U12924 ( .A1(n11859), .A2(n19175), .ZN(\pe6/poht [10]) );
  XOR2HSV2 U12925 ( .A1(n19173), .A2(n19174), .Z(n11859) );
  CLKNAND2HSV2 U12926 ( .A1(n26030), .A2(\pe6/got [6]), .ZN(n25975) );
  XNOR2HSV1 U12927 ( .A1(n25974), .A2(n25975), .ZN(n25976) );
  NOR2HSV4 U12928 ( .A1(n11861), .A2(n11860), .ZN(n14529) );
  CLKNAND2HSV2 U12929 ( .A1(n22097), .A2(n14526), .ZN(n11860) );
  CLKNHSV2 U12930 ( .I(n22094), .ZN(n11861) );
  INHSV4 U12931 ( .I(n18275), .ZN(n18204) );
  XOR2HSV2 U12932 ( .A1(n19608), .A2(n19607), .Z(n12122) );
  NAND2HSV2 U12933 ( .A1(n25980), .A2(n25420), .ZN(n23057) );
  CLKNAND2HSV2 U12934 ( .A1(\pe7/bq[15] ), .A2(\pe7/aot [16]), .ZN(n19192) );
  NAND2HSV2 U12935 ( .A1(n24377), .A2(n20977), .ZN(n21627) );
  CLKNAND2HSV4 U12936 ( .A1(n18275), .A2(n12361), .ZN(n18334) );
  XOR2HSV0 U12937 ( .A1(n23056), .A2(n23057), .Z(\pe6/poht [1]) );
  CLKNAND2HSV4 U12938 ( .A1(n25950), .A2(n26083), .ZN(n26088) );
  CLKXOR2HSV2 U12939 ( .A1(n26088), .A2(n26087), .Z(n26089) );
  BUFHSV6 U12940 ( .I(n12434), .Z(n12433) );
  CLKNAND2HSV2 U12941 ( .A1(n20984), .A2(n14045), .ZN(n20986) );
  NAND2HSV2 U12942 ( .A1(n28703), .A2(n24214), .ZN(n24215) );
  CLKNAND2HSV4 U12943 ( .A1(n18541), .A2(n18611), .ZN(n12724) );
  INHSV2 U12944 ( .I(n21102), .ZN(n17855) );
  XNOR2HSV4 U12945 ( .A1(n14541), .A2(n11862), .ZN(n14543) );
  XOR2HSV2 U12946 ( .A1(n14540), .A2(n14539), .Z(n11862) );
  CLKNAND2HSV2 U12947 ( .A1(n24377), .A2(\pe5/got [3]), .ZN(n21583) );
  CLKNAND2HSV4 U12948 ( .A1(n21571), .A2(n23275), .ZN(n28436) );
  CLKNAND2HSV2 U12949 ( .A1(n21222), .A2(n21223), .ZN(n21170) );
  NAND2HSV4 U12950 ( .A1(n17923), .A2(n17922), .ZN(n17924) );
  NOR2HSV4 U12951 ( .A1(n27277), .A2(n21645), .ZN(n21689) );
  CLKNAND2HSV2 U12952 ( .A1(n28707), .A2(n15242), .ZN(n15908) );
  NAND2HSV4 U12953 ( .A1(\pe10/aot [15]), .A2(\pe10/bq[12] ), .ZN(n16899) );
  XNOR2HSV4 U12954 ( .A1(n15107), .A2(n15106), .ZN(n15116) );
  DELHS1 U12955 ( .I(n28470), .Z(n11863) );
  CLKNAND2HSV4 U12956 ( .A1(n22692), .A2(n17121), .ZN(n17132) );
  OAI21HSV4 U12957 ( .A1(n12892), .A2(n23442), .B(n16178), .ZN(n23417) );
  CLKNAND2HSV4 U12958 ( .A1(n16111), .A2(n16110), .ZN(n26291) );
  CLKNAND2HSV2 U12959 ( .A1(n26291), .A2(n28930), .ZN(n16174) );
  INHSV2 U12960 ( .I(n22914), .ZN(n22900) );
  INHSV4 U12961 ( .I(n18270), .ZN(n18268) );
  CLKNAND2HSV4 U12962 ( .A1(n18268), .A2(n18267), .ZN(n18272) );
  CLKNAND2HSV2 U12963 ( .A1(n17893), .A2(n17892), .ZN(n17889) );
  CLKNAND2HSV4 U12964 ( .A1(n19522), .A2(n19523), .ZN(n25665) );
  NAND2HSV4 U12965 ( .A1(n19511), .A2(n19623), .ZN(n19522) );
  XOR2HSV2 U12966 ( .A1(n11865), .A2(n11864), .Z(n14313) );
  CLKNAND2HSV2 U12967 ( .A1(\pe6/aot [12]), .A2(\pe6/bq[14] ), .ZN(n11864) );
  CLKNAND2HSV2 U12968 ( .A1(\pe6/bq[10] ), .A2(\pe6/aot [16]), .ZN(n11865) );
  AND2HSV4 U12969 ( .A1(n21222), .A2(n21221), .Z(n21228) );
  NAND2HSV2 U12970 ( .A1(n15640), .A2(n13994), .ZN(n15537) );
  NOR2HSV2 U12971 ( .A1(n15426), .A2(n13078), .ZN(n15448) );
  INHSV2 U12972 ( .I(n19577), .ZN(n19576) );
  XNOR2HSV4 U12973 ( .A1(n17879), .A2(n11866), .ZN(n17880) );
  XNOR2HSV4 U12974 ( .A1(n17878), .A2(\pe9/phq [5]), .ZN(n11866) );
  INHSV2 U12975 ( .I(n11867), .ZN(n13969) );
  NAND2HSV0 U12976 ( .A1(n14181), .A2(n18847), .ZN(n11867) );
  INHSV6 U12977 ( .I(n22718), .ZN(n27195) );
  CLKNAND2HSV2 U12978 ( .A1(n28966), .A2(n19069), .ZN(n14340) );
  XNOR2HSV4 U12979 ( .A1(n11869), .A2(n11868), .ZN(n13287) );
  CLKNHSV2 U12980 ( .I(n13286), .ZN(n11868) );
  CLKNHSV2 U12981 ( .I(n13285), .ZN(n11869) );
  INHSV2 U12982 ( .I(\pe3/aot [16]), .ZN(n15108) );
  INHSV2 U12983 ( .I(n16553), .ZN(n12249) );
  XOR2HSV0 U12984 ( .A1(n25872), .A2(n25873), .Z(\pe6/poht [2]) );
  CLKNAND2HSV4 U12985 ( .A1(n21785), .A2(\pe11/ti_7t [14]), .ZN(n25053) );
  XOR2HSV0 U12986 ( .A1(n26028), .A2(n26029), .Z(\pe6/poht [5]) );
  NAND2HSV2 U12987 ( .A1(n29031), .A2(n22905), .ZN(n23059) );
  NAND2HSV0 U12988 ( .A1(n23059), .A2(n23058), .ZN(n21994) );
  NAND2HSV4 U12989 ( .A1(n15041), .A2(n11870), .ZN(n15043) );
  NAND3HSV2 U12990 ( .A1(n15040), .A2(\pe3/aot [16]), .A3(\pe3/bq[15] ), .ZN(
        n11870) );
  CLKNHSV0 U12991 ( .I(\pe5/ctrq ), .ZN(n14777) );
  NAND2HSV0 U12992 ( .A1(n26221), .A2(\pe10/got [2]), .ZN(n25066) );
  CLKNAND2HSV4 U12993 ( .A1(n11871), .A2(n25029), .ZN(n23438) );
  CLKNAND2HSV4 U12994 ( .A1(n23437), .A2(n23436), .ZN(n11871) );
  XOR2HSV2 U12995 ( .A1(n26079), .A2(n11872), .Z(n26080) );
  XOR2HSV2 U12996 ( .A1(n26077), .A2(n26078), .Z(n11872) );
  NAND2HSV4 U12997 ( .A1(n18706), .A2(n16554), .ZN(n18714) );
  NAND2HSV2 U12998 ( .A1(n16553), .A2(n16551), .ZN(n18706) );
  XOR2HSV4 U12999 ( .A1(n21965), .A2(n21964), .Z(\pe11/poht [2]) );
  XNOR2HSV4 U13000 ( .A1(n11873), .A2(n25487), .ZN(po6) );
  XOR2HSV2 U13001 ( .A1(n25486), .A2(n25485), .Z(n11873) );
  OR2HSV1 U13002 ( .A1(n20978), .A2(n20869), .Z(n20924) );
  NAND2HSV4 U13003 ( .A1(n12771), .A2(n12772), .ZN(n12774) );
  INHSV4 U13004 ( .I(n20849), .ZN(n20851) );
  NAND2HSV4 U13005 ( .A1(n20851), .A2(n20850), .ZN(n20919) );
  NAND2HSV2 U13006 ( .A1(\pe3/bq[16] ), .A2(\pe3/aot [14]), .ZN(n15018) );
  NAND2HSV4 U13007 ( .A1(n11874), .A2(n18843), .ZN(n19901) );
  CLKNAND2HSV4 U13008 ( .A1(n18842), .A2(n18841), .ZN(n11874) );
  NAND3HSV4 U13009 ( .A1(n19840), .A2(n19838), .A3(n19839), .ZN(n12241) );
  CLKNAND2HSV4 U13010 ( .A1(n20843), .A2(n11875), .ZN(n23320) );
  AOI22HSV2 U13011 ( .A1(n24884), .A2(n20770), .B1(n24881), .B2(n20769), .ZN(
        n11875) );
  NAND2HSV2 U13012 ( .A1(\pe8/bq[13] ), .A2(\pe8/aot [16]), .ZN(n16340) );
  XOR2HSV4 U13013 ( .A1(n16341), .A2(n16340), .Z(n12530) );
  CLKNAND2HSV4 U13014 ( .A1(n15478), .A2(n15484), .ZN(n15489) );
  INHSV4 U13015 ( .I(n15489), .ZN(n15565) );
  INHSV4 U13016 ( .I(n16809), .ZN(n12599) );
  NAND2HSV4 U13017 ( .A1(n12599), .A2(\pe10/aot [14]), .ZN(n16636) );
  OAI21HSV4 U13018 ( .A1(n12187), .A2(\pe5/phq [1]), .B(n11876), .ZN(n12192)
         );
  CLKNAND2HSV2 U13019 ( .A1(n12186), .A2(\pe5/phq [1]), .ZN(n11876) );
  CLKNAND2HSV2 U13020 ( .A1(n15126), .A2(n15189), .ZN(n15127) );
  CLKNHSV6 U13021 ( .I(n16976), .ZN(n14002) );
  NAND2HSV0 U13022 ( .A1(n16430), .A2(n16535), .ZN(n16421) );
  INAND2HSV4 U13023 ( .A1(n25668), .B1(n12678), .ZN(n12677) );
  INHSV4 U13024 ( .I(n18093), .ZN(n18094) );
  NAND2HSV4 U13025 ( .A1(n23320), .A2(n23319), .ZN(n25182) );
  CLKNAND2HSV4 U13026 ( .A1(n19179), .A2(n19180), .ZN(n19206) );
  XOR2HSV2 U13027 ( .A1(n11877), .A2(n17852), .Z(n17853) );
  XOR3HSV2 U13028 ( .A1(n17851), .A2(n17850), .A3(n17849), .Z(n11877) );
  NAND2HSV2 U13029 ( .A1(n23219), .A2(\pe10/got [3]), .ZN(n23228) );
  NAND2HSV2 U13030 ( .A1(n17991), .A2(n17992), .ZN(n17952) );
  NAND2HSV4 U13031 ( .A1(n26481), .A2(n26482), .ZN(n27000) );
  CLKNAND2HSV4 U13032 ( .A1(n17621), .A2(n11878), .ZN(n26482) );
  NAND2HSV4 U13033 ( .A1(n11880), .A2(n11879), .ZN(n11878) );
  INHSV2 U13034 ( .I(n17622), .ZN(n11879) );
  INHSV4 U13035 ( .I(n13962), .ZN(n11880) );
  CLKNAND2HSV4 U13036 ( .A1(n12698), .A2(n13338), .ZN(n29021) );
  NAND2HSV4 U13037 ( .A1(n29021), .A2(n19160), .ZN(n21743) );
  NAND2HSV4 U13038 ( .A1(n13200), .A2(n16420), .ZN(n13201) );
  CLKNAND2HSV2 U13039 ( .A1(n22063), .A2(n22062), .ZN(n22064) );
  XOR2HSV4 U13040 ( .A1(n21961), .A2(n21960), .Z(n21962) );
  XOR2HSV4 U13041 ( .A1(n24921), .A2(n24920), .Z(n24922) );
  CLKNAND2HSV2 U13042 ( .A1(n15895), .A2(n15894), .ZN(n15896) );
  CLKXOR2HSV4 U13043 ( .A1(n22557), .A2(n22556), .Z(n22559) );
  CLKNAND2HSV4 U13044 ( .A1(n26682), .A2(n26642), .ZN(n16098) );
  XOR3HSV2 U13045 ( .A1(n16099), .A2(n16098), .A3(n16097), .Z(n16100) );
  NAND2HSV2 U13046 ( .A1(n18021), .A2(n18022), .ZN(n28470) );
  AOI21HSV4 U13047 ( .A1(n17914), .A2(n17913), .B(n17912), .ZN(n18021) );
  NOR2HSV4 U13048 ( .A1(n18042), .A2(n22375), .ZN(n18090) );
  XNOR2HSV4 U13049 ( .A1(n24450), .A2(n11881), .ZN(n13757) );
  XOR2HSV2 U13050 ( .A1(n24449), .A2(n11882), .Z(n11881) );
  CLKNHSV2 U13051 ( .I(n24448), .ZN(n11882) );
  NAND2HSV2 U13052 ( .A1(n15281), .A2(n15280), .ZN(n15282) );
  XNOR2HSV4 U13053 ( .A1(n24847), .A2(n24846), .ZN(n24848) );
  CLKXOR2HSV4 U13054 ( .A1(n24849), .A2(n24848), .Z(n24852) );
  CLKXOR2HSV2 U13055 ( .A1(n16409), .A2(\pe8/phq [5]), .Z(n16410) );
  NAND2HSV2 U13056 ( .A1(\pe10/got [9]), .A2(n25060), .ZN(n22756) );
  NAND2HSV4 U13057 ( .A1(n23327), .A2(n28628), .ZN(n11887) );
  XNOR2HSV4 U13058 ( .A1(n15891), .A2(n11883), .ZN(n15893) );
  XNOR2HSV4 U13059 ( .A1(n15889), .A2(n15890), .ZN(n11883) );
  MUX2NHSV2 U13060 ( .I0(n17770), .I1(n14044), .S(n17818), .ZN(n11938) );
  CLKXOR2HSV4 U13061 ( .A1(n28256), .A2(n28255), .Z(n28258) );
  CLKXOR2HSV4 U13062 ( .A1(n28136), .A2(n28135), .Z(n28139) );
  CLKXOR2HSV4 U13063 ( .A1(n28181), .A2(n28180), .Z(n28183) );
  CLKNAND2HSV2 U13064 ( .A1(n28922), .A2(\pe11/got [9]), .ZN(n25179) );
  CLKXOR2HSV4 U13065 ( .A1(n26295), .A2(n26294), .Z(n13157) );
  NAND2HSV2 U13066 ( .A1(n13158), .A2(n13157), .ZN(n13159) );
  CLKNAND2HSV4 U13067 ( .A1(n28588), .A2(n26642), .ZN(n23369) );
  XNOR2HSV2 U13068 ( .A1(n23369), .A2(n23368), .ZN(n23370) );
  NAND2HSV2 U13069 ( .A1(n28110), .A2(n18078), .ZN(n17921) );
  CLKNAND2HSV4 U13070 ( .A1(n18673), .A2(\pe8/pvq [6]), .ZN(n16367) );
  INHSV4 U13071 ( .I(n25517), .ZN(n25521) );
  NAND2HSV4 U13072 ( .A1(n16511), .A2(\pe8/got [13]), .ZN(n11921) );
  CLKXOR2HSV4 U13073 ( .A1(n21690), .A2(n21691), .Z(n12595) );
  CLKNAND2HSV2 U13074 ( .A1(n22505), .A2(n22506), .ZN(n11884) );
  XNOR2HSV4 U13075 ( .A1(n25746), .A2(n11885), .ZN(n25747) );
  XOR2HSV2 U13076 ( .A1(n25744), .A2(n25745), .Z(n11885) );
  XNOR2HSV4 U13077 ( .A1(n12391), .A2(n12387), .ZN(n22714) );
  NAND2HSV4 U13078 ( .A1(n12129), .A2(\pe11/got [8]), .ZN(n12308) );
  AND2HSV2 U13079 ( .A1(n22624), .A2(\pe10/got [7]), .Z(n22625) );
  DELHS1 U13080 ( .I(n17554), .Z(n11886) );
  CLKNAND2HSV4 U13081 ( .A1(n28471), .A2(\pe11/got [9]), .ZN(n20749) );
  CLKXOR2HSV2 U13082 ( .A1(n20749), .A2(n20748), .Z(n20750) );
  CLKNAND2HSV8 U13083 ( .A1(n25370), .A2(n22919), .ZN(n22921) );
  NOR2HSV8 U13084 ( .A1(n22921), .A2(n22920), .ZN(n22923) );
  XNOR2HSV4 U13085 ( .A1(n15959), .A2(n11887), .ZN(n15970) );
  INHSV2 U13086 ( .I(n28432), .ZN(n26714) );
  NAND3HSV3 U13087 ( .A1(n19676), .A2(n19674), .A3(n19675), .ZN(n19706) );
  INHSV4 U13088 ( .I(n18167), .ZN(n27092) );
  XNOR2HSV4 U13089 ( .A1(n12633), .A2(n11888), .ZN(n14853) );
  XNOR2HSV4 U13090 ( .A1(n12627), .A2(n12631), .ZN(n11888) );
  XNOR2HSV4 U13091 ( .A1(n11889), .A2(n25783), .ZN(\pe6/poht [7]) );
  XNOR2HSV4 U13092 ( .A1(n25781), .A2(n25782), .ZN(n11889) );
  XNOR2HSV4 U13093 ( .A1(n11890), .A2(n12016), .ZN(n12015) );
  NOR2HSV4 U13094 ( .A1(n24045), .A2(n25338), .ZN(n11890) );
  NOR2HSV4 U13095 ( .A1(n12123), .A2(n14105), .ZN(n25476) );
  DELHS1 U13096 ( .I(\pe3/got [12]), .Z(n11891) );
  INHSV4 U13097 ( .I(n16346), .ZN(n16349) );
  INAND2HSV4 U13098 ( .A1(n20760), .B1(n20761), .ZN(n28919) );
  CLKNAND2HSV8 U13099 ( .A1(n18197), .A2(n12460), .ZN(n18210) );
  INHSV2 U13100 ( .I(n18210), .ZN(n25662) );
  INHSV4 U13101 ( .I(n15280), .ZN(n15278) );
  NAND2HSV4 U13102 ( .A1(n14497), .A2(n14965), .ZN(n13191) );
  CLKNAND2HSV4 U13103 ( .A1(n18310), .A2(n18398), .ZN(n12479) );
  CLKNAND2HSV1 U13104 ( .A1(n12377), .A2(n27228), .ZN(n15495) );
  XNOR2HSV4 U13105 ( .A1(n16299), .A2(\pe8/phq [3]), .ZN(n16300) );
  CLKNAND2HSV2 U13106 ( .A1(n15687), .A2(n15621), .ZN(n15689) );
  CLKNAND2HSV2 U13107 ( .A1(n18284), .A2(n18283), .ZN(n18322) );
  XNOR2HSV4 U13108 ( .A1(n23216), .A2(n23215), .ZN(n23217) );
  XNOR2HSV4 U13109 ( .A1(n11892), .A2(n24035), .ZN(n12275) );
  XNOR2HSV4 U13110 ( .A1(n24033), .A2(n11893), .ZN(n11892) );
  CLKNHSV2 U13111 ( .I(n24034), .ZN(n11893) );
  XNOR2HSV1 U13112 ( .A1(n11895), .A2(n11894), .ZN(n25872) );
  XOR2HSV0 U13113 ( .A1(n25870), .A2(n25871), .Z(n11894) );
  NAND2HSV0 U13114 ( .A1(n25950), .A2(\pe6/got [13]), .ZN(n11895) );
  CLKAND2HSV4 U13115 ( .A1(n21973), .A2(n22905), .Z(n13970) );
  NAND2HSV0 U13116 ( .A1(n21312), .A2(n23396), .ZN(n12892) );
  CLKNAND2HSV4 U13117 ( .A1(\pe8/pvq [2]), .A2(\pe8/ctrq ), .ZN(n16313) );
  MUX2NHSV4 U13118 ( .I0(\pe8/phq [2]), .I1(n16314), .S(n16313), .ZN(n16315)
         );
  CLKNAND2HSV4 U13119 ( .A1(n25500), .A2(n28610), .ZN(n23110) );
  CLKNAND2HSV2 U13120 ( .A1(n17292), .A2(n17291), .ZN(n17298) );
  CLKNAND2HSV2 U13121 ( .A1(n17299), .A2(n17298), .ZN(n17293) );
  MUX2NHSV4 U13122 ( .I0(n19529), .I1(n27213), .S(n19381), .ZN(n19383) );
  INHSV4 U13123 ( .I(n19684), .ZN(n11896) );
  NAND2HSV4 U13124 ( .A1(n12140), .A2(n21106), .ZN(n28942) );
  NAND2HSV4 U13125 ( .A1(n28942), .A2(n12013), .ZN(n12012) );
  NAND2HSV0 U13126 ( .A1(n13332), .A2(n13331), .ZN(n13333) );
  CLKNAND2HSV2 U13127 ( .A1(n13330), .A2(n11897), .ZN(n13331) );
  CLKNAND2HSV2 U13128 ( .A1(n11899), .A2(n11898), .ZN(n11897) );
  CLKNHSV2 U13129 ( .I(n13329), .ZN(n11898) );
  CLKNHSV2 U13130 ( .I(n13328), .ZN(n11899) );
  XNOR2HSV4 U13131 ( .A1(n21782), .A2(n21783), .ZN(\pe6/poht [11]) );
  CLKNAND2HSV2 U13132 ( .A1(n27485), .A2(n21692), .ZN(n21017) );
  CLKXOR2HSV4 U13133 ( .A1(n26347), .A2(n26346), .Z(n13063) );
  AOI22HSV4 U13134 ( .A1(\pe6/ti_7t [9]), .A2(n19138), .B1(n11900), .B2(n14696), .ZN(n18846) );
  NOR2HSV4 U13135 ( .A1(n25059), .A2(n14406), .ZN(n11900) );
  INHSV2 U13136 ( .I(n20254), .ZN(n11965) );
  INHSV2 U13137 ( .I(n16608), .ZN(n13597) );
  NAND2HSV4 U13138 ( .A1(n18690), .A2(n11901), .ZN(n16608) );
  INHSV2 U13139 ( .I(n12251), .ZN(n11901) );
  BUFHSV8 U13140 ( .I(\pe3/ctrq ), .Z(n23345) );
  INHSV4 U13141 ( .I(n11902), .ZN(n27284) );
  NAND2HSV4 U13142 ( .A1(n21632), .A2(n11903), .ZN(n11902) );
  INHSV4 U13143 ( .I(n25362), .ZN(n11903) );
  CLKNAND2HSV4 U13144 ( .A1(n21879), .A2(n21881), .ZN(n21632) );
  NOR2HSV4 U13145 ( .A1(n21167), .A2(n21217), .ZN(n21172) );
  NOR2HSV8 U13146 ( .A1(n21172), .A2(n21171), .ZN(n21640) );
  CLKNAND2HSV4 U13147 ( .A1(n19277), .A2(n19276), .ZN(n19322) );
  NAND2HSV4 U13148 ( .A1(n19322), .A2(n19321), .ZN(n19324) );
  OAI21HSV2 U13149 ( .A1(n12922), .A2(n12923), .B(n12924), .ZN(n22222) );
  XNOR2HSV2 U13150 ( .A1(n22223), .A2(n22222), .ZN(n22225) );
  INHSV24 U13151 ( .I(n20989), .ZN(n11904) );
  INHSV2 U13152 ( .I(pov5[10]), .ZN(n11905) );
  AOI21HSV4 U13153 ( .A1(n11905), .A2(n21422), .B(n11904), .ZN(n20990) );
  XNOR2HSV4 U13154 ( .A1(n11906), .A2(n16238), .ZN(n25653) );
  XNOR2HSV4 U13155 ( .A1(n16208), .A2(n16207), .ZN(n11906) );
  CLKXOR2HSV4 U13156 ( .A1(n21781), .A2(n21780), .Z(n21782) );
  CLKNAND2HSV4 U13157 ( .A1(n11908), .A2(n11907), .ZN(n28969) );
  CLKNAND2HSV2 U13158 ( .A1(n20927), .A2(n12309), .ZN(n11907) );
  OAI21HSV2 U13159 ( .A1(n28973), .A2(n21423), .B(n21414), .ZN(n21415) );
  OR2HSV8 U13160 ( .A1(n19684), .A2(n24220), .Z(n24276) );
  CLKXOR2HSV2 U13161 ( .A1(n24276), .A2(n24275), .Z(\pe7/poht [1]) );
  XNOR2HSV4 U13162 ( .A1(n12315), .A2(n19124), .ZN(n12314) );
  CLKNAND2HSV2 U13163 ( .A1(n29000), .A2(n18338), .ZN(n18340) );
  AOI21HSV2 U13164 ( .A1(n28662), .A2(\pe6/got [4]), .B(n25771), .ZN(n25772)
         );
  CLKXOR2HSV4 U13165 ( .A1(n24625), .A2(n24624), .Z(n24627) );
  INHSV2 U13166 ( .I(n14862), .ZN(n24634) );
  CLKNAND2HSV2 U13167 ( .A1(n18828), .A2(\pe8/got [12]), .ZN(n18753) );
  NAND2HSV4 U13168 ( .A1(n12395), .A2(n12394), .ZN(n16310) );
  CLKXOR2HSV4 U13169 ( .A1(n21022), .A2(n21021), .Z(n29041) );
  NAND2HSV4 U13170 ( .A1(n25660), .A2(n12478), .ZN(n18216) );
  CLKNAND2HSV2 U13171 ( .A1(n24322), .A2(n28645), .ZN(n12982) );
  XNOR2HSV4 U13172 ( .A1(n11910), .A2(n11909), .ZN(n16419) );
  CLKNHSV2 U13173 ( .I(n16417), .ZN(n11909) );
  XNOR2HSV4 U13174 ( .A1(n16413), .A2(n16412), .ZN(n11910) );
  CLKNAND2HSV2 U13175 ( .A1(\pe8/ctrq ), .A2(\pe8/pvq [1]), .ZN(n16292) );
  NOR2HSV4 U13176 ( .A1(n20050), .A2(n22138), .ZN(n25607) );
  NAND2HSV4 U13177 ( .A1(n11911), .A2(n18843), .ZN(n19831) );
  INHSV4 U13178 ( .I(n19062), .ZN(n19065) );
  CLKNAND2HSV2 U13179 ( .A1(n21241), .A2(n22085), .ZN(n12569) );
  CLKNAND2HSV2 U13180 ( .A1(n19239), .A2(n19190), .ZN(n19266) );
  AOI21HSV2 U13181 ( .A1(n21239), .A2(n21703), .B(n21238), .ZN(n21240) );
  XOR2HSV2 U13182 ( .A1(n11912), .A2(n22888), .Z(n22890) );
  XNOR2HSV4 U13183 ( .A1(n22878), .A2(n22879), .ZN(n11912) );
  OAI21HSV4 U13184 ( .A1(n19126), .A2(n19128), .B(n11913), .ZN(n12606) );
  AOI21HSV4 U13185 ( .A1(n12601), .A2(n12602), .B(n12600), .ZN(n11913) );
  XNOR2HSV4 U13186 ( .A1(n27819), .A2(n27818), .ZN(n27820) );
  CLKNAND2HSV4 U13187 ( .A1(n25622), .A2(\pe7/got [12]), .ZN(n12360) );
  CLKNAND2HSV8 U13188 ( .A1(n21421), .A2(\pe5/ti_7t [15]), .ZN(n23275) );
  CLKNAND2HSV3 U13189 ( .A1(\pe8/ti_1 ), .A2(\pe8/got [14]), .ZN(n16298) );
  CLKNAND2HSV4 U13190 ( .A1(n22084), .A2(n17767), .ZN(n21216) );
  CLKNAND2HSV4 U13191 ( .A1(\pe1/aot [14]), .A2(n26431), .ZN(n16222) );
  NAND2HSV2 U13192 ( .A1(n18648), .A2(n23717), .ZN(n28344) );
  NAND2HSV2 U13193 ( .A1(n14748), .A2(n14746), .ZN(n14751) );
  AOI21HSV4 U13194 ( .A1(n16167), .A2(n16166), .B(n16165), .ZN(n16171) );
  XNOR2HSV4 U13195 ( .A1(n21520), .A2(n21519), .ZN(po5) );
  AND3HSV8 U13196 ( .A1(n25653), .A2(n17215), .A3(n17602), .Z(n17199) );
  CLKXOR2HSV4 U13197 ( .A1(n22367), .A2(n22366), .Z(n22369) );
  CLKXOR2HSV4 U13198 ( .A1(n18666), .A2(n18665), .Z(n18670) );
  CLKXOR2HSV2 U13199 ( .A1(n18670), .A2(n18669), .Z(n18671) );
  AOI21HSV4 U13200 ( .A1(n20867), .A2(n14526), .B(n20866), .ZN(n20927) );
  INHSV4 U13201 ( .I(n16734), .ZN(n16848) );
  INHSV4 U13202 ( .I(n21157), .ZN(n13658) );
  CLKNAND2HSV4 U13203 ( .A1(n28706), .A2(n19837), .ZN(n19839) );
  INHSV6 U13204 ( .I(n14630), .ZN(n28664) );
  CLKNAND2HSV2 U13205 ( .A1(n15755), .A2(n11917), .ZN(n15756) );
  CLKNAND2HSV2 U13206 ( .A1(n15756), .A2(n15757), .ZN(n15808) );
  XNOR2HSV4 U13207 ( .A1(n26152), .A2(n26151), .ZN(n26155) );
  CLKNAND2HSV2 U13208 ( .A1(n21642), .A2(n21714), .ZN(n13308) );
  BUFHSV8 U13209 ( .I(n21422), .Z(n21346) );
  NAND2HSV4 U13210 ( .A1(n21230), .A2(n21229), .ZN(n21297) );
  INHSV4 U13211 ( .I(n21297), .ZN(n21298) );
  INHSV4 U13212 ( .I(n20393), .ZN(n13788) );
  CLKNHSV6 U13213 ( .I(n17023), .ZN(n28630) );
  BUFHSV4 U13214 ( .I(n16781), .Z(n16850) );
  XOR3HSV2 U13215 ( .A1(n16687), .A2(n16688), .A3(n16690), .Z(n16691) );
  CLKXOR2HSV4 U13216 ( .A1(n16652), .A2(n16651), .Z(n16654) );
  INHSV4 U13217 ( .I(n16654), .ZN(n16655) );
  XOR3HSV2 U13218 ( .A1(\pe7/phq [4]), .A2(n19241), .A3(n11961), .Z(n11960) );
  XNOR2HSV4 U13219 ( .A1(n23952), .A2(n23951), .ZN(n23953) );
  XNOR2HSV4 U13220 ( .A1(n17816), .A2(n17815), .ZN(n17818) );
  XNOR2HSV4 U13221 ( .A1(n11914), .A2(n17765), .ZN(n17816) );
  CLKNHSV2 U13222 ( .I(n17766), .ZN(n11914) );
  XNOR2HSV4 U13223 ( .A1(n15384), .A2(n15383), .ZN(n15385) );
  CLKNHSV2 U13224 ( .I(n22562), .ZN(n22561) );
  CLKNAND2HSV4 U13225 ( .A1(n25637), .A2(n17962), .ZN(n17992) );
  INHSV2 U13226 ( .I(\pe11/bq[16] ), .ZN(n20326) );
  AND2HSV2 U13227 ( .A1(n12517), .A2(\pe5/got [3]), .Z(n11973) );
  CLKNAND2HSV2 U13228 ( .A1(n21993), .A2(n25128), .ZN(n21996) );
  CLKNAND2HSV4 U13229 ( .A1(n15102), .A2(n15101), .ZN(n15144) );
  NAND2HSV2 U13230 ( .A1(n14992), .A2(n14993), .ZN(n14997) );
  CLKNAND2HSV2 U13231 ( .A1(n16245), .A2(\pe1/got [13]), .ZN(n16249) );
  NAND2HSV4 U13232 ( .A1(n14080), .A2(n28592), .ZN(n15834) );
  NAND2HSV4 U13233 ( .A1(n22916), .A2(n11915), .ZN(n25370) );
  INHSV2 U13234 ( .I(n22917), .ZN(n11915) );
  NOR2HSV4 U13235 ( .A1(n18190), .A2(n18207), .ZN(n18196) );
  NAND2HSV4 U13236 ( .A1(n18196), .A2(n18197), .ZN(n18275) );
  CLKNAND2HSV2 U13237 ( .A1(n12517), .A2(n28645), .ZN(n21551) );
  CLKXOR2HSV2 U13238 ( .A1(n21551), .A2(n21550), .Z(n21552) );
  XNOR2HSV4 U13239 ( .A1(n11916), .A2(n20688), .ZN(n20697) );
  XOR2HSV2 U13240 ( .A1(n20683), .A2(n20684), .Z(n11916) );
  CLKAND2HSV4 U13241 ( .A1(n22886), .A2(n21987), .Z(n13963) );
  CLKXOR2HSV4 U13242 ( .A1(n23712), .A2(n23711), .Z(n23713) );
  XNOR2HSV4 U13243 ( .A1(n23714), .A2(n23713), .ZN(\pe6/poht [12]) );
  NAND2HSV2 U13244 ( .A1(n24322), .A2(n14071), .ZN(n13313) );
  NAND2HSV2 U13245 ( .A1(n13312), .A2(n13313), .ZN(n13314) );
  INHSV2 U13246 ( .I(n15753), .ZN(n11917) );
  NAND2HSV4 U13247 ( .A1(n15844), .A2(n25131), .ZN(n15753) );
  XNOR2HSV4 U13248 ( .A1(n11918), .A2(n15172), .ZN(n12098) );
  XNOR2HSV4 U13249 ( .A1(n11919), .A2(n15165), .ZN(n11918) );
  XNOR2HSV4 U13250 ( .A1(n15166), .A2(n15167), .ZN(n11919) );
  NAND2HSV8 U13251 ( .A1(n21966), .A2(n21570), .ZN(n27112) );
  INHSV4 U13252 ( .I(n18703), .ZN(n18701) );
  NAND2HSV4 U13253 ( .A1(n18701), .A2(n18700), .ZN(n18705) );
  OAI21HSV4 U13254 ( .A1(n19829), .A2(n19840), .B(n11920), .ZN(n19975) );
  NOR2HSV4 U13255 ( .A1(n19827), .A2(n19828), .ZN(n11920) );
  CLKNAND2HSV2 U13256 ( .A1(n28946), .A2(n14072), .ZN(n24450) );
  CLKNAND2HSV4 U13257 ( .A1(n16343), .A2(n16307), .ZN(n16296) );
  XNOR2HSV4 U13258 ( .A1(n11921), .A2(n16342), .ZN(n12531) );
  NAND2HSV4 U13259 ( .A1(n18673), .A2(\pe8/pvq [5]), .ZN(n16409) );
  CLKNHSV2 U13260 ( .I(n23466), .ZN(n12056) );
  XNOR2HSV4 U13261 ( .A1(n18085), .A2(n18084), .ZN(n23466) );
  NAND2HSV4 U13262 ( .A1(n17908), .A2(n17907), .ZN(n17909) );
  CLKNAND2HSV4 U13263 ( .A1(n20983), .A2(n14757), .ZN(n20849) );
  NAND2HSV2 U13264 ( .A1(n17916), .A2(n17915), .ZN(n17946) );
  NAND2HSV2 U13265 ( .A1(n17889), .A2(n17890), .ZN(n17916) );
  INHSV4 U13266 ( .I(n15028), .ZN(n15026) );
  NAND3HSV4 U13267 ( .A1(n12446), .A2(n12447), .A3(n12444), .ZN(n25054) );
  INAND2HSV4 U13268 ( .A1(n11922), .B1(n12445), .ZN(n12444) );
  CLKNHSV2 U13269 ( .I(n25045), .ZN(n11922) );
  INHSV2 U13270 ( .I(n20983), .ZN(n20984) );
  CLKNAND2HSV4 U13271 ( .A1(n19474), .A2(n19472), .ZN(n19458) );
  CLKNAND2HSV4 U13272 ( .A1(n20272), .A2(\pe11/got [16]), .ZN(n14748) );
  CLKNAND2HSV8 U13273 ( .A1(n22993), .A2(n22992), .ZN(n18989) );
  CLKNHSV6 U13274 ( .I(n18989), .ZN(n18987) );
  XOR2HSV4 U13275 ( .A1(n15962), .A2(n15961), .Z(n23373) );
  INHSV4 U13276 ( .I(n21004), .ZN(n28426) );
  NAND2HSV0 U13277 ( .A1(n28426), .A2(\pe8/got [6]), .ZN(n25207) );
  INHSV4 U13278 ( .I(\pe1/bq[16] ), .ZN(n17302) );
  CLKNAND2HSV4 U13279 ( .A1(\pe7/bq[16] ), .A2(\pe7/aot [16]), .ZN(n12694) );
  AOI21HSV4 U13280 ( .A1(n20188), .A2(n20255), .B(n20620), .ZN(n20163) );
  NAND2HSV4 U13281 ( .A1(n20163), .A2(n20162), .ZN(n20219) );
  NAND2HSV2 U13282 ( .A1(\pe11/aot [16]), .A2(\pe11/bq[16] ), .ZN(n14753) );
  BUFHSV6 U13283 ( .I(\pe8/ctrq ), .Z(n18673) );
  CLKNAND2HSV2 U13284 ( .A1(n17215), .A2(n17617), .ZN(n16287) );
  INHSV2 U13285 ( .I(n14397), .ZN(n26033) );
  NOR2HSV4 U13286 ( .A1(n16749), .A2(n22503), .ZN(n22504) );
  CLKNAND2HSV2 U13287 ( .A1(n25692), .A2(n25691), .ZN(n28390) );
  INOR2HSV4 U13288 ( .A1(\pe3/ti_7t [8]), .B1(n21722), .ZN(n15236) );
  NAND3HSV3 U13289 ( .A1(n21868), .A2(n21866), .A3(n21163), .ZN(n27344) );
  NAND2HSV4 U13290 ( .A1(n11923), .A2(n21166), .ZN(n21868) );
  NOR2HSV4 U13291 ( .A1(n21218), .A2(n11924), .ZN(n11923) );
  INHSV4 U13292 ( .I(n21165), .ZN(n11924) );
  CLKNAND2HSV4 U13293 ( .A1(n11925), .A2(n16330), .ZN(n16381) );
  CLKNAND2HSV4 U13294 ( .A1(n16329), .A2(n16328), .ZN(n11925) );
  NAND2HSV4 U13295 ( .A1(n14138), .A2(n14137), .ZN(n14142) );
  NAND2HSV2 U13296 ( .A1(n25648), .A2(n25420), .ZN(n14185) );
  INHSV4 U13297 ( .I(n14185), .ZN(n14197) );
  CLKNAND2HSV2 U13298 ( .A1(n19576), .A2(n12178), .ZN(n12114) );
  INHSV4 U13299 ( .I(n14268), .ZN(n14269) );
  NAND2HSV4 U13300 ( .A1(\pe3/pvq [1]), .A2(\pe3/phq [1]), .ZN(n15004) );
  OAI22HSV2 U13301 ( .A1(n15936), .A2(n15004), .B1(\pe3/phq [1]), .B2(
        \pe3/pvq [1]), .ZN(n15006) );
  NAND2HSV2 U13302 ( .A1(n15754), .A2(n15753), .ZN(n15757) );
  NAND2HSV2 U13303 ( .A1(n17207), .A2(n17206), .ZN(n17208) );
  INHSV4 U13304 ( .I(n17208), .ZN(n17211) );
  INHSV6 U13305 ( .I(n22680), .ZN(n28603) );
  NAND2HSV2 U13306 ( .A1(n28603), .A2(n28479), .ZN(n26151) );
  CLKNAND2HSV2 U13307 ( .A1(n13321), .A2(n13322), .ZN(n13323) );
  CLKNAND2HSV2 U13308 ( .A1(n13320), .A2(n11926), .ZN(n13321) );
  CLKNAND2HSV2 U13309 ( .A1(n11928), .A2(n11927), .ZN(n11926) );
  CLKNHSV2 U13310 ( .I(n13318), .ZN(n11927) );
  CLKNHSV2 U13311 ( .I(n13319), .ZN(n11928) );
  CLKXOR2HSV4 U13312 ( .A1(n26217), .A2(n26216), .Z(n13485) );
  CLKXOR2HSV4 U13313 ( .A1(n26219), .A2(n13485), .Z(n13486) );
  CLKXOR2HSV4 U13314 ( .A1(n12830), .A2(n12831), .Z(n12832) );
  CLKNAND2HSV2 U13315 ( .A1(n12833), .A2(n12832), .ZN(n12834) );
  OAI31HSV2 U13316 ( .A1(n28368), .A2(n28367), .A3(n28286), .B(n28366), .ZN(
        n28372) );
  CLKNAND2HSV4 U13317 ( .A1(n12727), .A2(n20930), .ZN(n20998) );
  INHSV4 U13318 ( .I(n15014), .ZN(n15012) );
  NAND2HSV4 U13319 ( .A1(n15012), .A2(n15011), .ZN(n15016) );
  NAND2HSV2 U13320 ( .A1(\pe3/aot [10]), .A2(n23336), .ZN(n15112) );
  CLKNHSV2 U13321 ( .I(\pe3/ctrq ), .ZN(n15936) );
  CLKXOR2HSV4 U13322 ( .A1(n21627), .A2(n21626), .Z(n13060) );
  CLKXOR2HSV4 U13323 ( .A1(n21553), .A2(n21552), .Z(n13312) );
  XOR2HSV0 U13324 ( .A1(n25978), .A2(n25979), .Z(\pe6/poht [8]) );
  NAND2HSV2 U13325 ( .A1(n22431), .A2(n22430), .ZN(n22433) );
  XNOR2HSV4 U13326 ( .A1(n18134), .A2(n18133), .ZN(n18135) );
  CLKNAND2HSV4 U13327 ( .A1(n18399), .A2(n28134), .ZN(n18136) );
  XOR2HSV4 U13328 ( .A1(n18136), .A2(n18135), .Z(n18137) );
  NAND2HSV4 U13329 ( .A1(n28969), .A2(n14926), .ZN(n12727) );
  CLKNAND2HSV4 U13330 ( .A1(n28988), .A2(n22418), .ZN(n22690) );
  NAND2HSV4 U13331 ( .A1(n12323), .A2(n18280), .ZN(n12321) );
  CLKNAND2HSV4 U13332 ( .A1(n21299), .A2(n21300), .ZN(n25357) );
  CLKNAND2HSV4 U13333 ( .A1(\pe6/bq[15] ), .A2(\pe6/aot [16]), .ZN(n14112) );
  XOR2HSV4 U13334 ( .A1(n14113), .A2(n14112), .Z(n14144) );
  DELHS1 U13335 ( .I(\pe7/got [14]), .Z(n11929) );
  INHSV4 U13336 ( .I(n12481), .ZN(n22081) );
  NOR2HSV8 U13337 ( .A1(n22081), .A2(n16536), .ZN(n18833) );
  NAND2HSV4 U13338 ( .A1(n11930), .A2(n12491), .ZN(n18467) );
  INHSV2 U13339 ( .I(n12490), .ZN(n11930) );
  NOR2HSV2 U13340 ( .A1(n13673), .A2(n18336), .ZN(n12490) );
  INHSV4 U13341 ( .I(\pe3/ti_1 ), .ZN(n15162) );
  INHSV4 U13342 ( .I(n15162), .ZN(n15044) );
  CLKNAND2HSV4 U13343 ( .A1(n22499), .A2(n22498), .ZN(n22502) );
  CLKXOR2HSV4 U13344 ( .A1(n22755), .A2(n22754), .Z(n22757) );
  XNOR2HSV2 U13345 ( .A1(n22757), .A2(n22756), .ZN(n22760) );
  CLKNAND2HSV4 U13346 ( .A1(n17745), .A2(n17744), .ZN(n17859) );
  INHSV2 U13347 ( .I(n14621), .ZN(n14619) );
  DELHS1 U13348 ( .I(n24378), .Z(n11931) );
  NAND2HSV2 U13349 ( .A1(\pe2/bq[15] ), .A2(\pe2/aot [16]), .ZN(n17635) );
  NAND2HSV4 U13350 ( .A1(n21421), .A2(\pe5/ti_7t [13]), .ZN(n21338) );
  BUFHSV6 U13351 ( .I(\pe5/got [8]), .Z(n24340) );
  INHSV4 U13352 ( .I(n21109), .ZN(n21006) );
  INHSV4 U13353 ( .I(n17692), .ZN(n17695) );
  NAND2HSV4 U13354 ( .A1(n17695), .A2(n17694), .ZN(n11939) );
  BUFHSV2 U13355 ( .I(\pe3/aot [13]), .Z(n11932) );
  CLKNAND2HSV2 U13356 ( .A1(n19834), .A2(n19833), .ZN(n12242) );
  CLKNAND2HSV2 U13357 ( .A1(n24075), .A2(n23180), .ZN(n23181) );
  CLKNAND2HSV4 U13358 ( .A1(n12767), .A2(n12768), .ZN(n12770) );
  INHSV4 U13359 ( .I(n20457), .ZN(n23460) );
  INHSV4 U13360 ( .I(n28016), .ZN(n28134) );
  NOR2HSV8 U13361 ( .A1(n16285), .A2(n17287), .ZN(n17225) );
  INHSV2 U13362 ( .I(n21222), .ZN(n11933) );
  CLKNAND2HSV2 U13363 ( .A1(n11933), .A2(n28693), .ZN(n21167) );
  CLKNAND2HSV4 U13364 ( .A1(n14642), .A2(\pe5/got [15]), .ZN(n14675) );
  NAND2HSV2 U13365 ( .A1(n13487), .A2(n13486), .ZN(n13488) );
  CLKNAND2HSV2 U13366 ( .A1(n17648), .A2(n17647), .ZN(n17671) );
  XNOR2HSV4 U13367 ( .A1(n11934), .A2(n14533), .ZN(n14541) );
  XNOR2HSV4 U13368 ( .A1(n12174), .A2(n14534), .ZN(n11934) );
  INHSV4 U13369 ( .I(n28080), .ZN(n28373) );
  NOR2HSV2 U13370 ( .A1(n26916), .A2(n13030), .ZN(n22791) );
  CLKNAND2HSV2 U13371 ( .A1(n17800), .A2(n17799), .ZN(n17801) );
  XNOR2HSV2 U13372 ( .A1(n17719), .A2(n17718), .ZN(n17723) );
  NAND2HSV4 U13373 ( .A1(n19354), .A2(n19353), .ZN(n19355) );
  NAND2HSV4 U13374 ( .A1(n19356), .A2(n19355), .ZN(n19364) );
  CLKXOR2HSV4 U13375 ( .A1(n26644), .A2(n26643), .Z(n26647) );
  INHSV4 U13376 ( .I(n19900), .ZN(n28706) );
  CLKNAND2HSV2 U13377 ( .A1(n28706), .A2(n22136), .ZN(n20044) );
  CLKNAND2HSV2 U13378 ( .A1(n22375), .A2(n28669), .ZN(n13502) );
  CLKNHSV6 U13379 ( .I(n20999), .ZN(n12441) );
  OAI21HSV4 U13380 ( .A1(n16738), .A2(n23473), .B(n16737), .ZN(n16742) );
  CLKNAND2HSV4 U13381 ( .A1(n12364), .A2(n16641), .ZN(n16816) );
  CLKNAND2HSV2 U13382 ( .A1(n16816), .A2(n16759), .ZN(n16769) );
  CLKNAND2HSV2 U13383 ( .A1(n16511), .A2(\pe8/got [11]), .ZN(n16366) );
  XNOR2HSV2 U13384 ( .A1(n16366), .A2(n16365), .ZN(n16378) );
  XNOR2HSV4 U13385 ( .A1(n20209), .A2(n20208), .ZN(n20211) );
  XOR3HSV2 U13386 ( .A1(n16830), .A2(n16829), .A3(n16828), .Z(n16832) );
  CLKXOR2HSV4 U13387 ( .A1(n24432), .A2(n24431), .Z(n24433) );
  XNOR2HSV4 U13388 ( .A1(n24434), .A2(n24433), .ZN(n24435) );
  BUFHSV8 U13389 ( .I(\pe8/bq[15] ), .Z(n16400) );
  OAI21HSV4 U13390 ( .A1(pov5[15]), .A2(n23277), .B(n23276), .ZN(n13882) );
  NAND2HSV2 U13391 ( .A1(\pe1/aot [14]), .A2(n14991), .ZN(n14992) );
  DELHS1 U13392 ( .I(n25270), .Z(n11935) );
  DELHS1 U13393 ( .I(n21326), .Z(n11936) );
  NAND2HSV2 U13394 ( .A1(\pe2/aot [15]), .A2(\pe2/bq[14] ), .ZN(n17719) );
  INHSV4 U13395 ( .I(n11937), .ZN(n21005) );
  INHSV2 U13396 ( .I(n22199), .ZN(n23757) );
  INHSV4 U13397 ( .I(n15093), .ZN(n15036) );
  CLKNAND2HSV2 U13398 ( .A1(n15037), .A2(n15036), .ZN(n15038) );
  NAND3HSV3 U13399 ( .A1(n24075), .A2(n24074), .A3(n24073), .ZN(n25408) );
  NAND2HSV2 U13400 ( .A1(n25408), .A2(n24271), .ZN(n24272) );
  CLKNAND2HSV4 U13401 ( .A1(n11939), .A2(n12701), .ZN(n23471) );
  INHSV4 U13402 ( .I(n14764), .ZN(n14931) );
  CLKNHSV2 U13403 ( .I(n11940), .ZN(n25659) );
  CLKNAND2HSV2 U13404 ( .A1(n14764), .A2(n11941), .ZN(n11940) );
  CLKNHSV2 U13405 ( .I(n14684), .ZN(n11941) );
  NAND2HSV4 U13406 ( .A1(n14625), .A2(n14624), .ZN(n14764) );
  NOR2HSV4 U13407 ( .A1(n16439), .A2(n16438), .ZN(n16450) );
  NAND2HSV4 U13408 ( .A1(n11942), .A2(n16657), .ZN(n16662) );
  CLKNAND2HSV4 U13409 ( .A1(n16656), .A2(n16655), .ZN(n11942) );
  CLKNAND2HSV4 U13410 ( .A1(n16670), .A2(n25255), .ZN(n16625) );
  NAND2HSV0 U13411 ( .A1(n28584), .A2(n26603), .ZN(n24606) );
  OAI21HSV4 U13412 ( .A1(n15428), .A2(n21979), .B(n15420), .ZN(n15421) );
  INHSV2 U13413 ( .I(n14607), .ZN(n14610) );
  NAND2HSV2 U13414 ( .A1(n24411), .A2(n24635), .ZN(n14607) );
  INHSV6 U13415 ( .I(\pe7/ti_1 ), .ZN(n19243) );
  INHSV2 U13416 ( .I(n19243), .ZN(n25622) );
  XNOR2HSV4 U13417 ( .A1(n12716), .A2(n11943), .ZN(n23115) );
  NAND3HSV4 U13418 ( .A1(n12715), .A2(n12713), .A3(n12714), .ZN(n11943) );
  XNOR2HSV4 U13419 ( .A1(n19747), .A2(n19746), .ZN(n19748) );
  NAND2HSV4 U13420 ( .A1(n15415), .A2(n15414), .ZN(n15422) );
  CLKNAND2HSV2 U13421 ( .A1(n21065), .A2(n27231), .ZN(n17691) );
  CLKNAND2HSV4 U13422 ( .A1(n28690), .A2(n18765), .ZN(n18771) );
  INHSV4 U13423 ( .I(n18269), .ZN(n18267) );
  XNOR2HSV4 U13424 ( .A1(n13063), .A2(n13064), .ZN(n13065) );
  NAND2HSV2 U13425 ( .A1(n25060), .A2(n14070), .ZN(n22558) );
  INHSV4 U13426 ( .I(n25260), .ZN(n22499) );
  INHSV2 U13427 ( .I(n17414), .ZN(n17411) );
  CLKNAND2HSV4 U13428 ( .A1(n13125), .A2(n11944), .ZN(n17414) );
  NAND2HSV4 U13429 ( .A1(n11946), .A2(n11945), .ZN(n11944) );
  INHSV4 U13430 ( .I(n13123), .ZN(n11945) );
  INHSV2 U13431 ( .I(n13124), .ZN(n11946) );
  XNOR2HSV2 U13432 ( .A1(n26756), .A2(n26755), .ZN(n26757) );
  OAI22HSV4 U13433 ( .A1(n11948), .A2(n11947), .B1(n14007), .B2(n17346), .ZN(
        n17358) );
  CLKNAND2HSV2 U13434 ( .A1(n13957), .A2(n17351), .ZN(n11947) );
  CLKNHSV2 U13435 ( .I(n17352), .ZN(n11948) );
  CLKNAND2HSV2 U13436 ( .A1(n12039), .A2(n12037), .ZN(n12036) );
  INAND2HSV4 U13437 ( .A1(n17274), .B1(n11949), .ZN(n17276) );
  CLKNAND2HSV2 U13438 ( .A1(n17275), .A2(n26595), .ZN(n11949) );
  NAND2HSV2 U13439 ( .A1(n12396), .A2(n22507), .ZN(n11950) );
  CLKNAND2HSV2 U13440 ( .A1(n25597), .A2(n25602), .ZN(n19832) );
  INHSV4 U13441 ( .I(n19832), .ZN(n19833) );
  BUFHSV8 U13442 ( .I(n29052), .Z(n12023) );
  AOI21HSV2 U13443 ( .A1(n18456), .A2(n18455), .B(n11951), .ZN(n18523) );
  CLKNHSV2 U13444 ( .I(n18468), .ZN(n11951) );
  XNOR2HSV4 U13445 ( .A1(n11952), .A2(n22800), .ZN(n29028) );
  CLKNAND2HSV2 U13446 ( .A1(n27980), .A2(n15813), .ZN(n11952) );
  DELHS1 U13447 ( .I(n17785), .Z(n11953) );
  CLKNAND2HSV1 U13448 ( .A1(n13042), .A2(n13043), .ZN(n13044) );
  INHSV4 U13449 ( .I(n25490), .ZN(n20178) );
  XOR2HSV4 U13450 ( .A1(n23226), .A2(n23225), .Z(n23227) );
  CLKXOR2HSV4 U13451 ( .A1(n12607), .A2(n19144), .Z(n25517) );
  NAND2HSV4 U13452 ( .A1(n27284), .A2(n27283), .ZN(n28702) );
  NAND2HSV2 U13453 ( .A1(n26444), .A2(n27184), .ZN(n17178) );
  AOI31HSV2 U13454 ( .A1(n16798), .A2(n16797), .A3(n16796), .B(n16795), .ZN(
        n16799) );
  NAND3HSV4 U13455 ( .A1(n20312), .A2(n20311), .A3(n20310), .ZN(n20401) );
  NAND2HSV4 U13456 ( .A1(n16237), .A2(n11954), .ZN(n16281) );
  CLKNAND2HSV4 U13457 ( .A1(n16236), .A2(n16235), .ZN(n11954) );
  CLKNAND2HSV4 U13458 ( .A1(n28952), .A2(n28134), .ZN(n18437) );
  NAND2HSV4 U13459 ( .A1(n18340), .A2(n18339), .ZN(n28952) );
  CLKNAND2HSV4 U13460 ( .A1(n28809), .A2(n22085), .ZN(n27121) );
  CLKXOR2HSV4 U13461 ( .A1(n27897), .A2(n27896), .Z(n27898) );
  CLKXOR2HSV4 U13462 ( .A1(n27868), .A2(n27867), .Z(n27869) );
  INHSV8 U13463 ( .I(n26929), .ZN(n11955) );
  NOR2HSV4 U13464 ( .A1(n11955), .A2(n22796), .ZN(n12507) );
  OAI21HSV2 U13465 ( .A1(n14975), .A2(n14974), .B(n14978), .ZN(n14976) );
  NOR2HSV4 U13466 ( .A1(n29052), .A2(ctro1), .ZN(n14978) );
  CLKNAND2HSV8 U13467 ( .A1(n21000), .A2(n20999), .ZN(n21001) );
  CLKNAND2HSV4 U13468 ( .A1(n20132), .A2(n17117), .ZN(n20130) );
  CLKNAND2HSV4 U13469 ( .A1(n17118), .A2(n20130), .ZN(n22692) );
  NAND2HSV4 U13470 ( .A1(n12378), .A2(n21461), .ZN(n21462) );
  NAND3HSV4 U13471 ( .A1(n17930), .A2(\pe9/ti_1 ), .A3(\pe9/got [14]), .ZN(
        n17931) );
  INHSV4 U13472 ( .I(n20765), .ZN(n20764) );
  NAND2HSV4 U13473 ( .A1(n20764), .A2(n20763), .ZN(n12201) );
  XNOR2HSV4 U13474 ( .A1(n20845), .A2(n20846), .ZN(n24883) );
  XNOR2HSV4 U13475 ( .A1(n20842), .A2(n11956), .ZN(n20845) );
  CLKNHSV2 U13476 ( .I(n20841), .ZN(n11956) );
  NAND2HSV4 U13477 ( .A1(n27485), .A2(n28429), .ZN(n21057) );
  INHSV4 U13478 ( .I(n21057), .ZN(n13873) );
  XNOR2HSV4 U13479 ( .A1(n11957), .A2(n23950), .ZN(n23951) );
  XNOR2HSV4 U13480 ( .A1(n23948), .A2(n23949), .ZN(n11957) );
  NAND2HSV2 U13481 ( .A1(\pe7/aot [15]), .A2(\pe7/bq[16] ), .ZN(n19198) );
  NAND2HSV4 U13482 ( .A1(n27112), .A2(n24637), .ZN(n13222) );
  CLKNAND2HSV4 U13483 ( .A1(n14111), .A2(n11958), .ZN(n14145) );
  NAND2HSV4 U13484 ( .A1(n11959), .A2(n12435), .ZN(n11958) );
  NAND2HSV2 U13485 ( .A1(n12115), .A2(n12114), .ZN(n12117) );
  AND2HSV8 U13486 ( .A1(n23803), .A2(n23802), .Z(n23676) );
  CLKNAND2HSV4 U13487 ( .A1(n23677), .A2(n23676), .ZN(n26679) );
  AOI22HSV4 U13488 ( .A1(n24634), .A2(n20868), .B1(n28971), .B2(n21347), .ZN(
        n20926) );
  XNOR2HSV4 U13489 ( .A1(n12232), .A2(n12236), .ZN(n20865) );
  BUFHSV4 U13490 ( .I(n23266), .Z(n21452) );
  CLKNAND2HSV2 U13491 ( .A1(n14608), .A2(n14607), .ZN(n14612) );
  CLKNAND2HSV2 U13492 ( .A1(n17666), .A2(n21696), .ZN(n17644) );
  CLKNAND2HSV2 U13493 ( .A1(n17642), .A2(n17643), .ZN(n17666) );
  NAND2HSV2 U13494 ( .A1(\pe6/bq[16] ), .A2(\pe6/aot [13]), .ZN(n13634) );
  INHSV6 U13495 ( .I(n14674), .ZN(n14685) );
  NOR2HSV4 U13496 ( .A1(n12362), .A2(n12328), .ZN(n12316) );
  INHSV4 U13497 ( .I(n27121), .ZN(n17770) );
  CLKNHSV2 U13498 ( .I(n19494), .ZN(n11961) );
  NAND2HSV4 U13499 ( .A1(n11963), .A2(n11962), .ZN(n19179) );
  INHSV2 U13500 ( .I(n19178), .ZN(n11962) );
  INHSV2 U13501 ( .I(n19177), .ZN(n11963) );
  NAND2HSV2 U13502 ( .A1(n25950), .A2(\pe6/got [3]), .ZN(n23712) );
  MUX2NHSV2 U13503 ( .I0(n12879), .I1(n20314), .S(n11964), .ZN(n25513) );
  NOR2HSV4 U13504 ( .A1(n11966), .A2(n11965), .ZN(n11964) );
  CLKNAND2HSV2 U13505 ( .A1(n20253), .A2(n11967), .ZN(n11966) );
  CLKNAND2HSV2 U13506 ( .A1(n11969), .A2(n11968), .ZN(n11967) );
  CLKNHSV2 U13507 ( .I(n20619), .ZN(n11968) );
  CLKNHSV2 U13508 ( .I(n20348), .ZN(n11969) );
  NAND2HSV2 U13509 ( .A1(n25060), .A2(n14065), .ZN(n23226) );
  NAND2HSV4 U13510 ( .A1(n17731), .A2(n12765), .ZN(n17732) );
  NAND2HSV4 U13511 ( .A1(n17733), .A2(n17732), .ZN(n17738) );
  CLKNAND2HSV4 U13512 ( .A1(n17925), .A2(n17924), .ZN(n17960) );
  NAND2HSV2 U13513 ( .A1(n28927), .A2(n25030), .ZN(n21964) );
  INHSV2 U13514 ( .I(n19263), .ZN(n23137) );
  NOR2HSV4 U13515 ( .A1(n23137), .A2(n19267), .ZN(n19265) );
  INHSV4 U13516 ( .I(n14786), .ZN(n24406) );
  NOR2HSV4 U13517 ( .A1(n27942), .A2(n26932), .ZN(n22041) );
  NAND2HSV4 U13518 ( .A1(n21253), .A2(\pe2/pvq [5]), .ZN(n17677) );
  XOR3HSV4 U13519 ( .A1(\pe2/phq [5]), .A2(n17677), .A3(n17676), .Z(n17685) );
  CLKNAND2HSV2 U13520 ( .A1(n14040), .A2(\pe3/bq[10] ), .ZN(n15110) );
  CLKXOR2HSV2 U13521 ( .A1(n15110), .A2(n15109), .Z(n15114) );
  INHSV4 U13522 ( .I(n17628), .ZN(n17630) );
  XNOR2HSV4 U13523 ( .A1(n11970), .A2(n12074), .ZN(n12073) );
  XNOR2HSV4 U13524 ( .A1(n18261), .A2(n18230), .ZN(n11970) );
  NOR2HSV4 U13525 ( .A1(n18955), .A2(n14123), .ZN(n14125) );
  CLKNHSV2 U13526 ( .I(\pe6/got [14]), .ZN(n14123) );
  INHSV4 U13527 ( .I(n22566), .ZN(n25216) );
  NAND2HSV2 U13528 ( .A1(n25216), .A2(n27196), .ZN(n22580) );
  NAND2HSV4 U13529 ( .A1(n12544), .A2(n12543), .ZN(n16623) );
  NOR2HSV4 U13530 ( .A1(n22909), .A2(n22821), .ZN(n22889) );
  CLKNAND2HSV2 U13531 ( .A1(n22915), .A2(n26925), .ZN(n22909) );
  CLKNHSV6 U13532 ( .I(n18211), .ZN(n18195) );
  CLKNAND2HSV8 U13533 ( .A1(n18195), .A2(n18330), .ZN(n18197) );
  NAND2HSV4 U13534 ( .A1(n18324), .A2(n11971), .ZN(n18456) );
  INHSV4 U13535 ( .I(n18323), .ZN(n11971) );
  MUX2NHSV4 U13536 ( .I0(n18321), .I1(n18320), .S(n18319), .ZN(n18323) );
  AOI21HSV2 U13537 ( .A1(n20207), .A2(n25502), .B(n20206), .ZN(n20208) );
  CLKNAND2HSV4 U13538 ( .A1(\pe11/aot [15]), .A2(\pe11/bq[13] ), .ZN(n20268)
         );
  XOR3HSV2 U13539 ( .A1(n11972), .A2(n27546), .A3(n27545), .Z(\pe2/poht [4])
         );
  XNOR2HSV4 U13540 ( .A1(n27542), .A2(n27541), .ZN(n11972) );
  AOI22HSV2 U13541 ( .A1(n21423), .A2(n24634), .B1(n28973), .B2(n21347), .ZN(
        n20997) );
  NAND2HSV4 U13542 ( .A1(n22765), .A2(n22764), .ZN(n23219) );
  AO22HSV4 U13543 ( .A1(n14070), .A2(n16663), .B1(n28704), .B2(n16755), .Z(
        n16664) );
  CLKNHSV6 U13544 ( .I(n17960), .ZN(n12684) );
  INHSV4 U13545 ( .I(n17961), .ZN(n12685) );
  CLKNAND2HSV8 U13546 ( .A1(n12685), .A2(n12684), .ZN(n18044) );
  CLKNAND2HSV4 U13547 ( .A1(n15094), .A2(n15053), .ZN(n15097) );
  XNOR2HSV4 U13548 ( .A1(n11973), .A2(n24337), .ZN(n24338) );
  NOR2HSV2 U13549 ( .A1(n21009), .A2(n21014), .ZN(n21010) );
  NOR2HSV4 U13550 ( .A1(n11975), .A2(n11974), .ZN(n21009) );
  CLKNAND2HSV2 U13551 ( .A1(n17861), .A2(n27354), .ZN(n11974) );
  CLKNHSV2 U13552 ( .I(n14044), .ZN(n11975) );
  CLKXOR2HSV4 U13553 ( .A1(n12842), .A2(n12843), .Z(n12844) );
  NAND2HSV8 U13554 ( .A1(n21339), .A2(n21338), .ZN(n21718) );
  NAND2HSV4 U13555 ( .A1(n28790), .A2(n28134), .ZN(n18520) );
  NOR2HSV4 U13556 ( .A1(n26602), .A2(n26624), .ZN(n23813) );
  CLKNAND2HSV2 U13557 ( .A1(n12517), .A2(n28647), .ZN(n23272) );
  CLKXOR2HSV2 U13558 ( .A1(n23272), .A2(n23271), .Z(n23273) );
  XOR2HSV0 U13559 ( .A1(n21581), .A2(n21580), .Z(n21582) );
  NAND2HSV2 U13560 ( .A1(n21108), .A2(n21107), .ZN(n21110) );
  INHSV4 U13561 ( .I(n11976), .ZN(n16741) );
  NAND3HSV2 U13562 ( .A1(n16754), .A2(n23473), .A3(n16844), .ZN(n11976) );
  NOR2HSV2 U13563 ( .A1(n11977), .A2(n15496), .ZN(n15529) );
  CLKNHSV2 U13564 ( .I(n15495), .ZN(n11977) );
  INHSV4 U13565 ( .I(n14226), .ZN(n12153) );
  CLKBUFHSV12 U13566 ( .I(n28587), .Z(n11978) );
  NAND2HSV2 U13567 ( .A1(n12517), .A2(n24637), .ZN(n21625) );
  NAND2HSV2 U13568 ( .A1(n19274), .A2(n21326), .ZN(n19278) );
  CLKNAND2HSV4 U13569 ( .A1(n23458), .A2(n20456), .ZN(n20399) );
  CLKNAND2HSV4 U13570 ( .A1(n20396), .A2(n20397), .ZN(n23458) );
  NAND2HSV4 U13571 ( .A1(n21002), .A2(n21001), .ZN(n28965) );
  NAND2HSV4 U13572 ( .A1(n23444), .A2(n19964), .ZN(n19971) );
  XNOR4HSV4 U13573 ( .A1(\pe7/phq [3]), .A2(n19185), .A3(n11979), .A4(n19184), 
        .ZN(n19214) );
  NAND2HSV4 U13574 ( .A1(\pe7/ti_1 ), .A2(\pe7/got [14]), .ZN(n11979) );
  CLKNAND2HSV2 U13575 ( .A1(n13073), .A2(n13074), .ZN(n13075) );
  NOR2HSV2 U13576 ( .A1(n18383), .A2(n18469), .ZN(n18440) );
  INHSV4 U13577 ( .I(n17650), .ZN(n17648) );
  CLKNAND2HSV2 U13578 ( .A1(n16601), .A2(n16602), .ZN(n16603) );
  AOI21HSV4 U13579 ( .A1(n16598), .A2(n16597), .B(n16596), .ZN(n16601) );
  CLKNAND2HSV4 U13580 ( .A1(n12688), .A2(\pe7/pvq [1]), .ZN(n12689) );
  CLKNAND2HSV4 U13581 ( .A1(n15853), .A2(n28612), .ZN(n15668) );
  INHSV4 U13582 ( .I(n15668), .ZN(n15671) );
  NOR2HSV4 U13583 ( .A1(n20186), .A2(n11980), .ZN(n20193) );
  CLKNAND2HSV2 U13584 ( .A1(n11982), .A2(n11981), .ZN(n11980) );
  CLKNHSV2 U13585 ( .I(n20619), .ZN(n11981) );
  CLKNHSV2 U13586 ( .I(n20221), .ZN(n11982) );
  CLKNAND2HSV2 U13587 ( .A1(n19529), .A2(n24214), .ZN(n19531) );
  BUFHSV8 U13588 ( .I(\pe9/got [15]), .Z(n17940) );
  NAND2HSV2 U13589 ( .A1(n12311), .A2(n11983), .ZN(n20153) );
  CLKNAND2HSV2 U13590 ( .A1(n12310), .A2(n20150), .ZN(n11983) );
  NAND2HSV4 U13591 ( .A1(n15906), .A2(n15905), .ZN(n23327) );
  INHSV4 U13592 ( .I(n11994), .ZN(n14181) );
  NAND2HSV4 U13593 ( .A1(n15576), .A2(n15575), .ZN(n15577) );
  INHSV2 U13594 ( .I(n17729), .ZN(n17731) );
  XNOR2HSV4 U13595 ( .A1(n14314), .A2(n11984), .ZN(n14320) );
  XNOR2HSV4 U13596 ( .A1(n14312), .A2(n14313), .ZN(n11984) );
  CLKAND2HSV4 U13597 ( .A1(n28949), .A2(n18046), .Z(n18047) );
  XNOR2HSV4 U13598 ( .A1(n27043), .A2(n27042), .ZN(n27045) );
  CLKNAND2HSV2 U13599 ( .A1(n12955), .A2(\pe7/bq[15] ), .ZN(n19194) );
  NAND2HSV2 U13600 ( .A1(\pe7/bq[15] ), .A2(\pe7/aot [14]), .ZN(n19248) );
  INHSV4 U13601 ( .I(n17975), .ZN(n17976) );
  CLKNAND2HSV2 U13602 ( .A1(n11985), .A2(n13525), .ZN(n17975) );
  CLKNAND2HSV2 U13603 ( .A1(n11987), .A2(n11986), .ZN(n11985) );
  CLKNHSV2 U13604 ( .I(n13524), .ZN(n11986) );
  CLKNHSV2 U13605 ( .I(n13523), .ZN(n11987) );
  NAND2HSV2 U13606 ( .A1(\pe7/got [12]), .A2(n28587), .ZN(n13460) );
  NOR2HSV4 U13607 ( .A1(n12018), .A2(n22047), .ZN(n12017) );
  INAND2HSV2 U13608 ( .A1(n17901), .B1(n17900), .ZN(n17904) );
  INHSV2 U13609 ( .I(n14158), .ZN(n11988) );
  CLKNAND2HSV2 U13610 ( .A1(n11988), .A2(n27211), .ZN(n14187) );
  INHSV2 U13611 ( .I(n15473), .ZN(n11989) );
  NAND2HSV4 U13612 ( .A1(n11989), .A2(n12338), .ZN(n15479) );
  NAND2HSV2 U13613 ( .A1(\pe9/bq[13] ), .A2(\pe9/aot [16]), .ZN(n18302) );
  XNOR2HSV4 U13614 ( .A1(n11991), .A2(n11990), .ZN(n15669) );
  CLKNAND2HSV2 U13615 ( .A1(n28696), .A2(n25131), .ZN(n11990) );
  XNOR2HSV4 U13616 ( .A1(n11992), .A2(n15665), .ZN(n11991) );
  XNOR2HSV4 U13617 ( .A1(n15666), .A2(n15667), .ZN(n11992) );
  CLKXOR2HSV4 U13618 ( .A1(n21717), .A2(n21716), .Z(pov5[15]) );
  INHSV4 U13619 ( .I(n21992), .ZN(n27877) );
  AOI31HSV2 U13620 ( .A1(n19991), .A2(n19990), .A3(n22137), .B(n19989), .ZN(
        n20048) );
  CLKNAND2HSV2 U13621 ( .A1(n18844), .A2(n19831), .ZN(n19991) );
  OAI21HSV2 U13622 ( .A1(n19900), .A2(n13989), .B(n13959), .ZN(n19828) );
  CLKNAND2HSV4 U13623 ( .A1(n28920), .A2(n15245), .ZN(n15227) );
  INHSV2 U13624 ( .I(n22245), .ZN(n13324) );
  NAND2HSV0 U13625 ( .A1(n26229), .A2(\pe8/got [5]), .ZN(n22245) );
  NAND2HSV4 U13626 ( .A1(n16757), .A2(n26220), .ZN(n16754) );
  XNOR2HSV4 U13627 ( .A1(n15477), .A2(n11993), .ZN(n15532) );
  AOI21HSV4 U13628 ( .A1(n15567), .A2(n13503), .B(n15748), .ZN(n11993) );
  INHSV6 U13629 ( .I(n25914), .ZN(n26909) );
  AOI21HSV2 U13630 ( .A1(n24516), .A2(n21730), .B(n21727), .ZN(n16161) );
  INAND2HSV4 U13631 ( .A1(n16029), .B1(n21312), .ZN(n16175) );
  INHSV4 U13632 ( .I(n16175), .ZN(n16109) );
  CLKNAND2HSV2 U13633 ( .A1(n14119), .A2(n14396), .ZN(n11994) );
  NAND2HSV2 U13634 ( .A1(n13809), .A2(n11995), .ZN(\pe8/poht [9]) );
  CLKNAND2HSV2 U13635 ( .A1(n11997), .A2(n11996), .ZN(n11995) );
  CLKNHSV2 U13636 ( .I(n13807), .ZN(n11996) );
  CLKNHSV2 U13637 ( .I(n13808), .ZN(n11997) );
  CLKXOR2HSV4 U13638 ( .A1(n24742), .A2(n24741), .Z(n24743) );
  CLKXOR2HSV4 U13639 ( .A1(n24804), .A2(n24803), .Z(n24807) );
  XNOR2HSV4 U13640 ( .A1(n12615), .A2(n13592), .ZN(n12614) );
  CLKXOR2HSV4 U13641 ( .A1(n21806), .A2(n21805), .Z(n21807) );
  AOI21HSV4 U13642 ( .A1(n25045), .A2(n11998), .B(n20777), .ZN(n20780) );
  CLKNHSV2 U13643 ( .I(n11999), .ZN(n11998) );
  CLKNAND2HSV2 U13644 ( .A1(n20779), .A2(n20778), .ZN(n11999) );
  OAI21HSV2 U13645 ( .A1(n14390), .A2(n13539), .B(n13540), .ZN(n13541) );
  NAND2HSV2 U13646 ( .A1(n12000), .A2(\pe4/pvq [3]), .ZN(n15348) );
  INHSV2 U13647 ( .I(n15502), .ZN(n12000) );
  AOI21HSV4 U13648 ( .A1(n17982), .A2(n18481), .B(n12001), .ZN(n17984) );
  MUX2NHSV2 U13649 ( .I0(n18005), .I1(n17981), .S(n17980), .ZN(n12001) );
  IOA21HSV2 U13650 ( .A1(\pe9/ti_1 ), .A2(\pe9/got [14]), .B(\pe9/phq [3]), 
        .ZN(n17932) );
  XNOR2HSV2 U13651 ( .A1(n19040), .A2(n19039), .ZN(n19041) );
  BUFHSV6 U13652 ( .I(n16557), .Z(n28796) );
  CLKNAND2HSV2 U13653 ( .A1(n25377), .A2(n25334), .ZN(n19753) );
  NOR2HSV2 U13654 ( .A1(n17713), .A2(n17863), .ZN(n13638) );
  INHSV2 U13655 ( .I(n15808), .ZN(n15806) );
  XOR4HSV4 U13656 ( .A1(n26165), .A2(n12002), .A3(n16636), .A4(n16637), .Z(
        n16643) );
  AOI21HSV4 U13657 ( .A1(n16635), .A2(n16634), .B(n16633), .ZN(n12002) );
  CLKXOR2HSV4 U13658 ( .A1(n24609), .A2(n24608), .Z(n13224) );
  NAND2HSV2 U13659 ( .A1(n13225), .A2(n13224), .ZN(n13226) );
  CLKXOR2HSV4 U13660 ( .A1(n26758), .A2(n26757), .Z(n13402) );
  NAND2HSV2 U13661 ( .A1(n13403), .A2(n13402), .ZN(n13404) );
  INHSV4 U13662 ( .I(\pe11/got [13]), .ZN(n20201) );
  CLKNHSV6 U13663 ( .I(n20201), .ZN(n20707) );
  CLKNAND2HSV2 U13664 ( .A1(n17155), .A2(n17154), .ZN(n28622) );
  XNOR2HSV4 U13665 ( .A1(n12003), .A2(n24571), .ZN(n24572) );
  XNOR2HSV4 U13666 ( .A1(n24570), .A2(n24569), .ZN(n12003) );
  NAND2HSV4 U13667 ( .A1(\pe9/aot [16]), .A2(\pe9/bq[16] ), .ZN(n17884) );
  CLKXOR2HSV4 U13668 ( .A1(n25942), .A2(n25941), .Z(n25944) );
  AOI21HSV4 U13669 ( .A1(n19418), .A2(n28466), .B(n25499), .ZN(n19419) );
  XNOR2HSV4 U13670 ( .A1(n26412), .A2(n12004), .ZN(n12984) );
  CLKNHSV2 U13671 ( .I(n12005), .ZN(n12004) );
  CLKNAND2HSV2 U13672 ( .A1(n28652), .A2(n28930), .ZN(n12005) );
  INHSV4 U13673 ( .I(n16601), .ZN(n16599) );
  NAND2HSV4 U13674 ( .A1(n16600), .A2(n16599), .ZN(n16604) );
  CLKNAND2HSV4 U13675 ( .A1(\pe8/bq[10] ), .A2(\pe8/aot [16]), .ZN(n16468) );
  NAND2HSV2 U13676 ( .A1(n24377), .A2(n28645), .ZN(n23274) );
  NAND2HSV4 U13677 ( .A1(n12153), .A2(n12006), .ZN(n14227) );
  INHSV4 U13678 ( .I(n14225), .ZN(n12006) );
  DELHS1 U13679 ( .I(n25529), .Z(n12007) );
  CLKXOR2HSV4 U13680 ( .A1(n24876), .A2(n24875), .Z(n24877) );
  NAND2HSV2 U13681 ( .A1(n28603), .A2(n27196), .ZN(n25064) );
  XNOR2HSV4 U13682 ( .A1(n12008), .A2(n17764), .ZN(n17765) );
  XNOR2HSV4 U13683 ( .A1(n17762), .A2(n17763), .ZN(n12008) );
  NAND2HSV4 U13684 ( .A1(n25055), .A2(n25053), .ZN(n24902) );
  NAND2HSV2 U13685 ( .A1(\pe8/aot [16]), .A2(\pe8/bq[12] ), .ZN(n16407) );
  XNOR2HSV4 U13686 ( .A1(n25412), .A2(n25411), .ZN(\pe7/poht [7]) );
  NAND3HSV4 U13687 ( .A1(n15457), .A2(n15487), .A3(n15456), .ZN(n15500) );
  OAI21HSV2 U13688 ( .A1(n27678), .A2(n27677), .B(n13476), .ZN(n13477) );
  OAI31HSV2 U13689 ( .A1(n27678), .A2(n13476), .A3(n27677), .B(n13477), .ZN(
        n13478) );
  AOI21HSV2 U13690 ( .A1(n20187), .A2(n20188), .B(n20620), .ZN(n20191) );
  NOR2HSV4 U13691 ( .A1(n12010), .A2(n12009), .ZN(n20187) );
  CLKNHSV2 U13692 ( .I(n20171), .ZN(n12009) );
  CLKNHSV2 U13693 ( .I(n20181), .ZN(n12010) );
  CLKNAND2HSV2 U13694 ( .A1(n27106), .A2(n24637), .ZN(n21460) );
  NAND2HSV4 U13695 ( .A1(n14611), .A2(n14612), .ZN(n14629) );
  CLKNAND2HSV4 U13696 ( .A1(n14271), .A2(n14270), .ZN(n14391) );
  NOR2HSV4 U13697 ( .A1(n21732), .A2(n21720), .ZN(n16170) );
  NAND2HSV4 U13698 ( .A1(n12127), .A2(n12126), .ZN(n21239) );
  NOR2HSV4 U13699 ( .A1(n25502), .A2(n20689), .ZN(n20176) );
  DELHS1 U13700 ( .I(\pe11/aot [13]), .Z(n12011) );
  CLKNHSV2 U13701 ( .I(n21645), .ZN(n12013) );
  NAND2HSV2 U13702 ( .A1(n27106), .A2(n24635), .ZN(n24698) );
  XNOR2HSV4 U13703 ( .A1(n25343), .A2(n12014), .ZN(po7) );
  CLKNHSV2 U13704 ( .I(n25342), .ZN(n12016) );
  CLKXOR2HSV2 U13705 ( .A1(n16404), .A2(n16403), .Z(n16405) );
  CLKNAND2HSV2 U13706 ( .A1(n14031), .A2(\pe5/bq[11] ), .ZN(n14594) );
  CLKXOR2HSV2 U13707 ( .A1(n14595), .A2(n14594), .Z(n14596) );
  NOR2HSV4 U13708 ( .A1(n16327), .A2(n16353), .ZN(n16328) );
  XOR2HSV4 U13709 ( .A1(n12597), .A2(n12595), .Z(n21892) );
  CLKNAND2HSV4 U13710 ( .A1(n21815), .A2(n21144), .ZN(n12597) );
  XNOR2HSV4 U13711 ( .A1(n23371), .A2(n23370), .ZN(n23377) );
  XNOR2HSV2 U13712 ( .A1(n23377), .A2(n23376), .ZN(n23378) );
  NAND2HSV4 U13713 ( .A1(n28707), .A2(n26240), .ZN(n15235) );
  INHSV2 U13714 ( .I(n20151), .ZN(n20329) );
  CLKNAND2HSV4 U13715 ( .A1(n14207), .A2(n14206), .ZN(n14211) );
  CLKNAND2HSV4 U13716 ( .A1(n14211), .A2(n14210), .ZN(n14278) );
  CLKNAND2HSV4 U13717 ( .A1(n12065), .A2(n12064), .ZN(n14273) );
  NAND2HSV4 U13718 ( .A1(n16893), .A2(n22508), .ZN(n16882) );
  NAND2HSV4 U13719 ( .A1(n21145), .A2(n21144), .ZN(n21157) );
  NAND2HSV4 U13720 ( .A1(\pe2/got [14]), .A2(\pe2/ti_1 ), .ZN(n17657) );
  MUX2NHSV4 U13721 ( .I0(n12271), .I1(n13816), .S(n12017), .ZN(n13962) );
  NAND2HSV4 U13722 ( .A1(n12020), .A2(n12019), .ZN(n12018) );
  INHSV2 U13723 ( .I(n22054), .ZN(n12019) );
  INHSV4 U13724 ( .I(n26825), .ZN(n12020) );
  CLKNAND2HSV4 U13725 ( .A1(n17910), .A2(n17909), .ZN(n17914) );
  NAND2HSV4 U13726 ( .A1(n17831), .A2(\pe2/pvq [4]), .ZN(n17721) );
  CLKNAND2HSV2 U13727 ( .A1(n15190), .A2(n15189), .ZN(n15193) );
  NAND2HSV4 U13728 ( .A1(n15193), .A2(n15192), .ZN(n15199) );
  MUX2NHSV4 U13729 ( .I0(n12303), .I1(n13596), .S(n12021), .ZN(n28997) );
  BUFHSV8 U13730 ( .I(\pe4/bq[15] ), .Z(n26958) );
  NAND2HSV2 U13731 ( .A1(n15201), .A2(n15200), .ZN(n15204) );
  CLKNAND2HSV2 U13732 ( .A1(n15204), .A2(n15203), .ZN(n15206) );
  INHSV4 U13733 ( .I(n27322), .ZN(n21842) );
  NAND2HSV4 U13734 ( .A1(\pe2/aot [16]), .A2(\pe2/bq[14] ), .ZN(n17659) );
  XNOR2HSV4 U13735 ( .A1(n20753), .A2(n20752), .ZN(n20755) );
  CLKNAND2HSV4 U13736 ( .A1(n15282), .A2(n12022), .ZN(n15975) );
  CLKNAND2HSV4 U13737 ( .A1(n15279), .A2(n15278), .ZN(n12022) );
  CLKAND2HSV8 U13738 ( .A1(\pe10/ctrq ), .A2(\pe10/pvq [3]), .Z(n16634) );
  CLKXOR2HSV2 U13739 ( .A1(n26027), .A2(n26026), .Z(n26028) );
  XNOR2HSV4 U13740 ( .A1(n12537), .A2(n12540), .ZN(n12536) );
  XOR3HSV2 U13741 ( .A1(n18435), .A2(n12641), .A3(n18434), .Z(n18436) );
  XNOR2HSV4 U13742 ( .A1(n16783), .A2(n16782), .ZN(n16784) );
  NAND2HSV2 U13743 ( .A1(n26231), .A2(n26230), .ZN(n26235) );
  BUFHSV8 U13744 ( .I(\pe11/got [15]), .Z(n20171) );
  INHSV2 U13745 ( .I(n12024), .ZN(n13978) );
  NAND2HSV2 U13746 ( .A1(n15284), .A2(n15285), .ZN(n12024) );
  BUFHSV6 U13747 ( .I(n22078), .Z(n28467) );
  XOR2HSV4 U13748 ( .A1(n22877), .A2(n22876), .Z(n22878) );
  CLKNAND2HSV2 U13749 ( .A1(n13195), .A2(n13196), .ZN(n13197) );
  CLKNAND2HSV2 U13750 ( .A1(n13194), .A2(n12025), .ZN(n13195) );
  CLKNAND2HSV2 U13751 ( .A1(n12027), .A2(n12026), .ZN(n12025) );
  CLKNHSV2 U13752 ( .I(n13193), .ZN(n12026) );
  NOR2HSV4 U13753 ( .A1(n17068), .A2(n26091), .ZN(n12027) );
  INHSV8 U13754 ( .I(n14763), .ZN(n14526) );
  NAND2HSV2 U13755 ( .A1(n14484), .A2(\pe5/got [15]), .ZN(n14485) );
  CLKNAND2HSV4 U13756 ( .A1(n14477), .A2(n12028), .ZN(n14491) );
  INHSV4 U13757 ( .I(n12029), .ZN(n12028) );
  CLKNAND2HSV4 U13758 ( .A1(n14476), .A2(n14475), .ZN(n12029) );
  CLKXOR2HSV4 U13759 ( .A1(n24744), .A2(n24743), .Z(n24747) );
  INHSV2 U13760 ( .I(n16935), .ZN(n12030) );
  INHSV2 U13761 ( .I(n12032), .ZN(n12031) );
  OAI21HSV2 U13762 ( .A1(n16942), .A2(n17112), .B(n16740), .ZN(n12032) );
  NAND2HSV2 U13763 ( .A1(n23375), .A2(\pe3/got [11]), .ZN(n23376) );
  CLKXOR2HSV4 U13764 ( .A1(n14901), .A2(n14900), .Z(n14904) );
  NAND2HSV2 U13765 ( .A1(n28936), .A2(\pe11/got [2]), .ZN(n12452) );
  INHSV4 U13766 ( .I(n18210), .ZN(n12363) );
  INHSV4 U13767 ( .I(n16734), .ZN(n16757) );
  CLKNAND2HSV4 U13768 ( .A1(n19815), .A2(n23245), .ZN(n18636) );
  NAND2HSV4 U13769 ( .A1(n18632), .A2(n18633), .ZN(n19815) );
  CLKNAND2HSV2 U13770 ( .A1(n13069), .A2(n13068), .ZN(n13070) );
  CLKNAND2HSV2 U13771 ( .A1(n13164), .A2(n13163), .ZN(n13165) );
  XNOR2HSV4 U13772 ( .A1(n16253), .A2(n12033), .ZN(n16258) );
  XNOR2HSV4 U13773 ( .A1(n12034), .A2(n16250), .ZN(n12033) );
  XNOR2HSV4 U13774 ( .A1(n16251), .A2(n16252), .ZN(n12034) );
  OAI21HSV4 U13775 ( .A1(n12244), .A2(n12190), .B(n12035), .ZN(n12191) );
  CLKNAND2HSV2 U13776 ( .A1(n12188), .A2(n12190), .ZN(n12035) );
  NAND2HSV4 U13777 ( .A1(n16499), .A2(n16498), .ZN(n16503) );
  CLKNAND2HSV4 U13778 ( .A1(n16503), .A2(n16502), .ZN(n16506) );
  NAND2HSV0 U13779 ( .A1(n13336), .A2(n12036), .ZN(\pe3/poht [4]) );
  INHSV2 U13780 ( .I(n13335), .ZN(n12037) );
  INAND2HSV2 U13781 ( .A1(n12038), .B1(n26679), .ZN(n13335) );
  INHSV2 U13782 ( .I(n15245), .ZN(n12038) );
  CLKNHSV2 U13783 ( .I(n13334), .ZN(n12039) );
  NAND2HSV4 U13784 ( .A1(n21743), .A2(n21742), .ZN(n25952) );
  INHSV2 U13785 ( .I(n19266), .ZN(n19211) );
  CLKNAND2HSV4 U13786 ( .A1(n12720), .A2(n12719), .ZN(n21321) );
  NAND2HSV4 U13787 ( .A1(n23328), .A2(\pe3/got [11]), .ZN(n16153) );
  CLKNAND2HSV2 U13788 ( .A1(n19058), .A2(n19070), .ZN(n19157) );
  CLKNHSV12 U13789 ( .I(n15963), .ZN(n28931) );
  NAND2HSV4 U13790 ( .A1(n12040), .A2(n20156), .ZN(n20161) );
  CLKNAND2HSV2 U13791 ( .A1(n20154), .A2(n20155), .ZN(n12040) );
  BUFHSV8 U13792 ( .I(n19422), .Z(n19579) );
  NAND2HSV0 U13793 ( .A1(\pe7/got [12]), .A2(n19579), .ZN(n19608) );
  OAI21HSV4 U13794 ( .A1(n19137), .A2(n25519), .B(n19136), .ZN(n19140) );
  NAND2HSV2 U13795 ( .A1(n14398), .A2(\pe6/got [14]), .ZN(n14394) );
  CLKNAND2HSV4 U13796 ( .A1(n14894), .A2(n14852), .ZN(n14604) );
  INHSV4 U13797 ( .I(n14911), .ZN(n14762) );
  XNOR2HSV4 U13798 ( .A1(n15909), .A2(n15908), .ZN(n16018) );
  INHSV2 U13799 ( .I(n21765), .ZN(n26084) );
  BUFHSV8 U13800 ( .I(n16848), .Z(n28679) );
  INHSV2 U13801 ( .I(n12404), .ZN(n22310) );
  INHSV6 U13802 ( .I(n23717), .ZN(n28394) );
  XOR3HSV2 U13803 ( .A1(n12041), .A2(n22040), .A3(n22041), .Z(n22045) );
  CLKNHSV2 U13804 ( .I(n22039), .ZN(n12041) );
  CLKNHSV6 U13805 ( .I(n14761), .ZN(n14911) );
  XNOR2HSV4 U13806 ( .A1(n20762), .A2(n12042), .ZN(n20766) );
  CLKNAND2HSV2 U13807 ( .A1(n12434), .A2(n25504), .ZN(n12042) );
  INHSV4 U13808 ( .I(n13337), .ZN(n12697) );
  CLKNHSV0 U13809 ( .I(n19708), .ZN(n28656) );
  INHSV2 U13810 ( .I(n19614), .ZN(n19514) );
  OAI21HSV4 U13811 ( .A1(n19513), .A2(n19514), .B(n13990), .ZN(n12119) );
  XNOR2HSV4 U13812 ( .A1(n27815), .A2(n27814), .ZN(n27817) );
  XNOR2HSV2 U13813 ( .A1(n27817), .A2(n27816), .ZN(n27818) );
  NAND2HSV4 U13814 ( .A1(n25657), .A2(n12505), .ZN(n14759) );
  NAND3HSV4 U13815 ( .A1(n19132), .A2(n19131), .A3(n18921), .ZN(n12603) );
  INHSV2 U13816 ( .I(n16444), .ZN(n25651) );
  NAND2HSV4 U13817 ( .A1(n16425), .A2(n16445), .ZN(n16444) );
  XNOR2HSV4 U13818 ( .A1(n20200), .A2(n12043), .ZN(n20205) );
  XOR2HSV2 U13819 ( .A1(n20199), .A2(n20198), .Z(n12043) );
  CLKNAND2HSV2 U13820 ( .A1(n12877), .A2(n12044), .ZN(n12878) );
  CLKNAND2HSV2 U13821 ( .A1(n12046), .A2(n12045), .ZN(n12044) );
  CLKNHSV2 U13822 ( .I(n12876), .ZN(n12045) );
  CLKNAND2HSV2 U13823 ( .A1(n19507), .A2(n24181), .ZN(n12876) );
  CLKNHSV2 U13824 ( .I(n19508), .ZN(n12046) );
  INHSV2 U13825 ( .I(n12047), .ZN(n21166) );
  CLKNAND2HSV4 U13826 ( .A1(n13337), .A2(n12432), .ZN(n13338) );
  INHSV4 U13827 ( .I(n26625), .ZN(n28432) );
  XOR3HSV2 U13828 ( .A1(n20468), .A2(n12049), .A3(n12048), .Z(n20490) );
  CLKNHSV2 U13829 ( .I(n20488), .ZN(n12048) );
  CLKNHSV2 U13830 ( .I(n20469), .ZN(n12049) );
  CLKNAND2HSV2 U13831 ( .A1(n19579), .A2(n25334), .ZN(n19414) );
  XNOR2HSV4 U13832 ( .A1(n16827), .A2(n16826), .ZN(n16828) );
  NAND2HSV2 U13833 ( .A1(\pe4/bq[15] ), .A2(\pe4/aot [14]), .ZN(n13787) );
  INHSV6 U13834 ( .I(n14397), .ZN(n14398) );
  NAND3HSV2 U13835 ( .A1(n12050), .A2(n19704), .A3(n19703), .ZN(n12611) );
  CLKNHSV2 U13836 ( .I(n25674), .ZN(n12050) );
  NOR2HSV4 U13837 ( .A1(n19688), .A2(n12613), .ZN(n25674) );
  NAND2HSV4 U13838 ( .A1(n12051), .A2(n12077), .ZN(n19671) );
  INHSV4 U13839 ( .I(n19574), .ZN(n12051) );
  INAND2HSV4 U13840 ( .A1(n19617), .B1(n13399), .ZN(n25346) );
  CLKNAND2HSV2 U13841 ( .A1(n25347), .A2(n25346), .ZN(n12709) );
  XNOR2HSV4 U13842 ( .A1(n14740), .A2(n14741), .ZN(n19124) );
  NAND2HSV4 U13843 ( .A1(n14748), .A2(n14747), .ZN(n14750) );
  XNOR2HSV4 U13844 ( .A1(n12052), .A2(n16014), .ZN(n16020) );
  XNOR2HSV4 U13845 ( .A1(n12053), .A2(n16012), .ZN(n12052) );
  CLKNHSV2 U13846 ( .I(n16013), .ZN(n12053) );
  INHSV4 U13847 ( .I(n14484), .ZN(n14495) );
  CLKNHSV6 U13848 ( .I(n27192), .ZN(n12247) );
  CLKNHSV6 U13849 ( .I(n27494), .ZN(n27736) );
  NAND2HSV2 U13850 ( .A1(n27727), .A2(n27543), .ZN(n27395) );
  INHSV4 U13851 ( .I(n28703), .ZN(n25340) );
  NOR2HSV4 U13852 ( .A1(n25340), .A2(n19532), .ZN(n23215) );
  INHSV4 U13853 ( .I(n14333), .ZN(n12768) );
  XNOR2HSV4 U13854 ( .A1(n12054), .A2(n12149), .ZN(n12148) );
  XNOR2HSV4 U13855 ( .A1(n12152), .A2(n12874), .ZN(n12054) );
  NAND2HSV4 U13856 ( .A1(n14553), .A2(n14473), .ZN(n14476) );
  CLKNAND2HSV2 U13857 ( .A1(n15970), .A2(n15969), .ZN(n15971) );
  NAND2HSV2 U13858 ( .A1(n23409), .A2(n23408), .ZN(n23410) );
  NAND3HSV4 U13859 ( .A1(n14500), .A2(n14499), .A3(n14555), .ZN(n22094) );
  INHSV2 U13860 ( .I(n14673), .ZN(n13118) );
  INHSV2 U13861 ( .I(n25658), .ZN(n14613) );
  AOI22HSV4 U13862 ( .A1(n14616), .A2(\pe5/ti_7t [7]), .B1(n25658), .B2(n14615), .ZN(n12496) );
  AND2HSV4 U13863 ( .A1(n14611), .A2(n14612), .Z(n25658) );
  CLKNAND2HSV2 U13864 ( .A1(n18440), .A2(n18441), .ZN(n18442) );
  NAND2HSV2 U13865 ( .A1(n21223), .A2(n21702), .ZN(n21224) );
  INHSV4 U13866 ( .I(n21224), .ZN(n21227) );
  INHSV4 U13867 ( .I(n14231), .ZN(n12459) );
  CLKNAND2HSV2 U13868 ( .A1(n17926), .A2(n12055), .ZN(n17929) );
  CLKNAND2HSV2 U13869 ( .A1(\pe9/bq[15] ), .A2(\pe9/aot [15]), .ZN(n12055) );
  NOR2HSV4 U13870 ( .A1(n19129), .A2(n14745), .ZN(n18853) );
  AOI21HSV2 U13871 ( .A1(n22085), .A2(n25362), .B(n12594), .ZN(n12593) );
  NAND2HSV2 U13872 ( .A1(n12593), .A2(n21711), .ZN(n21891) );
  INHSV4 U13873 ( .I(n20979), .ZN(n24636) );
  NAND2HSV3 U13874 ( .A1(n17974), .A2(n17975), .ZN(n17979) );
  NAND2HSV4 U13875 ( .A1(n15026), .A2(n15025), .ZN(n15030) );
  NAND2HSV4 U13876 ( .A1(n15030), .A2(n15029), .ZN(n15034) );
  CLKNHSV6 U13877 ( .I(n27223), .ZN(n17479) );
  NAND2HSV4 U13878 ( .A1(n16495), .A2(n16494), .ZN(n16583) );
  INHSV4 U13879 ( .I(\pe3/ti_1 ), .ZN(n15007) );
  XNOR2HSV2 U13880 ( .A1(n19461), .A2(n19460), .ZN(n19467) );
  INHSV4 U13881 ( .I(n17064), .ZN(n17061) );
  NAND2HSV4 U13882 ( .A1(n17061), .A2(n17062), .ZN(n12059) );
  CLKNAND2HSV2 U13883 ( .A1(n20068), .A2(n20067), .ZN(n20069) );
  NAND2HSV2 U13884 ( .A1(n13357), .A2(n13356), .ZN(n13358) );
  NAND3HSV4 U13885 ( .A1(n12056), .A2(n18094), .A3(n23465), .ZN(n18095) );
  OAI21HSV4 U13886 ( .A1(n14638), .A2(n14924), .B(n14633), .ZN(n14634) );
  AOI21HSV4 U13887 ( .A1(n14635), .A2(n14636), .B(n14634), .ZN(n14641) );
  INHSV4 U13888 ( .I(n18280), .ZN(n12327) );
  NAND2HSV4 U13889 ( .A1(n12057), .A2(n19261), .ZN(n23844) );
  CLKNAND2HSV4 U13890 ( .A1(n19260), .A2(n19259), .ZN(n12057) );
  NAND2HSV4 U13891 ( .A1(\pe8/got [12]), .A2(n16511), .ZN(n16404) );
  NAND2HSV2 U13892 ( .A1(n25784), .A2(\pe6/got [4]), .ZN(n23714) );
  XNOR2HSV4 U13893 ( .A1(n23214), .A2(n23213), .ZN(n23216) );
  CLKNAND2HSV4 U13894 ( .A1(n12059), .A2(n12058), .ZN(n17131) );
  NAND3HSV4 U13895 ( .A1(n17064), .A2(n20070), .A3(n17063), .ZN(n12058) );
  CLKNAND2HSV4 U13896 ( .A1(n14571), .A2(n14570), .ZN(n23467) );
  NAND2HSV4 U13897 ( .A1(n23467), .A2(n12498), .ZN(n12497) );
  NAND3HSV3 U13898 ( .A1(n18143), .A2(n18144), .A3(n18028), .ZN(n18107) );
  NAND3HSV3 U13899 ( .A1(n25517), .A2(n19150), .A3(n19149), .ZN(n19153) );
  CLKNAND2HSV4 U13900 ( .A1(n12060), .A2(n16620), .ZN(n23484) );
  NAND2HSV4 U13901 ( .A1(n16619), .A2(n16618), .ZN(n12060) );
  CLKNAND2HSV4 U13902 ( .A1(n12111), .A2(n19146), .ZN(n25518) );
  CLKNAND2HSV2 U13903 ( .A1(n23467), .A2(n14628), .ZN(n25657) );
  INHSV2 U13904 ( .I(n26131), .ZN(n26200) );
  CLKNAND2HSV4 U13905 ( .A1(n27212), .A2(n14189), .ZN(n14190) );
  INHSV6 U13906 ( .I(n14190), .ZN(n14289) );
  NOR2HSV8 U13907 ( .A1(n14447), .A2(n14446), .ZN(n14445) );
  INHSV6 U13908 ( .I(n14448), .ZN(n27050) );
  CLKNAND2HSV4 U13909 ( .A1(n27050), .A2(n14445), .ZN(n14450) );
  NAND2HSV2 U13910 ( .A1(n27727), .A2(n27544), .ZN(n27545) );
  NAND3HSV3 U13911 ( .A1(n18185), .A2(n18184), .A3(n18183), .ZN(n18186) );
  NAND2HSV2 U13912 ( .A1(n12062), .A2(n12061), .ZN(n16294) );
  NAND2HSV2 U13913 ( .A1(n16464), .A2(\pe8/aot [16]), .ZN(n12061) );
  INHSV2 U13914 ( .I(n16292), .ZN(n12062) );
  XNOR2HSV2 U13915 ( .A1(n18437), .A2(n18436), .ZN(n18438) );
  XNOR2HSV4 U13916 ( .A1(n16297), .A2(n16298), .ZN(n16301) );
  CLKNAND2HSV4 U13917 ( .A1(n12560), .A2(n12559), .ZN(n12558) );
  NAND2HSV4 U13918 ( .A1(n14902), .A2(n24635), .ZN(n14810) );
  CLKXOR2HSV4 U13919 ( .A1(n13076), .A2(n13077), .Z(n18313) );
  CLKXOR2HSV4 U13920 ( .A1(n17875), .A2(n17874), .Z(n17881) );
  XOR2HSV4 U13921 ( .A1(n17881), .A2(n17880), .Z(n17920) );
  CLKNAND2HSV4 U13922 ( .A1(n12723), .A2(n12722), .ZN(n18541) );
  CLKNAND2HSV4 U13923 ( .A1(n14809), .A2(n14808), .ZN(n12635) );
  CLKNAND2HSV4 U13924 ( .A1(n12635), .A2(n12634), .ZN(n14902) );
  CLKAND2HSV4 U13925 ( .A1(n14054), .A2(n16030), .Z(n16033) );
  CLKNAND2HSV2 U13926 ( .A1(n14552), .A2(n14852), .ZN(n14545) );
  XNOR2HSV4 U13927 ( .A1(n21687), .A2(n21686), .ZN(n21688) );
  NAND2HSV4 U13928 ( .A1(n24378), .A2(\pe5/got [13]), .ZN(n14906) );
  NAND2HSV4 U13929 ( .A1(n14582), .A2(n14581), .ZN(n14894) );
  XNOR2HSV4 U13930 ( .A1(n12063), .A2(n15141), .ZN(n15143) );
  XNOR2HSV4 U13931 ( .A1(n15138), .A2(n15139), .ZN(n12063) );
  INAND2HSV4 U13932 ( .A1(n13992), .B1(n28664), .ZN(n14803) );
  INHSV4 U13933 ( .I(n14265), .ZN(n12064) );
  NAND2HSV4 U13934 ( .A1(n12191), .A2(n12192), .ZN(n12189) );
  CLKNAND2HSV2 U13935 ( .A1(n12066), .A2(n14294), .ZN(n14298) );
  CLKNAND2HSV2 U13936 ( .A1(n12068), .A2(n12067), .ZN(n12066) );
  CLKNHSV2 U13937 ( .I(n14296), .ZN(n12067) );
  CLKNHSV2 U13938 ( .I(n14295), .ZN(n12068) );
  NAND3HSV4 U13939 ( .A1(n12611), .A2(n12608), .A3(n12818), .ZN(n12069) );
  CLKNHSV2 U13940 ( .I(n12069), .ZN(n23871) );
  CLKNAND2HSV2 U13941 ( .A1(n12069), .A2(n24271), .ZN(n19755) );
  AOI31HSV2 U13942 ( .A1(n18218), .A2(n18217), .A3(n18216), .B(n12462), .ZN(
        n12070) );
  INHSV2 U13943 ( .I(n18264), .ZN(n12075) );
  NAND2HSV2 U13944 ( .A1(n12071), .A2(n12070), .ZN(n18264) );
  CLKNAND2HSV3 U13945 ( .A1(n25662), .A2(n18221), .ZN(n12071) );
  XNOR2HSV4 U13946 ( .A1(n12073), .A2(n12072), .ZN(n18262) );
  OAI21HSV4 U13947 ( .A1(n29000), .A2(n18194), .B(n18226), .ZN(n12072) );
  XNOR2HSV4 U13948 ( .A1(n18224), .A2(n18223), .ZN(n29000) );
  CLKNAND2HSV2 U13949 ( .A1(n19794), .A2(n28137), .ZN(n12074) );
  CLKNHSV4 U13950 ( .I(n12076), .ZN(n16026) );
  XNOR2HSV4 U13951 ( .A1(n16020), .A2(n16019), .ZN(n12076) );
  CLKNAND2HSV2 U13952 ( .A1(n12076), .A2(n16024), .ZN(n16028) );
  CLKNHSV2 U13953 ( .I(n19574), .ZN(n12081) );
  OAI22HSV4 U13954 ( .A1(n12081), .A2(n12080), .B1(n12079), .B2(n12078), .ZN(
        n19618) );
  CLKNAND2HSV2 U13955 ( .A1(n27131), .A2(n12082), .ZN(n12078) );
  CLKNHSV2 U13956 ( .I(n19575), .ZN(n12079) );
  CLKNHSV2 U13957 ( .I(n12082), .ZN(n12080) );
  CLKNHSV2 U13958 ( .I(n12121), .ZN(n12082) );
  XOR2HSV2 U13959 ( .A1(n13715), .A2(n12083), .Z(n13716) );
  XNOR2HSV4 U13960 ( .A1(n12086), .A2(n12084), .ZN(n12083) );
  XNOR2HSV4 U13961 ( .A1(n25970), .A2(n12085), .ZN(n12084) );
  CLKNHSV2 U13962 ( .I(n25971), .ZN(n12085) );
  CLKNAND2HSV2 U13963 ( .A1(n23041), .A2(n26083), .ZN(n12086) );
  CLKNHSV2 U13964 ( .I(n15244), .ZN(n15283) );
  XNOR2HSV1 U13965 ( .A1(n12087), .A2(n13450), .ZN(n15276) );
  CLKXOR2HSV4 U13966 ( .A1(n12088), .A2(n13449), .Z(n12087) );
  NOR2HSV3 U13967 ( .A1(n15244), .A2(n12089), .ZN(n12088) );
  INHSV2 U13968 ( .I(n15245), .ZN(n12089) );
  BUFHSV8 U13969 ( .I(\pe5/ti_1 ), .Z(n12090) );
  CLKNAND2HSV2 U13970 ( .A1(\pe5/ti_1 ), .A2(\pe5/got [15]), .ZN(n14451) );
  CLKNAND2HSV2 U13971 ( .A1(n12090), .A2(\pe5/got [3]), .ZN(n20939) );
  CLKNAND2HSV2 U13972 ( .A1(\pe5/got [11]), .A2(n12090), .ZN(n14536) );
  CLKNAND2HSV2 U13973 ( .A1(\pe5/got [12]), .A2(n12090), .ZN(n14436) );
  CLKNAND2HSV2 U13974 ( .A1(\pe5/got [9]), .A2(n12090), .ZN(n14645) );
  CLKNAND2HSV2 U13975 ( .A1(\pe5/got [5]), .A2(n25626), .ZN(n14942) );
  CLKNAND2HSV2 U13976 ( .A1(n28640), .A2(n12090), .ZN(n21477) );
  CLKNAND2HSV2 U13977 ( .A1(n14503), .A2(n12090), .ZN(n12152) );
  CLKNAND2HSV0 U13978 ( .A1(n12093), .A2(n12091), .ZN(n19360) );
  INHSV2 U13979 ( .I(n12092), .ZN(n12091) );
  CLKNAND2HSV3 U13980 ( .A1(n19366), .A2(n24271), .ZN(n12092) );
  NAND3HSV3 U13981 ( .A1(n12093), .A2(n23844), .A3(n19366), .ZN(n19370) );
  NAND2HSV2 U13982 ( .A1(n19284), .A2(n19281), .ZN(n12093) );
  XNOR2HSV4 U13983 ( .A1(n12095), .A2(n12094), .ZN(n15174) );
  NOR2HSV4 U13984 ( .A1(n15160), .A2(n23383), .ZN(n12094) );
  AOI21HSV4 U13985 ( .A1(n15145), .A2(n25635), .B(n15144), .ZN(n15160) );
  CLKNAND2HSV1 U13986 ( .A1(n13793), .A2(n15097), .ZN(n25635) );
  NOR2HSV4 U13987 ( .A1(n25636), .A2(n15238), .ZN(n15145) );
  XOR2HSV2 U13988 ( .A1(n15173), .A2(n12096), .Z(n12095) );
  XNOR2HSV4 U13989 ( .A1(n12098), .A2(n12097), .ZN(n12096) );
  CLKNAND2HSV2 U13990 ( .A1(n23480), .A2(n15245), .ZN(n12097) );
  XNOR2HSV4 U13991 ( .A1(n12105), .A2(n12099), .ZN(n13290) );
  AOI21HSV4 U13992 ( .A1(n12104), .A2(n12103), .B(n12100), .ZN(n12099) );
  CLKNHSV2 U13993 ( .I(n12101), .ZN(n12100) );
  AOI21HSV4 U13994 ( .A1(n16669), .A2(n12102), .B(n20065), .ZN(n12101) );
  CLKNHSV2 U13995 ( .I(\pe10/ti_7t [6]), .ZN(n12102) );
  CLKNHSV2 U13996 ( .I(n16669), .ZN(n12103) );
  CLKNHSV2 U13997 ( .I(n28997), .ZN(n12104) );
  XNOR2HSV4 U13998 ( .A1(n12106), .A2(n16881), .ZN(n12105) );
  CLKNAND2HSV2 U13999 ( .A1(n12108), .A2(n12107), .ZN(n12106) );
  CLKNAND2HSV2 U14000 ( .A1(n16879), .A2(n28794), .ZN(n12107) );
  CLKNAND2HSV2 U14001 ( .A1(n16878), .A2(n16877), .ZN(n12108) );
  CLKNAND2HSV3 U14002 ( .A1(n19139), .A2(n12111), .ZN(n12110) );
  CLKNAND2HSV4 U14003 ( .A1(n19067), .A2(n22993), .ZN(n12111) );
  CLKNAND2HSV2 U14004 ( .A1(n12111), .A2(n19135), .ZN(n19137) );
  NAND2HSV2 U14005 ( .A1(n12112), .A2(n20977), .ZN(n14602) );
  INHSV2 U14006 ( .I(n14583), .ZN(n12112) );
  CLKBUFHSV2 U14007 ( .I(n14583), .Z(n12113) );
  INAND2HSV4 U14008 ( .A1(n14583), .B1(\pe5/got [10]), .ZN(n14664) );
  INAND2HSV4 U14009 ( .A1(n12113), .B1(n14069), .ZN(n14788) );
  INAND2HSV4 U14010 ( .A1(n12113), .B1(n28645), .ZN(n14866) );
  INAND2HSV4 U14011 ( .A1(n12113), .B1(n28647), .ZN(n14932) );
  INAND2HSV4 U14012 ( .A1(n12113), .B1(n14072), .ZN(n20873) );
  INAND2HSV4 U14013 ( .A1(n12113), .B1(\pe5/got [3]), .ZN(n21389) );
  CLKNHSV4 U14014 ( .I(n19949), .ZN(n28690) );
  CLKNAND2HSV2 U14015 ( .A1(n28690), .A2(n19943), .ZN(n12196) );
  CLKNAND2HSV0 U14016 ( .A1(n19578), .A2(n19577), .ZN(n12115) );
  XNOR2HSV4 U14017 ( .A1(n12116), .A2(n12117), .ZN(n25347) );
  NOR2HSV4 U14018 ( .A1(n12119), .A2(n12118), .ZN(n12116) );
  NOR2HSV4 U14019 ( .A1(n12508), .A2(n12120), .ZN(n12118) );
  OAI21HSV4 U14020 ( .A1(n25347), .A2(n19695), .B(n19694), .ZN(n12710) );
  CLKNHSV2 U14021 ( .I(n19526), .ZN(n12120) );
  CLKNHSV2 U14022 ( .I(n19618), .ZN(n25672) );
  CLKNAND2HSV2 U14023 ( .A1(n19618), .A2(n25673), .ZN(n19675) );
  CLKNHSV2 U14024 ( .I(n19365), .ZN(n12121) );
  INAND2HSV4 U14025 ( .A1(n25673), .B1(n25339), .ZN(n19676) );
  XNOR2HSV4 U14026 ( .A1(n19611), .A2(n19612), .ZN(n25673) );
  NAND2HSV2 U14027 ( .A1(n19610), .A2(n24271), .ZN(n19612) );
  XNOR2HSV4 U14028 ( .A1(n19609), .A2(n12122), .ZN(n19611) );
  BUFHSV8 U14029 ( .I(n25818), .Z(n12123) );
  CLKNHSV8 U14030 ( .I(n23455), .ZN(n25818) );
  CLKNAND2HSV4 U14031 ( .A1(n12124), .A2(n19159), .ZN(n23455) );
  CLKNAND2HSV4 U14032 ( .A1(pov6[11]), .A2(n19127), .ZN(n12124) );
  XNOR2HSV4 U14033 ( .A1(n19044), .A2(n12125), .ZN(pov6[11]) );
  CLKNHSV2 U14034 ( .I(n19043), .ZN(n12125) );
  CLKNAND2HSV2 U14035 ( .A1(n21061), .A2(n21060), .ZN(n12126) );
  INHSV2 U14036 ( .I(n12128), .ZN(n12740) );
  CLKNAND2HSV2 U14037 ( .A1(n21239), .A2(n28693), .ZN(n12128) );
  BUFHSV8 U14038 ( .I(n24893), .Z(n12129) );
  CLKNAND2HSV4 U14039 ( .A1(n12130), .A2(n21786), .ZN(n21909) );
  CLKNAND2HSV3 U14040 ( .A1(n23437), .A2(n23436), .ZN(n12130) );
  XNOR2HSV4 U14041 ( .A1(n25034), .A2(n21734), .ZN(n23437) );
  CLKNAND2HSV2 U14042 ( .A1(\pe5/aot [15]), .A2(\pe5/bq[16] ), .ZN(n14453) );
  XNOR2HSV4 U14043 ( .A1(n12131), .A2(n18018), .ZN(n18020) );
  XOR3HSV2 U14044 ( .A1(n18009), .A2(n12133), .A3(n12132), .Z(n12131) );
  CLKNHSV2 U14045 ( .I(n18011), .ZN(n12132) );
  XOR2HSV2 U14046 ( .A1(n18008), .A2(\pe9/phq [7]), .Z(n12133) );
  OAI21HSV4 U14047 ( .A1(n18918), .A2(n19068), .B(n18917), .ZN(n12489) );
  XNOR2HSV4 U14048 ( .A1(n19043), .A2(n12134), .ZN(n18918) );
  XNOR2HSV4 U14049 ( .A1(n12136), .A2(n12135), .ZN(n12134) );
  NAND3HSV4 U14050 ( .A1(n12137), .A2(n18910), .A3(n13985), .ZN(n19043) );
  CLKNAND2HSV3 U14051 ( .A1(n14743), .A2(n18908), .ZN(n12137) );
  XNOR2HSV4 U14052 ( .A1(n19124), .A2(n18845), .ZN(n12135) );
  CLKNAND2HSV2 U14053 ( .A1(n18851), .A2(n18850), .ZN(n12136) );
  CLKNAND2HSV2 U14054 ( .A1(n12430), .A2(n14744), .ZN(n18910) );
  XOR2HSV2 U14055 ( .A1(n21286), .A2(n12138), .Z(n21288) );
  CLKNAND2HSV2 U14056 ( .A1(n28942), .A2(n12139), .ZN(n12138) );
  CLKNHSV2 U14057 ( .I(n17781), .ZN(n12139) );
  CLKNAND2HSV2 U14058 ( .A1(n29041), .A2(n21714), .ZN(n12140) );
  NAND2HSV3 U14059 ( .A1(n12141), .A2(n19066), .ZN(n12225) );
  CLKNAND2HSV0 U14060 ( .A1(\pe5/bq[15] ), .A2(\pe5/aot [16]), .ZN(n14454) );
  CLKNHSV2 U14061 ( .I(n23438), .ZN(n28922) );
  INAND2HSV4 U14062 ( .A1(n23438), .B1(\pe11/got [11]), .ZN(n24744) );
  INAND2HSV4 U14063 ( .A1(n23438), .B1(\pe11/got [10]), .ZN(n24849) );
  INAND2HSV4 U14064 ( .A1(n23438), .B1(n20227), .ZN(n24804) );
  INAND2HSV4 U14065 ( .A1(n23438), .B1(\pe11/got [6]), .ZN(n24878) );
  INAND2HSV4 U14066 ( .A1(n23438), .B1(\pe11/got [7]), .ZN(n24954) );
  CLKNHSV2 U14067 ( .I(\pe5/aot [15]), .ZN(n28687) );
  CLKNHSV2 U14068 ( .I(n14474), .ZN(n27191) );
  CLKNHSV0 U14069 ( .I(n12142), .ZN(n14475) );
  NOR2HSV1 U14070 ( .A1(n14484), .A2(n12143), .ZN(n12142) );
  CLKNAND2HSV3 U14071 ( .A1(n14474), .A2(n14473), .ZN(n12143) );
  CLKNAND2HSV4 U14072 ( .A1(n14442), .A2(n14441), .ZN(n14474) );
  CLKNAND2HSV0 U14073 ( .A1(\pe6/bq[15] ), .A2(\pe6/aot [13]), .ZN(n14219) );
  XNOR2HSV4 U14074 ( .A1(n12148), .A2(n12144), .ZN(n14507) );
  XOR2HSV2 U14075 ( .A1(n12145), .A2(n20953), .Z(n12144) );
  XOR2HSV2 U14076 ( .A1(n12147), .A2(n12146), .Z(n12145) );
  CLKNAND2HSV2 U14077 ( .A1(\pe5/bq[15] ), .A2(\pe5/aot [14]), .ZN(n12146) );
  CLKNAND2HSV0 U14078 ( .A1(\pe5/aot [13]), .A2(\pe5/bq[16] ), .ZN(n12147) );
  MUX2NHSV2 U14079 ( .I0(n14504), .I1(n12151), .S(n12150), .ZN(n12149) );
  CLKNHSV2 U14080 ( .I(\pe5/phq [4]), .ZN(n12150) );
  CLKNHSV2 U14081 ( .I(n14505), .ZN(n12151) );
  CLKNAND2HSV2 U14082 ( .A1(\pe5/aot [15]), .A2(\pe5/bq[14] ), .ZN(n14505) );
  XNOR2HSV4 U14083 ( .A1(n12156), .A2(n12154), .ZN(n14226) );
  XNOR2HSV4 U14084 ( .A1(n12155), .A2(n14218), .ZN(n12154) );
  XOR2HSV2 U14085 ( .A1(n14219), .A2(n14216), .Z(n12156) );
  XNOR2HSV4 U14086 ( .A1(n12157), .A2(n14224), .ZN(n14225) );
  XNOR2HSV4 U14087 ( .A1(n14222), .A2(n14221), .ZN(n12157) );
  INHSV2 U14088 ( .I(n16885), .ZN(n12158) );
  CLKNAND2HSV4 U14089 ( .A1(n12492), .A2(n16884), .ZN(n12159) );
  NAND3HSV4 U14090 ( .A1(n12492), .A2(n16885), .A3(n16884), .ZN(n12160) );
  CLKNAND2HSV2 U14091 ( .A1(n12367), .A2(n16999), .ZN(n16937) );
  INHSV2 U14092 ( .I(n12161), .ZN(n19199) );
  XNOR2HSV4 U14093 ( .A1(n19197), .A2(n19198), .ZN(n12161) );
  NAND3HSV2 U14094 ( .A1(n12161), .A2(n19202), .A3(n19201), .ZN(n19203) );
  XNOR2HSV4 U14095 ( .A1(n12164), .A2(n12162), .ZN(n12173) );
  XNOR2HSV4 U14096 ( .A1(n12163), .A2(\pe5/phq [5]), .ZN(n12162) );
  CLKNHSV2 U14097 ( .I(n14434), .ZN(n12163) );
  CLKNAND2HSV2 U14098 ( .A1(n12165), .A2(n14440), .ZN(n12164) );
  CLKNAND2HSV2 U14099 ( .A1(n12167), .A2(n12166), .ZN(n12165) );
  CLKNHSV2 U14100 ( .I(n14534), .ZN(n12166) );
  CLKNHSV2 U14101 ( .I(n14505), .ZN(n12167) );
  INHSV2 U14102 ( .I(n14474), .ZN(n14583) );
  XOR3HSV2 U14103 ( .A1(n12173), .A2(n12170), .A3(n12168), .Z(n14462) );
  CLKNAND2HSV2 U14104 ( .A1(n14474), .A2(n12169), .ZN(n12168) );
  CLKNHSV2 U14105 ( .I(n20869), .ZN(n12169) );
  XNOR2HSV4 U14106 ( .A1(n12172), .A2(n12171), .ZN(n12170) );
  XOR2HSV2 U14107 ( .A1(n14436), .A2(n14437), .Z(n12171) );
  XOR2HSV2 U14108 ( .A1(n14435), .A2(n14438), .Z(n12172) );
  NOR2HSV4 U14109 ( .A1(n12176), .A2(n12175), .ZN(n12174) );
  AOI22HSV4 U14110 ( .A1(\pe5/aot [16]), .A2(\pe5/bq[11] ), .B1(\pe5/bq[14] ), 
        .B2(\pe5/aot [13]), .ZN(n12175) );
  NOR2HSV4 U14111 ( .A1(n14835), .A2(n14765), .ZN(n12176) );
  CLKNAND2HSV2 U14112 ( .A1(\pe5/aot [13]), .A2(\pe5/bq[11] ), .ZN(n14765) );
  CLKNAND2HSV2 U14113 ( .A1(\pe5/bq[14] ), .A2(\pe5/aot [16]), .ZN(n14835) );
  INHSV2 U14114 ( .I(n12178), .ZN(n19578) );
  CLKNAND2HSV2 U14115 ( .A1(n19671), .A2(n12177), .ZN(n12178) );
  CLKNHSV2 U14116 ( .I(n12179), .ZN(n12177) );
  CLKNHSV2 U14117 ( .I(n24271), .ZN(n12179) );
  INHSV2 U14118 ( .I(n12180), .ZN(n12185) );
  AOI21HSV4 U14119 ( .A1(n28678), .A2(n14369), .B(n14368), .ZN(n22995) );
  OAI21HSV4 U14120 ( .A1(n28678), .A2(n14368), .B(n12181), .ZN(n14393) );
  AOI21HSV4 U14121 ( .A1(n12184), .A2(n12183), .B(n12182), .ZN(n12181) );
  CLKNHSV2 U14122 ( .I(n14236), .ZN(n12182) );
  CLKNHSV2 U14123 ( .I(n14369), .ZN(n12183) );
  CLKNHSV2 U14124 ( .I(n14368), .ZN(n12184) );
  CLKNHSV2 U14125 ( .I(n22995), .ZN(n12180) );
  CLKNAND2HSV1 U14126 ( .A1(\pe5/got [16]), .A2(\pe5/ti_1 ), .ZN(n12186) );
  CLKNAND2HSV2 U14127 ( .A1(\pe5/got [16]), .A2(\pe5/ti_1 ), .ZN(n12187) );
  CLKNAND2HSV2 U14128 ( .A1(\pe5/bq[16] ), .A2(\pe5/aot [16]), .ZN(n12188) );
  CLKNAND2HSV2 U14129 ( .A1(\pe5/ctrq ), .A2(\pe5/pvq [1]), .ZN(n12190) );
  CLKNHSV4 U14130 ( .I(n12189), .ZN(n14444) );
  OAI21HSV4 U14131 ( .A1(n14444), .A2(n14443), .B(n21346), .ZN(n14442) );
  NOR2HSV4 U14132 ( .A1(n12191), .A2(n12192), .ZN(n14443) );
  NAND2HSV4 U14133 ( .A1(\pe6/bq[16] ), .A2(\pe6/aot [16]), .ZN(n14091) );
  CLKNAND2HSV2 U14134 ( .A1(n28406), .A2(n28137), .ZN(n19818) );
  CLKNAND2HSV4 U14135 ( .A1(n28582), .A2(n14070), .ZN(n16838) );
  XOR2HSV4 U14136 ( .A1(n16838), .A2(n16839), .Z(n16840) );
  NAND2HSV2 U14137 ( .A1(\pe5/bq[14] ), .A2(\pe5/aot [12]), .ZN(n14586) );
  CLKNAND2HSV4 U14138 ( .A1(n14683), .A2(n14685), .ZN(n14566) );
  CLKNAND2HSV2 U14139 ( .A1(n14057), .A2(n14558), .ZN(n14494) );
  INHSV4 U14140 ( .I(n14494), .ZN(n14500) );
  OAI21HSV4 U14141 ( .A1(n14576), .A2(n14684), .B(n14473), .ZN(n14479) );
  INHSV4 U14142 ( .I(n14479), .ZN(n14490) );
  INHSV4 U14143 ( .I(n19133), .ZN(n19134) );
  CLKNAND2HSV4 U14144 ( .A1(n22434), .A2(n22696), .ZN(n22675) );
  CLKNAND2HSV4 U14145 ( .A1(n15016), .A2(n15015), .ZN(n15089) );
  NAND2HSV4 U14146 ( .A1(n15089), .A2(n23414), .ZN(n12456) );
  INHSV4 U14147 ( .I(\pe5/bq[15] ), .ZN(n14433) );
  NAND2HSV4 U14148 ( .A1(n12773), .A2(n12774), .ZN(n14333) );
  NAND2HSV4 U14149 ( .A1(n20505), .A2(\pe11/got [12]), .ZN(n20323) );
  OAI211HSV1 U14150 ( .A1(n28343), .A2(n13126), .B(n28347), .C(n18330), .ZN(
        n28352) );
  NAND3HSV3 U14151 ( .A1(n28352), .A2(n28351), .A3(n28350), .ZN(n28353) );
  NAND2HSV2 U14152 ( .A1(n24966), .A2(\pe11/got [11]), .ZN(n20434) );
  CLKNAND2HSV4 U14153 ( .A1(n21741), .A2(n14070), .ZN(n12958) );
  CLKXOR2HSV2 U14154 ( .A1(n25179), .A2(n25178), .Z(n25180) );
  AOI31HSV2 U14155 ( .A1(n27119), .A2(n15289), .A3(n15242), .B(n16015), .ZN(
        n15290) );
  INHSV2 U14156 ( .I(n15290), .ZN(n15293) );
  OAI21HSV4 U14157 ( .A1(n18154), .A2(n12287), .B(n18152), .ZN(n18177) );
  NOR2HSV4 U14158 ( .A1(n14931), .A2(n20869), .ZN(n14801) );
  CLKNAND2HSV4 U14159 ( .A1(n14512), .A2(n14511), .ZN(n14528) );
  NAND2HSV4 U14160 ( .A1(n14610), .A2(n14609), .ZN(n14611) );
  CLKXOR2HSV4 U14161 ( .A1(n19937), .A2(n19936), .Z(n19939) );
  XOR2HSV4 U14162 ( .A1(n19939), .A2(n19938), .Z(n19942) );
  NAND2HSV2 U14163 ( .A1(n28658), .A2(n28390), .ZN(n25693) );
  NAND3HSV4 U14164 ( .A1(n14273), .A2(n14271), .A3(n14267), .ZN(n14268) );
  NAND3HSV2 U14165 ( .A1(\pe11/phq [1]), .A2(\pe11/bq[16] ), .A3(
        \pe11/aot [16]), .ZN(n14754) );
  NOR2HSV4 U14166 ( .A1(n15206), .A2(n15205), .ZN(n15233) );
  NAND2HSV2 U14167 ( .A1(n28702), .A2(n14052), .ZN(n27658) );
  NAND2HSV2 U14168 ( .A1(\pe9/bq[16] ), .A2(\pe9/aot [13]), .ZN(n13520) );
  NAND2HSV4 U14169 ( .A1(n14552), .A2(n24635), .ZN(n14461) );
  CLKNAND2HSV4 U14170 ( .A1(n14495), .A2(n27191), .ZN(n14501) );
  CLKAND2HSV2 U14171 ( .A1(n14501), .A2(n14631), .Z(n14502) );
  CLKNAND2HSV2 U14172 ( .A1(n23388), .A2(n23387), .ZN(n23409) );
  AOI21HSV4 U14173 ( .A1(n20369), .A2(n20368), .B(n20372), .ZN(n20362) );
  OAI22HSV4 U14174 ( .A1(n23404), .A2(n27127), .B1(n23403), .B2(n23402), .ZN(
        n23405) );
  CLKNAND2HSV2 U14175 ( .A1(n28793), .A2(n14236), .ZN(n14331) );
  NAND2HSV4 U14176 ( .A1(n12470), .A2(n21346), .ZN(n14681) );
  INHSV4 U14177 ( .I(n25642), .ZN(n19268) );
  NOR2HSV4 U14178 ( .A1(n19268), .A2(n19466), .ZN(n19270) );
  NAND2HSV2 U14179 ( .A1(\pe3/bq[16] ), .A2(\pe3/aot [16]), .ZN(n15008) );
  NAND2HSV2 U14180 ( .A1(n27106), .A2(n28640), .ZN(n27110) );
  CLKNAND2HSV4 U14181 ( .A1(n25648), .A2(n14257), .ZN(n14258) );
  CLKNAND2HSV4 U14182 ( .A1(n28798), .A2(n14236), .ZN(n14120) );
  NAND2HSV4 U14183 ( .A1(n14286), .A2(n14284), .ZN(n14259) );
  NAND2HSV2 U14184 ( .A1(n14193), .A2(n19160), .ZN(n14194) );
  OAI21HSV4 U14185 ( .A1(n14195), .A2(n14194), .B(n18907), .ZN(n14196) );
  NAND2HSV2 U14186 ( .A1(n14552), .A2(n14463), .ZN(n14477) );
  NAND2HSV2 U14187 ( .A1(n20052), .A2(n13998), .ZN(n23867) );
  NAND2HSV4 U14188 ( .A1(n13120), .A2(n13119), .ZN(n13121) );
  OAI21HSV4 U14189 ( .A1(n28919), .A2(n20781), .B(n20703), .ZN(n20765) );
  NAND2HSV2 U14190 ( .A1(n28420), .A2(\pe8/got [3]), .ZN(n13590) );
  NAND2HSV2 U14191 ( .A1(n13590), .A2(n13589), .ZN(n13591) );
  CLKNAND2HSV2 U14192 ( .A1(\pe5/aot [15]), .A2(n23909), .ZN(n14537) );
  XOR2HSV0 U14193 ( .A1(n14537), .A2(n14536), .Z(n14540) );
  INHSV2 U14194 ( .I(n19158), .ZN(n22078) );
  NOR2HSV4 U14195 ( .A1(n14485), .A2(n14583), .ZN(n14487) );
  INHSV4 U14196 ( .I(\pe5/ctrq ), .ZN(n14448) );
  CLKNAND2HSV3 U14197 ( .A1(n12196), .A2(n12195), .ZN(n12194) );
  INHSV2 U14198 ( .I(n19946), .ZN(n12195) );
  CLKNAND2HSV0 U14199 ( .A1(n14755), .A2(n14754), .ZN(n12197) );
  CLKNHSV2 U14200 ( .I(n25502), .ZN(n20181) );
  XNOR2HSV4 U14201 ( .A1(n12198), .A2(n12197), .ZN(n25502) );
  NAND3HSV4 U14202 ( .A1(n14751), .A2(n14750), .A3(n14749), .ZN(n12198) );
  CLKNAND2HSV3 U14203 ( .A1(n12199), .A2(n25656), .ZN(n12504) );
  CLKNAND2HSV4 U14204 ( .A1(n14566), .A2(n14567), .ZN(n12199) );
  NOR2HSV4 U14205 ( .A1(n12199), .A2(n14568), .ZN(n14569) );
  NOR2HSV4 U14206 ( .A1(n12199), .A2(n14617), .ZN(n14618) );
  CLKNAND2HSV2 U14207 ( .A1(n12471), .A2(n12199), .ZN(n14571) );
  CLKNAND2HSV4 U14208 ( .A1(n24881), .A2(n20466), .ZN(n25055) );
  CLKNAND2HSV4 U14209 ( .A1(n12201), .A2(n12200), .ZN(n24881) );
  CLKNAND2HSV2 U14210 ( .A1(n20765), .A2(n20766), .ZN(n12200) );
  CLKNAND2HSV3 U14211 ( .A1(n25055), .A2(n25053), .ZN(n25414) );
  AOI22HSV4 U14212 ( .A1(n14631), .A2(n20868), .B1(n28971), .B2(n14926), .ZN(
        n13414) );
  XNOR2HSV4 U14213 ( .A1(n14923), .A2(n20860), .ZN(n28971) );
  CLKNAND2HSV3 U14214 ( .A1(n25050), .A2(n12202), .ZN(n12207) );
  CLKNHSV4 U14215 ( .I(n25055), .ZN(n12202) );
  CLKNAND2HSV4 U14216 ( .A1(n24957), .A2(n20561), .ZN(n12203) );
  XOR3HSV2 U14217 ( .A1(n12214), .A2(n12204), .A3(n12203), .Z(po11) );
  AOI21HSV4 U14218 ( .A1(n12207), .A2(n12206), .B(n12205), .ZN(n12204) );
  MUX2NHSV2 U14219 ( .I0(n12213), .I1(n12212), .S(n25054), .ZN(n12205) );
  CLKNAND2HSV2 U14220 ( .A1(n25055), .A2(n12208), .ZN(n12206) );
  NAND3HSV2 U14221 ( .A1(n12446), .A2(n12444), .A3(n12209), .ZN(n12208) );
  INHSV2 U14222 ( .I(n12210), .ZN(n12209) );
  INHSV2 U14223 ( .I(n25053), .ZN(n12211) );
  CLKNHSV0 U14224 ( .I(n25051), .ZN(n12212) );
  INHSV2 U14225 ( .I(n25052), .ZN(n12213) );
  INHSV1 U14226 ( .I(n25056), .ZN(n12214) );
  CLKNAND2HSV0 U14227 ( .A1(n12216), .A2(n12215), .ZN(n21716) );
  NAND3HSV4 U14228 ( .A1(n12216), .A2(n14628), .A3(n12215), .ZN(n12476) );
  CLKNHSV4 U14229 ( .I(n12399), .ZN(n12216) );
  NOR2HSV4 U14230 ( .A1(n25605), .A2(n12217), .ZN(n12221) );
  CLKNAND2HSV2 U14231 ( .A1(n12218), .A2(n12219), .ZN(n12222) );
  CLKNHSV2 U14232 ( .I(n23867), .ZN(n12218) );
  CLKNHSV2 U14233 ( .I(n12222), .ZN(n25605) );
  CLKNHSV2 U14234 ( .I(n20055), .ZN(n12219) );
  CLKNAND2HSV3 U14235 ( .A1(n12220), .A2(n20053), .ZN(n20064) );
  CLKNAND2HSV3 U14236 ( .A1(n12221), .A2(n25613), .ZN(n12220) );
  CLKNAND2HSV3 U14237 ( .A1(n12223), .A2(n20057), .ZN(n25613) );
  CLKNAND2HSV1 U14238 ( .A1(n19985), .A2(n20052), .ZN(n20057) );
  INHSV2 U14239 ( .I(n20054), .ZN(n12223) );
  CLKNAND2HSV3 U14240 ( .A1(n12226), .A2(n12225), .ZN(n12224) );
  CLKNAND2HSV3 U14241 ( .A1(pov6[15]), .A2(n19141), .ZN(n12227) );
  OAI21HSV4 U14242 ( .A1(n12226), .A2(n12225), .B(n12224), .ZN(pov6[15]) );
  CLKNAND2HSV3 U14243 ( .A1(n12227), .A2(n19143), .ZN(n28925) );
  NOR2HSV4 U14244 ( .A1(n12228), .A2(n20619), .ZN(n20183) );
  NOR2HSV4 U14245 ( .A1(n20219), .A2(n12228), .ZN(n20344) );
  NOR2HSV4 U14246 ( .A1(n25505), .A2(n20185), .ZN(n12228) );
  XNOR2HSV4 U14247 ( .A1(n12229), .A2(n20239), .ZN(n20241) );
  XNOR2HSV4 U14248 ( .A1(n12230), .A2(n20236), .ZN(n12229) );
  XNOR2HSV4 U14249 ( .A1(n12231), .A2(\pe11/phq [6]), .ZN(n12230) );
  CLKNAND2HSV2 U14250 ( .A1(n20587), .A2(\pe11/got [11]), .ZN(n12231) );
  CLKNHSV2 U14251 ( .I(n20865), .ZN(n13413) );
  XNOR2HSV4 U14252 ( .A1(n12235), .A2(n12233), .ZN(n12232) );
  XNOR2HSV4 U14253 ( .A1(n14968), .A2(n12234), .ZN(n12233) );
  XNOR2HSV4 U14254 ( .A1(n14969), .A2(n14970), .ZN(n12234) );
  NOR2HSV2 U14255 ( .A1(n20983), .A2(n21411), .ZN(n12235) );
  OAI211HSV2 U14256 ( .A1(n20849), .A2(n20985), .B(n12238), .C(n12237), .ZN(
        n12236) );
  NOR2HSV4 U14257 ( .A1(n20917), .A2(n13639), .ZN(n12237) );
  CLKNHSV2 U14258 ( .I(n20920), .ZN(n12238) );
  CLKNHSV2 U14259 ( .I(n19980), .ZN(n19977) );
  CLKNAND2HSV0 U14260 ( .A1(n12239), .A2(n19830), .ZN(n19978) );
  CLKNAND2HSV1 U14261 ( .A1(n19980), .A2(n12240), .ZN(n12239) );
  INHSV2 U14262 ( .I(n19976), .ZN(n12240) );
  CLKNAND2HSV4 U14263 ( .A1(n12242), .A2(n12241), .ZN(n19980) );
  NOR2HSV4 U14264 ( .A1(n14908), .A2(n13191), .ZN(n12243) );
  NAND2HSV3 U14265 ( .A1(n12243), .A2(n14816), .ZN(n14864) );
  NAND3HSV4 U14266 ( .A1(n12243), .A2(n14816), .A3(n14628), .ZN(n14818) );
  CLKNAND2HSV2 U14267 ( .A1(\pe5/bq[16] ), .A2(\pe5/aot [16]), .ZN(n12244) );
  NOR2HSV4 U14268 ( .A1(n12245), .A2(n18658), .ZN(n18694) );
  NOR2HSV3 U14269 ( .A1(n12245), .A2(n18717), .ZN(n18756) );
  NOR2HSV4 U14270 ( .A1(n29007), .A2(n18657), .ZN(n12245) );
  NOR2HSV8 U14271 ( .A1(n12247), .A2(n12246), .ZN(n14481) );
  CLKNAND2HSV4 U14272 ( .A1(n14519), .A2(n21346), .ZN(n12246) );
  CLKNAND2HSV2 U14273 ( .A1(n14460), .A2(n14909), .ZN(n14514) );
  NOR2HSV2 U14274 ( .A1(n14058), .A2(n14483), .ZN(n14488) );
  NOR2HSV4 U14275 ( .A1(n14480), .A2(n14481), .ZN(n14058) );
  OAI21HSV4 U14276 ( .A1(n14513), .A2(n14514), .B(n14518), .ZN(n14480) );
  XNOR2HSV4 U14277 ( .A1(n14456), .A2(n14455), .ZN(n14513) );
  CLKNAND2HSV2 U14278 ( .A1(n14042), .A2(\pe8/got [9]), .ZN(n19886) );
  CLKNAND2HSV2 U14279 ( .A1(n14042), .A2(n23605), .ZN(n20036) );
  CLKNAND2HSV2 U14280 ( .A1(n14042), .A2(\pe8/got [5]), .ZN(n22174) );
  CLKNAND2HSV2 U14281 ( .A1(n14042), .A2(n25577), .ZN(n22312) );
  CLKNAND2HSV2 U14282 ( .A1(n14042), .A2(\pe8/got [2]), .ZN(n22267) );
  CLKNAND2HSV2 U14283 ( .A1(n14042), .A2(\pe8/got [3]), .ZN(n23585) );
  CLKNAND2HSV0 U14284 ( .A1(n14042), .A2(\pe8/got [6]), .ZN(n23646) );
  CLKNAND2HSV2 U14285 ( .A1(n14042), .A2(n26230), .ZN(n23743) );
  CLKNAND2HSV2 U14286 ( .A1(n14042), .A2(n14060), .ZN(n25587) );
  OAI21HSV2 U14287 ( .A1(n19884), .A2(n19883), .B(n19885), .ZN(n14042) );
  NOR2HSV4 U14288 ( .A1(n12248), .A2(n18656), .ZN(n18703) );
  NOR2HSV4 U14289 ( .A1(n12248), .A2(n16555), .ZN(n16605) );
  NOR2HSV4 U14290 ( .A1(n16552), .A2(n12249), .ZN(n12248) );
  CLKNAND2HSV2 U14291 ( .A1(n12250), .A2(n16587), .ZN(n16597) );
  CLKNHSV2 U14292 ( .I(n16608), .ZN(n12250) );
  OAI21HSV4 U14293 ( .A1(n19883), .A2(n19884), .B(n19885), .ZN(n18690) );
  CLKNHSV2 U14294 ( .I(n19835), .ZN(n12251) );
  CLKNAND2HSV4 U14295 ( .A1(n28965), .A2(n14526), .ZN(n21464) );
  INHSV8 U14296 ( .I(n12252), .ZN(n24377) );
  NOR2HSV4 U14297 ( .A1(n12254), .A2(n12253), .ZN(n12252) );
  NOR2HSV4 U14298 ( .A1(n21002), .A2(n12255), .ZN(n12253) );
  OAI21HSV4 U14299 ( .A1(n21001), .A2(n12255), .B(n21463), .ZN(n12254) );
  CLKNHSV2 U14300 ( .I(n14526), .ZN(n12255) );
  CLKNAND2HSV2 U14301 ( .A1(n24377), .A2(\pe5/got [2]), .ZN(n12914) );
  XNOR2HSV4 U14302 ( .A1(n12259), .A2(n12256), .ZN(n12975) );
  XNOR2HSV4 U14303 ( .A1(n12258), .A2(n12257), .ZN(n12256) );
  XOR2HSV2 U14304 ( .A1(n25201), .A2(n25202), .Z(n12257) );
  CLKNAND2HSV2 U14305 ( .A1(n28616), .A2(n26230), .ZN(n12258) );
  CLKNHSV2 U14306 ( .I(n12974), .ZN(n12259) );
  NAND2HSV4 U14307 ( .A1(n15003), .A2(n15002), .ZN(n29050) );
  INHSV2 U14308 ( .I(n27220), .ZN(n27221) );
  CLKNAND2HSV2 U14309 ( .A1(n21897), .A2(n28590), .ZN(n21903) );
  INOR2HSV2 U14310 ( .A1(n25681), .B1(n25682), .ZN(n13600) );
  CLKNAND2HSV2 U14311 ( .A1(n14982), .A2(n14987), .ZN(n14983) );
  NAND3HSV3 U14312 ( .A1(n28814), .A2(n15001), .A3(n17617), .ZN(n15002) );
  BUFHSV4 U14313 ( .I(n16535), .Z(n18823) );
  CLKXOR2HSV4 U14314 ( .A1(n18754), .A2(n18753), .Z(n18755) );
  INHSV2 U14315 ( .I(n15704), .ZN(n15620) );
  NAND2HSV4 U14316 ( .A1(n22690), .A2(n22689), .ZN(n22718) );
  NAND2HSV2 U14317 ( .A1(n22690), .A2(n22689), .ZN(n22624) );
  INHSV2 U14318 ( .I(n22624), .ZN(n24451) );
  CLKXOR2HSV4 U14319 ( .A1(n21735), .A2(poh11[13]), .Z(po[14]) );
  AND2HSV2 U14320 ( .A1(n28703), .A2(n14022), .Z(n23904) );
  INHSV2 U14321 ( .I(n25520), .ZN(n12260) );
  NAND2HSV2 U14322 ( .A1(n17692), .A2(n17693), .ZN(n12701) );
  MOAI22HSV4 U14323 ( .A1(n22091), .A2(n19368), .B1(n19466), .B2(
        \pe7/ti_7t [5]), .ZN(n19369) );
  INHSV4 U14324 ( .I(n19617), .ZN(n19708) );
  NAND2HSV0 U14325 ( .A1(n13499), .A2(n23424), .ZN(n13500) );
  OAI21HSV0 U14326 ( .A1(n13499), .A2(n23424), .B(n13500), .ZN(pov8[14]) );
  CLKNAND2HSV2 U14327 ( .A1(n16047), .A2(n16046), .ZN(n16048) );
  CLKNAND2HSV2 U14328 ( .A1(n21312), .A2(n23382), .ZN(n21314) );
  INOR2HSV1 U14329 ( .A1(n26349), .B1(n24313), .ZN(n26411) );
  NOR2HSV2 U14330 ( .A1(n17349), .A2(n17348), .ZN(n17352) );
  CLKNAND2HSV4 U14331 ( .A1(n17804), .A2(n17774), .ZN(n17807) );
  NAND2HSV2 U14332 ( .A1(n20143), .A2(n20144), .ZN(n20147) );
  INHSV2 U14333 ( .I(n28347), .ZN(n13810) );
  MUX2NHSV1 U14334 ( .I0(n28347), .I1(n13810), .S(n13813), .ZN(pov9[15]) );
  NAND2HSV0 U14335 ( .A1(n28421), .A2(n28590), .ZN(n13886) );
  OAI31HSV2 U14336 ( .A1(n23717), .A2(n23719), .A3(n13811), .B(n13812), .ZN(
        n13813) );
  NAND2HSV4 U14337 ( .A1(n15810), .A2(n15809), .ZN(n15830) );
  INHSV4 U14338 ( .I(n19044), .ZN(n19047) );
  INHSV4 U14339 ( .I(n23997), .ZN(n25784) );
  NAND2HSV2 U14340 ( .A1(n28940), .A2(n22992), .ZN(n12315) );
  XOR3HSV2 U14341 ( .A1(n12591), .A2(n12261), .A3(n12588), .Z(n26999) );
  XNOR2HSV4 U14342 ( .A1(n26997), .A2(n26996), .ZN(n12261) );
  CLKNHSV6 U14343 ( .I(n27941), .ZN(n25079) );
  NAND2HSV0 U14344 ( .A1(n28012), .A2(\pe4/got [4]), .ZN(n28013) );
  NAND2HSV0 U14345 ( .A1(n28012), .A2(\pe4/got [16]), .ZN(n26998) );
  NAND2HSV0 U14346 ( .A1(n28012), .A2(n25134), .ZN(n25135) );
  MUX2NHSV2 U14347 ( .I0(n13087), .I1(n19125), .S(n13089), .ZN(n19128) );
  INAND2HSV2 U14348 ( .A1(n27223), .B1(n27220), .ZN(n26414) );
  NOR2HSV0 U14349 ( .A1(n27217), .A2(n27220), .ZN(n22077) );
  XNOR2HSV4 U14350 ( .A1(n17466), .A2(n17465), .ZN(n17467) );
  NAND2HSV0 U14351 ( .A1(n25901), .A2(n28425), .ZN(n12753) );
  INHSV4 U14352 ( .I(n21981), .ZN(n21984) );
  NAND2HSV4 U14353 ( .A1(n15897), .A2(n15896), .ZN(n21981) );
  INHSV4 U14354 ( .I(n21980), .ZN(n21983) );
  CLKNAND2HSV2 U14355 ( .A1(n16675), .A2(n12369), .ZN(n16676) );
  INHSV4 U14356 ( .I(n16994), .ZN(n21738) );
  NAND3HSV4 U14357 ( .A1(n23476), .A2(n16710), .A3(n16709), .ZN(n16797) );
  XNOR2HSV4 U14358 ( .A1(n20122), .A2(n20121), .ZN(n20124) );
  XOR2HSV0 U14359 ( .A1(n27187), .A2(n27186), .Z(n27188) );
  NAND2HSV4 U14360 ( .A1(n28704), .A2(n16995), .ZN(n12364) );
  CLKNAND2HSV2 U14361 ( .A1(n13755), .A2(n13754), .ZN(n13756) );
  OAI21HSV0 U14362 ( .A1(n13754), .A2(n13755), .B(n13756), .ZN(\pe10/poht [5])
         );
  CLKNHSV0 U14363 ( .I(n25690), .ZN(n13674) );
  CLKXOR2HSV4 U14364 ( .A1(n25127), .A2(n25126), .Z(n25130) );
  CLKNAND2HSV2 U14365 ( .A1(n18673), .A2(\pe8/pvq [4]), .ZN(n13438) );
  XNOR2HSV1 U14366 ( .A1(n23868), .A2(n25613), .ZN(n29004) );
  NAND2HSV0 U14367 ( .A1(n26909), .A2(\pe1/got [5]), .ZN(n26848) );
  NAND2HSV4 U14368 ( .A1(n17534), .A2(n17360), .ZN(n17413) );
  NAND2HSV4 U14369 ( .A1(n17361), .A2(n12742), .ZN(n17534) );
  XOR2HSV0 U14370 ( .A1(n26814), .A2(n12262), .Z(n26816) );
  XOR2HSV0 U14371 ( .A1(n26813), .A2(n26812), .Z(n12262) );
  INHSV6 U14372 ( .I(n22680), .ZN(n25060) );
  NOR2HSV2 U14373 ( .A1(n17342), .A2(n17341), .ZN(n17344) );
  INHSV4 U14374 ( .I(n17276), .ZN(n12331) );
  INHSV6 U14375 ( .I(n25680), .ZN(n17471) );
  AOI21HSV2 U14376 ( .A1(n21629), .A2(n21628), .B(n21631), .ZN(n21638) );
  INHSV6 U14377 ( .I(n21323), .ZN(n25901) );
  INHSV4 U14378 ( .I(n17402), .ZN(n21323) );
  XOR2HSV1 U14379 ( .A1(n27207), .A2(n27206), .Z(n27208) );
  XOR3HSV2 U14380 ( .A1(n23106), .A2(n23105), .A3(n23104), .Z(\pe4/poht [3])
         );
  XOR2HSV0 U14381 ( .A1(n23103), .A2(n23102), .Z(n23105) );
  NOR2HSV0 U14382 ( .A1(n21218), .A2(n17863), .ZN(n21219) );
  CLKNHSV0 U14383 ( .I(n20144), .ZN(n12263) );
  XNOR2HSV4 U14384 ( .A1(n12264), .A2(n12795), .ZN(n18614) );
  XNOR2HSV4 U14385 ( .A1(n18521), .A2(n18520), .ZN(n12264) );
  INHSV2 U14386 ( .I(n15705), .ZN(n12265) );
  INHSV4 U14387 ( .I(n15711), .ZN(n15705) );
  NAND2HSV4 U14388 ( .A1(n12340), .A2(n15475), .ZN(n12339) );
  NAND2HSV2 U14389 ( .A1(n17210), .A2(n17207), .ZN(n17223) );
  CLKNAND2HSV4 U14390 ( .A1(n28974), .A2(n15839), .ZN(n12340) );
  CLKNAND2HSV2 U14391 ( .A1(n17604), .A2(n28460), .ZN(n26824) );
  INHSV4 U14392 ( .I(n16642), .ZN(n22103) );
  OAI21HSV4 U14393 ( .A1(n16670), .A2(n16663), .B(n12819), .ZN(n16642) );
  NOR2HSV2 U14394 ( .A1(n26540), .A2(n26417), .ZN(n12733) );
  INHSV2 U14395 ( .I(n26540), .ZN(n26418) );
  NOR2HSV2 U14396 ( .A1(n26540), .A2(n17364), .ZN(n17538) );
  NAND2HSV2 U14397 ( .A1(\pe10/got [16]), .A2(\pe10/ti_1 ), .ZN(n16610) );
  XOR2HSV4 U14398 ( .A1(n22629), .A2(n22628), .Z(n22633) );
  CLKNAND2HSV2 U14399 ( .A1(n12286), .A2(n22630), .ZN(n22635) );
  INHSV2 U14400 ( .I(n22632), .ZN(n12286) );
  CLKNHSV0 U14401 ( .I(n21745), .ZN(n12266) );
  INHSV2 U14402 ( .I(n12266), .ZN(n12267) );
  NAND2HSV4 U14403 ( .A1(n17155), .A2(n17154), .ZN(n26426) );
  CLKNAND2HSV2 U14404 ( .A1(n16185), .A2(\pe1/ti_7t [1]), .ZN(n17154) );
  NAND3HSV3 U14405 ( .A1(n22795), .A2(n22794), .A3(n22793), .ZN(n22799) );
  NAND2HSV2 U14406 ( .A1(n22197), .A2(n22196), .ZN(\pe8/poht [2]) );
  NOR2HSV4 U14407 ( .A1(n16219), .A2(n16233), .ZN(n23478) );
  NOR2HSV2 U14408 ( .A1(n15490), .A2(n15489), .ZN(n12377) );
  INHSV4 U14409 ( .I(n19815), .ZN(n12268) );
  NAND2HSV2 U14410 ( .A1(n23115), .A2(n14030), .ZN(n25498) );
  NAND2HSV2 U14411 ( .A1(n23114), .A2(n23115), .ZN(n23119) );
  OAI21HSV2 U14412 ( .A1(n13578), .A2(n13579), .B(n13580), .ZN(n13581) );
  CLKXOR2HSV2 U14413 ( .A1(n24498), .A2(n24497), .Z(n13578) );
  NAND2HSV2 U14414 ( .A1(n13579), .A2(n13578), .ZN(n13580) );
  NAND2HSV2 U14415 ( .A1(n13582), .A2(n13581), .ZN(n13583) );
  NAND2HSV4 U14416 ( .A1(n22104), .A2(n16640), .ZN(n12419) );
  AOI21HSV4 U14417 ( .A1(n22103), .A2(n13915), .B(n16639), .ZN(n16640) );
  XOR3HSV2 U14418 ( .A1(n24130), .A2(n12269), .A3(n24129), .Z(n24131) );
  CLKNAND2HSV4 U14419 ( .A1(n22502), .A2(n22501), .ZN(n12626) );
  CLKNAND2HSV4 U14420 ( .A1(n12313), .A2(n17000), .ZN(n21741) );
  XNOR2HSV4 U14421 ( .A1(n15537), .A2(n15536), .ZN(n15559) );
  XNOR2HSV4 U14422 ( .A1(n15559), .A2(n15558), .ZN(n15560) );
  INHSV4 U14423 ( .I(n22102), .ZN(n13915) );
  INHSV4 U14424 ( .I(n15490), .ZN(n15564) );
  XNOR2HSV4 U14425 ( .A1(n17163), .A2(n17162), .ZN(n17164) );
  XNOR2HSV4 U14426 ( .A1(n17161), .A2(n17160), .ZN(n17163) );
  INAND2HSV2 U14427 ( .A1(n16809), .B1(\pe10/aot [7]), .ZN(n16909) );
  INAND2HSV2 U14428 ( .A1(n16809), .B1(\pe10/aot [8]), .ZN(n16851) );
  INAND2HSV2 U14429 ( .A1(n16809), .B1(\pe10/aot [12]), .ZN(n16688) );
  NAND2HSV2 U14430 ( .A1(n12609), .A2(n25674), .ZN(n12608) );
  CLKNHSV0 U14431 ( .I(n25674), .ZN(n19690) );
  CLKNHSV3 U14432 ( .I(n23871), .ZN(n24287) );
  NAND2HSV2 U14433 ( .A1(n18644), .A2(n18643), .ZN(n18653) );
  NOR2HSV0 U14434 ( .A1(n22084), .A2(n21242), .ZN(n12270) );
  NOR2HSV2 U14435 ( .A1(n22084), .A2(n21242), .ZN(n21153) );
  INHSV2 U14436 ( .I(n12597), .ZN(n12596) );
  AOI22HSV0 U14437 ( .A1(n21901), .A2(\pe2/ti_7t [15]), .B1(n23435), .B2(
        n21900), .ZN(n21902) );
  CLKNAND2HSV2 U14438 ( .A1(n21903), .A2(n21902), .ZN(n21908) );
  INAND2HSV4 U14439 ( .A1(n12729), .B1(n12731), .ZN(n17419) );
  INHSV2 U14440 ( .I(n22066), .ZN(n12271) );
  OAI21HSV4 U14441 ( .A1(n22066), .A2(n22065), .B(n22064), .ZN(n22067) );
  NAND2HSV2 U14442 ( .A1(n16648), .A2(n12418), .ZN(n16704) );
  INHSV2 U14443 ( .I(n21012), .ZN(n21013) );
  CLKXOR2HSV4 U14444 ( .A1(n15461), .A2(n15460), .Z(n15464) );
  XOR2HSV4 U14445 ( .A1(n15464), .A2(n15463), .Z(n15465) );
  XNOR2HSV4 U14446 ( .A1(n17464), .A2(n17463), .ZN(n17466) );
  CLKNAND2HSV4 U14447 ( .A1(n17473), .A2(n17426), .ZN(n17472) );
  INHSV2 U14448 ( .I(n18438), .ZN(n18441) );
  CLKXOR2HSV4 U14449 ( .A1(n16929), .A2(n16928), .Z(n16931) );
  OAI31HSV2 U14450 ( .A1(n27438), .A2(n21306), .A3(n21305), .B(n13204), .ZN(
        n13205) );
  AOI21HSV4 U14451 ( .A1(n28956), .A2(n12739), .B(n12737), .ZN(n27438) );
  XNOR2HSV4 U14452 ( .A1(n21307), .A2(n21306), .ZN(n21309) );
  INHSV4 U14453 ( .I(n22598), .ZN(n27197) );
  CLKNAND2HSV2 U14454 ( .A1(n13389), .A2(n15705), .ZN(n15852) );
  NOR2HSV2 U14455 ( .A1(n19158), .A2(n13469), .ZN(n12607) );
  CLKNAND2HSV2 U14456 ( .A1(n13593), .A2(n13594), .ZN(n13595) );
  OAI21HSV2 U14457 ( .A1(n13593), .A2(n13594), .B(n13595), .ZN(\pe11/poht [12]) );
  XNOR2HSV4 U14458 ( .A1(n12616), .A2(n12614), .ZN(n13593) );
  CLKNAND2HSV4 U14459 ( .A1(n15488), .A2(n13981), .ZN(n15496) );
  NAND2HSV4 U14460 ( .A1(n27229), .A2(n15486), .ZN(n15488) );
  INHSV4 U14461 ( .I(n19157), .ZN(n19057) );
  CLKNHSV0 U14462 ( .I(n15852), .ZN(n12272) );
  INHSV2 U14463 ( .I(n12272), .ZN(n12273) );
  CLKNAND2HSV4 U14464 ( .A1(n18459), .A2(n18458), .ZN(n18534) );
  NAND3HSV4 U14465 ( .A1(n15566), .A2(n15565), .A3(n15564), .ZN(n13503) );
  NAND2HSV4 U14466 ( .A1(n22043), .A2(n22042), .ZN(n14080) );
  XOR2HSV0 U14467 ( .A1(n24036), .A2(n12275), .Z(\pe7/poht [8]) );
  NOR2HSV2 U14468 ( .A1(n18335), .A2(n18334), .ZN(n18383) );
  INHSV4 U14469 ( .I(n22802), .ZN(n27942) );
  INOR2HSV4 U14470 ( .A1(n22802), .B1(n22880), .ZN(n13360) );
  INHSV4 U14471 ( .I(n22802), .ZN(n27876) );
  NAND2HSV4 U14472 ( .A1(n15829), .A2(n15828), .ZN(n22802) );
  NAND2HSV2 U14473 ( .A1(n18471), .A2(n18472), .ZN(n12795) );
  XNOR2HSV4 U14474 ( .A1(n21971), .A2(n21974), .ZN(pov4[13]) );
  NOR2HSV4 U14475 ( .A1(n21750), .A2(n21749), .ZN(n17234) );
  CLKNAND2HSV2 U14476 ( .A1(n12755), .A2(n12752), .ZN(n12751) );
  NAND3HSV2 U14477 ( .A1(n17363), .A2(n17407), .A3(n17346), .ZN(n12274) );
  NAND3HSV0 U14478 ( .A1(n17363), .A2(n17407), .A3(n17346), .ZN(n25879) );
  CLKXOR2HSV2 U14479 ( .A1(n21294), .A2(n21293), .Z(n12816) );
  BUFHSV2 U14480 ( .I(n25945), .Z(n28787) );
  INHSV4 U14481 ( .I(n25945), .ZN(n21765) );
  CLKXOR2HSV2 U14482 ( .A1(n25743), .A2(n25742), .Z(n25744) );
  BUFHSV4 U14483 ( .I(n22078), .Z(n26031) );
  CLKNHSV0 U14484 ( .I(n22071), .ZN(n12276) );
  INHSV2 U14485 ( .I(n12276), .ZN(n12277) );
  INHSV4 U14486 ( .I(n17521), .ZN(n16260) );
  INHSV2 U14487 ( .I(n12617), .ZN(n12616) );
  NAND2HSV4 U14488 ( .A1(n21975), .A2(n21973), .ZN(n21971) );
  XOR2HSV4 U14489 ( .A1(n16767), .A2(n16766), .Z(n16768) );
  CLKXOR2HSV4 U14490 ( .A1(n16765), .A2(n16764), .Z(n16766) );
  CLKNAND2HSV8 U14491 ( .A1(n12392), .A2(n22599), .ZN(n26215) );
  IAO21HSV2 U14492 ( .A1(n28996), .A2(n22442), .B(n12279), .ZN(n12278) );
  AO21HSV1 U14493 ( .A1(n22442), .A2(n16992), .B(n17065), .Z(n12279) );
  NAND2HSV2 U14494 ( .A1(n26082), .A2(n25419), .ZN(n25487) );
  MUX2NHSV4 U14495 ( .I0(n15447), .I1(n15448), .S(n12280), .ZN(n15449) );
  XNOR2HSV4 U14496 ( .A1(n15446), .A2(n13973), .ZN(n12280) );
  OAI21HSV4 U14497 ( .A1(n23420), .A2(n23419), .B(n23418), .ZN(n24628) );
  INHSV4 U14498 ( .I(n20131), .ZN(n23716) );
  CLKNAND2HSV2 U14499 ( .A1(n17125), .A2(n17124), .ZN(n22432) );
  XNOR2HSV4 U14500 ( .A1(n22187), .A2(n22186), .ZN(n22188) );
  XNOR2HSV4 U14501 ( .A1(n22191), .A2(n22190), .ZN(n22194) );
  XOR2HSV4 U14502 ( .A1(n22189), .A2(n22188), .Z(n22190) );
  NAND2HSV4 U14503 ( .A1(n15403), .A2(n15404), .ZN(n12573) );
  INHSV4 U14504 ( .I(n21765), .ZN(n25950) );
  NAND2HSV4 U14505 ( .A1(n18203), .A2(n18216), .ZN(n12362) );
  CLKNAND2HSV4 U14506 ( .A1(n15899), .A2(n15898), .ZN(n21977) );
  NAND2HSV4 U14507 ( .A1(n12403), .A2(n12402), .ZN(n23454) );
  CLKNAND2HSV2 U14508 ( .A1(n20632), .A2(n20567), .ZN(n12403) );
  NOR2HSV4 U14509 ( .A1(n25660), .A2(n12479), .ZN(n18207) );
  CLKNAND2HSV4 U14510 ( .A1(n15199), .A2(n15198), .ZN(n15332) );
  CLKXOR2HSV4 U14511 ( .A1(n20127), .A2(n20126), .Z(n13127) );
  XOR3HSV2 U14512 ( .A1(n12281), .A2(n19819), .A3(n19818), .Z(\pe9/poht [3])
         );
  XNOR2HSV1 U14513 ( .A1(n19813), .A2(n19812), .ZN(n12281) );
  BUFHSV8 U14514 ( .I(n12729), .Z(n12329) );
  NOR2HSV0 U14515 ( .A1(n17222), .A2(n17221), .ZN(n17228) );
  CLKNHSV0 U14516 ( .I(n13770), .ZN(n12282) );
  OR2HSV2 U14517 ( .A1(n21744), .A2(n12267), .Z(n21748) );
  NAND2HSV2 U14518 ( .A1(n21745), .A2(n21968), .ZN(n15842) );
  XOR2HSV0 U14519 ( .A1(n23954), .A2(n23953), .Z(\pe5/poht [3]) );
  NAND3HSV3 U14520 ( .A1(n15677), .A2(n15676), .A3(n15852), .ZN(n15678) );
  NAND2HSV4 U14521 ( .A1(n23320), .A2(n23319), .ZN(n28927) );
  NAND2HSV2 U14522 ( .A1(n13460), .A2(n13459), .ZN(n13461) );
  MUX2NHSV1 U14523 ( .I0(n13768), .I1(n15007), .S(n23517), .ZN(\pe3/ti_1t ) );
  NOR2HSV0 U14524 ( .A1(n15007), .A2(n26680), .ZN(n15209) );
  NOR2HSV0 U14525 ( .A1(n26241), .A2(n15007), .ZN(n15129) );
  NAND2HSV4 U14526 ( .A1(n15580), .A2(n15579), .ZN(n15853) );
  INHSV4 U14527 ( .I(n15637), .ZN(n15697) );
  CLKNAND2HSV4 U14528 ( .A1(n12441), .A2(n20998), .ZN(n21002) );
  INHSV4 U14529 ( .I(n18090), .ZN(n18184) );
  NAND2HSV4 U14530 ( .A1(n19769), .A2(n19768), .ZN(n22375) );
  INHSV2 U14531 ( .I(n18631), .ZN(n12283) );
  INHSV4 U14532 ( .I(n12283), .ZN(n12284) );
  CLKNAND2HSV2 U14533 ( .A1(n19816), .A2(n19815), .ZN(n23242) );
  NAND2HSV2 U14534 ( .A1(n18222), .A2(n28081), .ZN(n18224) );
  BUFHSV4 U14535 ( .I(n18222), .Z(n18310) );
  NAND3HSV4 U14536 ( .A1(n12656), .A2(n12658), .A3(n12659), .ZN(n18624) );
  NAND3HSV4 U14537 ( .A1(n23243), .A2(n23242), .A3(n19817), .ZN(n28140) );
  NAND2HSV2 U14538 ( .A1(n13673), .A2(n18336), .ZN(n12491) );
  NOR2HSV4 U14539 ( .A1(n18626), .A2(n12284), .ZN(n18627) );
  XOR2HSV0 U14540 ( .A1(n12596), .A2(n12595), .Z(n12285) );
  CLKNAND2HSV4 U14541 ( .A1(n23522), .A2(\pe7/pvq [3]), .ZN(n19184) );
  CLKNAND2HSV4 U14542 ( .A1(n20071), .A2(n20070), .ZN(n13128) );
  CLKNAND2HSV2 U14543 ( .A1(n15573), .A2(n15574), .ZN(n15578) );
  INHSV2 U14544 ( .I(n22631), .ZN(n22632) );
  NAND2HSV0 U14545 ( .A1(n28059), .A2(\pe9/got [11]), .ZN(n18260) );
  BUFHSV4 U14546 ( .I(n18231), .Z(n28059) );
  CLKNAND2HSV2 U14547 ( .A1(n18231), .A2(n18005), .ZN(n18035) );
  INHSV6 U14548 ( .I(n19158), .ZN(n22993) );
  NAND2HSV2 U14549 ( .A1(n22911), .A2(n25371), .ZN(n22912) );
  INHSV0 U14550 ( .I(n15481), .ZN(n12571) );
  NAND2HSV0 U14551 ( .A1(n18144), .A2(n18143), .ZN(n12287) );
  CLKXOR2HSV2 U14552 ( .A1(n25177), .A2(n25176), .Z(n25178) );
  CLKNAND2HSV2 U14553 ( .A1(n19328), .A2(n19327), .ZN(n12288) );
  INHSV4 U14554 ( .I(n17199), .ZN(n17207) );
  INHSV4 U14555 ( .I(n23328), .ZN(n23459) );
  NAND2HSV4 U14556 ( .A1(n16057), .A2(n16016), .ZN(n23328) );
  INAND3HSV2 U14557 ( .A1(n12490), .B1(n12491), .B2(n18468), .ZN(n18337) );
  CLKNAND2HSV2 U14558 ( .A1(n12803), .A2(n12802), .ZN(n12804) );
  OAI21HSV2 U14559 ( .A1(n13493), .A2(n13494), .B(n13495), .ZN(n13496) );
  NAND2HSV2 U14560 ( .A1(n28943), .A2(n14039), .ZN(n28143) );
  NAND2HSV2 U14561 ( .A1(n28943), .A2(n28423), .ZN(n28185) );
  NAND2HSV2 U14562 ( .A1(n28943), .A2(n28227), .ZN(n28228) );
  NAND2HSV2 U14563 ( .A1(n28943), .A2(\pe9/got [8]), .ZN(n28259) );
  INAND2HSV2 U14564 ( .A1(n28431), .B1(n17117), .ZN(n20073) );
  NAND2HSV2 U14565 ( .A1(n28431), .A2(n12371), .ZN(n12370) );
  XOR2HSV4 U14566 ( .A1(n16955), .A2(n16954), .Z(n28431) );
  MUX2NHSV2 U14567 ( .I0(n15974), .I1(n12820), .S(n15975), .ZN(n16106) );
  AOI22HSV2 U14568 ( .A1(n12688), .A2(n12690), .B1(n12689), .B2(n19176), .ZN(
        n12289) );
  INHSV4 U14569 ( .I(n15970), .ZN(n15968) );
  OAI21HSV4 U14570 ( .A1(n15177), .A2(n15239), .B(n15056), .ZN(n15180) );
  NOR2HSV2 U14571 ( .A1(n15178), .A2(n15243), .ZN(n15179) );
  NAND2HSV0 U14572 ( .A1(n23327), .A2(\pe3/got [11]), .ZN(n16103) );
  NOR2HSV2 U14573 ( .A1(n19311), .A2(n19310), .ZN(n19326) );
  OAI21HSV2 U14574 ( .A1(n27214), .A2(n23120), .B(n19215), .ZN(n19382) );
  CLKNAND2HSV2 U14575 ( .A1(n27214), .A2(n19380), .ZN(n19377) );
  INHSV6 U14576 ( .I(n27687), .ZN(n27494) );
  NAND2HSV2 U14577 ( .A1(n27687), .A2(n14046), .ZN(n27689) );
  OAI21HSV4 U14578 ( .A1(n18545), .A2(n28961), .B(n18052), .ZN(n18085) );
  NOR2HSV4 U14579 ( .A1(n18335), .A2(n18334), .ZN(n18439) );
  CLKNAND2HSV2 U14580 ( .A1(n14575), .A2(n14574), .ZN(n14582) );
  NAND2HSV2 U14581 ( .A1(n18396), .A2(n18397), .ZN(n12963) );
  NOR2HSV4 U14582 ( .A1(n18550), .A2(n28343), .ZN(n28346) );
  AOI21HSV4 U14583 ( .A1(n14525), .A2(n14524), .B(n14523), .ZN(n12290) );
  CLKNAND2HSV4 U14584 ( .A1(n20501), .A2(n20502), .ZN(n20503) );
  NAND2HSV2 U14585 ( .A1(n18523), .A2(n18522), .ZN(n18527) );
  CLKNHSV0 U14586 ( .I(n18522), .ZN(n12495) );
  CLKNAND2HSV2 U14587 ( .A1(n17407), .A2(n17406), .ZN(n12756) );
  NAND2HSV4 U14588 ( .A1(n16259), .A2(n17207), .ZN(n17521) );
  CLKNAND2HSV2 U14589 ( .A1(n23483), .A2(n15394), .ZN(n15397) );
  NAND2HSV4 U14590 ( .A1(n15968), .A2(n15967), .ZN(n15972) );
  INHSV4 U14591 ( .I(n15969), .ZN(n15967) );
  CLKNAND2HSV4 U14592 ( .A1(n19616), .A2(n19615), .ZN(n12508) );
  NOR2HSV8 U14593 ( .A1(n19521), .A2(n19520), .ZN(n19616) );
  XOR2HSV4 U14594 ( .A1(n19755), .A2(n19754), .Z(n19763) );
  CLKNHSV6 U14595 ( .I(n27494), .ZN(n27727) );
  NAND2HSV4 U14596 ( .A1(n23229), .A2(n23230), .ZN(n27687) );
  NAND2HSV2 U14597 ( .A1(n19257), .A2(n19258), .ZN(n19261) );
  NOR2HSV2 U14598 ( .A1(n19706), .A2(n12610), .ZN(n12609) );
  CLKNAND2HSV2 U14599 ( .A1(n20191), .A2(n20190), .ZN(n20222) );
  NAND2HSV2 U14600 ( .A1(n14764), .A2(n12632), .ZN(n12631) );
  INHSV2 U14601 ( .I(n14263), .ZN(n13436) );
  NAND2HSV4 U14602 ( .A1(n14273), .A2(n14272), .ZN(n14297) );
  XNOR2HSV4 U14603 ( .A1(n20175), .A2(n20174), .ZN(n12291) );
  CLKNAND2HSV2 U14604 ( .A1(n20178), .A2(n20177), .ZN(n12292) );
  NAND2HSV0 U14605 ( .A1(n20177), .A2(n20178), .ZN(n12293) );
  CLKNAND2HSV2 U14606 ( .A1(n20178), .A2(n20177), .ZN(n20288) );
  INHSV4 U14607 ( .I(n12709), .ZN(n19693) );
  CLKNHSV0 U14608 ( .I(n14495), .ZN(n12294) );
  INHSV6 U14609 ( .I(n22439), .ZN(n22680) );
  NAND3HSV4 U14610 ( .A1(n14391), .A2(n14297), .A3(n18920), .ZN(n14274) );
  CLKNAND2HSV4 U14611 ( .A1(n12497), .A2(n12496), .ZN(n12502) );
  NAND2HSV4 U14612 ( .A1(n15085), .A2(n15084), .ZN(n14041) );
  CLKNHSV4 U14613 ( .I(n12296), .ZN(n12297) );
  NAND2HSV4 U14614 ( .A1(n16787), .A2(n16786), .ZN(n16790) );
  NAND2HSV4 U14615 ( .A1(n16893), .A2(n16892), .ZN(n16955) );
  CLKNAND2HSV4 U14616 ( .A1(n16888), .A2(n16845), .ZN(n16893) );
  CLKNAND2HSV2 U14617 ( .A1(n12459), .A2(n14239), .ZN(n28798) );
  CLKNAND2HSV4 U14618 ( .A1(n14450), .A2(n14449), .ZN(n14452) );
  INHSV4 U14619 ( .I(n15675), .ZN(n15677) );
  NOR2HSV8 U14620 ( .A1(n16742), .A2(n16741), .ZN(n16744) );
  NAND2HSV0 U14621 ( .A1(n22136), .A2(n28420), .ZN(n13895) );
  OAI21HSV2 U14622 ( .A1(n22328), .A2(n22329), .B(n13893), .ZN(n13894) );
  BUFHSV4 U14623 ( .I(n19794), .Z(n12295) );
  CLKNAND2HSV2 U14624 ( .A1(n18443), .A2(n18442), .ZN(n18447) );
  OAI21HSV0 U14625 ( .A1(n18439), .A2(n18469), .B(n18438), .ZN(n18443) );
  CLKNAND2HSV2 U14626 ( .A1(n18322), .A2(n18323), .ZN(n18455) );
  INHSV4 U14627 ( .I(n15281), .ZN(n15279) );
  INHSV4 U14628 ( .I(n25059), .ZN(n12296) );
  INHSV4 U14629 ( .I(n14278), .ZN(n14276) );
  NAND2HSV4 U14630 ( .A1(n27126), .A2(n16170), .ZN(n23440) );
  IOA22HSV4 U14631 ( .B1(n28801), .B2(n23667), .A1(n23664), .A2(n16031), .ZN(
        n23665) );
  XNOR2HSV4 U14632 ( .A1(n23598), .A2(n23597), .ZN(n23599) );
  XNOR2HSV4 U14633 ( .A1(n23596), .A2(n23595), .ZN(n23597) );
  XNOR2HSV4 U14634 ( .A1(n23657), .A2(n23656), .ZN(n23658) );
  INHSV2 U14635 ( .I(n18560), .ZN(n18564) );
  OAI21HSV0 U14636 ( .A1(n18560), .A2(n28016), .B(n18389), .ZN(n18390) );
  NAND2HSV4 U14637 ( .A1(n20395), .A2(n20448), .ZN(n20396) );
  MUX2NHSV2 U14638 ( .I0(n13873), .I1(n21057), .S(n13874), .ZN(n21058) );
  IOA21HSV2 U14639 ( .A1(n21053), .A2(n21052), .B(n21056), .ZN(n13874) );
  BUFHSV2 U14640 ( .I(n24961), .Z(n12298) );
  NOR2HSV4 U14641 ( .A1(n17611), .A2(n23432), .ZN(n17612) );
  INHSV4 U14642 ( .I(n19243), .ZN(n23138) );
  AOI21HSV4 U14643 ( .A1(n19266), .A2(n19265), .B(n19372), .ZN(n19272) );
  CLKNHSV6 U14644 ( .I(n14157), .ZN(n27212) );
  CLKXOR2HSV4 U14645 ( .A1(n20173), .A2(n20172), .Z(n20174) );
  NAND2HSV4 U14646 ( .A1(n17637), .A2(n17636), .ZN(n17654) );
  CLKNAND2HSV2 U14647 ( .A1(n13124), .A2(n13123), .ZN(n13125) );
  INHSV2 U14648 ( .I(n19460), .ZN(n13294) );
  XOR2HSV4 U14649 ( .A1(n19414), .A2(n19413), .Z(n19461) );
  NAND2HSV2 U14650 ( .A1(n17824), .A2(n17825), .ZN(n13714) );
  NAND2HSV2 U14651 ( .A1(n20691), .A2(n20692), .ZN(n12721) );
  AOI21HSV2 U14652 ( .A1(n20631), .A2(n12385), .B(n12382), .ZN(n20616) );
  CLKNHSV0 U14653 ( .I(n15570), .ZN(n23985) );
  CLKNAND2HSV2 U14654 ( .A1(n14054), .A2(n23372), .ZN(n24500) );
  NAND2HSV0 U14655 ( .A1(n24500), .A2(n24499), .ZN(n23375) );
  NAND3HSV4 U14656 ( .A1(n14432), .A2(n14431), .A3(n14401), .ZN(n14402) );
  NAND2HSV2 U14657 ( .A1(n18848), .A2(n18847), .ZN(n18851) );
  CLKNAND2HSV2 U14658 ( .A1(n12740), .A2(n21241), .ZN(n21642) );
  OAI21HSV4 U14659 ( .A1(n19956), .A2(n18773), .B(n18772), .ZN(n18779) );
  NAND2HSV4 U14660 ( .A1(n18779), .A2(n18778), .ZN(n18780) );
  CLKNHSV0 U14661 ( .I(n18615), .ZN(n12299) );
  INHSV2 U14662 ( .I(n12299), .ZN(n12300) );
  NAND2HSV2 U14663 ( .A1(n16616), .A2(n16617), .ZN(n16620) );
  OAI21HSV2 U14664 ( .A1(n13042), .A2(n13043), .B(n13044), .ZN(n26216) );
  CLKXOR2HSV4 U14665 ( .A1(n16984), .A2(n13192), .Z(n13193) );
  NAND2HSV4 U14666 ( .A1(n15972), .A2(n15971), .ZN(n15978) );
  CLKXOR2HSV4 U14667 ( .A1(n24954), .A2(n24953), .Z(n24955) );
  CLKNAND2HSV4 U14668 ( .A1(n14606), .A2(n14605), .ZN(n14642) );
  NAND2HSV4 U14669 ( .A1(n12290), .A2(n14605), .ZN(n24411) );
  INHSV4 U14670 ( .I(n14902), .ZN(n21325) );
  NAND2HSV2 U14671 ( .A1(\pe5/bq[16] ), .A2(\pe5/aot [14]), .ZN(n12426) );
  CLKNAND2HSV4 U14672 ( .A1(n15187), .A2(n15291), .ZN(n28707) );
  CLKBUFHSV2 U14673 ( .I(n12274), .Z(n26854) );
  AOI21HSV4 U14674 ( .A1(n20702), .A2(n25026), .B(n20701), .ZN(n20703) );
  INHSV2 U14675 ( .I(n26929), .ZN(n26928) );
  AOI21HSV4 U14676 ( .A1(n23184), .A2(n23186), .B(n23183), .ZN(n23185) );
  AOI21HSV4 U14677 ( .A1(n19739), .A2(n22091), .B(n19320), .ZN(n19321) );
  CLKNAND2HSV4 U14678 ( .A1(n19619), .A2(n23901), .ZN(n19705) );
  CLKNAND2HSV2 U14679 ( .A1(n23112), .A2(n23111), .ZN(n23113) );
  NOR2HSV2 U14680 ( .A1(n23181), .A2(n12663), .ZN(n23184) );
  NOR2HSV2 U14681 ( .A1(n23427), .A2(n12663), .ZN(n23428) );
  CLKNAND2HSV4 U14682 ( .A1(n20772), .A2(n20771), .ZN(n20761) );
  NAND2HSV4 U14683 ( .A1(n23454), .A2(n20635), .ZN(n20771) );
  NAND2HSV4 U14684 ( .A1(n25055), .A2(n25053), .ZN(n28936) );
  NAND3HSV2 U14685 ( .A1(n21222), .A2(n21223), .A3(n21221), .ZN(n21866) );
  CLKNAND2HSV8 U14686 ( .A1(n12510), .A2(n12405), .ZN(n25529) );
  XNOR2HSV4 U14687 ( .A1(n18689), .A2(n18688), .ZN(n18693) );
  CLKXOR2HSV4 U14688 ( .A1(n19172), .A2(n19171), .Z(n19173) );
  NAND2HSV2 U14689 ( .A1(n28936), .A2(\pe11/got [3]), .ZN(n12617) );
  NAND3HSV4 U14690 ( .A1(n16463), .A2(n16462), .A3(n16461), .ZN(n28799) );
  INAND2HSV4 U14691 ( .A1(n16308), .B1(n21330), .ZN(n16462) );
  AOI21HSV4 U14692 ( .A1(n16053), .A2(n16045), .B(n16044), .ZN(n16046) );
  CLKXOR2HSV4 U14693 ( .A1(n26641), .A2(n26640), .Z(n26644) );
  NAND2HSV2 U14694 ( .A1(n25054), .A2(n25504), .ZN(n25050) );
  NAND2HSV4 U14695 ( .A1(n27284), .A2(n27283), .ZN(n27640) );
  NAND2HSV2 U14696 ( .A1(n13670), .A2(n13669), .ZN(n13671) );
  AOI21HSV2 U14697 ( .A1(n23407), .A2(n23406), .B(n23405), .ZN(n12301) );
  NAND2HSV2 U14698 ( .A1(n13744), .A2(n13743), .ZN(n13745) );
  AOI22HSV2 U14699 ( .A1(n28967), .A2(n27354), .B1(\pe2/ti_7t [14]), .B2(
        n27571), .ZN(n12302) );
  INHSV2 U14700 ( .I(n16310), .ZN(n13746) );
  CLKNAND2HSV4 U14701 ( .A1(n16356), .A2(n16355), .ZN(n16454) );
  INAND2HSV4 U14702 ( .A1(n19708), .B1(n13657), .ZN(n25345) );
  CLKNAND2HSV2 U14703 ( .A1(n20776), .A2(n20698), .ZN(n20781) );
  CLKXOR2HSV4 U14704 ( .A1(n24878), .A2(n24877), .Z(n24879) );
  BUFHSV8 U14705 ( .I(n18690), .Z(n18828) );
  CLKXOR2HSV2 U14706 ( .A1(n24919), .A2(n24918), .Z(n24920) );
  OAI21HSV4 U14707 ( .A1(n15412), .A2(n12573), .B(n15411), .ZN(n28923) );
  NAND2HSV2 U14708 ( .A1(n15481), .A2(n15487), .ZN(n15412) );
  NOR2HSV4 U14709 ( .A1(n21991), .A2(n21990), .ZN(n22046) );
  MUX2NHSV4 U14710 ( .I0(n16744), .I1(n13656), .S(n16743), .ZN(n12303) );
  INHSV2 U14711 ( .I(n22718), .ZN(n12304) );
  MUX2NHSV1 U14712 ( .I0(n16744), .I1(n13656), .S(n16743), .ZN(n16803) );
  INHSV2 U14713 ( .I(n19620), .ZN(n19619) );
  NAND2HSV0 U14714 ( .A1(n19620), .A2(n25339), .ZN(n19682) );
  MUX2NHSV2 U14715 ( .I0(n19612), .I1(n12852), .S(n19611), .ZN(n19620) );
  NOR2HSV2 U14716 ( .A1(n14910), .A2(n14763), .ZN(n14825) );
  CLKXOR2HSV2 U14717 ( .A1(n21959), .A2(n21958), .Z(n21960) );
  XOR2HSV4 U14718 ( .A1(n21808), .A2(n21807), .Z(n21809) );
  CLKNAND2HSV2 U14719 ( .A1(n28973), .A2(n21422), .ZN(n21522) );
  CLKNAND2HSV2 U14720 ( .A1(n28973), .A2(n24634), .ZN(n21337) );
  MUX2NHSV4 U14721 ( .I0(n20865), .I1(n13413), .S(n13414), .ZN(n28973) );
  XNOR2HSV4 U14722 ( .A1(n12306), .A2(n12305), .ZN(n13817) );
  XNOR2HSV4 U14723 ( .A1(n12308), .A2(n12307), .ZN(n12306) );
  XOR2HSV2 U14724 ( .A1(n23308), .A2(n23307), .Z(n12307) );
  XNOR2HSV4 U14725 ( .A1(n20926), .A2(n20925), .ZN(n12309) );
  CLKNHSV2 U14726 ( .I(n20587), .ZN(n12310) );
  MUX2NHSV1 U14727 ( .I0(n20150), .I1(n12312), .S(n20613), .ZN(n12311) );
  NOR2HSV0 U14728 ( .A1(n12477), .A2(n20151), .ZN(n12312) );
  CLKNHSV2 U14729 ( .I(n20153), .ZN(n20154) );
  CLKNAND2HSV2 U14730 ( .A1(n16999), .A2(n16998), .ZN(n12313) );
  XNOR2HSV4 U14731 ( .A1(n12314), .A2(n19125), .ZN(n19044) );
  CLKNAND2HSV1 U14732 ( .A1(n28938), .A2(n25420), .ZN(n19125) );
  NAND2HSV3 U14733 ( .A1(n18210), .A2(n12316), .ZN(n12317) );
  CLKNAND2HSV3 U14734 ( .A1(n12318), .A2(n12317), .ZN(n12323) );
  CLKNAND2HSV3 U14735 ( .A1(n18204), .A2(n12324), .ZN(n12318) );
  NAND3HSV4 U14736 ( .A1(n12322), .A2(n12321), .A3(n12320), .ZN(n12319) );
  CLKNHSV2 U14737 ( .I(n18205), .ZN(n12320) );
  NAND3HSV4 U14738 ( .A1(n12327), .A2(n12325), .A3(n12326), .ZN(n12322) );
  NOR2HSV4 U14739 ( .A1(n12363), .A2(n12362), .ZN(n18335) );
  CLKNHSV2 U14740 ( .I(n12328), .ZN(n12324) );
  CLKNHSV2 U14741 ( .I(n12453), .ZN(n12325) );
  NOR2HSV4 U14742 ( .A1(n18204), .A2(n12328), .ZN(n12326) );
  CLKNHSV2 U14743 ( .I(n18330), .ZN(n12328) );
  XNOR2HSV4 U14744 ( .A1(n12455), .A2(n12454), .ZN(n18280) );
  CLKNAND2HSV4 U14745 ( .A1(n12332), .A2(n12330), .ZN(n12729) );
  OAI21HSV4 U14746 ( .A1(n12331), .A2(n12730), .B(n12335), .ZN(n12330) );
  CLKNAND2HSV2 U14747 ( .A1(n12334), .A2(n12333), .ZN(n12332) );
  CLKNHSV2 U14748 ( .I(n12331), .ZN(n12333) );
  NOR2HSV4 U14749 ( .A1(n12335), .A2(n12730), .ZN(n12334) );
  CLKNHSV2 U14750 ( .I(n12729), .ZN(n12750) );
  CLKNAND2HSV4 U14751 ( .A1(n17293), .A2(n14056), .ZN(n12335) );
  AOI22HSV4 U14752 ( .A1(n24634), .A2(n14865), .B1(pov5[9]), .B2(n21347), .ZN(
        n14922) );
  XNOR2HSV4 U14753 ( .A1(n14864), .A2(n14863), .ZN(pov5[9]) );
  NAND3HSV1 U14754 ( .A1(n15479), .A2(n15478), .A3(n12337), .ZN(n12336) );
  CLKNHSV2 U14755 ( .I(n15476), .ZN(n12337) );
  NOR2HSV4 U14756 ( .A1(n15472), .A2(n15474), .ZN(n12338) );
  XNOR2HSV4 U14757 ( .A1(n12341), .A2(n12573), .ZN(n28974) );
  CLKNHSV2 U14758 ( .I(n15481), .ZN(n12341) );
  XNOR2HSV4 U14759 ( .A1(n18610), .A2(n12342), .ZN(n18634) );
  XOR2HSV2 U14760 ( .A1(n12343), .A2(n18609), .Z(n12342) );
  NOR2HSV4 U14761 ( .A1(n18560), .A2(n12344), .ZN(n12343) );
  CLKNHSV2 U14762 ( .I(n28137), .ZN(n12344) );
  CLKNAND2HSV2 U14763 ( .A1(n28959), .A2(n16995), .ZN(n16847) );
  CLKNHSV2 U14764 ( .I(n16807), .ZN(n12345) );
  NOR2HSV4 U14765 ( .A1(n28959), .A2(n16808), .ZN(n16788) );
  XNOR2HSV4 U14766 ( .A1(n16754), .A2(n16753), .ZN(n28959) );
  CLKNHSV4 U14767 ( .I(n18645), .ZN(n23717) );
  CLKNAND2HSV4 U14768 ( .A1(n12347), .A2(n12346), .ZN(n18645) );
  NAND3HSV3 U14769 ( .A1(n25681), .A2(n25683), .A3(n18544), .ZN(n12346) );
  CLKNAND2HSV3 U14770 ( .A1(n12349), .A2(n12348), .ZN(n12347) );
  AOI21HSV4 U14771 ( .A1(n28705), .A2(n13988), .B(n18540), .ZN(n12348) );
  CLKNAND2HSV4 U14772 ( .A1(n25683), .A2(n18538), .ZN(n12349) );
  CLKNAND2HSV3 U14773 ( .A1(n18542), .A2(n18463), .ZN(n25681) );
  NOR2HSV4 U14774 ( .A1(n16877), .A2(n12350), .ZN(n16879) );
  CLKNHSV2 U14775 ( .I(n16876), .ZN(n12350) );
  XNOR2HSV4 U14776 ( .A1(n12351), .A2(n16875), .ZN(n16877) );
  CLKNHSV2 U14777 ( .I(n16874), .ZN(n12351) );
  XNOR2HSV4 U14778 ( .A1(n12358), .A2(n12352), .ZN(n19228) );
  XNOR2HSV4 U14779 ( .A1(n12355), .A2(n12353), .ZN(n12352) );
  XNOR2HSV4 U14780 ( .A1(n12354), .A2(\pe7/phq [5]), .ZN(n12353) );
  CLKNAND2HSV2 U14781 ( .A1(\pe7/aot [15]), .A2(\pe7/bq[13] ), .ZN(n12354) );
  XNOR2HSV4 U14782 ( .A1(n12357), .A2(n12356), .ZN(n12355) );
  CLKNAND2HSV2 U14783 ( .A1(n25273), .A2(\pe7/aot [12]), .ZN(n12356) );
  CLKNAND2HSV2 U14784 ( .A1(n27104), .A2(\pe7/pvq [5]), .ZN(n12357) );
  XNOR2HSV4 U14785 ( .A1(n19223), .A2(n12359), .ZN(n12358) );
  XNOR2HSV4 U14786 ( .A1(n19225), .A2(n12360), .ZN(n12359) );
  CLKNHSV3 U14787 ( .I(n18280), .ZN(n18336) );
  OAI21HSV2 U14788 ( .A1(n18335), .A2(n18334), .B(n13672), .ZN(n13673) );
  INHSV2 U14789 ( .I(n18274), .ZN(n12361) );
  CLKNHSV1 U14790 ( .I(n16816), .ZN(n16907) );
  CLKNAND2HSV3 U14791 ( .A1(n12366), .A2(n12365), .ZN(n16942) );
  AOI21HSV4 U14792 ( .A1(n12705), .A2(n16890), .B(n16889), .ZN(n12365) );
  CLKNAND2HSV2 U14793 ( .A1(n16894), .A2(n16955), .ZN(n12366) );
  CLKNHSV2 U14794 ( .I(n12368), .ZN(n12367) );
  CLKNAND2HSV2 U14795 ( .A1(n16942), .A2(n17120), .ZN(n12368) );
  CLKNHSV4 U14796 ( .I(n17067), .ZN(n12371) );
  CLKNAND2HSV2 U14797 ( .A1(n12374), .A2(n12372), .ZN(n17010) );
  CLKNAND2HSV2 U14798 ( .A1(n12373), .A2(n28431), .ZN(n12372) );
  CLKNHSV2 U14799 ( .I(n17005), .ZN(n12373) );
  CLKNAND2HSV2 U14800 ( .A1(n17004), .A2(n12744), .ZN(n12374) );
  NAND3HSV2 U14801 ( .A1(n12376), .A2(n15493), .A3(n12375), .ZN(n27228) );
  INHSV2 U14802 ( .I(n13982), .ZN(n12375) );
  CLKNHSV4 U14803 ( .I(n15492), .ZN(n12376) );
  CLKNHSV4 U14804 ( .I(n15479), .ZN(n15490) );
  CLKNAND2HSV3 U14805 ( .A1(n21343), .A2(n21342), .ZN(n12378) );
  CLKNAND2HSV2 U14806 ( .A1(n12378), .A2(n21715), .ZN(n21717) );
  CLKNHSV2 U14807 ( .I(n12380), .ZN(n16997) );
  CLKNHSV2 U14808 ( .I(n12381), .ZN(n12379) );
  CLKNAND2HSV2 U14809 ( .A1(n12380), .A2(n21738), .ZN(n21739) );
  CLKNHSV2 U14810 ( .I(n17120), .ZN(n12381) );
  CLKNHSV2 U14811 ( .I(n23451), .ZN(n20566) );
  CLKNHSV2 U14812 ( .I(n20631), .ZN(n20567) );
  CLKNAND2HSV2 U14813 ( .A1(n12383), .A2(n23436), .ZN(n12382) );
  CLKNAND2HSV2 U14814 ( .A1(n23451), .A2(n12384), .ZN(n12383) );
  CLKNHSV2 U14815 ( .I(n25488), .ZN(n12384) );
  NOR2HSV4 U14816 ( .A1(n23451), .A2(n12386), .ZN(n12385) );
  CLKNHSV2 U14817 ( .I(n20565), .ZN(n12386) );
  CLKNAND2HSV2 U14818 ( .A1(n20564), .A2(n20563), .ZN(n23451) );
  XNOR2HSV4 U14819 ( .A1(n20558), .A2(n20557), .ZN(n20631) );
  CLKNHSV0 U14820 ( .I(n22714), .ZN(n22713) );
  OAI21HSV2 U14821 ( .A1(n12390), .A2(n12389), .B(n12388), .ZN(n12387) );
  CLKNAND2HSV3 U14822 ( .A1(n12390), .A2(n12389), .ZN(n12388) );
  XNOR2HSV2 U14823 ( .A1(n22710), .A2(n22711), .ZN(n12389) );
  NOR2HSV3 U14824 ( .A1(n12304), .A2(n24453), .ZN(n12390) );
  INHSV2 U14825 ( .I(n13390), .ZN(n12391) );
  CLKNAND2HSV4 U14826 ( .A1(n28996), .A2(n22418), .ZN(n12392) );
  INHSV24 U14827 ( .I(\pe8/phq [1]), .ZN(n12393) );
  NAND3HSV4 U14828 ( .A1(\pe8/phq [1]), .A2(\pe8/ti_1 ), .A3(\pe8/got [16]), 
        .ZN(n12394) );
  IOA21HSV4 U14829 ( .A1(\pe8/ti_1 ), .A2(\pe8/got [16]), .B(n12393), .ZN(
        n12395) );
  CLKNHSV2 U14830 ( .I(n22506), .ZN(n12396) );
  XNOR2HSV4 U14831 ( .A1(n12398), .A2(n12397), .ZN(n22506) );
  XNOR2HSV4 U14832 ( .A1(n22437), .A2(n22438), .ZN(n12398) );
  NOR2HSV4 U14833 ( .A1(n21420), .A2(n12400), .ZN(n12399) );
  CLKNAND2HSV2 U14834 ( .A1(n21418), .A2(n21417), .ZN(n12400) );
  CLKNAND2HSV1 U14835 ( .A1(n20771), .A2(n20772), .ZN(n20773) );
  OAI21HSV2 U14836 ( .A1(n23452), .A2(n12401), .B(n20633), .ZN(n20772) );
  AOI21HSV2 U14837 ( .A1(n20631), .A2(n20778), .B(n20627), .ZN(n12401) );
  CLKNAND2HSV0 U14838 ( .A1(n20628), .A2(n20631), .ZN(n12402) );
  BUFHSV8 U14839 ( .I(n25529), .Z(n12404) );
  CLKNAND2HSV3 U14840 ( .A1(n12406), .A2(n12407), .ZN(n12405) );
  INHSV2 U14841 ( .I(n12515), .ZN(n12406) );
  CLKNAND2HSV0 U14842 ( .A1(n12404), .A2(\pe8/got [12]), .ZN(n18689) );
  CLKNHSV2 U14843 ( .I(n12513), .ZN(n12407) );
  NOR2HSV8 U14844 ( .A1(n16023), .A2(n15960), .ZN(n15962) );
  NOR2HSV8 U14845 ( .A1(n12408), .A2(n15236), .ZN(n16023) );
  XNOR2HSV4 U14846 ( .A1(n15332), .A2(n15331), .ZN(n12408) );
  XNOR2HSV4 U14847 ( .A1(n15235), .A2(n15234), .ZN(n15331) );
  XNOR2HSV4 U14848 ( .A1(n12415), .A2(n12409), .ZN(n18908) );
  XNOR2HSV4 U14849 ( .A1(n12411), .A2(n12410), .ZN(n12409) );
  NAND3HSV1 U14850 ( .A1(n14431), .A2(n14432), .A3(n13526), .ZN(n12410) );
  XOR3HSV2 U14851 ( .A1(n14430), .A2(n12413), .A3(n12412), .Z(n12411) );
  CLKNAND2HSV2 U14852 ( .A1(n26033), .A2(n14236), .ZN(n12412) );
  NOR2HSV4 U14853 ( .A1(n12185), .A2(n12414), .ZN(n12413) );
  CLKNHSV2 U14854 ( .I(n28593), .ZN(n12414) );
  OAI21HSV4 U14855 ( .A1(n28676), .A2(n19142), .B(n14410), .ZN(n12415) );
  XNOR2HSV4 U14856 ( .A1(n14409), .A2(n14408), .ZN(n28676) );
  XNOR2HSV4 U14857 ( .A1(n14366), .A2(n14365), .ZN(n14408) );
  AOI21HSV4 U14858 ( .A1(n12655), .A2(n19069), .B(n13792), .ZN(n14409) );
  AOI21HSV4 U14859 ( .A1(n16901), .A2(n12416), .B(n16771), .ZN(n16772) );
  CLKNHSV2 U14860 ( .I(n12417), .ZN(n12416) );
  XNOR2HSV4 U14861 ( .A1(n16660), .A2(n12417), .ZN(n16661) );
  CLKNAND2HSV2 U14862 ( .A1(n16897), .A2(\pe10/aot [14]), .ZN(n12417) );
  CLKNHSV2 U14863 ( .I(n16795), .ZN(n12418) );
  NAND3HSV4 U14864 ( .A1(n12419), .A2(n16680), .A3(n16679), .ZN(n16648) );
  XNOR2HSV4 U14865 ( .A1(n23650), .A2(n12420), .ZN(n23652) );
  XOR2HSV2 U14866 ( .A1(n23649), .A2(n12421), .Z(n12420) );
  XNOR2HSV4 U14867 ( .A1(n23648), .A2(n12422), .ZN(n12421) );
  XNOR2HSV4 U14868 ( .A1(n12424), .A2(n12423), .ZN(n12422) );
  XOR2HSV2 U14869 ( .A1(n23647), .A2(n23645), .Z(n12423) );
  CLKNHSV2 U14870 ( .I(n23646), .ZN(n12424) );
  OAI21HSV2 U14871 ( .A1(n25644), .A2(\pe5/got [15]), .B(n14815), .ZN(n14486)
         );
  XNOR2HSV4 U14872 ( .A1(n14471), .A2(n14470), .ZN(n25644) );
  XNOR2HSV4 U14873 ( .A1(n14835), .A2(n12425), .ZN(n14470) );
  CLKNHSV2 U14874 ( .I(n12426), .ZN(n12425) );
  XNOR2HSV4 U14875 ( .A1(n12428), .A2(n12427), .ZN(n14471) );
  OAI21HSV4 U14876 ( .A1(\pe5/phq [3]), .A2(n14468), .B(n14467), .ZN(n12427)
         );
  XNOR2HSV4 U14877 ( .A1(n14464), .A2(n14465), .ZN(n12428) );
  CLKNAND2HSV3 U14878 ( .A1(n12429), .A2(n18856), .ZN(n28940) );
  CLKNAND2HSV2 U14879 ( .A1(n14696), .A2(n18927), .ZN(n12429) );
  XNOR2HSV4 U14880 ( .A1(n14409), .A2(n14408), .ZN(n14696) );
  CLKNHSV4 U14881 ( .I(n18908), .ZN(n12430) );
  INHSV2 U14882 ( .I(n12431), .ZN(n12432) );
  CLKNHSV2 U14883 ( .I(n18908), .ZN(n12431) );
  CLKNAND2HSV2 U14884 ( .A1(n12433), .A2(n14049), .ZN(n24801) );
  CLKNAND2HSV2 U14885 ( .A1(n12433), .A2(\pe11/got [4]), .ZN(n21805) );
  CLKNAND2HSV2 U14886 ( .A1(n12433), .A2(\pe11/got [11]), .ZN(n21958) );
  CLKNAND2HSV2 U14887 ( .A1(n12433), .A2(\pe11/got [9]), .ZN(n24846) );
  CLKNAND2HSV2 U14888 ( .A1(n12433), .A2(\pe11/got [5]), .ZN(n24875) );
  CLKNAND2HSV2 U14889 ( .A1(n12433), .A2(\pe11/got [8]), .ZN(n25176) );
  CLKNAND2HSV2 U14890 ( .A1(n12433), .A2(\pe11/got [2]), .ZN(n12670) );
  CLKNAND2HSV4 U14891 ( .A1(n20774), .A2(n20761), .ZN(n12434) );
  INHSV2 U14892 ( .I(n14109), .ZN(n12435) );
  NAND3HSV4 U14893 ( .A1(n12437), .A2(n12436), .A3(\pe6/pvq [2]), .ZN(n12440)
         );
  CLKNHSV2 U14894 ( .I(n14108), .ZN(n12436) );
  INHSV2 U14895 ( .I(\pe6/ctrq ), .ZN(n14047) );
  CLKNAND2HSV2 U14896 ( .A1(\pe6/aot [15]), .A2(\pe6/bq[16] ), .ZN(n14109) );
  CLKNAND2HSV2 U14897 ( .A1(n12439), .A2(n14108), .ZN(n12438) );
  CLKNAND2HSV2 U14898 ( .A1(\pe6/ctrq ), .A2(\pe6/pvq [2]), .ZN(n12439) );
  XNOR2HSV4 U14899 ( .A1(n12442), .A2(n21336), .ZN(n20999) );
  CLKNHSV2 U14900 ( .I(n20997), .ZN(n12442) );
  AOI21HSV4 U14901 ( .A1(n12448), .A2(n12449), .B(n12443), .ZN(n12446) );
  CLKNHSV2 U14902 ( .I(n25049), .ZN(n12443) );
  CLKNAND2HSV2 U14903 ( .A1(n25044), .A2(n25043), .ZN(n12445) );
  CLKNHSV2 U14904 ( .I(n25039), .ZN(n12448) );
  CLKNHSV2 U14905 ( .I(n25038), .ZN(n12449) );
  CLKNHSV2 U14906 ( .I(n25036), .ZN(n12450) );
  CLKNHSV2 U14907 ( .I(n25037), .ZN(n12451) );
  CLKNHSV2 U14908 ( .I(n18202), .ZN(n12453) );
  XNOR2HSV4 U14909 ( .A1(n18140), .A2(n18139), .ZN(n12454) );
  NOR2HSV4 U14910 ( .A1(n18102), .A2(n18103), .ZN(n12455) );
  CLKNAND2HSV0 U14911 ( .A1(n12456), .A2(n15285), .ZN(n15095) );
  AOI31HSV2 U14912 ( .A1(n23481), .A2(n12456), .A3(n15973), .B(n15096), .ZN(
        n15054) );
  CLKNAND2HSV4 U14913 ( .A1(n14179), .A2(n12457), .ZN(n14239) );
  CLKNHSV3 U14914 ( .I(n12458), .ZN(n12457) );
  CLKNAND2HSV1 U14915 ( .A1(n14178), .A2(n18920), .ZN(n12458) );
  CLKNHSV2 U14916 ( .I(n14117), .ZN(n14179) );
  CLKNAND2HSV4 U14917 ( .A1(n14116), .A2(n14148), .ZN(n14231) );
  CLKNHSV2 U14918 ( .I(n12461), .ZN(n12460) );
  CLKNHSV4 U14919 ( .I(n18212), .ZN(n12461) );
  CLKNHSV1 U14920 ( .I(n18220), .ZN(n12462) );
  XNOR2HSV4 U14921 ( .A1(n12463), .A2(n21157), .ZN(n21160) );
  XNOR2HSV4 U14922 ( .A1(n21158), .A2(n12464), .ZN(n12463) );
  CLKNHSV2 U14923 ( .I(n21155), .ZN(n12464) );
  XNOR2HSV4 U14924 ( .A1(n12466), .A2(n12465), .ZN(n21155) );
  CLKNAND2HSV2 U14925 ( .A1(n27524), .A2(n27544), .ZN(n12465) );
  XOR2HSV2 U14926 ( .A1(n21142), .A2(n12467), .Z(n12466) );
  CLKNHSV2 U14927 ( .I(n21143), .ZN(n12467) );
  INHSV2 U14928 ( .I(n12468), .ZN(n20186) );
  CLKNAND2HSV2 U14929 ( .A1(n12469), .A2(n20227), .ZN(n20245) );
  CLKNAND2HSV2 U14930 ( .A1(n12469), .A2(\pe11/got [9]), .ZN(n20406) );
  CLKNHSV2 U14931 ( .I(n20186), .ZN(n12469) );
  CLKNAND2HSV2 U14932 ( .A1(n12292), .A2(n20180), .ZN(n12468) );
  XNOR2HSV4 U14933 ( .A1(n14620), .A2(n24411), .ZN(n12470) );
  CLKNAND2HSV2 U14934 ( .A1(n14681), .A2(n14680), .ZN(n12471) );
  CLKNHSV2 U14935 ( .I(n15074), .ZN(n15077) );
  XNOR2HSV4 U14936 ( .A1(n12473), .A2(n12472), .ZN(n15074) );
  CLKNAND2HSV2 U14937 ( .A1(n15118), .A2(n28930), .ZN(n12472) );
  CLKNAND2HSV2 U14938 ( .A1(n15061), .A2(n13977), .ZN(n15118) );
  XNOR2HSV4 U14939 ( .A1(n12475), .A2(n12474), .ZN(n12473) );
  XNOR2HSV4 U14940 ( .A1(n15070), .A2(n15072), .ZN(n12474) );
  XNOR2HSV4 U14941 ( .A1(n15073), .A2(n15071), .ZN(n12475) );
  XNOR2HSV4 U14942 ( .A1(n21462), .A2(n12476), .ZN(n21571) );
  XNOR2HSV4 U14943 ( .A1(n21462), .A2(n12476), .ZN(n21966) );
  CLKNHSV2 U14944 ( .I(n20151), .ZN(n20587) );
  CLKNHSV4 U14945 ( .I(\pe11/phq [3]), .ZN(n12477) );
  CLKNHSV2 U14946 ( .I(n12479), .ZN(n12478) );
  XOR2HSV2 U14947 ( .A1(n25660), .A2(n12479), .Z(n25661) );
  CLKNAND2HSV3 U14948 ( .A1(n18714), .A2(n12480), .ZN(n12481) );
  CLKNHSV2 U14949 ( .I(n18715), .ZN(n12480) );
  CLKNAND2HSV2 U14950 ( .A1(n12481), .A2(n28599), .ZN(n18759) );
  CLKNHSV2 U14951 ( .I(n15919), .ZN(n15240) );
  MUX2NHSV2 U14952 ( .I0(n29036), .I1(\pe3/ti_7t [5]), .S(n21313), .ZN(n15244)
         );
  OAI22HSV4 U14953 ( .A1(n15919), .A2(n12486), .B1(n12483), .B2(n12482), .ZN(
        n29036) );
  CLKNHSV2 U14954 ( .I(n15243), .ZN(n12482) );
  NOR2HSV4 U14955 ( .A1(n12485), .A2(n12484), .ZN(n12483) );
  CLKNHSV2 U14956 ( .I(n15242), .ZN(n12484) );
  CLKNHSV2 U14957 ( .I(n15241), .ZN(n12485) );
  CLKNAND2HSV2 U14958 ( .A1(n15239), .A2(n26413), .ZN(n12486) );
  CLKNAND2HSV3 U14959 ( .A1(n28964), .A2(n18454), .ZN(n12487) );
  CLKNAND2HSV4 U14960 ( .A1(n18272), .A2(n18271), .ZN(n28964) );
  CLKNAND2HSV0 U14961 ( .A1(n28795), .A2(n18005), .ZN(n18615) );
  CLKNAND2HSV4 U14962 ( .A1(n12487), .A2(n18273), .ZN(n28795) );
  CLKNAND2HSV2 U14963 ( .A1(n28436), .A2(\pe5/got [2]), .ZN(n27111) );
  CLKNAND2HSV2 U14964 ( .A1(n28436), .A2(\pe5/got [3]), .ZN(n23239) );
  CLKNHSV2 U14965 ( .I(n18467), .ZN(pov9[9]) );
  CLKNAND2HSV2 U14966 ( .A1(n18444), .A2(pov9[9]), .ZN(n18451) );
  CLKNAND2HSV4 U14967 ( .A1(n16842), .A2(n20142), .ZN(n12492) );
  CLKNAND2HSV1 U14968 ( .A1(n18525), .A2(n12493), .ZN(n18526) );
  NOR2HSV2 U14969 ( .A1(n18522), .A2(n12494), .ZN(n12493) );
  INHSV2 U14970 ( .I(n18558), .ZN(n12494) );
  AOI21HSV4 U14971 ( .A1(n12495), .A2(n18525), .B(n18457), .ZN(n18458) );
  NAND2HSV2 U14972 ( .A1(n28964), .A2(n18454), .ZN(n18522) );
  INHSV2 U14973 ( .I(n12506), .ZN(n12498) );
  NOR2HSV8 U14974 ( .A1(n12500), .A2(n12499), .ZN(n12501) );
  CLKNAND2HSV4 U14975 ( .A1(n14931), .A2(n14628), .ZN(n12499) );
  CLKXOR2HSV4 U14976 ( .A1(n14618), .A2(n14629), .Z(n12500) );
  NOR2HSV8 U14977 ( .A1(n12502), .A2(n12501), .ZN(n14760) );
  NAND3HSV4 U14978 ( .A1(n14760), .A2(n14759), .A3(n14758), .ZN(n14905) );
  NAND3HSV4 U14979 ( .A1(n12503), .A2(n25659), .A3(n14628), .ZN(n14758) );
  XNOR2HSV4 U14980 ( .A1(n12504), .A2(n14629), .ZN(n12503) );
  NOR2HSV4 U14981 ( .A1(n25658), .A2(n14627), .ZN(n12505) );
  CLKNHSV2 U14982 ( .I(n13967), .ZN(n12506) );
  CLKNHSV2 U14983 ( .I(\pe11/got [16]), .ZN(n20179) );
  CLKNAND2HSV2 U14984 ( .A1(n12507), .A2(n22797), .ZN(n22798) );
  MUX2NHSV4 U14985 ( .I0(n22046), .I1(n22903), .S(n22904), .ZN(n26929) );
  INHSV2 U14986 ( .I(n12508), .ZN(n12613) );
  NAND3HSV4 U14987 ( .A1(n12509), .A2(n19705), .A3(n19702), .ZN(n19677) );
  CLKNHSV2 U14988 ( .I(n12613), .ZN(n12509) );
  CLKNHSV3 U14989 ( .I(n12514), .ZN(n12512) );
  CLKNAND2HSV2 U14990 ( .A1(n16458), .A2(n16459), .ZN(n12514) );
  CLKNAND2HSV4 U14991 ( .A1(n12515), .A2(n12514), .ZN(n28984) );
  CLKNAND2HSV3 U14992 ( .A1(n16456), .A2(n16457), .ZN(n12515) );
  AOI21HSV4 U14993 ( .A1(n12512), .A2(n19830), .B(n12511), .ZN(n12510) );
  CLKNHSV2 U14994 ( .I(n16556), .ZN(n12511) );
  CLKNHSV2 U14995 ( .I(n19830), .ZN(n12513) );
  OAI21HSV4 U14996 ( .A1(n29021), .A2(n14281), .B(n18998), .ZN(n19042) );
  CLKNAND2HSV4 U14997 ( .A1(n28969), .A2(n21342), .ZN(n21339) );
  CLKNHSV2 U14998 ( .I(n12516), .ZN(n12622) );
  CLKNAND2HSV2 U14999 ( .A1(n12516), .A2(n12523), .ZN(n23476) );
  CLKNAND2HSV2 U15000 ( .A1(n16707), .A2(n16706), .ZN(n12516) );
  BUFHSV8 U15001 ( .I(n21718), .Z(n12517) );
  XNOR2HSV4 U15002 ( .A1(n12522), .A2(n12518), .ZN(n21519) );
  XNOR2HSV4 U15003 ( .A1(n12520), .A2(n12519), .ZN(n12518) );
  CLKNAND2HSV2 U15004 ( .A1(n12517), .A2(n24635), .ZN(n12519) );
  XNOR2HSV4 U15005 ( .A1(n21518), .A2(n12521), .ZN(n12520) );
  XOR2HSV2 U15006 ( .A1(n21517), .A2(n21516), .Z(n12521) );
  CLKNAND2HSV2 U15007 ( .A1(n24377), .A2(\pe5/got [15]), .ZN(n12522) );
  CLKNAND2HSV2 U15008 ( .A1(n12523), .A2(n12623), .ZN(n12621) );
  NAND2HSV2 U15009 ( .A1(n16704), .A2(n16705), .ZN(n12523) );
  CLKNAND2HSV4 U15010 ( .A1(n12525), .A2(n12524), .ZN(n16781) );
  NOR2HSV4 U15011 ( .A1(n16668), .A2(n16667), .ZN(n12525) );
  OAI21HSV2 U15012 ( .A1(n16672), .A2(n16671), .B(n23484), .ZN(n12524) );
  XNOR2HSV4 U15013 ( .A1(n12526), .A2(n16345), .ZN(n16346) );
  XNOR2HSV4 U15014 ( .A1(n12528), .A2(n12527), .ZN(n12526) );
  XNOR2HSV4 U15015 ( .A1(n12529), .A2(n19921), .ZN(n12527) );
  XNOR2HSV4 U15016 ( .A1(n12531), .A2(n12530), .ZN(n12528) );
  CLKNAND2HSV2 U15017 ( .A1(n28641), .A2(n23627), .ZN(n19921) );
  MUX2NHSV2 U15018 ( .I0(\pe8/phq [4]), .I1(n13437), .S(n13438), .ZN(n12529)
         );
  CLKNHSV2 U15019 ( .I(n16530), .ZN(n28788) );
  INAND2HSV4 U15020 ( .A1(n16530), .B1(n16418), .ZN(n12854) );
  INAND2HSV4 U15021 ( .A1(n16530), .B1(\pe8/got [13]), .ZN(n16382) );
  CLKNAND2HSV3 U15022 ( .A1(n28945), .A2(n15086), .ZN(n12538) );
  CLKNAND2HSV3 U15023 ( .A1(n16108), .A2(n16107), .ZN(n28945) );
  CLKNAND2HSV3 U15024 ( .A1(n16053), .A2(n12539), .ZN(n16110) );
  MUX2NHSV4 U15025 ( .I0(n16052), .I1(n16038), .S(n28708), .ZN(n16053) );
  CLKNAND2HSV3 U15026 ( .A1(n16037), .A2(n16036), .ZN(n16049) );
  XNOR2HSV4 U15027 ( .A1(n12535), .A2(n12532), .ZN(n21732) );
  CLKNAND2HSV2 U15028 ( .A1(n12534), .A2(n12533), .ZN(n12532) );
  CLKNHSV2 U15029 ( .I(n23402), .ZN(n12533) );
  CLKNAND2HSV2 U15030 ( .A1(n16111), .A2(n16110), .ZN(n12534) );
  AOI22HSV4 U15031 ( .A1(\pe3/ti_7t [11]), .A2(n16054), .B1(n16050), .B2(
        n16049), .ZN(n16111) );
  XNOR2HSV4 U15032 ( .A1(n12538), .A2(n12536), .ZN(n12535) );
  XOR2HSV2 U15033 ( .A1(n16156), .A2(n16155), .Z(n12537) );
  AOI21HSV4 U15034 ( .A1(n21719), .A2(n16052), .B(n16051), .ZN(n12539) );
  AOI21HSV4 U15035 ( .A1(n16035), .A2(n28708), .B(n16034), .ZN(n16050) );
  OAI21HSV4 U15036 ( .A1(n14054), .A2(n23374), .B(n16158), .ZN(n12540) );
  XNOR2HSV4 U15037 ( .A1(n12541), .A2(\pe4/phq [5]), .ZN(n13702) );
  CLKNAND2HSV2 U15038 ( .A1(\pe4/got [12]), .A2(\pe4/ti_1 ), .ZN(n12541) );
  CLKNAND2HSV2 U15039 ( .A1(n12542), .A2(\pe3/phq [2]), .ZN(n15041) );
  CLKNAND2HSV2 U15040 ( .A1(\pe3/aot [16]), .A2(\pe3/bq[15] ), .ZN(n12542) );
  CLKNAND2HSV2 U15041 ( .A1(n21632), .A2(n25364), .ZN(n21628) );
  XNOR2HSV4 U15042 ( .A1(n21311), .A2(n21310), .ZN(n21629) );
  IOA21HSV4 U15043 ( .A1(\pe10/pvq [1]), .A2(\pe10/ctrq ), .B(\pe10/phq [1]), 
        .ZN(n12543) );
  NAND3HSV4 U15044 ( .A1(n12545), .A2(\pe10/ctrq ), .A3(\pe10/pvq [1]), .ZN(
        n12544) );
  CLKNHSV2 U15045 ( .I(\pe10/phq [1]), .ZN(n12545) );
  CLKNHSV2 U15046 ( .I(n28795), .ZN(n18560) );
  CLKNAND2HSV2 U15047 ( .A1(n28795), .A2(n14039), .ZN(n13482) );
  XNOR2HSV4 U15048 ( .A1(n16174), .A2(n16173), .ZN(n16167) );
  XNOR2HSV4 U15049 ( .A1(n12547), .A2(n12546), .ZN(n16173) );
  CLKNAND2HSV2 U15050 ( .A1(n28945), .A2(\pe3/got [13]), .ZN(n12546) );
  XNOR2HSV4 U15051 ( .A1(n16104), .A2(n16105), .ZN(n12547) );
  CLKNAND2HSV1 U15052 ( .A1(n12548), .A2(n20992), .ZN(n20996) );
  CLKNHSV2 U15053 ( .I(n12549), .ZN(n27574) );
  CLKNAND2HSV2 U15054 ( .A1(n12558), .A2(n12550), .ZN(n12549) );
  CLKNHSV2 U15055 ( .I(n27572), .ZN(n12550) );
  CLKNHSV2 U15056 ( .I(n12551), .ZN(n27665) );
  CLKNAND2HSV2 U15057 ( .A1(n12558), .A2(n12552), .ZN(n12551) );
  CLKNHSV2 U15058 ( .I(n27663), .ZN(n12552) );
  CLKNHSV2 U15059 ( .I(n12553), .ZN(n27721) );
  CLKNAND2HSV2 U15060 ( .A1(n12558), .A2(n12554), .ZN(n12553) );
  CLKNHSV2 U15061 ( .I(n27718), .ZN(n12554) );
  OAI21HSV1 U15062 ( .A1(n12562), .A2(n12557), .B(n12555), .ZN(n13735) );
  CLKNAND2HSV3 U15063 ( .A1(n12556), .A2(n13734), .ZN(n12555) );
  CLKNAND2HSV4 U15064 ( .A1(n12558), .A2(n12563), .ZN(n12556) );
  INHSV2 U15065 ( .I(n12558), .ZN(n12557) );
  CLKNAND2HSV3 U15066 ( .A1(n27571), .A2(\pe2/ti_7t [14]), .ZN(n12559) );
  NAND2HSV2 U15067 ( .A1(n28967), .A2(n12561), .ZN(n12560) );
  INHSV2 U15068 ( .I(n27571), .ZN(n12561) );
  CLKNAND2HSV1 U15069 ( .A1(n12564), .A2(n12563), .ZN(n12562) );
  CLKNHSV4 U15070 ( .I(n27735), .ZN(n12563) );
  CLKNHSV1 U15071 ( .I(n13734), .ZN(n12564) );
  XOR2HSV2 U15072 ( .A1(n12566), .A2(n12565), .Z(n20152) );
  CLKNAND2HSV2 U15073 ( .A1(\pe11/aot [14]), .A2(\pe11/bq[16] ), .ZN(n12565)
         );
  CLKNAND2HSV2 U15074 ( .A1(\pe11/aot [15]), .A2(\pe11/bq[15] ), .ZN(n12566)
         );
  CLKNHSV2 U15075 ( .I(n18223), .ZN(n18100) );
  NOR2HSV4 U15076 ( .A1(n12567), .A2(n18098), .ZN(n18099) );
  NOR2HSV4 U15077 ( .A1(n18223), .A2(n12568), .ZN(n12567) );
  CLKNHSV2 U15078 ( .I(n18529), .ZN(n12568) );
  CLKNAND2HSV4 U15079 ( .A1(n21149), .A2(n21148), .ZN(n21241) );
  CLKNAND2HSV4 U15080 ( .A1(n29039), .A2(n21714), .ZN(n21149) );
  CLKNAND2HSV2 U15081 ( .A1(n15399), .A2(n15400), .ZN(n15404) );
  CLKNAND2HSV4 U15082 ( .A1(n15402), .A2(n15401), .ZN(n15403) );
  NAND3HSV4 U15083 ( .A1(n12572), .A2(n15405), .A3(n12575), .ZN(n15481) );
  CLKNHSV3 U15084 ( .I(n15480), .ZN(n12574) );
  CLKNHSV3 U15085 ( .I(n15374), .ZN(n12575) );
  CLKNAND2HSV2 U15086 ( .A1(\pe10/bq[14] ), .A2(\pe10/aot [14]), .ZN(n16689)
         );
  CLKNAND2HSV2 U15087 ( .A1(n17985), .A2(n12576), .ZN(n17986) );
  CLKNHSV2 U15088 ( .I(n17983), .ZN(n12576) );
  CLKNAND2HSV2 U15089 ( .A1(n12578), .A2(n12577), .ZN(n17983) );
  CLKNHSV2 U15090 ( .I(n18530), .ZN(n12577) );
  CLKNAND2HSV2 U15091 ( .A1(n18021), .A2(n18022), .ZN(n12578) );
  XNOR2HSV4 U15092 ( .A1(n12878), .A2(n12579), .ZN(n19566) );
  CLKNAND2HSV2 U15093 ( .A1(n25270), .A2(n24271), .ZN(n12579) );
  CLKNAND2HSV4 U15094 ( .A1(n12603), .A2(n18922), .ZN(n19158) );
  INHSV4 U15095 ( .I(n16336), .ZN(n12580) );
  CLKNAND2HSV4 U15096 ( .A1(n16557), .A2(n12583), .ZN(n16336) );
  CLKNAND2HSV2 U15097 ( .A1(n16388), .A2(n12581), .ZN(n16308) );
  CLKNAND2HSV2 U15098 ( .A1(n12582), .A2(n12584), .ZN(n12581) );
  CLKNAND2HSV2 U15099 ( .A1(n16334), .A2(n16307), .ZN(n12582) );
  CLKNAND2HSV2 U15100 ( .A1(n12580), .A2(n21328), .ZN(n16388) );
  CLKNHSV2 U15101 ( .I(n16336), .ZN(n21329) );
  CLKNHSV2 U15102 ( .I(n12587), .ZN(n12583) );
  CLKNHSV0 U15103 ( .I(n16557), .ZN(n16385) );
  CLKNAND2HSV2 U15104 ( .A1(n16557), .A2(n12585), .ZN(n12584) );
  CLKNHSV2 U15105 ( .I(n12908), .ZN(n12585) );
  XNOR2HSV4 U15106 ( .A1(n16306), .A2(n16305), .ZN(n16334) );
  XNOR2HSV4 U15107 ( .A1(n12586), .A2(n16303), .ZN(n16305) );
  CLKNHSV2 U15108 ( .I(n16302), .ZN(n12586) );
  XNOR2HSV4 U15109 ( .A1(n16301), .A2(n16300), .ZN(n16306) );
  CLKNHSV2 U15110 ( .I(n28695), .ZN(n12587) );
  AOI21HSV4 U15111 ( .A1(n26921), .A2(n26922), .B(n12589), .ZN(n12588) );
  CLKNAND2HSV2 U15112 ( .A1(n12590), .A2(n26931), .ZN(n12589) );
  CLKNAND2HSV2 U15113 ( .A1(n26927), .A2(n26928), .ZN(n12590) );
  CLKNAND2HSV2 U15114 ( .A1(n27940), .A2(n28612), .ZN(n12591) );
  INAND2HSV4 U15115 ( .A1(n12592), .B1(n22928), .ZN(n27940) );
  CLKNHSV2 U15116 ( .I(n22927), .ZN(n12592) );
  NOR2HSV4 U15117 ( .A1(n21814), .A2(n23434), .ZN(n21886) );
  XNOR2HSV4 U15118 ( .A1(n21892), .A2(n21891), .ZN(n21814) );
  INHSV2 U15119 ( .I(n16809), .ZN(n12598) );
  CLKNAND2HSV2 U15120 ( .A1(n16615), .A2(n16614), .ZN(n16613) );
  CLKNAND2HSV2 U15121 ( .A1(n12598), .A2(\pe10/aot [15]), .ZN(n16614) );
  INHSV2 U15122 ( .I(n19130), .ZN(n12601) );
  CLKNHSV2 U15123 ( .I(n12851), .ZN(n12600) );
  CLKNHSV2 U15124 ( .I(n12850), .ZN(n12602) );
  XNOR2HSV4 U15125 ( .A1(n12606), .A2(n12604), .ZN(n19144) );
  XOR3HSV2 U15126 ( .A1(n19122), .A2(n19123), .A3(n12605), .Z(n12604) );
  CLKNAND2HSV2 U15127 ( .A1(n19075), .A2(n19074), .ZN(n12605) );
  CLKNHSV2 U15128 ( .I(n19705), .ZN(n12610) );
  INOR2HSV4 U15129 ( .A1(n19683), .B1(n12612), .ZN(n19704) );
  CLKNAND2HSV2 U15130 ( .A1(n19682), .A2(n19699), .ZN(n12612) );
  CLKNAND2HSV2 U15131 ( .A1(n19618), .A2(n19619), .ZN(n19683) );
  AOI21HSV4 U15132 ( .A1(n19679), .A2(n19678), .B(n25628), .ZN(n19688) );
  CLKNAND2HSV4 U15133 ( .A1(n25182), .A2(\pe11/got [4]), .ZN(n13594) );
  CLKNAND2HSV4 U15134 ( .A1(n20847), .A2(n25415), .ZN(n23319) );
  CLKBUFHSV2 U15135 ( .I(\pe9/aot [16]), .Z(n12618) );
  CLKNAND2HSV2 U15136 ( .A1(\pe9/aot [16]), .A2(\pe9/bq[12] ), .ZN(n17876) );
  CLKNAND2HSV2 U15137 ( .A1(n12618), .A2(\pe9/bq[5] ), .ZN(n18414) );
  CLKNAND2HSV2 U15138 ( .A1(n12618), .A2(\pe9/bq[7] ), .ZN(n18232) );
  CLKNAND2HSV2 U15139 ( .A1(n12618), .A2(\pe9/bq[3] ), .ZN(n18583) );
  CLKNAND2HSV2 U15140 ( .A1(n12618), .A2(\pe9/bq[1] ), .ZN(n28036) );
  NOR2HSV3 U15141 ( .A1(n12622), .A2(n12621), .ZN(n12619) );
  CLKNAND2HSV3 U15142 ( .A1(n16710), .A2(n16678), .ZN(n12620) );
  XOR2HSV4 U15143 ( .A1(n16848), .A2(n16753), .Z(n16710) );
  CLKNHSV3 U15144 ( .I(n16708), .ZN(n12623) );
  BUFHSV8 U15145 ( .I(n22084), .Z(n12624) );
  CLKNAND2HSV4 U15146 ( .A1(n21149), .A2(n21148), .ZN(n22084) );
  NAND3HSV4 U15147 ( .A1(n25687), .A2(n12626), .A3(n16844), .ZN(n22764) );
  NOR2HSV4 U15148 ( .A1(n12625), .A2(n22504), .ZN(n22765) );
  NOR2HSV4 U15149 ( .A1(n25687), .A2(n12626), .ZN(n12625) );
  CLKNAND2HSV4 U15150 ( .A1(n22441), .A2(n16892), .ZN(n25687) );
  XNOR2HSV4 U15151 ( .A1(n14851), .A2(n12628), .ZN(n12627) );
  XOR2HSV2 U15152 ( .A1(n12630), .A2(n12629), .Z(n12628) );
  CLKNAND2HSV2 U15153 ( .A1(n14848), .A2(n24637), .ZN(n12629) );
  XNOR2HSV4 U15154 ( .A1(n14849), .A2(n14850), .ZN(n12630) );
  CLKNHSV2 U15155 ( .I(n20979), .ZN(n12632) );
  CLKNAND2HSV2 U15156 ( .A1(n14902), .A2(n14852), .ZN(n12633) );
  AOI21HSV4 U15157 ( .A1(n14806), .A2(n14807), .B(n14805), .ZN(n12634) );
  NAND2HSV2 U15158 ( .A1(n14905), .A2(n12639), .ZN(n12636) );
  INHSV2 U15159 ( .I(n12636), .ZN(n14824) );
  OAI22HSV4 U15160 ( .A1(n14822), .A2(n14821), .B1(n12638), .B2(n12637), .ZN(
        n14823) );
  INAND2HSV4 U15161 ( .A1(n14821), .B1(n12639), .ZN(n12637) );
  CLKNHSV2 U15162 ( .I(n14905), .ZN(n12638) );
  CLKNHSV2 U15163 ( .I(n12640), .ZN(n12639) );
  CLKNHSV8 U15164 ( .I(n14497), .ZN(n12640) );
  AOI21HSV4 U15165 ( .A1(n18048), .A2(n18049), .B(n18047), .ZN(n18096) );
  CLKNAND2HSV2 U15166 ( .A1(n19794), .A2(n28423), .ZN(n12641) );
  OAI21HSV4 U15167 ( .A1(n18096), .A2(n18097), .B(n12642), .ZN(n19794) );
  CLKNAND2HSV2 U15168 ( .A1(n18091), .A2(n23465), .ZN(n12642) );
  AOI21HSV4 U15169 ( .A1(n23466), .A2(n18338), .B(n18086), .ZN(n18097) );
  OAI21HSV4 U15170 ( .A1(n29041), .A2(n12646), .B(n12643), .ZN(n21156) );
  AOI21HSV4 U15171 ( .A1(n21106), .A2(n12645), .B(n12644), .ZN(n12643) );
  CLKNHSV2 U15172 ( .I(n28429), .ZN(n12644) );
  CLKNHSV2 U15173 ( .I(n21714), .ZN(n12645) );
  CLKNHSV2 U15174 ( .I(n21106), .ZN(n12646) );
  XNOR2HSV4 U15175 ( .A1(n12650), .A2(n12647), .ZN(n14352) );
  XNOR2HSV4 U15176 ( .A1(n12649), .A2(n12648), .ZN(n12647) );
  CLKNAND2HSV2 U15177 ( .A1(n27072), .A2(\pe6/pvq [8]), .ZN(n12648) );
  XOR2HSV2 U15178 ( .A1(n23021), .A2(\pe6/phq [8]), .Z(n12649) );
  XOR2HSV2 U15179 ( .A1(n14344), .A2(n12651), .Z(n12650) );
  XOR2HSV2 U15180 ( .A1(n12652), .A2(n14341), .Z(n12651) );
  CLKNAND2HSV2 U15181 ( .A1(n25701), .A2(\pe6/aot [13]), .ZN(n12652) );
  XNOR2HSV4 U15182 ( .A1(n24690), .A2(n12653), .ZN(n24692) );
  CLKNAND2HSV2 U15183 ( .A1(\pe5/ti_7[10] ), .A2(n24637), .ZN(n12653) );
  CLKNAND2HSV2 U15184 ( .A1(pov5[10]), .A2(n14815), .ZN(n12654) );
  XNOR2HSV4 U15185 ( .A1(n20986), .A2(n20985), .ZN(pov5[10]) );
  MUX2NHSV1 U15186 ( .I0(n14398), .I1(n14397), .S(n14736), .ZN(n12655) );
  AOI21HSV2 U15187 ( .A1(n12662), .A2(n12657), .B(n18623), .ZN(n12656) );
  INHSV2 U15188 ( .I(n18622), .ZN(n12657) );
  INAND2HSV2 U15189 ( .A1(n12660), .B1(n18614), .ZN(n12658) );
  NAND3HSV2 U15190 ( .A1(n12661), .A2(n12660), .A3(n18622), .ZN(n12659) );
  OAI21HSV2 U15191 ( .A1(n18620), .A2(n18616), .B(n12300), .ZN(n12660) );
  INHSV2 U15192 ( .I(n12662), .ZN(n12661) );
  NOR2HSV2 U15193 ( .A1(n18620), .A2(n18621), .ZN(n12662) );
  OAI21HSV1 U15194 ( .A1(pov4[14]), .A2(n27976), .B(n27975), .ZN(n27997) );
  NAND2HSV2 U15195 ( .A1(n13602), .A2(n12664), .ZN(pov4[14]) );
  CLKNAND2HSV1 U15196 ( .A1(n12666), .A2(n12665), .ZN(n12664) );
  NOR2HSV3 U15197 ( .A1(n22796), .A2(n26930), .ZN(n12665) );
  CLKNHSV0 U15198 ( .I(n26928), .ZN(n12666) );
  XNOR2HSV4 U15199 ( .A1(n12673), .A2(n12667), .ZN(n23317) );
  MUX2NHSV2 U15200 ( .I0(n12671), .I1(n12670), .S(n12668), .ZN(n12667) );
  XNOR2HSV4 U15201 ( .A1(n12669), .A2(n23316), .ZN(n12668) );
  CLKNAND2HSV2 U15202 ( .A1(n24965), .A2(\pe11/got [1]), .ZN(n12669) );
  CLKNHSV2 U15203 ( .I(n12672), .ZN(n12671) );
  CLKNAND2HSV2 U15204 ( .A1(n28919), .A2(\pe11/got [2]), .ZN(n12672) );
  CLKNAND2HSV2 U15205 ( .A1(n24903), .A2(\pe11/got [3]), .ZN(n12673) );
  INHSV2 U15206 ( .I(n22043), .ZN(n12674) );
  CLKNAND2HSV0 U15207 ( .A1(n22043), .A2(n22042), .ZN(n27980) );
  NOR2HSV4 U15208 ( .A1(n12674), .A2(n12675), .ZN(n15904) );
  CLKNAND2HSV2 U15209 ( .A1(n22042), .A2(n12676), .ZN(n12675) );
  CLKNHSV2 U15210 ( .I(n22801), .ZN(n12676) );
  CLKNAND2HSV4 U15211 ( .A1(n12679), .A2(n12677), .ZN(n22043) );
  CLKNAND2HSV2 U15212 ( .A1(n12683), .A2(n12682), .ZN(n12678) );
  AOI21HSV4 U15213 ( .A1(n25666), .A2(n25668), .B(n22801), .ZN(n12679) );
  XNOR2HSV4 U15214 ( .A1(n15750), .A2(n15749), .ZN(n25668) );
  NOR2HSV4 U15215 ( .A1(n12681), .A2(n12680), .ZN(n25667) );
  CLKNHSV2 U15216 ( .I(n12682), .ZN(n12680) );
  CLKNHSV2 U15217 ( .I(n12683), .ZN(n12681) );
  CLKNAND2HSV2 U15218 ( .A1(n21993), .A2(n15699), .ZN(n12682) );
  CLKNAND2HSV2 U15219 ( .A1(n15751), .A2(n15842), .ZN(n12683) );
  CLKNAND2HSV3 U15220 ( .A1(n18104), .A2(n18325), .ZN(n18042) );
  CLKNAND2HSV4 U15221 ( .A1(n18044), .A2(n18043), .ZN(n18104) );
  CLKNAND2HSV2 U15222 ( .A1(n17961), .A2(n17960), .ZN(n18043) );
  NOR2HSV4 U15223 ( .A1(n12687), .A2(n12686), .ZN(n12692) );
  CLKNAND2HSV2 U15224 ( .A1(\pe7/ti_1 ), .A2(\pe7/got [16]), .ZN(n12686) );
  CLKNHSV2 U15225 ( .I(n12694), .ZN(n12687) );
  BUFHSV8 U15226 ( .I(\pe7/ctrq ), .Z(n12688) );
  AOI22HSV4 U15227 ( .A1(n12688), .A2(n12690), .B1(n12689), .B2(n19176), .ZN(
        n19178) );
  CLKNHSV2 U15228 ( .I(n12691), .ZN(n12690) );
  CLKNAND2HSV2 U15229 ( .A1(\pe7/phq [1]), .A2(\pe7/pvq [1]), .ZN(n12691) );
  AOI21HSV4 U15230 ( .A1(n12695), .A2(n12693), .B(n12692), .ZN(n19177) );
  CLKNHSV2 U15231 ( .I(n12694), .ZN(n12693) );
  CLKNAND2HSV2 U15232 ( .A1(n23138), .A2(\pe7/got [16]), .ZN(n12695) );
  CLKNAND2HSV2 U15233 ( .A1(n29023), .A2(n18927), .ZN(n18929) );
  OAI21HSV4 U15234 ( .A1(n29023), .A2(n18992), .B(n14739), .ZN(n14740) );
  OAI21HSV1 U15235 ( .A1(n29023), .A2(n18859), .B(n18858), .ZN(n18898) );
  XNOR2HSV2 U15236 ( .A1(n14737), .A2(n14736), .ZN(n29023) );
  CLKNAND2HSV4 U15237 ( .A1(n12697), .A2(n12696), .ZN(n12698) );
  CLKNHSV4 U15238 ( .I(n12432), .ZN(n12696) );
  NAND3HSV4 U15239 ( .A1(n12698), .A2(n13338), .A3(n12699), .ZN(n19075) );
  INHSV2 U15240 ( .I(n18925), .ZN(n12699) );
  CLKNAND2HSV2 U15241 ( .A1(\pe9/aot [16]), .A2(\pe9/bq[14] ), .ZN(n17939) );
  XOR2HSV2 U15242 ( .A1(n17939), .A2(n12700), .Z(n17941) );
  CLKNAND2HSV2 U15243 ( .A1(\pe9/bq[16] ), .A2(\pe9/aot [14]), .ZN(n12700) );
  CLKNAND2HSV3 U15244 ( .A1(n17771), .A2(n21696), .ZN(n12703) );
  XNOR2HSV4 U15245 ( .A1(n17747), .A2(n17746), .ZN(n17771) );
  INHSV2 U15246 ( .I(n12702), .ZN(n17858) );
  NOR2HSV4 U15247 ( .A1(n23471), .A2(n12703), .ZN(n12702) );
  CLKBUFHSV2 U15248 ( .I(n12705), .Z(n12704) );
  CLKNHSV2 U15249 ( .I(n12705), .ZN(n12746) );
  CLKNAND2HSV2 U15250 ( .A1(n12705), .A2(\pe10/got [13]), .ZN(n13196) );
  CLKNAND2HSV2 U15251 ( .A1(n12704), .A2(\pe10/got [9]), .ZN(n22487) );
  CLKNAND2HSV2 U15252 ( .A1(n12704), .A2(n14065), .ZN(n22743) );
  CLKNAND2HSV2 U15253 ( .A1(n12704), .A2(\pe10/got [5]), .ZN(n22668) );
  CLKNAND2HSV2 U15254 ( .A1(n12704), .A2(\pe10/got [4]), .ZN(n24486) );
  INAND2HSV4 U15255 ( .A1(n12706), .B1(n16896), .ZN(n12705) );
  CLKNHSV2 U15256 ( .I(n16895), .ZN(n12706) );
  INHSV24 U15257 ( .I(n19622), .ZN(n12707) );
  INHSV2 U15258 ( .I(n25345), .ZN(n12708) );
  CLKNAND2HSV2 U15259 ( .A1(n19698), .A2(n23112), .ZN(n14030) );
  OAI21HSV4 U15260 ( .A1(n12712), .A2(n12711), .B(n12710), .ZN(n23112) );
  CLKNHSV2 U15261 ( .I(n25345), .ZN(n12711) );
  CLKNAND2HSV2 U15262 ( .A1(n25346), .A2(n19697), .ZN(n12712) );
  CLKNAND2HSV2 U15263 ( .A1(n19693), .A2(n19692), .ZN(n19698) );
  NOR2HSV4 U15264 ( .A1(n12708), .A2(n12707), .ZN(n19692) );
  CLKNAND2HSV2 U15265 ( .A1(n19681), .A2(n19680), .ZN(n12713) );
  CLKNHSV2 U15266 ( .I(n13986), .ZN(n12714) );
  CLKNAND2HSV2 U15267 ( .A1(n19691), .A2(n19690), .ZN(n12715) );
  XNOR2HSV4 U15268 ( .A1(n12718), .A2(n12717), .ZN(n12716) );
  XNOR2HSV4 U15269 ( .A1(n19673), .A2(n19672), .ZN(n12717) );
  CLKNAND2HSV2 U15270 ( .A1(n25377), .A2(n24271), .ZN(n12718) );
  CLKNAND2HSV2 U15271 ( .A1(n21321), .A2(n20227), .ZN(n20757) );
  CLKNHSV2 U15272 ( .I(n20706), .ZN(n12719) );
  CLKNAND2HSV2 U15273 ( .A1(n25352), .A2(n23436), .ZN(n12720) );
  XNOR2HSV4 U15274 ( .A1(n12721), .A2(n20693), .ZN(n25352) );
  XNOR2HSV4 U15275 ( .A1(n20445), .A2(n20560), .ZN(n20693) );
  CLKNAND2HSV3 U15276 ( .A1(n18535), .A2(n18534), .ZN(n12722) );
  CLKNAND2HSV3 U15277 ( .A1(n18461), .A2(n18460), .ZN(n12723) );
  XOR2HSV2 U15278 ( .A1(n12726), .A2(n12725), .Z(n14167) );
  CLKNAND2HSV2 U15279 ( .A1(\pe6/aot [16]), .A2(\pe6/bq[13] ), .ZN(n12725) );
  CLKNAND2HSV2 U15280 ( .A1(\pe6/aot [15]), .A2(\pe6/bq[14] ), .ZN(n12726) );
  INHSV2 U15281 ( .I(n17407), .ZN(n12728) );
  NOR2HSV4 U15282 ( .A1(n17277), .A2(n17278), .ZN(n12730) );
  INOR2HSV4 U15283 ( .A1(n17363), .B1(n12728), .ZN(n12731) );
  CLKNAND2HSV2 U15284 ( .A1(n17404), .A2(n17403), .ZN(n17363) );
  CLKNAND2HSV2 U15285 ( .A1(n17240), .A2(n12732), .ZN(n17403) );
  CLKNHSV2 U15286 ( .I(n17241), .ZN(n12732) );
  NOR2HSV4 U15287 ( .A1(n17238), .A2(n17341), .ZN(n17404) );
  XOR2HSV2 U15288 ( .A1(n17595), .A2(n12733), .Z(n17596) );
  AOI21HSV4 U15289 ( .A1(n28968), .A2(n12735), .B(n12734), .ZN(n26540) );
  CLKNHSV2 U15290 ( .I(n17532), .ZN(n12734) );
  CLKNHSV2 U15291 ( .I(n17531), .ZN(n12735) );
  CLKNAND2HSV0 U15292 ( .A1(n28997), .A2(n12736), .ZN(n17020) );
  INHSV2 U15293 ( .I(n22442), .ZN(n12736) );
  OAI21HSV4 U15294 ( .A1(n28997), .A2(n16843), .B(n16806), .ZN(n16841) );
  CLKNAND2HSV2 U15295 ( .A1(n18645), .A2(n14039), .ZN(n18549) );
  NOR2HSV2 U15296 ( .A1(n27438), .A2(n21305), .ZN(n21307) );
  INHSV2 U15297 ( .I(n12738), .ZN(n12737) );
  CLKNAND2HSV3 U15298 ( .A1(n21643), .A2(\pe2/ti_7t [9]), .ZN(n12738) );
  INHSV2 U15299 ( .I(n21643), .ZN(n12739) );
  INAND2HSV2 U15300 ( .A1(n21644), .B1(n21642), .ZN(n28956) );
  AOI21HSV2 U15301 ( .A1(n22084), .A2(\pe2/got [16]), .B(n21064), .ZN(n21644)
         );
  NAND3HSV4 U15302 ( .A1(n12741), .A2(n17414), .A3(n17536), .ZN(n17415) );
  CLKNHSV2 U15303 ( .I(n17413), .ZN(n12741) );
  CLKNHSV2 U15304 ( .I(n12743), .ZN(n12742) );
  CLKNAND2HSV2 U15305 ( .A1(n22082), .A2(n17359), .ZN(n12743) );
  CLKNAND2HSV2 U15306 ( .A1(n13732), .A2(n13731), .ZN(n13733) );
  CLKNAND2HSV2 U15307 ( .A1(n28590), .A2(n14055), .ZN(n13732) );
  CLKNAND2HSV2 U15308 ( .A1(n27295), .A2(n27294), .ZN(n27731) );
  CLKNAND2HSV2 U15309 ( .A1(n21636), .A2(n21304), .ZN(n27294) );
  CLKNHSV2 U15310 ( .I(n17003), .ZN(n17007) );
  NAND3HSV4 U15311 ( .A1(n17003), .A2(n26212), .A3(n17002), .ZN(n12744) );
  NOR2HSV4 U15312 ( .A1(n12746), .A2(n12745), .ZN(n17003) );
  CLKNHSV2 U15313 ( .I(n16759), .ZN(n12745) );
  CLKNHSV4 U15314 ( .I(\pe9/ctrq ), .ZN(n18167) );
  CLKNHSV0 U15315 ( .I(n17408), .ZN(n12748) );
  OAI21HSV4 U15316 ( .A1(n12756), .A2(n12749), .B(n12747), .ZN(n28968) );
  OAI21HSV4 U15317 ( .A1(n12756), .A2(n12748), .B(n12329), .ZN(n12747) );
  CLKNAND2HSV2 U15318 ( .A1(n12750), .A2(n17408), .ZN(n12749) );
  OAI21HSV2 U15319 ( .A1(n12755), .A2(n12752), .B(n12751), .ZN(n13123) );
  XNOR2HSV1 U15320 ( .A1(n12754), .A2(n12753), .ZN(n12752) );
  XNOR2HSV2 U15321 ( .A1(n17401), .A2(n17400), .ZN(n12754) );
  INAND2HSV2 U15322 ( .A1(n17364), .B1(n12274), .ZN(n12755) );
  OAI21HSV2 U15323 ( .A1(n28968), .A2(n17410), .B(n17409), .ZN(n13124) );
  NOR2HSV0 U15324 ( .A1(n17706), .A2(n21159), .ZN(n17709) );
  INHSV4 U15325 ( .I(n17130), .ZN(n17133) );
  CLKNHSV6 U15326 ( .I(n15747), .ZN(n21992) );
  INHSV4 U15327 ( .I(n17914), .ZN(n25634) );
  NAND2HSV2 U15328 ( .A1(n17857), .A2(n17856), .ZN(n12759) );
  CLKNAND2HSV2 U15329 ( .A1(n12757), .A2(n12758), .ZN(n12760) );
  CLKNAND2HSV2 U15330 ( .A1(n12759), .A2(n12760), .ZN(n17868) );
  CLKNHSV2 U15331 ( .I(n17857), .ZN(n12757) );
  CLKNHSV2 U15332 ( .I(n17856), .ZN(n12758) );
  NAND2HSV4 U15333 ( .A1(n16702), .A2(n16703), .ZN(n16705) );
  CLKNAND2HSV4 U15334 ( .A1(n16701), .A2(n16700), .ZN(n16702) );
  NAND2HSV2 U15335 ( .A1(n24007), .A2(n24006), .ZN(n12763) );
  CLKNAND2HSV2 U15336 ( .A1(n12761), .A2(n12762), .ZN(n12764) );
  NAND2HSV2 U15337 ( .A1(n12763), .A2(n12764), .ZN(\pe6/poht [13]) );
  CLKNHSV2 U15338 ( .I(n24007), .ZN(n12761) );
  CLKNHSV2 U15339 ( .I(n24006), .ZN(n12762) );
  CLKXOR2HSV2 U15340 ( .A1(n24005), .A2(n24004), .Z(n24006) );
  CLKNAND2HSV2 U15341 ( .A1(n14580), .A2(n14561), .ZN(n14562) );
  NOR2HSV4 U15342 ( .A1(n25663), .A2(n15480), .ZN(n15680) );
  CLKNAND2HSV4 U15343 ( .A1(n13968), .A2(n14269), .ZN(n14275) );
  XOR2HSV4 U15344 ( .A1(n17728), .A2(n17727), .Z(n12765) );
  CKMUX2HSV2 U15345 ( .I0(bo6[15]), .I1(\pe6/bq[15] ), .S(n22109), .Z(n28868)
         );
  NAND2HSV4 U15346 ( .A1(n17687), .A2(n17686), .ZN(n17708) );
  NAND2HSV4 U15347 ( .A1(n14259), .A2(n18907), .ZN(n14260) );
  CLKNAND2HSV4 U15348 ( .A1(n14289), .A2(n14288), .ZN(n14286) );
  MOAI22HSV4 U15349 ( .A1(n24964), .A2(n14147), .B1(n25058), .B2(n14146), .ZN(
        n14150) );
  CLKXOR2HSV4 U15350 ( .A1(n22553), .A2(n22552), .Z(n22555) );
  INHSV4 U15351 ( .I(n26215), .ZN(n26093) );
  AND2HSV2 U15352 ( .A1(n26215), .A2(n26132), .Z(n22586) );
  INHSV2 U15353 ( .I(n22787), .ZN(n22785) );
  XNOR2HSV4 U15354 ( .A1(n22784), .A2(n22783), .ZN(n22787) );
  CLKXOR2HSV4 U15355 ( .A1(n22782), .A2(n22781), .Z(n22784) );
  OAI31HSV0 U15356 ( .A1(n22698), .A2(n27194), .A3(n22692), .B(n22697), .ZN(
        n22699) );
  XNOR2HSV4 U15357 ( .A1(n21996), .A2(n21995), .ZN(n22040) );
  CLKNAND2HSV4 U15358 ( .A1(n15679), .A2(n15678), .ZN(n25663) );
  CLKNAND2HSV4 U15359 ( .A1(n13130), .A2(n13131), .ZN(n13132) );
  INHSV2 U15360 ( .I(n14231), .ZN(n12766) );
  NAND2HSV4 U15361 ( .A1(n17827), .A2(n17826), .ZN(n17804) );
  CLKNAND2HSV4 U15362 ( .A1(n14261), .A2(n14260), .ZN(n14271) );
  INHSV4 U15363 ( .I(n14258), .ZN(n14261) );
  NAND2HSV4 U15364 ( .A1(n13128), .A2(n13127), .ZN(n13129) );
  CLKNAND2HSV2 U15365 ( .A1(n14197), .A2(n14196), .ZN(n14205) );
  NAND2HSV4 U15366 ( .A1(n14205), .A2(n14204), .ZN(n14208) );
  AND2HSV4 U15367 ( .A1(n14270), .A2(n14272), .Z(n13968) );
  INHSV4 U15368 ( .I(n14507), .ZN(n14510) );
  NAND2HSV2 U15369 ( .A1(n14333), .A2(n14334), .ZN(n12769) );
  NAND2HSV4 U15370 ( .A1(n12769), .A2(n12770), .ZN(n14335) );
  CLKNHSV2 U15371 ( .I(n14334), .ZN(n12767) );
  INHSV4 U15372 ( .I(n23471), .ZN(n17697) );
  XNOR2HSV4 U15373 ( .A1(n17056), .A2(n17055), .ZN(n17057) );
  INHSV6 U15374 ( .I(\pe6/phq [2]), .ZN(n14108) );
  NAND3HSV2 U15375 ( .A1(n18912), .A2(n18911), .A3(n18910), .ZN(n18913) );
  INHSV2 U15376 ( .I(n14200), .ZN(n12793) );
  NAND2HSV2 U15377 ( .A1(n14332), .A2(n14331), .ZN(n12773) );
  INHSV4 U15378 ( .I(n14332), .ZN(n12771) );
  CLKNHSV0 U15379 ( .I(n14331), .ZN(n12772) );
  NAND2HSV4 U15380 ( .A1(n14737), .A2(n14399), .ZN(n14431) );
  CLKNAND2HSV4 U15381 ( .A1(n17741), .A2(n17740), .ZN(n17746) );
  NAND2HSV4 U15382 ( .A1(n17827), .A2(n17826), .ZN(n21817) );
  CLKNAND2HSV4 U15383 ( .A1(n17771), .A2(n21641), .ZN(n17827) );
  XNOR2HSV4 U15384 ( .A1(n23224), .A2(n12775), .ZN(n23225) );
  XOR2HSV0 U15385 ( .A1(n23223), .A2(n26162), .Z(n12775) );
  NAND2HSV2 U15386 ( .A1(n23241), .A2(n23240), .ZN(\pe5/poht [13]) );
  CLKNAND2HSV2 U15387 ( .A1(n20994), .A2(n20993), .ZN(n20995) );
  MUX2NHSV4 U15388 ( .I0(n18453), .I1(n13481), .S(n13482), .ZN(n18535) );
  NAND2HSV0 U15389 ( .A1(n13725), .A2(n13724), .ZN(n13726) );
  NAND2HSV4 U15390 ( .A1(n20996), .A2(n20995), .ZN(n21336) );
  NOR2HSV4 U15391 ( .A1(n14577), .A2(n14576), .ZN(n14579) );
  MUX2NHSV4 U15392 ( .I0(n14673), .I1(n13118), .S(n14672), .ZN(n13119) );
  BUFHSV4 U15393 ( .I(n14894), .Z(n14848) );
  CLKNAND2HSV2 U15394 ( .A1(n14642), .A2(\pe5/got [16]), .ZN(n14621) );
  XNOR2HSV4 U15395 ( .A1(n14799), .A2(n14798), .ZN(n14800) );
  XNOR2HSV4 U15396 ( .A1(n14797), .A2(n14796), .ZN(n14799) );
  CLKNAND2HSV4 U15397 ( .A1(n21638), .A2(n21637), .ZN(n21712) );
  CLKNAND2HSV4 U15398 ( .A1(n17859), .A2(n17858), .ZN(n28809) );
  NAND3HSV4 U15399 ( .A1(n14760), .A2(n14759), .A3(n14758), .ZN(n14761) );
  CLKXOR2HSV4 U15400 ( .A1(n19120), .A2(n19119), .Z(n19123) );
  CLKAND2HSV4 U15401 ( .A1(n20068), .A2(n16993), .Z(n17063) );
  CLKNAND2HSV4 U15402 ( .A1(n17987), .A2(n17986), .ZN(n17997) );
  INHSV4 U15403 ( .I(n16643), .ZN(n22102) );
  CLKNAND2HSV4 U15404 ( .A1(n23117), .A2(n23116), .ZN(n23118) );
  CLKNAND2HSV2 U15405 ( .A1(n25665), .A2(n23120), .ZN(n19513) );
  NOR2HSV4 U15406 ( .A1(n21066), .A2(n21164), .ZN(n17689) );
  NAND2HSV4 U15407 ( .A1(n22765), .A2(n22764), .ZN(n26221) );
  OAI21HSV2 U15408 ( .A1(n13195), .A2(n13196), .B(n13197), .ZN(n16985) );
  CLKXOR2HSV2 U15409 ( .A1(n22709), .A2(n22708), .Z(n22710) );
  CLKXOR2HSV4 U15410 ( .A1(n17854), .A2(n17853), .Z(n17857) );
  CLKNAND2HSV4 U15411 ( .A1(n17135), .A2(n17134), .ZN(n28988) );
  NAND2HSV4 U15412 ( .A1(n22440), .A2(n25689), .ZN(n22439) );
  NAND2HSV4 U15413 ( .A1(n14398), .A2(n28472), .ZN(n14737) );
  NAND2HSV4 U15414 ( .A1(n17111), .A2(n17110), .ZN(n17124) );
  INHSV4 U15415 ( .I(n17123), .ZN(n17110) );
  MUX2NHSV2 U15416 ( .I0(n12957), .I1(n17109), .S(n12958), .ZN(n17123) );
  NAND2HSV4 U15417 ( .A1(n14407), .A2(n18846), .ZN(n28938) );
  CLKNHSV0 U15418 ( .I(n29039), .ZN(n14032) );
  CLKNAND2HSV2 U15419 ( .A1(n26541), .A2(n13971), .ZN(n17347) );
  NAND2HSV2 U15420 ( .A1(n17171), .A2(n17170), .ZN(n16288) );
  NAND2HSV4 U15421 ( .A1(n19462), .A2(n19455), .ZN(n19569) );
  NAND2HSV2 U15422 ( .A1(n27907), .A2(n28612), .ZN(n22044) );
  NAND2HSV2 U15423 ( .A1(n18285), .A2(n18464), .ZN(n18320) );
  CLKNAND2HSV2 U15424 ( .A1(n16647), .A2(n16646), .ZN(n16680) );
  INHSV6 U15425 ( .I(ctro9), .ZN(n17998) );
  NAND2HSV2 U15426 ( .A1(n25334), .A2(n19670), .ZN(n12803) );
  NAND2HSV0 U15427 ( .A1(n25325), .A2(n24214), .ZN(n23161) );
  INHSV4 U15428 ( .I(n19371), .ZN(n19362) );
  NAND2HSV4 U15429 ( .A1(n15832), .A2(n15831), .ZN(n21975) );
  NAND2HSV4 U15430 ( .A1(n19971), .A2(n19970), .ZN(n20052) );
  NAND2HSV2 U15431 ( .A1(n18708), .A2(n18707), .ZN(n18712) );
  INHSV2 U15432 ( .I(n18709), .ZN(n18708) );
  XNOR2HSV1 U15433 ( .A1(n14311), .A2(\pe6/phq [7]), .ZN(n14312) );
  XOR2HSV0 U15434 ( .A1(n15164), .A2(n15163), .Z(n15165) );
  NAND2HSV2 U15435 ( .A1(n14753), .A2(n14752), .ZN(n14755) );
  OAI21HSV2 U15436 ( .A1(n14429), .A2(n13100), .B(n13101), .ZN(n13102) );
  AOI21HSV2 U15437 ( .A1(n29012), .A2(n16311), .B(n16504), .ZN(n16326) );
  NOR2HSV2 U15438 ( .A1(n19243), .A2(n19242), .ZN(n19244) );
  CLKNAND2HSV2 U15439 ( .A1(n19518), .A2(n19517), .ZN(n19519) );
  INHSV4 U15440 ( .I(ctro4), .ZN(n15417) );
  NAND2HSV2 U15441 ( .A1(n20295), .A2(n20296), .ZN(n20300) );
  NAND2HSV2 U15442 ( .A1(n20262), .A2(n20261), .ZN(n20295) );
  INHSV4 U15443 ( .I(n17664), .ZN(n13451) );
  NAND3HSV2 U15444 ( .A1(n19156), .A2(n19155), .A3(n19059), .ZN(n19060) );
  NAND3HSV2 U15445 ( .A1(n23389), .A2(n26349), .A3(n26348), .ZN(n23408) );
  NAND2HSV2 U15446 ( .A1(n17482), .A2(n17481), .ZN(n22072) );
  NAND2HSV4 U15447 ( .A1(n17542), .A2(n26595), .ZN(n17599) );
  NOR2HSV2 U15448 ( .A1(n20860), .A2(n21003), .ZN(n20854) );
  NAND2HSV2 U15449 ( .A1(n17888), .A2(n17887), .ZN(n17892) );
  NAND2HSV2 U15450 ( .A1(n17884), .A2(\pe9/phq [1]), .ZN(n17891) );
  NAND2HSV4 U15451 ( .A1(n18455), .A2(n18456), .ZN(n18528) );
  CLKNAND2HSV2 U15452 ( .A1(n19200), .A2(n19199), .ZN(n19204) );
  INHSV2 U15453 ( .I(n19565), .ZN(n19570) );
  NAND2HSV2 U15454 ( .A1(n13964), .A2(n28526), .ZN(n14432) );
  NAND2HSV2 U15455 ( .A1(n15671), .A2(n15670), .ZN(n15672) );
  CLKNAND2HSV2 U15456 ( .A1(n17628), .A2(n17627), .ZN(n17632) );
  NOR2HSV4 U15457 ( .A1(n15180), .A2(n15179), .ZN(n15289) );
  CLKNAND2HSV2 U15458 ( .A1(n19897), .A2(n19977), .ZN(n19898) );
  NAND2HSV2 U15459 ( .A1(n25692), .A2(n25691), .ZN(n28406) );
  XNOR2HSV1 U15460 ( .A1(n23773), .A2(n23772), .ZN(n23774) );
  NAND2HSV4 U15461 ( .A1(n20288), .A2(n20279), .ZN(n20228) );
  NAND2HSV2 U15462 ( .A1(n19062), .A2(n19063), .ZN(n19066) );
  NAND2HSV2 U15463 ( .A1(n19139), .A2(n19135), .ZN(n19136) );
  NAND2HSV2 U15464 ( .A1(n22889), .A2(n22890), .ZN(n22894) );
  AND2HSV2 U15465 ( .A1(n23395), .A2(n23400), .Z(n27126) );
  NAND2HSV2 U15466 ( .A1(n22791), .A2(n22915), .ZN(n22794) );
  INHSV2 U15467 ( .I(n27940), .ZN(n27977) );
  CLKNAND2HSV2 U15468 ( .A1(n28795), .A2(n18326), .ZN(n23447) );
  NAND2HSV2 U15469 ( .A1(n19376), .A2(n23180), .ZN(n19231) );
  XOR2HSV0 U15470 ( .A1(n23602), .A2(n23601), .Z(n23603) );
  XNOR2HSV1 U15471 ( .A1(n24180), .A2(n24179), .ZN(n24184) );
  XNOR2HSV1 U15472 ( .A1(n24080), .A2(n24079), .ZN(\pe7/poht [6]) );
  NAND2HSV0 U15473 ( .A1(n26030), .A2(\pe6/got [10]), .ZN(n26078) );
  XOR2HSV0 U15474 ( .A1(n25977), .A2(n25976), .Z(n25978) );
  XNOR2HSV1 U15475 ( .A1(n16468), .A2(n16467), .ZN(n16469) );
  NAND2HSV2 U15476 ( .A1(n20264), .A2(\pe11/pvq [5]), .ZN(n20265) );
  NAND2HSV2 U15477 ( .A1(n14002), .A2(\pe10/pvq [4]), .ZN(n16652) );
  NOR2HSV2 U15478 ( .A1(n28431), .A2(n17008), .ZN(n17009) );
  NAND2HSV2 U15479 ( .A1(n18035), .A2(n18034), .ZN(n18036) );
  XNOR2HSV1 U15480 ( .A1(n18031), .A2(n18030), .ZN(n18034) );
  NOR2HSV4 U15481 ( .A1(n18182), .A2(n18003), .ZN(n18004) );
  NAND2HSV2 U15482 ( .A1(n15525), .A2(n15524), .ZN(n15526) );
  NAND2HSV2 U15483 ( .A1(n22694), .A2(n26218), .ZN(n20136) );
  NAND2HSV2 U15484 ( .A1(n18393), .A2(n18392), .ZN(n18397) );
  XNOR2HSV1 U15485 ( .A1(n21288), .A2(n21287), .ZN(n21294) );
  NAND2HSV2 U15486 ( .A1(n23177), .A2(n23430), .ZN(n23178) );
  NOR2HSV2 U15487 ( .A1(n14213), .A2(n14212), .ZN(n14214) );
  NAND3HSV3 U15488 ( .A1(n18100), .A2(n18200), .A3(n18543), .ZN(n18092) );
  OAI21HSV2 U15489 ( .A1(\pe9/phq [2]), .A2(n17897), .B(n17896), .ZN(n17899)
         );
  NAND2HSV2 U15490 ( .A1(n17897), .A2(\pe9/phq [2]), .ZN(n17896) );
  XNOR2HSV1 U15491 ( .A1(n14389), .A2(n14388), .ZN(n14390) );
  NAND2HSV2 U15492 ( .A1(n16837), .A2(n12303), .ZN(n16747) );
  NAND2HSV2 U15493 ( .A1(n16489), .A2(n16488), .ZN(n16491) );
  INHSV2 U15494 ( .I(n23481), .ZN(n15094) );
  NAND2HSV2 U15495 ( .A1(n16959), .A2(n16958), .ZN(n16986) );
  NAND3HSV2 U15496 ( .A1(n14918), .A2(n14917), .A3(n14916), .ZN(n14919) );
  NAND2HSV2 U15497 ( .A1(n21504), .A2(\pe5/got [11]), .ZN(n14963) );
  INHSV2 U15498 ( .I(n21060), .ZN(n21063) );
  NAND2HSV2 U15499 ( .A1(n21020), .A2(n21019), .ZN(n21060) );
  CLKNAND2HSV2 U15500 ( .A1(n21881), .A2(n21882), .ZN(n21885) );
  NAND2HSV2 U15501 ( .A1(n21522), .A2(n21521), .ZN(n24341) );
  MUX2NHSV1 U15502 ( .I0(n18449), .I1(n18448), .S(n18447), .ZN(n18450) );
  INHSV2 U15503 ( .I(n27226), .ZN(n16329) );
  NOR2HSV2 U15504 ( .A1(n16459), .A2(n18773), .ZN(n16425) );
  NOR2HSV2 U15505 ( .A1(n15363), .A2(n15871), .ZN(n15364) );
  NAND2HSV2 U15506 ( .A1(n20319), .A2(n20320), .ZN(n25489) );
  INHSV4 U15507 ( .I(n19711), .ZN(n28673) );
  NOR2HSV2 U15508 ( .A1(n25513), .A2(n20367), .ZN(n20301) );
  NAND2HSV4 U15509 ( .A1(n18337), .A2(n18470), .ZN(n19767) );
  NOR2HSV2 U15510 ( .A1(n26602), .A2(n26601), .ZN(n26641) );
  CLKXOR2HSV4 U15511 ( .A1(n19966), .A2(n19965), .Z(n23443) );
  NAND2HSV2 U15512 ( .A1(n17709), .A2(n17712), .ZN(n17710) );
  CLKNAND2HSV2 U15513 ( .A1(n17712), .A2(n17774), .ZN(n17735) );
  INHSV2 U15514 ( .I(n17738), .ZN(n17734) );
  NAND2HSV4 U15515 ( .A1(n25529), .A2(n13998), .ZN(n16607) );
  AOI22HSV2 U15516 ( .A1(n15976), .A2(n15017), .B1(n16106), .B2(n23396), .ZN(
        n15977) );
  NAND2HSV2 U15517 ( .A1(n19949), .A2(n19948), .ZN(n18770) );
  CLKNAND2HSV2 U15518 ( .A1(n23440), .A2(n16171), .ZN(n23420) );
  XNOR2HSV1 U15519 ( .A1(n25815), .A2(n25814), .ZN(n25816) );
  NAND2HSV0 U15520 ( .A1(n27640), .A2(n27647), .ZN(n27539) );
  NAND2HSV0 U15521 ( .A1(n27679), .A2(n14046), .ZN(n27535) );
  NAND2HSV2 U15522 ( .A1(n18522), .A2(n18523), .ZN(n18459) );
  INAND2HSV2 U15523 ( .A1(n16535), .B1(n28625), .ZN(n25650) );
  INHSV2 U15524 ( .I(n19257), .ZN(n19260) );
  NAND2HSV2 U15525 ( .A1(n19452), .A2(n19451), .ZN(n19453) );
  NAND2HSV2 U15526 ( .A1(n15674), .A2(n15675), .ZN(n15679) );
  NAND2HSV2 U15527 ( .A1(n23059), .A2(n23058), .ZN(n27957) );
  MUX2NHSV2 U15528 ( .I0(n13658), .I1(n21157), .S(n13660), .ZN(n22086) );
  XNOR2HSV2 U15529 ( .A1(n25416), .A2(n25415), .ZN(n25417) );
  CLKXOR2HSV2 U15530 ( .A1(n25133), .A2(n25132), .Z(n25136) );
  XOR2HSV0 U15531 ( .A1(n24436), .A2(n24435), .Z(\pe5/poht [2]) );
  NAND2HSV2 U15532 ( .A1(n28406), .A2(\pe9/got [6]), .ZN(n28374) );
  NAND2HSV2 U15533 ( .A1(n28406), .A2(n28405), .ZN(n28407) );
  NAND2HSV4 U15534 ( .A1(n15580), .A2(n15579), .ZN(n28933) );
  NAND2HSV2 U15535 ( .A1(n20344), .A2(n20345), .ZN(n20350) );
  INHSV6 U15536 ( .I(n18604), .ZN(n28790) );
  NAND2HSV2 U15537 ( .A1(n27290), .A2(n27289), .ZN(n28701) );
  CLKNAND2HSV2 U15538 ( .A1(n13753), .A2(n25269), .ZN(n13755) );
  XNOR2HSV1 U15539 ( .A1(n23903), .A2(n23902), .ZN(n23906) );
  INHSV4 U15540 ( .I(n19710), .ZN(n24214) );
  XNOR2HSV1 U15541 ( .A1(n27870), .A2(n27869), .ZN(n27873) );
  XNOR2HSV1 U15542 ( .A1(n27899), .A2(n27898), .ZN(n27902) );
  MUX2NHSV1 U15543 ( .I0(n13760), .I1(n23843), .S(n13761), .ZN(\pe7/poht [10])
         );
  NAND2HSV4 U15544 ( .A1(n17168), .A2(n17615), .ZN(n17240) );
  OAI21HSV2 U15545 ( .A1(n16206), .A2(n16204), .B(n16205), .ZN(n16207) );
  AOI21HSV2 U15546 ( .A1(n16201), .A2(n16200), .B(n16199), .ZN(n16202) );
  NAND2HSV2 U15547 ( .A1(n16232), .A2(n16231), .ZN(n16219) );
  CLKNHSV0 U15548 ( .I(\pe6/phq [14]), .ZN(n12776) );
  NAND2HSV0 U15549 ( .A1(\pe6/pvq [14]), .A2(n22109), .ZN(n12777) );
  MUX2NHSV1 U15550 ( .I0(\pe6/phq [14]), .I1(n12776), .S(n12777), .ZN(n19079)
         );
  XOR2HSV0 U15551 ( .A1(n18304), .A2(n18305), .Z(n12778) );
  XOR2HSV0 U15552 ( .A1(n18300), .A2(n18299), .Z(n12779) );
  XOR2HSV0 U15553 ( .A1(n12778), .A2(n12779), .Z(n12780) );
  NAND2HSV0 U15554 ( .A1(\pe9/got [8]), .A2(n28110), .ZN(n12781) );
  CLKNAND2HSV0 U15555 ( .A1(n12781), .A2(n12780), .ZN(n12782) );
  OAI21HSV0 U15556 ( .A1(n12780), .A2(n12781), .B(n12782), .ZN(n12783) );
  NAND2HSV0 U15557 ( .A1(n28688), .A2(\pe9/got [7]), .ZN(n12784) );
  CLKNAND2HSV0 U15558 ( .A1(n12784), .A2(n12783), .ZN(n12785) );
  OAI21HSV0 U15559 ( .A1(n12783), .A2(n12784), .B(n12785), .ZN(n12786) );
  NAND2HSV0 U15560 ( .A1(n28804), .A2(\pe9/got [9]), .ZN(n12787) );
  NAND2HSV0 U15561 ( .A1(n12787), .A2(n12786), .ZN(n12788) );
  OAI21HSV2 U15562 ( .A1(n12786), .A2(n12787), .B(n12788), .ZN(n18306) );
  CLKNHSV0 U15563 ( .I(n19714), .ZN(n12789) );
  NAND2HSV0 U15564 ( .A1(\pe7/pvq [14]), .A2(n27087), .ZN(n12790) );
  NAND2HSV0 U15565 ( .A1(n12790), .A2(\pe7/phq [14]), .ZN(n12791) );
  OAI21HSV2 U15566 ( .A1(\pe7/phq [14]), .A2(n12790), .B(n12791), .ZN(n12792)
         );
  MUX2NHSV1 U15567 ( .I0(n12789), .I1(n19714), .S(n12792), .ZN(n19722) );
  NAND2HSV0 U15568 ( .A1(n14199), .A2(n14198), .ZN(n12794) );
  MUX2NHSV2 U15569 ( .I0(n14200), .I1(n12793), .S(n12794), .ZN(n14213) );
  XOR2HSV0 U15570 ( .A1(n19564), .A2(n19563), .Z(n12796) );
  NAND2HSV0 U15571 ( .A1(n14022), .A2(n25270), .ZN(n12797) );
  CLKNAND2HSV0 U15572 ( .A1(n12797), .A2(n12796), .ZN(n12798) );
  OAI21HSV0 U15573 ( .A1(n12796), .A2(n12797), .B(n12798), .ZN(n12799) );
  NAND2HSV0 U15574 ( .A1(\pe7/got [12]), .A2(n19711), .ZN(n12800) );
  CLKNAND2HSV0 U15575 ( .A1(n12800), .A2(n12799), .ZN(n12801) );
  OAI21HSV2 U15576 ( .A1(n12799), .A2(n12800), .B(n12801), .ZN(n12802) );
  OAI21HSV2 U15577 ( .A1(n12802), .A2(n12803), .B(n12804), .ZN(n19577) );
  NAND3HSV0 U15578 ( .A1(n15688), .A2(n15370), .A3(n15628), .ZN(n12805) );
  NOR2HSV4 U15579 ( .A1(n12805), .A2(n15629), .ZN(n15698) );
  CLKNHSV0 U15580 ( .I(n24328), .ZN(n12806) );
  XOR2HSV0 U15581 ( .A1(n21561), .A2(n21559), .Z(n12807) );
  XOR2HSV0 U15582 ( .A1(n21556), .A2(n21555), .Z(n12808) );
  XOR2HSV0 U15583 ( .A1(n12807), .A2(n12808), .Z(n12809) );
  MUX2NHSV0 U15584 ( .I0(n12806), .I1(n24328), .S(n12809), .ZN(n12810) );
  OAI21HSV0 U15585 ( .A1(n24638), .A2(n24686), .B(n12810), .ZN(n12811) );
  OAI31HSV0 U15586 ( .A1(n24638), .A2(n12810), .A3(n24686), .B(n12811), .ZN(
        n12812) );
  NAND2HSV0 U15587 ( .A1(\pe5/got [2]), .A2(\pe5/ti_7[10] ), .ZN(n12813) );
  NAND2HSV0 U15588 ( .A1(n12813), .A2(n12812), .ZN(n12814) );
  OAI21HSV2 U15589 ( .A1(n12812), .A2(n12813), .B(n12814), .ZN(n21563) );
  INHSV2 U15590 ( .I(n21295), .ZN(n12815) );
  MUX2NHSV2 U15591 ( .I0(n12815), .I1(n21295), .S(n12816), .ZN(n21708) );
  CLKNHSV0 U15592 ( .I(n22128), .ZN(n12817) );
  AOI21HSV0 U15593 ( .A1(n18776), .A2(n29006), .B(n12817), .ZN(n18768) );
  CLKNHSV0 U15594 ( .I(n19707), .ZN(n12818) );
  AOI21HSV0 U15595 ( .A1(n16956), .A2(n16641), .B(n25256), .ZN(n12819) );
  NAND2HSV0 U15596 ( .A1(n23336), .A2(\pe3/aot [2]), .ZN(n12821) );
  OAI21HSV0 U15597 ( .A1(n24535), .A2(n24581), .B(n12821), .ZN(n12822) );
  OAI31HSV2 U15598 ( .A1(n24535), .A2(n12821), .A3(n24581), .B(n12822), .ZN(
        n12823) );
  NAND2HSV0 U15599 ( .A1(n14040), .A2(\pe3/bq[2] ), .ZN(n12824) );
  NAND2HSV0 U15600 ( .A1(n12824), .A2(n12823), .ZN(n12825) );
  OAI21HSV0 U15601 ( .A1(n12823), .A2(n12824), .B(n12825), .ZN(n12826) );
  NAND2HSV0 U15602 ( .A1(n11932), .A2(\pe3/bq[5] ), .ZN(n12827) );
  CLKNAND2HSV0 U15603 ( .A1(n12827), .A2(n12826), .ZN(n12828) );
  OAI21HSV0 U15604 ( .A1(n12826), .A2(n12827), .B(n12828), .ZN(n23337) );
  AOI21HSV0 U15605 ( .A1(n27082), .A2(\pe7/pvq [10]), .B(\pe7/phq [10]), .ZN(
        n12829) );
  AO31HSV2 U15606 ( .A1(n27082), .A2(\pe7/pvq [10]), .A3(\pe7/phq [10]), .B(
        n12829), .Z(n19398) );
  XOR2HSV0 U15607 ( .A1(n19722), .A2(n19723), .Z(n12830) );
  XOR2HSV0 U15608 ( .A1(n19738), .A2(n19721), .Z(n12831) );
  NAND2HSV0 U15609 ( .A1(n25292), .A2(n25375), .ZN(n12833) );
  OAI21HSV2 U15610 ( .A1(n12832), .A2(n12833), .B(n12834), .ZN(n12835) );
  XOR2HSV0 U15611 ( .A1(n19737), .A2(n19736), .Z(n12836) );
  CLKXOR2HSV2 U15612 ( .A1(n12835), .A2(n12836), .Z(n12837) );
  NAND2HSV0 U15613 ( .A1(n24250), .A2(\pe7/got [6]), .ZN(n12838) );
  NAND2HSV2 U15614 ( .A1(n12838), .A2(n12837), .ZN(n12839) );
  OAI21HSV2 U15615 ( .A1(n12837), .A2(n12838), .B(n12839), .ZN(n19741) );
  CLKNHSV0 U15616 ( .I(\pe6/pvq [9]), .ZN(n12840) );
  OAI21HSV2 U15617 ( .A1(n27074), .A2(n12840), .B(\pe6/phq [9]), .ZN(n12841)
         );
  OAI31HSV2 U15618 ( .A1(n27074), .A2(\pe6/phq [9]), .A3(n12840), .B(n12841), 
        .ZN(n14379) );
  XOR2HSV0 U15619 ( .A1(n20389), .A2(n20390), .Z(n12842) );
  XOR2HSV0 U15620 ( .A1(n20376), .A2(n20375), .Z(n12843) );
  NAND2HSV0 U15621 ( .A1(n28807), .A2(n14049), .ZN(n12845) );
  NAND2HSV2 U15622 ( .A1(n12845), .A2(n12844), .ZN(n12846) );
  OAI21HSV2 U15623 ( .A1(n12844), .A2(n12845), .B(n12846), .ZN(n12847) );
  NAND2HSV0 U15624 ( .A1(n20467), .A2(n20292), .ZN(n12848) );
  NAND2HSV2 U15625 ( .A1(n12848), .A2(n12847), .ZN(n12849) );
  OAI21HSV2 U15626 ( .A1(n12847), .A2(n12848), .B(n12849), .ZN(n20392) );
  INOR2HSV0 U15627 ( .A1(\pe9/ti_7t [6]), .B1(n17998), .ZN(n18086) );
  NAND2HSV0 U15628 ( .A1(n19127), .A2(n19128), .ZN(n12850) );
  NOR2HSV0 U15629 ( .A1(n19129), .A2(n14123), .ZN(n12851) );
  INOR2HSV1 U15630 ( .A1(n18538), .B1(n25682), .ZN(n13988) );
  CLKNHSV0 U15631 ( .I(n19612), .ZN(n12852) );
  INHSV2 U15632 ( .I(n16419), .ZN(n12853) );
  MUX2NHSV2 U15633 ( .I0(n16419), .I1(n12853), .S(n12854), .ZN(n16420) );
  CLKNHSV0 U15634 ( .I(n24443), .ZN(n12855) );
  XOR2HSV0 U15635 ( .A1(n24441), .A2(n24442), .Z(n12856) );
  XOR2HSV0 U15636 ( .A1(n24438), .A2(n24437), .Z(n12857) );
  XOR2HSV0 U15637 ( .A1(n12856), .A2(n12857), .Z(n12858) );
  NAND2HSV0 U15638 ( .A1(\pe5/aot [3]), .A2(\pe5/bq[4] ), .ZN(n12859) );
  CLKNAND2HSV0 U15639 ( .A1(n12859), .A2(n12858), .ZN(n12860) );
  OAI21HSV0 U15640 ( .A1(n12858), .A2(n12859), .B(n12860), .ZN(n12861) );
  MUX2NHSV0 U15641 ( .I0(n24443), .I1(n12855), .S(n12861), .ZN(n12862) );
  NAND2HSV0 U15642 ( .A1(n28640), .A2(\pe5/ti_7[10] ), .ZN(n12863) );
  NAND2HSV0 U15643 ( .A1(n12863), .A2(n12862), .ZN(n12864) );
  OAI21HSV2 U15644 ( .A1(n12862), .A2(n12863), .B(n12864), .ZN(n24445) );
  OA21HSV2 U15645 ( .A1(n25494), .A2(\pe7/ti_7t [5]), .B(n28610), .Z(n19319)
         );
  INOR2HSV0 U15646 ( .A1(\pe11/ti_7t [11]), .B1(n20636), .ZN(n23450) );
  NAND2HSV0 U15647 ( .A1(\pe9/bq[4] ), .A2(\pe9/aot [15]), .ZN(n12865) );
  AOI21HSV0 U15648 ( .A1(\pe9/got [3]), .A2(n28019), .B(n12865), .ZN(n12866)
         );
  AO31HSV0 U15649 ( .A1(\pe9/got [3]), .A2(n28019), .A3(n12865), .B(n12866), 
        .Z(n18572) );
  NAND2HSV0 U15650 ( .A1(n21335), .A2(\pe3/pvq [15]), .ZN(n12867) );
  NAND2HSV0 U15651 ( .A1(n12867), .A2(\pe3/phq [15]), .ZN(n12868) );
  OAI21HSV0 U15652 ( .A1(\pe3/phq [15]), .A2(n12867), .B(n12868), .ZN(n23346)
         );
  CLKNAND2HSV2 U15653 ( .A1(\pe8/pvq [8]), .A2(n14036), .ZN(n12869) );
  NAND2HSV2 U15654 ( .A1(n12869), .A2(\pe8/phq [8]), .ZN(n12870) );
  OAI21HSV2 U15655 ( .A1(\pe8/phq [8]), .A2(n12869), .B(n12870), .ZN(n12871)
         );
  NAND2HSV0 U15656 ( .A1(\pe8/aot [11]), .A2(n23627), .ZN(n12872) );
  NAND2HSV2 U15657 ( .A1(n12872), .A2(n12871), .ZN(n12873) );
  OAI21HSV2 U15658 ( .A1(n12871), .A2(n12872), .B(n12873), .ZN(n16525) );
  NAND2HSV2 U15659 ( .A1(\pe5/pvq [4]), .A2(n27050), .ZN(n12874) );
  NAND2HSV0 U15660 ( .A1(n18227), .A2(n18029), .ZN(n12875) );
  NOR2HSV4 U15661 ( .A1(n18229), .A2(n12875), .ZN(n18138) );
  INAND2HSV2 U15662 ( .A1(n19678), .B1(n19702), .ZN(n13990) );
  NOR2HSV4 U15663 ( .A1(n14676), .A2(n14616), .ZN(n21347) );
  CLKNAND2HSV0 U15664 ( .A1(n12876), .A2(n19508), .ZN(n12877) );
  INHSV2 U15665 ( .I(n20314), .ZN(n12879) );
  XOR2HSV0 U15666 ( .A1(n22274), .A2(n22273), .Z(n12880) );
  NAND2HSV0 U15667 ( .A1(\pe8/got [6]), .A2(n14059), .ZN(n12881) );
  CLKNAND2HSV0 U15668 ( .A1(n12881), .A2(n12880), .ZN(n12882) );
  OAI21HSV0 U15669 ( .A1(n12880), .A2(n12881), .B(n12882), .ZN(n12883) );
  NAND2HSV0 U15670 ( .A1(n14060), .A2(n28706), .ZN(n12884) );
  CLKNAND2HSV0 U15671 ( .A1(n12884), .A2(n12883), .ZN(n12885) );
  OAI21HSV0 U15672 ( .A1(n12883), .A2(n12884), .B(n12885), .ZN(n12886) );
  NAND2HSV0 U15673 ( .A1(\pe8/got [8]), .A2(n25185), .ZN(n12887) );
  CLKNAND2HSV0 U15674 ( .A1(n12887), .A2(n12886), .ZN(n12888) );
  OAI21HSV0 U15675 ( .A1(n12886), .A2(n12887), .B(n12888), .ZN(n12889) );
  NAND2HSV0 U15676 ( .A1(n23757), .A2(\pe8/got [9]), .ZN(n12890) );
  NAND2HSV0 U15677 ( .A1(n12889), .A2(n12890), .ZN(n12891) );
  OAI21HSV0 U15678 ( .A1(n12889), .A2(n12890), .B(n12891), .ZN(n22275) );
  NAND2HSV0 U15679 ( .A1(\pe9/aot [5]), .A2(\pe9/bq[16] ), .ZN(n12893) );
  OAI21HSV0 U15680 ( .A1(n18407), .A2(n27101), .B(n12893), .ZN(n12894) );
  OAI31HSV0 U15681 ( .A1(n18407), .A2(n12893), .A3(n27101), .B(n12894), .ZN(
        n18411) );
  CLKNHSV0 U15682 ( .I(\pe3/phq [7]), .ZN(n12895) );
  NAND2HSV4 U15683 ( .A1(\pe3/pvq [7]), .A2(n21335), .ZN(n12896) );
  MUX2NHSV2 U15684 ( .I0(\pe3/phq [7]), .I1(n12895), .S(n12896), .ZN(n15107)
         );
  NAND2HSV0 U15685 ( .A1(\pe2/pvq [12]), .A2(n21253), .ZN(n12897) );
  NAND2HSV0 U15686 ( .A1(n12897), .A2(\pe2/phq [12]), .ZN(n12898) );
  OAI21HSV2 U15687 ( .A1(\pe2/phq [12]), .A2(n12897), .B(n12898), .ZN(n21255)
         );
  NAND2HSV0 U15688 ( .A1(\pe7/aot [10]), .A2(\pe7/bq[8] ), .ZN(n12899) );
  NAND2HSV0 U15689 ( .A1(\pe7/bq[11] ), .A2(\pe7/aot [7]), .ZN(n12900) );
  NAND2HSV0 U15690 ( .A1(n12900), .A2(n12899), .ZN(n12901) );
  OAI21HSV2 U15691 ( .A1(n12899), .A2(n12900), .B(n12901), .ZN(n12902) );
  NAND2HSV0 U15692 ( .A1(\pe7/bq[14] ), .A2(\pe7/aot [4]), .ZN(n12903) );
  NAND2HSV2 U15693 ( .A1(n12903), .A2(n12902), .ZN(n12904) );
  OAI21HSV2 U15694 ( .A1(n12902), .A2(n12903), .B(n12904), .ZN(n12905) );
  NAND2HSV0 U15695 ( .A1(\pe7/aot [5]), .A2(\pe7/bq[13] ), .ZN(n12906) );
  CLKNAND2HSV0 U15696 ( .A1(n12906), .A2(n12905), .ZN(n12907) );
  OAI21HSV2 U15697 ( .A1(n12905), .A2(n12906), .B(n12907), .ZN(n23145) );
  NAND2HSV0 U15698 ( .A1(n22129), .A2(n18784), .ZN(n12908) );
  INHSV4 U15699 ( .I(n19054), .ZN(n12909) );
  MUX2NHSV4 U15700 ( .I0(n19054), .I1(n12909), .S(n19053), .ZN(n19070) );
  NAND2HSV2 U15701 ( .A1(n19615), .A2(n19616), .ZN(n12910) );
  CLKNHSV0 U15702 ( .I(n24329), .ZN(n12911) );
  MUX2NHSV0 U15703 ( .I0(n12911), .I1(n24329), .S(n23234), .ZN(n12912) );
  XOR2HSV0 U15704 ( .A1(n23235), .A2(n12912), .Z(n12913) );
  NAND2HSV2 U15705 ( .A1(n12914), .A2(n12913), .ZN(n12915) );
  OAI21HSV2 U15706 ( .A1(n12913), .A2(n12914), .B(n12915), .ZN(n23238) );
  XOR2HSV0 U15707 ( .A1(n22221), .A2(n22220), .Z(n12916) );
  NAND2HSV0 U15708 ( .A1(n25204), .A2(\pe8/got [5]), .ZN(n12917) );
  CLKNAND2HSV0 U15709 ( .A1(n12917), .A2(n12916), .ZN(n12918) );
  OAI21HSV0 U15710 ( .A1(n12916), .A2(n12917), .B(n12918), .ZN(n12919) );
  NAND2HSV0 U15711 ( .A1(\pe8/got [6]), .A2(n28698), .ZN(n12920) );
  NAND2HSV0 U15712 ( .A1(n12920), .A2(n12919), .ZN(n12921) );
  OAI21HSV0 U15713 ( .A1(n12919), .A2(n12920), .B(n12921), .ZN(n12922) );
  NAND2HSV0 U15714 ( .A1(n14060), .A2(n23757), .ZN(n12923) );
  NAND2HSV0 U15715 ( .A1(n12923), .A2(n12922), .ZN(n12924) );
  NAND2HSV0 U15716 ( .A1(n28652), .A2(n26751), .ZN(n12926) );
  CLKNAND2HSV0 U15717 ( .A1(n12926), .A2(n12925), .ZN(n12927) );
  OAI21HSV0 U15718 ( .A1(n12925), .A2(n12926), .B(n12927), .ZN(n12928) );
  NAND2HSV0 U15719 ( .A1(n26760), .A2(\pe3/got [4]), .ZN(n12929) );
  CLKNAND2HSV0 U15720 ( .A1(n12929), .A2(n12928), .ZN(n12930) );
  OAI21HSV0 U15721 ( .A1(n12928), .A2(n12929), .B(n12930), .ZN(n12931) );
  NAND2HSV0 U15722 ( .A1(\pe3/got [5]), .A2(n28661), .ZN(n12932) );
  NAND2HSV0 U15723 ( .A1(n12932), .A2(n12931), .ZN(n12933) );
  OAI21HSV0 U15724 ( .A1(n12931), .A2(n12932), .B(n12933), .ZN(\pe3/poht [11])
         );
  OAI21HSV0 U15725 ( .A1(n23546), .A2(n28199), .B(n18301), .ZN(n12934) );
  OAI21HSV0 U15726 ( .A1(n18302), .A2(n22377), .B(n12934), .ZN(n12935) );
  CLKNAND2HSV0 U15727 ( .A1(\pe9/pvq [11]), .A2(n27078), .ZN(n12936) );
  NAND2HSV2 U15728 ( .A1(n12936), .A2(\pe9/phq [11]), .ZN(n12937) );
  OAI21HSV2 U15729 ( .A1(\pe9/phq [11]), .A2(n12936), .B(n12937), .ZN(n12938)
         );
  NAND2HSV2 U15730 ( .A1(n12935), .A2(n12938), .ZN(n12939) );
  OAI21HSV2 U15731 ( .A1(n12935), .A2(n12938), .B(n12939), .ZN(n18305) );
  INOR2HSV1 U15732 ( .A1(n20953), .B1(n23255), .ZN(n20955) );
  CLKNHSV0 U15733 ( .I(\pe4/phq [7]), .ZN(n12940) );
  NAND2HSV4 U15734 ( .A1(\pe4/pvq [7]), .A2(n27105), .ZN(n12941) );
  MUX2NHSV2 U15735 ( .I0(\pe4/phq [7]), .I1(n12940), .S(n12941), .ZN(n15435)
         );
  CLKNHSV0 U15736 ( .I(\pe6/phq [10]), .ZN(n12942) );
  NAND2HSV2 U15737 ( .A1(\pe6/pvq [10]), .A2(n23498), .ZN(n12943) );
  MUX2NHSV2 U15738 ( .I0(\pe6/phq [10]), .I1(n12942), .S(n12943), .ZN(n14417)
         );
  NAND2HSV2 U15739 ( .A1(\pe2/pvq [14]), .A2(n23539), .ZN(n12944) );
  NAND2HSV2 U15740 ( .A1(n12944), .A2(\pe2/phq [14]), .ZN(n12945) );
  OAI21HSV2 U15741 ( .A1(\pe2/phq [14]), .A2(n12944), .B(n12945), .ZN(n12946)
         );
  NAND2HSV0 U15742 ( .A1(\pe2/aot [8]), .A2(\pe2/bq[11] ), .ZN(n12947) );
  NAND2HSV2 U15743 ( .A1(n12947), .A2(n12946), .ZN(n12948) );
  OAI21HSV2 U15744 ( .A1(n12946), .A2(n12947), .B(n12948), .ZN(n21655) );
  CLKNHSV0 U15745 ( .I(\pe7/phq [12]), .ZN(n12949) );
  NAND2HSV2 U15746 ( .A1(\pe7/pvq [12]), .A2(n27099), .ZN(n12950) );
  MUX2NHSV1 U15747 ( .I0(\pe7/phq [12]), .I1(n12949), .S(n12950), .ZN(n19553)
         );
  AOI22HSV0 U15748 ( .A1(\pe10/bq[2] ), .A2(\pe10/aot [14]), .B1(
        \pe10/aot [12]), .B2(\pe10/bq[4] ), .ZN(n12951) );
  IAO21HSV2 U15749 ( .A1(n22527), .A2(n24465), .B(n12951), .ZN(n12952) );
  NAND2HSV0 U15750 ( .A1(\pe10/bq[3] ), .A2(\pe10/aot [13]), .ZN(n12953) );
  CLKNAND2HSV0 U15751 ( .A1(n12953), .A2(n12952), .ZN(n12954) );
  OAI21HSV2 U15752 ( .A1(n12952), .A2(n12953), .B(n12954), .ZN(n22528) );
  NOR2HSV4 U15753 ( .A1(n14077), .A2(\pe7/phq [2]), .ZN(n12955) );
  INAND2HSV0 U15754 ( .A1(\pe11/ti_7t [10]), .B1(ctro11), .ZN(n20562) );
  INHSV2 U15755 ( .I(n18213), .ZN(n12956) );
  AOI21HSV0 U15756 ( .A1(n18212), .A2(n18211), .B(n12956), .ZN(n18218) );
  CLKNHSV0 U15757 ( .I(n17109), .ZN(n12957) );
  CLKNHSV0 U15758 ( .I(\pe5/ti_7t [1]), .ZN(n12959) );
  AOI21HSV0 U15759 ( .A1(n21412), .A2(n12959), .B(n21411), .ZN(n12960) );
  OAI21HSV0 U15760 ( .A1(n28455), .A2(n14616), .B(n12960), .ZN(n14508) );
  NAND2HSV0 U15761 ( .A1(n28812), .A2(n15423), .ZN(n12961) );
  OAI21HSV2 U15762 ( .A1(n29033), .A2(n28812), .B(n12961), .ZN(n15723) );
  NAND3HSV0 U15763 ( .A1(n26923), .A2(n26924), .A3(n26918), .ZN(n26926) );
  INHSV4 U15764 ( .I(n18465), .ZN(n12962) );
  MUX2NHSV4 U15765 ( .I0(n12962), .I1(n18465), .S(n12963), .ZN(n18648) );
  INOR2HSV1 U15766 ( .A1(n21898), .B1(n21899), .ZN(n21900) );
  CLKNHSV0 U15767 ( .I(n26683), .ZN(n12964) );
  NAND2HSV0 U15768 ( .A1(\pe3/aot [5]), .A2(\pe3/bq[1] ), .ZN(n12965) );
  CLKNAND2HSV0 U15769 ( .A1(n12965), .A2(n23673), .ZN(n12966) );
  OAI21HSV0 U15770 ( .A1(n23673), .A2(n12965), .B(n12966), .ZN(n12967) );
  NAND2HSV0 U15771 ( .A1(\pe3/aot [2]), .A2(\pe3/bq[4] ), .ZN(n12968) );
  CLKNAND2HSV0 U15772 ( .A1(n12968), .A2(n12967), .ZN(n12969) );
  OAI21HSV0 U15773 ( .A1(n12967), .A2(n12968), .B(n12969), .ZN(n12970) );
  MUX2NHSV0 U15774 ( .I0(n26683), .I1(n12964), .S(n12970), .ZN(n12971) );
  NAND2HSV0 U15775 ( .A1(\pe3/got [1]), .A2(n28584), .ZN(n12972) );
  NAND2HSV0 U15776 ( .A1(n12972), .A2(n12971), .ZN(n12973) );
  OAI21HSV0 U15777 ( .A1(n12971), .A2(n12972), .B(n12973), .ZN(n23674) );
  NAND2HSV0 U15778 ( .A1(n25186), .A2(\pe8/got [2]), .ZN(n12974) );
  NAND2HSV0 U15779 ( .A1(n14059), .A2(\pe8/got [3]), .ZN(n12976) );
  NAND2HSV0 U15780 ( .A1(n12976), .A2(n12975), .ZN(n12977) );
  OAI21HSV0 U15781 ( .A1(n12975), .A2(n12976), .B(n12977), .ZN(n12978) );
  NAND2HSV0 U15782 ( .A1(n25203), .A2(n25204), .ZN(n12979) );
  NAND2HSV0 U15783 ( .A1(n12979), .A2(n12978), .ZN(n12980) );
  OAI21HSV0 U15784 ( .A1(n12978), .A2(n12979), .B(n12980), .ZN(n25205) );
  CLKNAND2HSV0 U15785 ( .A1(n12982), .A2(n12981), .ZN(n12983) );
  OAI21HSV0 U15786 ( .A1(n12981), .A2(n12982), .B(n12983), .ZN(\pe5/poht [9])
         );
  NAND2HSV0 U15787 ( .A1(n26729), .A2(n15157), .ZN(n12985) );
  CLKNAND2HSV0 U15788 ( .A1(n12985), .A2(n12984), .ZN(n12986) );
  OAI21HSV0 U15789 ( .A1(n12984), .A2(n12985), .B(n12986), .ZN(n12987) );
  NAND2HSV0 U15790 ( .A1(n26600), .A2(n26413), .ZN(n12988) );
  CLKNAND2HSV0 U15791 ( .A1(n12988), .A2(n12987), .ZN(n12989) );
  OAI21HSV0 U15792 ( .A1(n12987), .A2(n12988), .B(n12989), .ZN(po3) );
  NAND2HSV0 U15793 ( .A1(\pe11/aot [5]), .A2(n24997), .ZN(n12990) );
  NAND2HSV0 U15794 ( .A1(\pe11/aot [11]), .A2(\pe11/bq[9] ), .ZN(n12991) );
  NAND2HSV0 U15795 ( .A1(n12991), .A2(n12990), .ZN(n12992) );
  OAI21HSV0 U15796 ( .A1(n12990), .A2(n12991), .B(n12992), .ZN(n20657) );
  XOR2HSV0 U15797 ( .A1(n19908), .A2(n19909), .Z(n12993) );
  XOR2HSV0 U15798 ( .A1(n19907), .A2(n19906), .Z(n12994) );
  XOR2HSV0 U15799 ( .A1(n12993), .A2(n12994), .Z(n12995) );
  XOR2HSV0 U15800 ( .A1(n19916), .A2(n19917), .Z(n12996) );
  XOR2HSV0 U15801 ( .A1(n19915), .A2(n19914), .Z(n12997) );
  XOR2HSV0 U15802 ( .A1(n12996), .A2(n12997), .Z(n12998) );
  XOR2HSV0 U15803 ( .A1(n19918), .A2(\pe8/phq [13]), .Z(n12999) );
  OAI21HSV0 U15804 ( .A1(n19921), .A2(n23731), .B(n19920), .ZN(n13000) );
  CLKNAND2HSV0 U15805 ( .A1(n13000), .A2(n12999), .ZN(n13001) );
  OAI21HSV2 U15806 ( .A1(n13000), .A2(n12999), .B(n13001), .ZN(n13002) );
  XOR2HSV0 U15807 ( .A1(n13002), .A2(n12998), .Z(n13003) );
  XOR2HSV0 U15808 ( .A1(n19913), .A2(n19912), .Z(n13004) );
  XOR2HSV0 U15809 ( .A1(n13003), .A2(n13004), .Z(n13005) );
  XOR2HSV0 U15810 ( .A1(n12995), .A2(n13005), .Z(n19922) );
  NAND2HSV0 U15811 ( .A1(\pe3/aot [14]), .A2(\pe3/bq[15] ), .ZN(n13006) );
  NAND2HSV2 U15812 ( .A1(n13006), .A2(\pe3/phq [4]), .ZN(n13007) );
  OAI21HSV2 U15813 ( .A1(\pe3/phq [4]), .A2(n13006), .B(n13007), .ZN(n15073)
         );
  CLKNHSV0 U15814 ( .I(\pe2/phq [13]), .ZN(n13008) );
  NAND2HSV0 U15815 ( .A1(n23539), .A2(\pe2/pvq [13]), .ZN(n13009) );
  MUX2NHSV1 U15816 ( .I0(n13008), .I1(\pe2/phq [13]), .S(n13009), .ZN(n21090)
         );
  XOR2HSV0 U15817 ( .A1(n17557), .A2(n17556), .Z(n13010) );
  XOR2HSV0 U15818 ( .A1(n27021), .A2(n26556), .Z(n13011) );
  XOR2HSV0 U15819 ( .A1(n13010), .A2(n13011), .Z(n17559) );
  AOI22HSV0 U15820 ( .A1(\pe10/aot [3]), .A2(\pe10/bq[13] ), .B1(\pe10/bq[14] ), .B2(\pe10/aot [2]), .ZN(n13012) );
  AOI21HSV0 U15821 ( .A1(n26106), .A2(n26164), .B(n13012), .ZN(n22530) );
  CLKNAND2HSV2 U15822 ( .A1(\pe7/pvq [8]), .A2(n27096), .ZN(n13013) );
  NAND2HSV2 U15823 ( .A1(n13013), .A2(\pe7/phq [8]), .ZN(n13014) );
  OAI21HSV2 U15824 ( .A1(\pe7/phq [8]), .A2(n13013), .B(n13014), .ZN(n13015)
         );
  NAND2HSV0 U15825 ( .A1(\pe7/aot [10]), .A2(\pe7/bq[15] ), .ZN(n13016) );
  NAND2HSV2 U15826 ( .A1(n13016), .A2(n13015), .ZN(n13017) );
  OAI21HSV2 U15827 ( .A1(n13015), .A2(n13016), .B(n13017), .ZN(n19434) );
  NAND2HSV0 U15828 ( .A1(\pe2/bq[8] ), .A2(\pe2/aot [15]), .ZN(n13018) );
  AOI21HSV2 U15829 ( .A1(\pe2/got [7]), .A2(n21269), .B(n13018), .ZN(n13019)
         );
  AO31HSV0 U15830 ( .A1(\pe2/got [7]), .A2(n21269), .A3(n13018), .B(n13019), 
        .Z(n21121) );
  INAND2HSV0 U15831 ( .A1(\pe4/ti_7t [7]), .B1(n15534), .ZN(n15638) );
  CLKNHSV0 U15832 ( .I(\pe3/phq [5]), .ZN(n13020) );
  NAND2HSV0 U15833 ( .A1(\pe3/pvq [5]), .A2(n23541), .ZN(n13021) );
  MUX2NHSV0 U15834 ( .I0(\pe3/phq [5]), .I1(n13020), .S(n13021), .ZN(n15130)
         );
  NAND2HSV0 U15835 ( .A1(\pe5/aot [14]), .A2(\pe5/bq[3] ), .ZN(n13022) );
  OAI21HSV0 U15836 ( .A1(n23923), .A2(n21493), .B(n13022), .ZN(n13023) );
  OAI31HSV0 U15837 ( .A1(n23923), .A2(n13022), .A3(n21493), .B(n13023), .ZN(
        n13024) );
  NAND2HSV0 U15838 ( .A1(\pe5/aot [10]), .A2(\pe5/bq[7] ), .ZN(n13025) );
  NAND2HSV0 U15839 ( .A1(n13025), .A2(n13024), .ZN(n13026) );
  OAI21HSV0 U15840 ( .A1(n13024), .A2(n13025), .B(n13026), .ZN(n13027) );
  NAND2HSV0 U15841 ( .A1(\pe5/aot [11]), .A2(\pe5/bq[6] ), .ZN(n13028) );
  CLKNAND2HSV0 U15842 ( .A1(n13028), .A2(n13027), .ZN(n13029) );
  OAI21HSV0 U15843 ( .A1(n13027), .A2(n13028), .B(n13029), .ZN(n21494) );
  INAND2HSV0 U15844 ( .A1(\pe9/ti_7t [7]), .B1(n18628), .ZN(n18225) );
  NAND2HSV0 U15845 ( .A1(n26924), .A2(n22792), .ZN(n13030) );
  INHSV4 U15846 ( .I(n16384), .ZN(n13031) );
  NOR2HSV4 U15847 ( .A1(n16364), .A2(n16363), .ZN(n13032) );
  MUX2NHSV4 U15848 ( .I0(n16384), .I1(n13031), .S(n13032), .ZN(n16430) );
  CLKNHSV0 U15849 ( .I(n18785), .ZN(n13033) );
  OAI21HSV4 U15850 ( .A1(n29006), .A2(n13033), .B(n18776), .ZN(n21315) );
  NOR2HSV0 U15851 ( .A1(n21116), .A2(n21236), .ZN(n13034) );
  OAI21HSV2 U15852 ( .A1(n21239), .A2(n21149), .B(n13034), .ZN(n21152) );
  XOR2HSV0 U15853 ( .A1(n26208), .A2(n26207), .Z(n13035) );
  NAND2HSV0 U15854 ( .A1(n28585), .A2(n28644), .ZN(n13036) );
  CLKNAND2HSV0 U15855 ( .A1(n13036), .A2(n13035), .ZN(n13037) );
  OAI21HSV2 U15856 ( .A1(n13035), .A2(n13036), .B(n13037), .ZN(n13038) );
  NAND2HSV0 U15857 ( .A1(n26214), .A2(n26215), .ZN(n13039) );
  NAND2HSV0 U15858 ( .A1(n27197), .A2(\pe10/got [13]), .ZN(n13043) );
  XOR2HSV0 U15859 ( .A1(n23900), .A2(n23899), .Z(n13045) );
  XOR2HSV0 U15860 ( .A1(n23898), .A2(n13045), .Z(n13046) );
  NAND2HSV0 U15861 ( .A1(\pe7/got [5]), .A2(n11978), .ZN(n13047) );
  CLKNAND2HSV0 U15862 ( .A1(n13047), .A2(n13046), .ZN(n13048) );
  OAI21HSV0 U15863 ( .A1(n13046), .A2(n13047), .B(n13048), .ZN(n13049) );
  NAND2HSV0 U15864 ( .A1(n25397), .A2(\pe7/got [6]), .ZN(n13050) );
  CLKNAND2HSV0 U15865 ( .A1(n13050), .A2(n13049), .ZN(n13051) );
  OAI21HSV0 U15866 ( .A1(n13049), .A2(n13050), .B(n13051), .ZN(n13052) );
  NAND2HSV0 U15867 ( .A1(\pe7/got [7]), .A2(n28656), .ZN(n13053) );
  CLKNAND2HSV0 U15868 ( .A1(n13053), .A2(n13052), .ZN(n13054) );
  OAI21HSV0 U15869 ( .A1(n13052), .A2(n13053), .B(n13054), .ZN(n13055) );
  NAND2HSV0 U15870 ( .A1(\pe7/got [8]), .A2(n25376), .ZN(n13056) );
  NAND2HSV0 U15871 ( .A1(n13056), .A2(n13055), .ZN(n13057) );
  OAI21HSV2 U15872 ( .A1(n13055), .A2(n13056), .B(n13057), .ZN(n23903) );
  NAND2HSV0 U15873 ( .A1(n20770), .A2(n24881), .ZN(n13058) );
  NAND2HSV0 U15874 ( .A1(n13058), .A2(poh11[14]), .ZN(n13059) );
  OAI21HSV2 U15875 ( .A1(poh11[14]), .A2(n13058), .B(n13059), .ZN(po[15]) );
  NAND2HSV0 U15876 ( .A1(n26759), .A2(n11891), .ZN(n13064) );
  NAND2HSV0 U15877 ( .A1(n26729), .A2(\pe3/got [13]), .ZN(n13066) );
  CLKNAND2HSV0 U15878 ( .A1(n13066), .A2(n13065), .ZN(n13067) );
  OAI21HSV0 U15879 ( .A1(n13065), .A2(n13066), .B(n13067), .ZN(n13068) );
  NAND2HSV0 U15880 ( .A1(n26348), .A2(n26600), .ZN(n13069) );
  OAI21HSV0 U15881 ( .A1(n13068), .A2(n13069), .B(n13070), .ZN(\pe3/poht [2])
         );
  CLKNAND2HSV2 U15882 ( .A1(\pe4/pvq [6]), .A2(n23508), .ZN(n13071) );
  NAND2HSV2 U15883 ( .A1(n13071), .A2(\pe4/phq [6]), .ZN(n13072) );
  OAI21HSV2 U15884 ( .A1(\pe4/phq [6]), .A2(n13071), .B(n13072), .ZN(n13073)
         );
  NAND2HSV0 U15885 ( .A1(n15784), .A2(\pe4/bq[12] ), .ZN(n13074) );
  OAI21HSV2 U15886 ( .A1(n13073), .A2(n13074), .B(n13075), .ZN(n15504) );
  NAND2HSV0 U15887 ( .A1(n28463), .A2(n15424), .ZN(n13078) );
  NAND2HSV0 U15888 ( .A1(n24771), .A2(\pe11/bq[11] ), .ZN(n13079) );
  AOI21HSV0 U15889 ( .A1(\pe11/pvq [8]), .A2(n20650), .B(n13079), .ZN(n13080)
         );
  AO31HSV0 U15890 ( .A1(\pe11/pvq [8]), .A2(n20650), .A3(n13079), .B(n13080), 
        .Z(n13081) );
  NAND2HSV0 U15891 ( .A1(\pe11/aot [10]), .A2(n24997), .ZN(n13082) );
  NAND2HSV2 U15892 ( .A1(n13082), .A2(n13081), .ZN(n13083) );
  OAI21HSV2 U15893 ( .A1(n13081), .A2(n13082), .B(n13083), .ZN(n13084) );
  NAND2HSV0 U15894 ( .A1(\pe11/bq[13] ), .A2(\pe11/aot [12]), .ZN(n13085) );
  NAND2HSV0 U15895 ( .A1(n13085), .A2(n13084), .ZN(n13086) );
  OAI21HSV0 U15896 ( .A1(n13084), .A2(n13085), .B(n13086), .ZN(n20389) );
  CLKNHSV0 U15897 ( .I(n19125), .ZN(n13087) );
  CLKNHSV0 U15898 ( .I(n19124), .ZN(n13088) );
  MUX2NHSV1 U15899 ( .I0(n13088), .I1(n19124), .S(n25764), .ZN(n13089) );
  NAND2HSV0 U15900 ( .A1(\pe10/bq[16] ), .A2(\pe10/aot [1]), .ZN(n13090) );
  OAI21HSV0 U15901 ( .A1(n26185), .A2(n26186), .B(n13090), .ZN(n13091) );
  OAI31HSV0 U15902 ( .A1(n26185), .A2(n13090), .A3(n26186), .B(n13091), .ZN(
        n13092) );
  NAND2HSV0 U15903 ( .A1(\pe10/aot [2]), .A2(\pe10/bq[15] ), .ZN(n13093) );
  NAND2HSV0 U15904 ( .A1(n13093), .A2(n13092), .ZN(n13094) );
  OAI21HSV0 U15905 ( .A1(n13092), .A2(n13093), .B(n13094), .ZN(n13095) );
  NAND2HSV0 U15906 ( .A1(\pe10/aot [5]), .A2(\pe10/bq[12] ), .ZN(n13096) );
  CLKNAND2HSV0 U15907 ( .A1(n13096), .A2(n13095), .ZN(n13097) );
  OAI21HSV0 U15908 ( .A1(n13095), .A2(n13096), .B(n13097), .ZN(n26187) );
  AOI22HSV0 U15909 ( .A1(\pe9/bq[2] ), .A2(\pe9/aot [14]), .B1(\pe9/bq[5] ), 
        .B2(\pe9/aot [11]), .ZN(n13098) );
  IAO21HSV2 U15910 ( .A1(n28089), .A2(n28088), .B(n13098), .ZN(n28093) );
  AOI22HSV0 U15911 ( .A1(\pe2/bq[9] ), .A2(\pe2/aot [8]), .B1(\pe2/aot [2]), 
        .B2(n27239), .ZN(n13099) );
  IAO21HSV2 U15912 ( .A1(n27299), .A2(n27576), .B(n13099), .ZN(n27300) );
  NAND2HSV0 U15913 ( .A1(\pe6/ti_7[1] ), .A2(\pe6/got [8]), .ZN(n13100) );
  NAND2HSV2 U15914 ( .A1(n13100), .A2(n14429), .ZN(n13101) );
  NAND2HSV0 U15915 ( .A1(n18930), .A2(\pe6/got [9]), .ZN(n13103) );
  NAND2HSV2 U15916 ( .A1(n13103), .A2(n13102), .ZN(n13104) );
  OAI21HSV2 U15917 ( .A1(n13102), .A2(n13103), .B(n13104), .ZN(n13105) );
  NAND2HSV0 U15918 ( .A1(n19076), .A2(\pe6/got [10]), .ZN(n13106) );
  NAND2HSV2 U15919 ( .A1(n13106), .A2(n13105), .ZN(n13107) );
  OAI21HSV2 U15920 ( .A1(n13105), .A2(n13106), .B(n13107), .ZN(n13108) );
  NAND2HSV0 U15921 ( .A1(n19109), .A2(\pe6/got [11]), .ZN(n13109) );
  NAND2HSV2 U15922 ( .A1(n13109), .A2(n13108), .ZN(n13110) );
  OAI21HSV2 U15923 ( .A1(n13108), .A2(n13109), .B(n13110), .ZN(n14430) );
  XOR2HSV0 U15924 ( .A1(n14957), .A2(n14958), .Z(n13111) );
  XOR2HSV0 U15925 ( .A1(n14947), .A2(n14946), .Z(n13112) );
  XOR2HSV0 U15926 ( .A1(n13111), .A2(n13112), .Z(n13113) );
  XOR2HSV0 U15927 ( .A1(n14933), .A2(n14932), .Z(n13114) );
  XOR2HSV0 U15928 ( .A1(n13113), .A2(n13114), .Z(n13115) );
  NAND2HSV0 U15929 ( .A1(n24340), .A2(n28614), .ZN(n13116) );
  NAND2HSV2 U15930 ( .A1(n13116), .A2(n13115), .ZN(n13117) );
  OAI21HSV2 U15931 ( .A1(n13115), .A2(n13116), .B(n13117), .ZN(n14960) );
  INAND2HSV0 U15932 ( .A1(\pe10/ti_7t [8]), .B1(n16843), .ZN(n17002) );
  INAND2HSV0 U15933 ( .A1(\pe2/ti_7t [6]), .B1(n21235), .ZN(n17864) );
  CLKNAND2HSV2 U15934 ( .A1(n14691), .A2(n14690), .ZN(n13120) );
  OAI21HSV4 U15935 ( .A1(n13119), .A2(n13120), .B(n13121), .ZN(n14910) );
  CLKNHSV0 U15936 ( .I(\pe6/ti_7t [14]), .ZN(n13122) );
  AOI21HSV0 U15937 ( .A1(n19068), .A2(n13122), .B(n24962), .ZN(n19135) );
  AO22HSV4 U15938 ( .A1(\pe8/ti_7t [7]), .A2(n18788), .B1(n29007), .B2(n18787), 
        .Z(n22141) );
  NAND2HSV0 U15939 ( .A1(n28345), .A2(n28344), .ZN(n13126) );
  INOR2HSV0 U15940 ( .A1(\pe2/ti_7t [13]), .B1(n21714), .ZN(n21630) );
  OAI21HSV4 U15941 ( .A1(n13127), .A2(n13128), .B(n13129), .ZN(n13130) );
  OAI21HSV4 U15942 ( .A1(n20141), .A2(n23716), .B(n20140), .ZN(n13131) );
  OAI21HSV4 U15943 ( .A1(n13130), .A2(n13131), .B(n13132), .ZN(n25685) );
  XOR2HSV0 U15944 ( .A1(n24210), .A2(n24209), .Z(n13133) );
  NAND2HSV0 U15945 ( .A1(n14067), .A2(\pe7/got [3]), .ZN(n13134) );
  CLKNAND2HSV0 U15946 ( .A1(n13134), .A2(n13133), .ZN(n13135) );
  OAI21HSV0 U15947 ( .A1(n13133), .A2(n13134), .B(n13135), .ZN(n13136) );
  NAND2HSV0 U15948 ( .A1(\pe7/got [4]), .A2(n11978), .ZN(n13137) );
  CLKNAND2HSV0 U15949 ( .A1(n13137), .A2(n13136), .ZN(n13138) );
  OAI21HSV0 U15950 ( .A1(n13136), .A2(n13137), .B(n13138), .ZN(n13139) );
  NAND2HSV0 U15951 ( .A1(n25397), .A2(n25375), .ZN(n13140) );
  CLKNAND2HSV0 U15952 ( .A1(n13140), .A2(n13139), .ZN(n13141) );
  OAI21HSV0 U15953 ( .A1(n13139), .A2(n13140), .B(n13141), .ZN(n13142) );
  NAND2HSV0 U15954 ( .A1(\pe7/got [6]), .A2(n25377), .ZN(n13143) );
  CLKNAND2HSV0 U15955 ( .A1(n13143), .A2(n13142), .ZN(n13144) );
  OAI21HSV0 U15956 ( .A1(n13142), .A2(n13143), .B(n13144), .ZN(n13145) );
  NAND2HSV0 U15957 ( .A1(n25271), .A2(n24287), .ZN(n13146) );
  NAND2HSV0 U15958 ( .A1(n13146), .A2(n13145), .ZN(n13147) );
  OAI21HSV2 U15959 ( .A1(n13145), .A2(n13146), .B(n13147), .ZN(n24212) );
  NAND2HSV0 U15960 ( .A1(n23450), .A2(n20775), .ZN(n13148) );
  NAND2HSV0 U15961 ( .A1(n13148), .A2(n23451), .ZN(n13149) );
  OAI21HSV0 U15962 ( .A1(n23451), .A2(n13148), .B(n13149), .ZN(n13150) );
  NAND2HSV0 U15963 ( .A1(n13150), .A2(n23452), .ZN(n13151) );
  OAI211HSV0 U15964 ( .A1(n23452), .A2(n13150), .B(n13151), .C(n20770), .ZN(
        n13152) );
  NAND2HSV0 U15965 ( .A1(n13152), .A2(poh11[12]), .ZN(n13153) );
  OAI21HSV2 U15966 ( .A1(poh11[12]), .A2(n13152), .B(n13153), .ZN(po[13]) );
  CLKNAND2HSV0 U15967 ( .A1(n13154), .A2(n13155), .ZN(n13156) );
  NAND2HSV0 U15968 ( .A1(n26759), .A2(\pe3/got [13]), .ZN(n13158) );
  OAI21HSV0 U15969 ( .A1(n13157), .A2(n13158), .B(n13159), .ZN(n13160) );
  NAND2HSV0 U15970 ( .A1(n26729), .A2(n26348), .ZN(n13161) );
  CLKNAND2HSV0 U15971 ( .A1(n13161), .A2(n13160), .ZN(n13162) );
  OAI21HSV0 U15972 ( .A1(n13160), .A2(n13161), .B(n13162), .ZN(n13163) );
  NAND2HSV0 U15973 ( .A1(n26240), .A2(n26600), .ZN(n13164) );
  OAI21HSV0 U15974 ( .A1(n13163), .A2(n13164), .B(n13165), .ZN(\pe3/poht [1])
         );
  AOI21HSV0 U15975 ( .A1(\pe6/pvq [13]), .A2(n23486), .B(\pe6/phq [13]), .ZN(
        n13166) );
  AO31HSV2 U15976 ( .A1(\pe6/pvq [13]), .A2(n23486), .A3(\pe6/phq [13]), .B(
        n13166), .Z(n13167) );
  NAND2HSV0 U15977 ( .A1(n19021), .A2(\pe6/got [4]), .ZN(n13168) );
  NAND2HSV2 U15978 ( .A1(n13168), .A2(n13167), .ZN(n13169) );
  OAI21HSV2 U15979 ( .A1(n13167), .A2(n13168), .B(n13169), .ZN(n13170) );
  NAND2HSV0 U15980 ( .A1(\pe6/bq[5] ), .A2(n28680), .ZN(n13171) );
  NAND2HSV2 U15981 ( .A1(n13171), .A2(n13170), .ZN(n13172) );
  OAI21HSV2 U15982 ( .A1(n13170), .A2(n13171), .B(n13172), .ZN(n19022) );
  CLKNHSV0 U15983 ( .I(\pe7/bq[13] ), .ZN(n13173) );
  OAI21HSV0 U15984 ( .A1(n19492), .A2(n13173), .B(n19491), .ZN(n19493) );
  AOI22HSV0 U15985 ( .A1(\pe6/bq[3] ), .A2(\pe6/aot [14]), .B1(\pe6/bq[4] ), 
        .B2(\pe6/aot [13]), .ZN(n13174) );
  IAO21HSV2 U15986 ( .A1(n25427), .A2(n25426), .B(n13174), .ZN(n25428) );
  NAND2HSV0 U15987 ( .A1(\pe3/bq[11] ), .A2(\pe3/aot [12]), .ZN(n13175) );
  OAI21HSV0 U15988 ( .A1(n15260), .A2(n26246), .B(n13175), .ZN(n13176) );
  OAI31HSV2 U15989 ( .A1(n15260), .A2(n13175), .A3(n26246), .B(n13176), .ZN(
        n15264) );
  INAND2HSV2 U15990 ( .A1(n16749), .B1(\pe10/ti_7t [2]), .ZN(n16666) );
  CLKNHSV0 U15991 ( .I(\pe7/phq [6]), .ZN(n13177) );
  NAND2HSV2 U15992 ( .A1(\pe7/pvq [6]), .A2(n27104), .ZN(n13178) );
  MUX2NHSV2 U15993 ( .I0(\pe7/phq [6]), .I1(n13177), .S(n13178), .ZN(n19288)
         );
  NAND2HSV0 U15994 ( .A1(\pe2/bq[10] ), .A2(\pe2/aot [16]), .ZN(n13179) );
  CLKNAND2HSV0 U15995 ( .A1(n13179), .A2(\pe2/phq [7]), .ZN(n13180) );
  OAI21HSV0 U15996 ( .A1(\pe2/phq [7]), .A2(n13179), .B(n13180), .ZN(n13181)
         );
  MUX2NHSV1 U15997 ( .I0(n27255), .I1(n17751), .S(n17750), .ZN(n13182) );
  CLKXOR2HSV4 U15998 ( .A1(n13181), .A2(n13182), .Z(n17760) );
  AO22HSV2 U15999 ( .A1(\pe11/bq[9] ), .A2(\pe11/aot [12]), .B1(\pe11/aot [9]), 
        .B2(\pe11/bq[12] ), .Z(n13183) );
  OAI21HSV2 U16000 ( .A1(n20711), .A2(n20786), .B(n13183), .ZN(n13184) );
  CLKNAND2HSV0 U16001 ( .A1(n13184), .A2(n24765), .ZN(n13185) );
  OAI21HSV0 U16002 ( .A1(n13184), .A2(n24765), .B(n13185), .ZN(n20591) );
  NAND2HSV0 U16003 ( .A1(n25029), .A2(n25030), .ZN(n13186) );
  NOR2HSV0 U16004 ( .A1(n25042), .A2(n13186), .ZN(n25039) );
  CLKNHSV0 U16005 ( .I(n19987), .ZN(n13187) );
  OAI21HSV0 U16006 ( .A1(n20058), .A2(n19988), .B(n13187), .ZN(n13989) );
  AOI22HSV0 U16007 ( .A1(\pe9/bq[5] ), .A2(\pe9/aot [8]), .B1(\pe9/aot [2]), 
        .B2(\pe9/bq[11] ), .ZN(n13188) );
  IAO21HSV2 U16008 ( .A1(n22333), .A2(n28363), .B(n13188), .ZN(n22334) );
  CLKNHSV0 U16009 ( .I(n27553), .ZN(n13189) );
  AOI22HSV0 U16010 ( .A1(\pe2/aot [8]), .A2(\pe2/bq[1] ), .B1(\pe2/bq[8] ), 
        .B2(\pe2/aot [1]), .ZN(n13190) );
  AOI21HSV2 U16011 ( .A1(n27672), .A2(n13189), .B(n13190), .ZN(n27557) );
  XOR2HSV0 U16012 ( .A1(n16983), .A2(n16982), .Z(n13192) );
  OAI21HSV0 U16013 ( .A1(n17068), .A2(n26091), .B(n13193), .ZN(n13194) );
  NOR2HSV0 U16014 ( .A1(n18075), .A2(n18552), .ZN(n13198) );
  NAND3HSV2 U16015 ( .A1(n13198), .A2(n18077), .A3(n18076), .ZN(n18080) );
  NOR2HSV0 U16016 ( .A1(n15483), .A2(n15482), .ZN(n13199) );
  CLKNAND2HSV4 U16017 ( .A1(n16398), .A2(n16399), .ZN(n13200) );
  OAI21HSV4 U16018 ( .A1(n16420), .A2(n13200), .B(n13201), .ZN(n16459) );
  CLKNHSV0 U16019 ( .I(n21308), .ZN(n13202) );
  CLKNHSV0 U16020 ( .I(\pe2/got [13]), .ZN(n13203) );
  OAI21HSV0 U16021 ( .A1(n27438), .A2(n13203), .B(n21306), .ZN(n13204) );
  MUX2NHSV1 U16022 ( .I0(n21308), .I1(n13202), .S(n13205), .ZN(n25361) );
  OAI21HSV0 U16023 ( .A1(n25256), .A2(n27195), .B(n25260), .ZN(n13206) );
  IOA21HSV2 U16024 ( .A1(n22624), .A2(n25264), .B(n13206), .ZN(n25690) );
  XOR2HSV0 U16025 ( .A1(n24070), .A2(n24069), .Z(n13207) );
  NAND2HSV0 U16026 ( .A1(\pe7/got [3]), .A2(n11978), .ZN(n13208) );
  CLKNAND2HSV0 U16027 ( .A1(n13208), .A2(n13207), .ZN(n13209) );
  OAI21HSV0 U16028 ( .A1(n13207), .A2(n13208), .B(n13209), .ZN(n13210) );
  NAND2HSV0 U16029 ( .A1(n25397), .A2(n25272), .ZN(n13211) );
  CLKNAND2HSV0 U16030 ( .A1(n13211), .A2(n13210), .ZN(n13212) );
  OAI21HSV0 U16031 ( .A1(n13210), .A2(n13211), .B(n13212), .ZN(n13213) );
  NAND2HSV0 U16032 ( .A1(\pe7/got [5]), .A2(n28656), .ZN(n13214) );
  CLKNAND2HSV0 U16033 ( .A1(n13214), .A2(n13213), .ZN(n13215) );
  OAI21HSV0 U16034 ( .A1(n13213), .A2(n13214), .B(n13215), .ZN(n13216) );
  NAND2HSV0 U16035 ( .A1(n28665), .A2(\pe7/got [6]), .ZN(n13217) );
  NAND2HSV0 U16036 ( .A1(n13217), .A2(n13216), .ZN(n13218) );
  OAI21HSV2 U16037 ( .A1(n13216), .A2(n13217), .B(n13218), .ZN(n24072) );
  NAND2HSV0 U16038 ( .A1(n20770), .A2(n23454), .ZN(n13219) );
  NAND2HSV0 U16039 ( .A1(n13219), .A2(poh11[11]), .ZN(n13220) );
  OAI21HSV2 U16040 ( .A1(poh11[11]), .A2(n13219), .B(n13220), .ZN(po[12]) );
  NAND2HSV0 U16041 ( .A1(n13222), .A2(n13221), .ZN(n13223) );
  OAI21HSV0 U16042 ( .A1(n13222), .A2(n13221), .B(n13223), .ZN(\pe5/poht [6])
         );
  NAND2HSV0 U16043 ( .A1(n28652), .A2(\pe3/got [7]), .ZN(n13225) );
  OAI21HSV0 U16044 ( .A1(n13224), .A2(n13225), .B(n13226), .ZN(n13227) );
  NAND2HSV0 U16045 ( .A1(n28648), .A2(n26760), .ZN(n13228) );
  CLKNAND2HSV0 U16046 ( .A1(n13228), .A2(n13227), .ZN(n13229) );
  OAI21HSV0 U16047 ( .A1(n13227), .A2(n13228), .B(n13229), .ZN(n13230) );
  NAND2HSV0 U16048 ( .A1(n26679), .A2(\pe3/got [9]), .ZN(n13231) );
  NAND2HSV0 U16049 ( .A1(n13231), .A2(n13230), .ZN(n13232) );
  OAI21HSV0 U16050 ( .A1(n13230), .A2(n13231), .B(n13232), .ZN(\pe3/poht [7])
         );
  CLKNHSV0 U16051 ( .I(\pe5/phq [8]), .ZN(n13233) );
  CLKNAND2HSV0 U16052 ( .A1(\pe5/pvq [8]), .A2(n14646), .ZN(n13234) );
  MUX2NHSV1 U16053 ( .I0(\pe5/phq [8]), .I1(n13233), .S(n13234), .ZN(n14647)
         );
  NAND2HSV0 U16054 ( .A1(\pe11/aot [6]), .A2(\pe11/bq[14] ), .ZN(n13235) );
  OAI21HSV0 U16055 ( .A1(n20267), .A2(n20811), .B(n13235), .ZN(n13236) );
  OAI31HSV2 U16056 ( .A1(n20267), .A2(n13235), .A3(n20811), .B(n13236), .ZN(
        n20658) );
  CLKNHSV0 U16057 ( .I(n19021), .ZN(n13237) );
  NAND2HSV0 U16058 ( .A1(\pe6/aot [14]), .A2(\pe6/bq[7] ), .ZN(n13238) );
  NAND2HSV0 U16059 ( .A1(\pe6/aot [7]), .A2(\pe6/bq[14] ), .ZN(n13239) );
  NAND2HSV0 U16060 ( .A1(n13239), .A2(n13238), .ZN(n13240) );
  OAI21HSV2 U16061 ( .A1(n13238), .A2(n13239), .B(n13240), .ZN(n13241) );
  NAND2HSV0 U16062 ( .A1(\pe6/aot [6]), .A2(\pe6/bq[15] ), .ZN(n13242) );
  NAND2HSV2 U16063 ( .A1(n13242), .A2(n13241), .ZN(n13243) );
  OAI21HSV2 U16064 ( .A1(n13241), .A2(n13242), .B(n13243), .ZN(n13244) );
  OAI21HSV0 U16065 ( .A1(n26014), .A2(n13237), .B(n13244), .ZN(n13245) );
  OAI31HSV2 U16066 ( .A1(n26014), .A2(n13244), .A3(n13237), .B(n13245), .ZN(
        n18869) );
  OAI21HSV0 U16067 ( .A1(n27846), .A2(n26940), .B(n22829), .ZN(n13246) );
  NAND2HSV0 U16068 ( .A1(\pe4/pvq [12]), .A2(n27129), .ZN(n13247) );
  CLKNAND2HSV0 U16069 ( .A1(n13247), .A2(\pe4/phq [12]), .ZN(n13248) );
  OAI21HSV0 U16070 ( .A1(\pe4/phq [12]), .A2(n13247), .B(n13248), .ZN(n13249)
         );
  OAI21HSV0 U16071 ( .A1(n22001), .A2(n26942), .B(n13246), .ZN(n13250) );
  NAND2HSV0 U16072 ( .A1(n13250), .A2(n13249), .ZN(n13251) );
  OAI21HSV2 U16073 ( .A1(n13250), .A2(n13249), .B(n13251), .ZN(n15877) );
  NAND2HSV0 U16074 ( .A1(n23519), .A2(\pe8/pvq [15]), .ZN(n13252) );
  NAND2HSV0 U16075 ( .A1(n13252), .A2(\pe8/phq [15]), .ZN(n13253) );
  OAI21HSV0 U16076 ( .A1(\pe8/phq [15]), .A2(n13252), .B(n13253), .ZN(n19998)
         );
  AOI22HSV0 U16077 ( .A1(\pe3/bq[11] ), .A2(\pe3/aot [16]), .B1(\pe3/aot [13]), 
        .B2(\pe3/bq[14] ), .ZN(n13254) );
  IAO21HSV2 U16078 ( .A1(n15161), .A2(n15304), .B(n13254), .ZN(n15166) );
  NAND2HSV0 U16079 ( .A1(n23541), .A2(\pe3/pvq [11]), .ZN(n13255) );
  NAND2HSV2 U16080 ( .A1(n13255), .A2(\pe3/phq [11]), .ZN(n13256) );
  OAI21HSV2 U16081 ( .A1(\pe3/phq [11]), .A2(n13255), .B(n13256), .ZN(n15998)
         );
  INOR2HSV0 U16082 ( .A1(\pe2/aot [10]), .B1(n27322), .ZN(n13257) );
  CLKNAND2HSV0 U16083 ( .A1(n22114), .A2(\pe2/pvq [7]), .ZN(n13258) );
  CLKNAND2HSV0 U16084 ( .A1(n13258), .A2(n13257), .ZN(n13259) );
  OAI21HSV0 U16085 ( .A1(n13257), .A2(n13258), .B(n13259), .ZN(n17761) );
  CLKNHSV0 U16086 ( .I(n26166), .ZN(n13260) );
  AOI22HSV0 U16087 ( .A1(\pe10/bq[6] ), .A2(\pe10/aot [11]), .B1(n16973), .B2(
        \pe10/bq[2] ), .ZN(n13261) );
  AOI21HSV0 U16088 ( .A1(n26167), .A2(n13260), .B(n13261), .ZN(n26168) );
  NAND2HSV0 U16089 ( .A1(\pe9/aot [6]), .A2(\pe9/bq[9] ), .ZN(n13262) );
  NAND2HSV0 U16090 ( .A1(\pe9/bq[8] ), .A2(\pe9/aot [7]), .ZN(n13263) );
  NAND2HSV0 U16091 ( .A1(n13263), .A2(n13262), .ZN(n13264) );
  OAI21HSV2 U16092 ( .A1(n13262), .A2(n13263), .B(n13264), .ZN(n13265) );
  NAND2HSV0 U16093 ( .A1(\pe9/bq[10] ), .A2(\pe9/aot [5]), .ZN(n13266) );
  NAND2HSV2 U16094 ( .A1(n13266), .A2(n13265), .ZN(n13267) );
  OAI21HSV2 U16095 ( .A1(n13265), .A2(n13266), .B(n13267), .ZN(n13268) );
  NAND2HSV0 U16096 ( .A1(\pe9/aot [8]), .A2(\pe9/bq[7] ), .ZN(n13269) );
  CLKNAND2HSV0 U16097 ( .A1(n13269), .A2(n13268), .ZN(n13270) );
  OAI21HSV2 U16098 ( .A1(n13268), .A2(n13269), .B(n13270), .ZN(n22395) );
  CLKNHSV0 U16099 ( .I(n17941), .ZN(n13271) );
  MUX2NHSV2 U16100 ( .I0(n17941), .I1(n13271), .S(n17942), .ZN(n17951) );
  CLKNHSV0 U16101 ( .I(\pe11/phq [4]), .ZN(n13272) );
  NAND2HSV0 U16102 ( .A1(\pe11/ti_1 ), .A2(n20707), .ZN(n13273) );
  MUX2NHSV1 U16103 ( .I0(\pe11/phq [4]), .I1(n13272), .S(n13273), .ZN(n20203)
         );
  AOI21HSV0 U16104 ( .A1(n18856), .A2(n19147), .B(n18855), .ZN(n13274) );
  OAI21HSV0 U16105 ( .A1(n18857), .A2(n28676), .B(n13274), .ZN(n18900) );
  INAND2HSV0 U16106 ( .A1(\pe5/ti_7t [8]), .B1(ctro5), .ZN(n14965) );
  INOR2HSV4 U16107 ( .A1(n25357), .B1(n21301), .ZN(n21881) );
  CLKNHSV0 U16108 ( .I(n25756), .ZN(n13275) );
  AOI22HSV0 U16109 ( .A1(\pe6/bq[5] ), .A2(\pe6/aot [9]), .B1(\pe6/aot [13]), 
        .B2(\pe6/bq[1] ), .ZN(n13276) );
  AOI21HSV2 U16110 ( .A1(n25716), .A2(n13275), .B(n13276), .ZN(n25720) );
  XOR2HSV0 U16111 ( .A1(n19603), .A2(n19604), .Z(n13277) );
  XOR2HSV0 U16112 ( .A1(n19590), .A2(n19589), .Z(n13278) );
  XOR2HSV0 U16113 ( .A1(n13277), .A2(n13278), .Z(n13279) );
  NAND2HSV0 U16114 ( .A1(n25271), .A2(n11858), .ZN(n13280) );
  NAND2HSV2 U16115 ( .A1(n13280), .A2(n13279), .ZN(n13281) );
  OAI21HSV2 U16116 ( .A1(n13279), .A2(n13280), .B(n13281), .ZN(n13282) );
  NAND2HSV0 U16117 ( .A1(n25292), .A2(\pe7/got [8]), .ZN(n13283) );
  NAND2HSV0 U16118 ( .A1(n13283), .A2(n13282), .ZN(n13284) );
  OAI21HSV0 U16119 ( .A1(n13282), .A2(n13283), .B(n13284), .ZN(n13285) );
  NAND2HSV0 U16120 ( .A1(\pe7/got [9]), .A2(n12288), .ZN(n13286) );
  NAND2HSV0 U16121 ( .A1(\pe7/got [10]), .A2(n19739), .ZN(n13288) );
  NAND2HSV2 U16122 ( .A1(n13288), .A2(n13287), .ZN(n13289) );
  OAI21HSV2 U16123 ( .A1(n13287), .A2(n13288), .B(n13289), .ZN(n19606) );
  MUX2NHSV4 U16124 ( .I0(n16883), .I1(n13290), .S(n16882), .ZN(n16885) );
  INOR2HSV2 U16125 ( .A1(n14573), .B1(n14549), .ZN(n14575) );
  AOI21HSV0 U16126 ( .A1(n16164), .A2(n16016), .B(n23383), .ZN(n13291) );
  OAI21HSV4 U16127 ( .A1(n16018), .A2(n16056), .B(n13291), .ZN(n15277) );
  INHSV4 U16128 ( .I(n17600), .ZN(n13292) );
  NOR2HSV2 U16129 ( .A1(n15413), .A2(n15752), .ZN(n13293) );
  MUX2NHSV2 U16130 ( .I0(n13294), .I1(n19460), .S(n19461), .ZN(n19517) );
  CLKNHSV0 U16131 ( .I(\pe2/aot [6]), .ZN(n13295) );
  IOA22HSV1 U16132 ( .B1(n27652), .B2(n13295), .A1(\pe2/aot [3]), .A2(
        \pe2/bq[4] ), .ZN(n13296) );
  OAI21HSV0 U16133 ( .A1(n27653), .A2(n27734), .B(n13296), .ZN(n13297) );
  CLKNHSV0 U16134 ( .I(\pe2/aot [4]), .ZN(n13298) );
  OAI21HSV0 U16135 ( .A1(n27710), .A2(n13298), .B(n27651), .ZN(n13299) );
  OAI21HSV0 U16136 ( .A1(n27708), .A2(n27711), .B(n13299), .ZN(n13300) );
  NAND2HSV0 U16137 ( .A1(n13300), .A2(n13297), .ZN(n13301) );
  OAI21HSV2 U16138 ( .A1(n13300), .A2(n13297), .B(n13301), .ZN(n13302) );
  NAND2HSV0 U16139 ( .A1(\pe2/aot [2]), .A2(\pe2/bq[5] ), .ZN(n13303) );
  NAND2HSV2 U16140 ( .A1(n13303), .A2(n13302), .ZN(n13304) );
  OAI21HSV2 U16141 ( .A1(n13302), .A2(n13303), .B(n13304), .ZN(n13305) );
  OAI21HSV0 U16142 ( .A1(n27654), .A2(n27693), .B(n13305), .ZN(n13306) );
  OAI31HSV0 U16143 ( .A1(n27654), .A2(n13305), .A3(n27693), .B(n13306), .ZN(
        n27655) );
  CLKNHSV0 U16144 ( .I(\pe7/ti_7t [13]), .ZN(n13307) );
  AOI21HSV0 U16145 ( .A1(n23188), .A2(n13307), .B(n27134), .ZN(n25496) );
  CLKNHSV0 U16146 ( .I(n21643), .ZN(n13309) );
  OAI22HSV2 U16147 ( .A1(n21644), .A2(n13308), .B1(\pe2/ti_7t [9]), .B2(n13309), .ZN(n27277) );
  AND2HSV2 U16148 ( .A1(n25255), .A2(n28603), .Z(n25257) );
  CLKNHSV0 U16149 ( .I(n25352), .ZN(n13310) );
  OAI21HSV0 U16150 ( .A1(n25515), .A2(n13310), .B(poh11[10]), .ZN(n13311) );
  OAI31HSV2 U16151 ( .A1(n25515), .A2(poh11[10]), .A3(n13310), .B(n13311), 
        .ZN(po[11]) );
  OAI21HSV0 U16152 ( .A1(n13312), .A2(n13313), .B(n13314), .ZN(\pe5/poht [7])
         );
  XOR2HSV0 U16153 ( .A1(n22417), .A2(n22416), .Z(n13315) );
  NAND2HSV0 U16154 ( .A1(n28394), .A2(\pe9/got [12]), .ZN(n13316) );
  CLKNAND2HSV0 U16155 ( .A1(n13316), .A2(n13315), .ZN(n13317) );
  OAI21HSV0 U16156 ( .A1(n13315), .A2(n13316), .B(n13317), .ZN(n13318) );
  NAND3HSV2 U16157 ( .A1(n28340), .A2(\pe9/got [13]), .A3(n28404), .ZN(n13319)
         );
  NAND2HSV0 U16158 ( .A1(n13319), .A2(n13318), .ZN(n13320) );
  NAND2HSV0 U16159 ( .A1(n28928), .A2(n28414), .ZN(n13322) );
  OAI21HSV0 U16160 ( .A1(n13321), .A2(n13322), .B(n13323), .ZN(\pe9/poht [2])
         );
  CLKNHSV0 U16161 ( .I(n22244), .ZN(n13325) );
  NAND2HSV0 U16162 ( .A1(n26231), .A2(n25577), .ZN(n13326) );
  MUX2NHSV0 U16163 ( .I0(n13325), .I1(n22244), .S(n13326), .ZN(n13327) );
  MUX2NHSV1 U16164 ( .I0(n22245), .I1(n13324), .S(n13327), .ZN(\pe8/poht [11])
         );
  XOR2HSV0 U16165 ( .A1(n26728), .A2(n26727), .Z(n13328) );
  NAND2HSV0 U16166 ( .A1(n26759), .A2(\pe3/got [10]), .ZN(n13329) );
  CLKNAND2HSV0 U16167 ( .A1(n13329), .A2(n13328), .ZN(n13330) );
  NAND2HSV0 U16168 ( .A1(\pe3/got [11]), .A2(n26729), .ZN(n13332) );
  OAI21HSV0 U16169 ( .A1(n13331), .A2(n13332), .B(n13333), .ZN(n13334) );
  NAND2HSV0 U16170 ( .A1(n13335), .A2(n13334), .ZN(n13336) );
  NAND2HSV4 U16171 ( .A1(n19121), .A2(n25647), .ZN(n13337) );
  CLKNHSV0 U16172 ( .I(\pe9/phq [12]), .ZN(n13339) );
  NAND2HSV0 U16173 ( .A1(\pe9/pvq [12]), .A2(n21760), .ZN(n13340) );
  MUX2NHSV0 U16174 ( .I0(\pe9/phq [12]), .I1(n13339), .S(n13340), .ZN(n18417)
         );
  CLKNHSV0 U16175 ( .I(\pe6/phq [6]), .ZN(n13341) );
  NAND2HSV4 U16176 ( .A1(\pe6/pvq [6]), .A2(n27073), .ZN(n13342) );
  MUX2NHSV2 U16177 ( .I0(\pe6/phq [6]), .I1(n13341), .S(n13342), .ZN(n14101)
         );
  CLKNHSV0 U16178 ( .I(\pe9/bq[6] ), .ZN(n13343) );
  IOA22HSV1 U16179 ( .B1(n22330), .B2(n13343), .A1(\pe9/aot [11]), .A2(
        \pe9/bq[1] ), .ZN(n28147) );
  NAND2HSV0 U16180 ( .A1(\pe8/bq[14] ), .A2(\pe8/aot [3]), .ZN(n13344) );
  OAI21HSV2 U16181 ( .A1(n25531), .A2(n25530), .B(n13344), .ZN(n13345) );
  OAI31HSV2 U16182 ( .A1(n25531), .A2(n13344), .A3(n25530), .B(n13345), .ZN(
        n25536) );
  XOR2HSV0 U16183 ( .A1(n16971), .A2(n16972), .Z(n13346) );
  XOR2HSV0 U16184 ( .A1(n16966), .A2(n16965), .Z(n13347) );
  XOR2HSV0 U16185 ( .A1(n13346), .A2(n13347), .Z(n13348) );
  NAND2HSV0 U16186 ( .A1(n28642), .A2(n16850), .ZN(n13349) );
  NAND2HSV0 U16187 ( .A1(n13349), .A2(n13348), .ZN(n13350) );
  OAI21HSV2 U16188 ( .A1(n13348), .A2(n13349), .B(n13350), .ZN(n13351) );
  NAND2HSV0 U16189 ( .A1(\pe10/got [7]), .A2(n28666), .ZN(n13352) );
  NAND2HSV2 U16190 ( .A1(n13351), .A2(n13352), .ZN(n13353) );
  OAI21HSV2 U16191 ( .A1(n13351), .A2(n13352), .B(n13353), .ZN(n13354) );
  XOR2HSV0 U16192 ( .A1(n16981), .A2(n16980), .Z(n13355) );
  CLKXOR2HSV4 U16193 ( .A1(n13354), .A2(n13355), .Z(n13356) );
  NAND2HSV0 U16194 ( .A1(\pe10/got [9]), .A2(n28679), .ZN(n13357) );
  OAI21HSV2 U16195 ( .A1(n13356), .A2(n13357), .B(n13358), .ZN(n16982) );
  INHSV2 U16196 ( .I(n15830), .ZN(n13359) );
  MUX2NHSV2 U16197 ( .I0(n13359), .I1(n15830), .S(n13360), .ZN(n15833) );
  AOI22HSV0 U16198 ( .A1(\pe7/bq[5] ), .A2(\pe7/aot [11]), .B1(\pe7/aot [5]), 
        .B2(\pe7/bq[11] ), .ZN(n13361) );
  IAO21HSV2 U16199 ( .A1(n24241), .A2(n25382), .B(n13361), .ZN(n24242) );
  NAND2HSV0 U16200 ( .A1(\pe6/bq[3] ), .A2(\pe6/aot [8]), .ZN(n13362) );
  AOI22HSV0 U16201 ( .A1(n25994), .A2(n25961), .B1(n25992), .B2(n13362), .ZN(
        n25791) );
  NAND2HSV0 U16202 ( .A1(\pe5/bq[7] ), .A2(\pe5/aot [7]), .ZN(n13363) );
  OAI21HSV0 U16203 ( .A1(n24440), .A2(n27049), .B(n13363), .ZN(n13364) );
  OAI31HSV0 U16204 ( .A1(n24440), .A2(n13363), .A3(n27049), .B(n13364), .ZN(
        n23914) );
  NAND2HSV0 U16205 ( .A1(\pe1/bq[4] ), .A2(\pe1/aot [12]), .ZN(n13365) );
  AOI22HSV0 U16206 ( .A1(n27022), .A2(n26556), .B1(n26557), .B2(n13365), .ZN(
        n26558) );
  CLKNHSV0 U16207 ( .I(\pe4/phq [2]), .ZN(n13366) );
  INAND2HSV2 U16208 ( .A1(n20372), .B1(n20562), .ZN(n20624) );
  NAND2HSV0 U16209 ( .A1(\pe3/aot [3]), .A2(\pe3/bq[8] ), .ZN(n13368) );
  CLKNAND2HSV0 U16210 ( .A1(n13368), .A2(n23689), .ZN(n13369) );
  OAI21HSV0 U16211 ( .A1(n23689), .A2(n13368), .B(n13369), .ZN(n13370) );
  NAND2HSV0 U16212 ( .A1(\pe3/aot [6]), .A2(\pe3/bq[5] ), .ZN(n13371) );
  CLKNAND2HSV0 U16213 ( .A1(n13371), .A2(n13370), .ZN(n13372) );
  OAI21HSV0 U16214 ( .A1(n13370), .A2(n13371), .B(n13372), .ZN(n13373) );
  CLKNHSV0 U16215 ( .I(n26610), .ZN(n13374) );
  XOR2HSV0 U16216 ( .A1(n23685), .A2(n23684), .Z(n13375) );
  OAI21HSV0 U16217 ( .A1(n23688), .A2(n23687), .B(n13375), .ZN(n13376) );
  OAI31HSV0 U16218 ( .A1(n23688), .A2(n13375), .A3(n23687), .B(n13376), .ZN(
        n13377) );
  NAND2HSV0 U16219 ( .A1(\pe3/bq[2] ), .A2(\pe3/aot [9]), .ZN(n13378) );
  CLKNAND2HSV0 U16220 ( .A1(n13378), .A2(n13377), .ZN(n13379) );
  OAI21HSV0 U16221 ( .A1(n13377), .A2(n13378), .B(n13379), .ZN(n13380) );
  MUX2NHSV0 U16222 ( .I0(n13374), .I1(n26610), .S(n13380), .ZN(n13381) );
  XOR2HSV0 U16223 ( .A1(n23690), .A2(n13373), .Z(n13382) );
  XOR2HSV0 U16224 ( .A1(n13381), .A2(n13382), .Z(n13383) );
  NAND2HSV0 U16225 ( .A1(\pe3/got [1]), .A2(n23683), .ZN(n13384) );
  CLKNAND2HSV0 U16226 ( .A1(n13384), .A2(n13383), .ZN(n13385) );
  OAI21HSV0 U16227 ( .A1(n13383), .A2(n13384), .B(n13385), .ZN(n13386) );
  NAND2HSV0 U16228 ( .A1(\pe3/got [2]), .A2(n23328), .ZN(n13387) );
  CLKNAND2HSV0 U16229 ( .A1(n13387), .A2(n13386), .ZN(n13388) );
  OAI21HSV2 U16230 ( .A1(n13386), .A2(n13387), .B(n13388), .ZN(n23691) );
  NOR2HSV0 U16231 ( .A1(n15704), .A2(n15900), .ZN(n13389) );
  IOA21HSV4 U16232 ( .A1(n17819), .A2(n28454), .B(n17715), .ZN(n21065) );
  NAND2HSV0 U16233 ( .A1(n26132), .A2(n22439), .ZN(n13390) );
  XOR2HSV0 U16234 ( .A1(n27038), .A2(n27037), .Z(n13391) );
  XOR2HSV0 U16235 ( .A1(n27039), .A2(n13391), .Z(n13392) );
  NAND2HSV0 U16236 ( .A1(\pe1/got [7]), .A2(n12274), .ZN(n13393) );
  CLKNAND2HSV0 U16237 ( .A1(n13393), .A2(n13392), .ZN(n13394) );
  OAI21HSV0 U16238 ( .A1(n13392), .A2(n13393), .B(n13394), .ZN(n13395) );
  OAI21HSV0 U16239 ( .A1(n27004), .A2(n27003), .B(n13395), .ZN(n13396) );
  OAI31HSV0 U16240 ( .A1(n27004), .A2(n13395), .A3(n27003), .B(n13396), .ZN(
        n13397) );
  OAI21HSV0 U16241 ( .A1(n27002), .A2(n27001), .B(n13397), .ZN(n13398) );
  OAI31HSV2 U16242 ( .A1(n27002), .A2(n13397), .A3(n27001), .B(n13398), .ZN(
        n27040) );
  INAND2HSV4 U16243 ( .A1(n16441), .B1(n16443), .ZN(n25652) );
  AOI31HSV2 U16244 ( .A1(n19676), .A2(n19705), .A3(n19675), .B(n19613), .ZN(
        n13399) );
  NAND2HSV0 U16245 ( .A1(n23457), .A2(n20770), .ZN(n13400) );
  NAND2HSV0 U16246 ( .A1(n13400), .A2(poh11[9]), .ZN(n13401) );
  OAI21HSV2 U16247 ( .A1(poh11[9]), .A2(n13400), .B(n13401), .ZN(po[10]) );
  NAND2HSV0 U16248 ( .A1(n26759), .A2(\pe3/got [6]), .ZN(n13403) );
  OAI21HSV0 U16249 ( .A1(n13402), .A2(n13403), .B(n13404), .ZN(n13405) );
  NAND2HSV0 U16250 ( .A1(\pe3/got [7]), .A2(n26760), .ZN(n13406) );
  CLKNAND2HSV0 U16251 ( .A1(n13406), .A2(n13405), .ZN(n13407) );
  OAI21HSV0 U16252 ( .A1(n13405), .A2(n13406), .B(n13407), .ZN(n13408) );
  NAND2HSV0 U16253 ( .A1(n28648), .A2(n28661), .ZN(n13409) );
  NAND2HSV0 U16254 ( .A1(n13409), .A2(n13408), .ZN(n13410) );
  OAI21HSV0 U16255 ( .A1(n13408), .A2(n13409), .B(n13410), .ZN(\pe3/poht [8])
         );
  INHSV4 U16256 ( .I(n17997), .ZN(n13411) );
  AOI21HSV2 U16257 ( .A1(n28110), .A2(n17996), .B(n17995), .ZN(n13412) );
  MUX2NHSV4 U16258 ( .I0(n17997), .I1(n13411), .S(n13412), .ZN(n28961) );
  AOI22HSV0 U16259 ( .A1(\pe11/aot [7]), .A2(\pe11/bq[12] ), .B1(\pe11/bq[7] ), 
        .B2(\pe11/aot [12]), .ZN(n13415) );
  IAO21HSV2 U16260 ( .A1(n20711), .A2(n24715), .B(n13415), .ZN(n13416) );
  CLKNAND2HSV0 U16261 ( .A1(n24980), .A2(\pe11/pvq [14]), .ZN(n13417) );
  NAND2HSV2 U16262 ( .A1(n13417), .A2(n13416), .ZN(n13418) );
  OAI21HSV2 U16263 ( .A1(n13416), .A2(n13417), .B(n13418), .ZN(n20720) );
  CLKNHSV0 U16264 ( .I(\pe5/bq[5] ), .ZN(n13419) );
  OAI21HSV0 U16265 ( .A1(n23789), .A2(n13419), .B(n14954), .ZN(n13420) );
  OAI21HSV0 U16266 ( .A1(n14955), .A2(n21470), .B(n13420), .ZN(n13421) );
  NOR2HSV0 U16267 ( .A1(n14956), .A2(n23923), .ZN(n13422) );
  NAND2HSV0 U16268 ( .A1(n13422), .A2(n13421), .ZN(n13423) );
  OAI21HSV0 U16269 ( .A1(n13422), .A2(n13421), .B(n13423), .ZN(n14957) );
  NAND2HSV0 U16270 ( .A1(n25273), .A2(\pe7/aot [8]), .ZN(n13424) );
  OAI21HSV0 U16271 ( .A1(n24105), .A2(n25278), .B(n13424), .ZN(n13425) );
  OAI31HSV0 U16272 ( .A1(n24105), .A2(n13424), .A3(n25278), .B(n13425), .ZN(
        n19483) );
  NAND2HSV0 U16273 ( .A1(\pe1/bq[2] ), .A2(\pe1/aot [11]), .ZN(n13426) );
  OAI21HSV0 U16274 ( .A1(n26764), .A2(n26763), .B(n13426), .ZN(n13427) );
  OAI31HSV0 U16275 ( .A1(n26764), .A2(n13426), .A3(n26763), .B(n13427), .ZN(
        n26765) );
  NOR2HSV0 U16276 ( .A1(n23723), .A2(n23760), .ZN(n13428) );
  OAI22HSV0 U16277 ( .A1(n23561), .A2(n13428), .B1(n26226), .B2(n22252), .ZN(
        n22256) );
  AOI22HSV0 U16278 ( .A1(\pe8/bq[7] ), .A2(\pe8/aot [6]), .B1(\pe8/aot [5]), 
        .B2(\pe8/bq[8] ), .ZN(n13429) );
  IAO21HSV2 U16279 ( .A1(n23563), .A2(n23562), .B(n13429), .ZN(n23564) );
  NAND2HSV0 U16280 ( .A1(\pe10/bq[9] ), .A2(\pe10/aot [3]), .ZN(n13430) );
  AOI22HSV0 U16281 ( .A1(n25223), .A2(n27199), .B1(n25224), .B2(n13430), .ZN(
        n13431) );
  NAND2HSV0 U16282 ( .A1(\pe10/bq[6] ), .A2(\pe10/aot [6]), .ZN(n13432) );
  NAND2HSV0 U16283 ( .A1(\pe10/bq[3] ), .A2(\pe10/aot [9]), .ZN(n13433) );
  CLKNAND2HSV0 U16284 ( .A1(n13433), .A2(n13432), .ZN(n13434) );
  OAI21HSV0 U16285 ( .A1(n13432), .A2(n13433), .B(n13434), .ZN(n13435) );
  XOR2HSV0 U16286 ( .A1(n13431), .A2(n13435), .Z(n25232) );
  IOA22HSV4 U16287 ( .B1(n14265), .B2(n13436), .A1(n14264), .A2(n14262), .ZN(
        n14272) );
  CLKNHSV0 U16288 ( .I(\pe8/phq [4]), .ZN(n13437) );
  AOI21HSV0 U16289 ( .A1(n27089), .A2(\pe4/pvq [11]), .B(\pe4/phq [11]), .ZN(
        n13439) );
  AO31HSV2 U16290 ( .A1(n27089), .A2(\pe4/pvq [11]), .A3(\pe4/phq [11]), .B(
        n13439), .Z(n13440) );
  NAND2HSV0 U16291 ( .A1(n15784), .A2(\pe4/bq[7] ), .ZN(n13441) );
  NAND2HSV2 U16292 ( .A1(n13441), .A2(n13440), .ZN(n13442) );
  OAI21HSV2 U16293 ( .A1(n13440), .A2(n13441), .B(n13442), .ZN(n13443) );
  NAND2HSV0 U16294 ( .A1(n23076), .A2(\pe4/aot [9]), .ZN(n13444) );
  NAND2HSV0 U16295 ( .A1(n13444), .A2(n13443), .ZN(n13445) );
  OAI21HSV0 U16296 ( .A1(n13443), .A2(n13444), .B(n13445), .ZN(n15739) );
  XOR2HSV0 U16297 ( .A1(n15274), .A2(n15273), .Z(n13446) );
  NAND2HSV0 U16298 ( .A1(n16112), .A2(\pe3/got [11]), .ZN(n13447) );
  CLKNAND2HSV0 U16299 ( .A1(n13447), .A2(n13446), .ZN(n13448) );
  OAI21HSV2 U16300 ( .A1(n13446), .A2(n13447), .B(n13448), .ZN(n13449) );
  NAND2HSV0 U16301 ( .A1(n28628), .A2(n23683), .ZN(n13450) );
  XOR2HSV0 U16302 ( .A1(n17663), .A2(n17662), .Z(n13452) );
  MUX2NHSV4 U16303 ( .I0(n17664), .I1(n13451), .S(n13452), .ZN(n17700) );
  XOR2HSV0 U16304 ( .A1(n19669), .A2(n19668), .Z(n13453) );
  NAND2HSV0 U16305 ( .A1(n24214), .A2(n28466), .ZN(n13454) );
  CLKNAND2HSV0 U16306 ( .A1(n13454), .A2(n13453), .ZN(n13455) );
  OAI21HSV0 U16307 ( .A1(n13453), .A2(n13454), .B(n13455), .ZN(n13456) );
  NAND2HSV0 U16308 ( .A1(n14022), .A2(n14066), .ZN(n13457) );
  CLKNAND2HSV0 U16309 ( .A1(n13457), .A2(n13456), .ZN(n13458) );
  OAI21HSV0 U16310 ( .A1(n13456), .A2(n13457), .B(n13458), .ZN(n13459) );
  OAI21HSV2 U16311 ( .A1(n13459), .A2(n13460), .B(n13461), .ZN(n19673) );
  INAND2HSV2 U16312 ( .A1(n22905), .B1(\pe4/ti_7t [14]), .ZN(n22792) );
  CLKNHSV0 U16313 ( .I(\pe7/ti_7t [9]), .ZN(n13462) );
  AOI21HSV0 U16314 ( .A1(n19695), .A2(n13462), .B(n27134), .ZN(n19523) );
  CLKNHSV0 U16315 ( .I(n26043), .ZN(n13463) );
  MUX2NHSV0 U16316 ( .I0(n13463), .I1(n26043), .S(n19167), .ZN(n13464) );
  XOR2HSV0 U16317 ( .A1(n19168), .A2(n13464), .Z(n13465) );
  NAND2HSV0 U16318 ( .A1(n25952), .A2(n26083), .ZN(n13466) );
  XOR2HSV0 U16319 ( .A1(n13465), .A2(n13466), .Z(n13467) );
  OAI21HSV0 U16320 ( .A1(n12123), .A2(n28651), .B(n13467), .ZN(n13468) );
  OAI31HSV0 U16321 ( .A1(n12123), .A2(n13467), .A3(n28651), .B(n13468), .ZN(
        n19169) );
  CLKNHSV0 U16322 ( .I(n25420), .ZN(n13469) );
  CLKNHSV0 U16323 ( .I(n27711), .ZN(n13470) );
  CLKNHSV0 U16324 ( .I(n27707), .ZN(n13471) );
  MUX2NHSV0 U16325 ( .I0(n13471), .I1(n27707), .S(n27671), .ZN(n13472) );
  XOR2HSV0 U16326 ( .A1(n27676), .A2(n13472), .Z(n13473) );
  XOR2HSV0 U16327 ( .A1(n27670), .A2(n27669), .Z(n13474) );
  XOR2HSV0 U16328 ( .A1(n13473), .A2(n13474), .Z(n13475) );
  MUX2NHSV0 U16329 ( .I0(n13470), .I1(n27711), .S(n13475), .ZN(n13476) );
  NAND2HSV0 U16330 ( .A1(n27679), .A2(\pe2/got [2]), .ZN(n13479) );
  NAND2HSV0 U16331 ( .A1(n13479), .A2(n13478), .ZN(n13480) );
  OAI21HSV2 U16332 ( .A1(n13478), .A2(n13479), .B(n13480), .ZN(n27680) );
  NAND2HSV0 U16333 ( .A1(n23458), .A2(n23470), .ZN(n13483) );
  NAND2HSV0 U16334 ( .A1(n13483), .A2(poh11[8]), .ZN(n13484) );
  OAI21HSV2 U16335 ( .A1(poh11[8]), .A2(n13483), .B(n13484), .ZN(po[9]) );
  NAND2HSV0 U16336 ( .A1(n26220), .A2(n26221), .ZN(n13487) );
  OAI21HSV0 U16337 ( .A1(n13486), .A2(n13487), .B(n13488), .ZN(po10) );
  CLKNHSV0 U16338 ( .I(n24049), .ZN(n13489) );
  NAND2HSV0 U16339 ( .A1(\pe7/got [4]), .A2(n28659), .ZN(n13490) );
  MUX2NHSV1 U16340 ( .I0(n13489), .I1(n24049), .S(n13490), .ZN(\pe7/poht [12])
         );
  NAND2HSV0 U16341 ( .A1(n26759), .A2(\pe3/got [5]), .ZN(n13491) );
  CLKNAND2HSV0 U16342 ( .A1(n13491), .A2(n24521), .ZN(n13492) );
  OAI21HSV0 U16343 ( .A1(n24521), .A2(n13491), .B(n13492), .ZN(n13493) );
  NAND2HSV0 U16344 ( .A1(n24522), .A2(\pe3/got [6]), .ZN(n13494) );
  CLKNAND2HSV0 U16345 ( .A1(n13494), .A2(n13493), .ZN(n13495) );
  NAND2HSV0 U16346 ( .A1(n26600), .A2(\pe3/got [7]), .ZN(n13497) );
  CLKNAND2HSV2 U16347 ( .A1(n13497), .A2(n13496), .ZN(n13498) );
  OAI21HSV0 U16348 ( .A1(n13496), .A2(n13497), .B(n13498), .ZN(\pe3/poht [9])
         );
  INOR2HSV0 U16349 ( .A1(n23421), .B1(n23422), .ZN(n13499) );
  CLKNHSV0 U16350 ( .I(n18002), .ZN(n13501) );
  MUX2NHSV4 U16351 ( .I0(n18002), .I1(n13501), .S(n13502), .ZN(n29001) );
  CLKNAND2HSV2 U16352 ( .A1(n13503), .A2(n15567), .ZN(n28696) );
  XOR2HSV0 U16353 ( .A1(n23432), .A2(n23431), .Z(n13504) );
  NAND2HSV0 U16354 ( .A1(n27218), .A2(n22067), .ZN(n13505) );
  NAND2HSV0 U16355 ( .A1(n13505), .A2(n13504), .ZN(n13506) );
  OAI21HSV0 U16356 ( .A1(n13504), .A2(n13505), .B(n13506), .ZN(n29046) );
  AOI21HSV0 U16357 ( .A1(n25624), .A2(n25203), .B(n22252), .ZN(n13507) );
  AO31HSV2 U16358 ( .A1(n25624), .A2(n25203), .A3(n22252), .B(n13507), .Z(
        n19912) );
  INOR2HSV2 U16359 ( .A1(n15643), .B1(n22115), .ZN(n13508) );
  NAND2HSV0 U16360 ( .A1(\pe4/aot [16]), .A2(\pe4/bq[11] ), .ZN(n13509) );
  NAND2HSV2 U16361 ( .A1(n13509), .A2(n13508), .ZN(n13510) );
  OAI21HSV2 U16362 ( .A1(n13508), .A2(n13509), .B(n13510), .ZN(n15503) );
  NAND2HSV0 U16363 ( .A1(n20157), .A2(\pe11/bq[10] ), .ZN(n13511) );
  OAI21HSV0 U16364 ( .A1(n24314), .A2(n20385), .B(n13511), .ZN(n13512) );
  OAI31HSV0 U16365 ( .A1(n24314), .A2(n13511), .A3(n20385), .B(n13512), .ZN(
        n20337) );
  NAND2HSV0 U16366 ( .A1(n28811), .A2(\pe10/pvq [15]), .ZN(n13513) );
  NAND2HSV2 U16367 ( .A1(n13513), .A2(\pe10/phq [15]), .ZN(n13514) );
  OAI21HSV2 U16368 ( .A1(\pe10/phq [15]), .A2(n13513), .B(n13514), .ZN(n22448)
         );
  NAND2HSV0 U16369 ( .A1(\pe7/bq[11] ), .A2(\pe7/aot [14]), .ZN(n13515) );
  OAI21HSV0 U16370 ( .A1(n19492), .A2(n25278), .B(n13515), .ZN(n13516) );
  OAI31HSV2 U16371 ( .A1(n19492), .A2(n13515), .A3(n25278), .B(n13516), .ZN(
        n19433) );
  INOR2HSV0 U16372 ( .A1(\pe2/aot [7]), .B1(n27322), .ZN(n13517) );
  NAND2HSV0 U16373 ( .A1(\pe2/aot [10]), .A2(\pe2/bq[13] ), .ZN(n13518) );
  NAND2HSV0 U16374 ( .A1(n13518), .A2(n13517), .ZN(n13519) );
  OAI21HSV0 U16375 ( .A1(n13517), .A2(n13518), .B(n13519), .ZN(n21125) );
  NAND2HSV0 U16376 ( .A1(\pe9/got [13]), .A2(\pe9/ti_1 ), .ZN(n13521) );
  NAND2HSV0 U16377 ( .A1(n13521), .A2(n13520), .ZN(n13522) );
  OAI21HSV2 U16378 ( .A1(n13520), .A2(n13521), .B(n13522), .ZN(n13523) );
  NAND2HSV0 U16379 ( .A1(n21761), .A2(\pe9/aot [14]), .ZN(n13524) );
  NAND2HSV2 U16380 ( .A1(n13524), .A2(n13523), .ZN(n13525) );
  NOR2HSV0 U16381 ( .A1(n14738), .A2(n18996), .ZN(n13526) );
  CLKNHSV0 U16382 ( .I(n26097), .ZN(n13527) );
  NAND2HSV0 U16383 ( .A1(\pe10/aot [3]), .A2(\pe10/bq[5] ), .ZN(n13528) );
  NAND2HSV0 U16384 ( .A1(n13528), .A2(n22766), .ZN(n13529) );
  OAI21HSV2 U16385 ( .A1(n22766), .A2(n13528), .B(n13529), .ZN(n13530) );
  OAI21HSV0 U16386 ( .A1(n26163), .A2(n26102), .B(n13530), .ZN(n13531) );
  OAI31HSV2 U16387 ( .A1(n26163), .A2(n13530), .A3(n26102), .B(n13531), .ZN(
        n13532) );
  MUX2NHSV1 U16388 ( .I0(n26097), .I1(n13527), .S(n13532), .ZN(n22772) );
  XOR2HSV0 U16389 ( .A1(n26051), .A2(n26052), .Z(n13533) );
  XOR2HSV0 U16390 ( .A1(n26053), .A2(n26054), .Z(n13534) );
  XOR2HSV0 U16391 ( .A1(n13533), .A2(n13534), .Z(n26055) );
  NAND2HSV0 U16392 ( .A1(\pe5/bq[6] ), .A2(\pe5/aot [8]), .ZN(n13535) );
  OAI21HSV0 U16393 ( .A1(n23924), .A2(n23923), .B(n13535), .ZN(n13536) );
  OAI31HSV0 U16394 ( .A1(n23924), .A2(n13535), .A3(n23923), .B(n13536), .ZN(
        n23925) );
  AOI22HSV0 U16395 ( .A1(\pe1/bq[1] ), .A2(n28468), .B1(\pe1/bq[5] ), .B2(
        \pe1/aot [11]), .ZN(n13537) );
  IAO21HSV2 U16396 ( .A1(n26542), .A2(n27150), .B(n13537), .ZN(n26543) );
  NOR2HSV4 U16397 ( .A1(n15704), .A2(n15900), .ZN(n13538) );
  NAND2HSV4 U16398 ( .A1(n22931), .A2(n13538), .ZN(n15685) );
  NAND2HSV0 U16399 ( .A1(\pe6/ti_7[1] ), .A2(\pe6/got [9]), .ZN(n13539) );
  CLKNAND2HSV0 U16400 ( .A1(n13539), .A2(n14390), .ZN(n13540) );
  NAND2HSV0 U16401 ( .A1(n18930), .A2(\pe6/got [10]), .ZN(n13542) );
  CLKNAND2HSV0 U16402 ( .A1(n13542), .A2(n13541), .ZN(n13543) );
  OAI21HSV2 U16403 ( .A1(n13541), .A2(n13542), .B(n13543), .ZN(n13544) );
  NAND2HSV0 U16404 ( .A1(n19076), .A2(n28586), .ZN(n13545) );
  CLKNAND2HSV0 U16405 ( .A1(n13545), .A2(n13544), .ZN(n13546) );
  OAI21HSV2 U16406 ( .A1(n13544), .A2(n13545), .B(n13546), .ZN(n13547) );
  CLKNAND2HSV0 U16407 ( .A1(n19109), .A2(n28593), .ZN(n13548) );
  NAND2HSV2 U16408 ( .A1(n13548), .A2(n13547), .ZN(n13549) );
  OAI21HSV2 U16409 ( .A1(n13547), .A2(n13548), .B(n13549), .ZN(n14392) );
  CLKNHSV0 U16410 ( .I(\pe2/aot [3]), .ZN(n13550) );
  OAI21HSV0 U16411 ( .A1(n27710), .A2(n13550), .B(n27709), .ZN(n13551) );
  NAND2HSV0 U16412 ( .A1(\pe2/aot [2]), .A2(n27706), .ZN(n13552) );
  CLKNHSV0 U16413 ( .I(n27707), .ZN(n13553) );
  AOI22HSV0 U16414 ( .A1(n27708), .A2(n13552), .B1(n27733), .B2(n13553), .ZN(
        n13554) );
  OAI21HSV0 U16415 ( .A1(n27711), .A2(n27734), .B(n13551), .ZN(n13555) );
  NAND2HSV0 U16416 ( .A1(n13555), .A2(n13554), .ZN(n13556) );
  OAI21HSV0 U16417 ( .A1(n13555), .A2(n13554), .B(n13556), .ZN(n13557) );
  NAND2HSV0 U16418 ( .A1(\pe2/aot [1]), .A2(\pe2/bq[5] ), .ZN(n13558) );
  CLKNAND2HSV0 U16419 ( .A1(n13558), .A2(n13557), .ZN(n13559) );
  OAI21HSV0 U16420 ( .A1(n13557), .A2(n13558), .B(n13559), .ZN(n27713) );
  AOI22HSV2 U16421 ( .A1(n28967), .A2(n27354), .B1(\pe2/ti_7t [14]), .B2(
        n27571), .ZN(n27646) );
  CLKNAND2HSV2 U16422 ( .A1(n23805), .A2(n23804), .ZN(n13560) );
  NAND3HSV2 U16423 ( .A1(n13560), .A2(n23802), .A3(n23803), .ZN(n26600) );
  XOR2HSV0 U16424 ( .A1(n27487), .A2(n27486), .Z(n13561) );
  OAI21HSV0 U16425 ( .A1(n27527), .A2(n27718), .B(n13561), .ZN(n13562) );
  OAI31HSV0 U16426 ( .A1(n27594), .A2(n13561), .A3(n27718), .B(n13562), .ZN(
        n13563) );
  OAI21HSV0 U16427 ( .A1(n27595), .A2(n27663), .B(n13563), .ZN(n13564) );
  OAI31HSV0 U16428 ( .A1(n27595), .A2(n13563), .A3(n27663), .B(n13564), .ZN(
        n13565) );
  NAND2HSV0 U16429 ( .A1(n27614), .A2(n14003), .ZN(n13566) );
  NAND2HSV0 U16430 ( .A1(n13566), .A2(n13565), .ZN(n13567) );
  OAI21HSV2 U16431 ( .A1(n13565), .A2(n13566), .B(n13567), .ZN(n13568) );
  OAI21HSV0 U16432 ( .A1(n27634), .A2(n27572), .B(n13568), .ZN(n13569) );
  OAI31HSV2 U16433 ( .A1(n27634), .A2(n13568), .A3(n27572), .B(n13569), .ZN(
        n13570) );
  NAND2HSV0 U16434 ( .A1(n28474), .A2(\pe2/got [8]), .ZN(n13571) );
  CLKNAND2HSV0 U16435 ( .A1(n13571), .A2(n13570), .ZN(n13572) );
  OAI21HSV0 U16436 ( .A1(n13570), .A2(n13571), .B(n13572), .ZN(n27488) );
  CLKNHSV0 U16437 ( .I(n17945), .ZN(n13573) );
  AOI21HSV2 U16438 ( .A1(n18650), .A2(n17945), .B(n17950), .ZN(n13574) );
  OAI21HSV4 U16439 ( .A1(n17946), .A2(n13573), .B(n13574), .ZN(n25638) );
  INHSV4 U16440 ( .I(n15051), .ZN(n13575) );
  CLKNAND2HSV0 U16441 ( .A1(n15049), .A2(n15050), .ZN(n13576) );
  MUX2NHSV4 U16442 ( .I0(n15051), .I1(n13575), .S(n13576), .ZN(n23481) );
  OAI21HSV0 U16443 ( .A1(n25515), .A2(n25516), .B(poh11[6]), .ZN(n13577) );
  OAI31HSV0 U16444 ( .A1(n25515), .A2(poh11[6]), .A3(n25516), .B(n13577), .ZN(
        po[7]) );
  NAND2HSV0 U16445 ( .A1(\pe10/got [11]), .A2(n25060), .ZN(n13579) );
  NAND2HSV0 U16446 ( .A1(n26212), .A2(n26221), .ZN(n13582) );
  OAI21HSV0 U16447 ( .A1(n13581), .A2(n13582), .B(n13583), .ZN(\pe10/poht [4])
         );
  CLKNHSV0 U16448 ( .I(n26226), .ZN(n13584) );
  MUX2NHSV0 U16449 ( .I0(n13584), .I1(n26226), .S(n26227), .ZN(n13585) );
  XOR2HSV0 U16450 ( .A1(n26228), .A2(n13585), .Z(n13586) );
  NAND2HSV0 U16451 ( .A1(n25525), .A2(\pe8/got [2]), .ZN(n13587) );
  CLKNAND2HSV0 U16452 ( .A1(n13587), .A2(n13586), .ZN(n13588) );
  OAI21HSV0 U16453 ( .A1(n13586), .A2(n13587), .B(n13588), .ZN(n13589) );
  OAI21HSV0 U16454 ( .A1(n13589), .A2(n13590), .B(n13591), .ZN(\pe8/poht [13])
         );
  XOR2HSV0 U16455 ( .A1(n24901), .A2(n24900), .Z(n13592) );
  CLKNHSV0 U16456 ( .I(n12303), .ZN(n13596) );
  INHSV2 U16457 ( .I(n16607), .ZN(n13598) );
  MUX2NHSV2 U16458 ( .I0(n13598), .I1(n16607), .S(n16606), .ZN(n13599) );
  MUX2NHSV4 U16459 ( .I0(n13597), .I1(n16608), .S(n13599), .ZN(n29007) );
  CLKNAND2HSV0 U16460 ( .A1(n13600), .A2(n25684), .ZN(n13601) );
  OAI21HSV0 U16461 ( .A1(n13600), .A2(n25684), .B(n13601), .ZN(pov9[13]) );
  AOI21HSV4 U16462 ( .A1(n19155), .A2(n19156), .B(n19057), .ZN(n29019) );
  OAI21HSV0 U16463 ( .A1(n22796), .A2(n26930), .B(n26928), .ZN(n13602) );
  NAND2HSV0 U16464 ( .A1(n27125), .A2(n27126), .ZN(n13603) );
  NAND2HSV0 U16465 ( .A1(n13603), .A2(n27127), .ZN(n13604) );
  OAI21HSV0 U16466 ( .A1(n27127), .A2(n13603), .B(n13604), .ZN(n28963) );
  AOI21HSV0 U16467 ( .A1(n26426), .A2(n27218), .B(n25627), .ZN(n13605) );
  AO31HSV2 U16468 ( .A1(n26426), .A2(n27218), .A3(n25627), .B(n13605), .Z(
        n29051) );
  INOR2HSV2 U16469 ( .A1(n20505), .B1(n20229), .ZN(n20244) );
  INOR2HSV2 U16470 ( .A1(n15146), .B1(n14041), .ZN(n15088) );
  INOR2HSV0 U16471 ( .A1(\pe2/aot [6]), .B1(n27322), .ZN(n13606) );
  NAND2HSV0 U16472 ( .A1(\pe2/aot [7]), .A2(\pe2/bq[15] ), .ZN(n13607) );
  CLKNAND2HSV0 U16473 ( .A1(n13607), .A2(n13606), .ZN(n13608) );
  OAI21HSV0 U16474 ( .A1(n13606), .A2(n13607), .B(n13608), .ZN(n21182) );
  INOR2HSV0 U16475 ( .A1(n28424), .B1(n26163), .ZN(n13609) );
  CLKNHSV0 U16476 ( .I(n26162), .ZN(n13610) );
  OAI22HSV0 U16477 ( .A1(n26164), .A2(n13609), .B1(n26165), .B2(n13610), .ZN(
        n26169) );
  AOI22HSV0 U16478 ( .A1(\pe7/aot [14]), .A2(\pe7/bq[3] ), .B1(\pe7/bq[6] ), 
        .B2(\pe7/aot [11]), .ZN(n13611) );
  IAO21HSV2 U16479 ( .A1(n25280), .A2(n25279), .B(n13611), .ZN(n25281) );
  NAND2HSV0 U16480 ( .A1(\pe2/bq[8] ), .A2(\pe2/aot [9]), .ZN(n13612) );
  OAI21HSV0 U16481 ( .A1(n27462), .A2(n27654), .B(n13612), .ZN(n13613) );
  OAI31HSV0 U16482 ( .A1(n27462), .A2(n13612), .A3(n27654), .B(n13613), .ZN(
        n27304) );
  XOR2HSV0 U16483 ( .A1(n16567), .A2(n16568), .Z(n13614) );
  XOR2HSV0 U16484 ( .A1(n16563), .A2(n16562), .Z(n13615) );
  CLKXOR2HSV4 U16485 ( .A1(n13614), .A2(n13615), .Z(n13616) );
  NAND2HSV0 U16486 ( .A1(\pe8/aot [12]), .A2(\pe8/bq[12] ), .ZN(n13617) );
  CLKNAND2HSV0 U16487 ( .A1(n13617), .A2(n16570), .ZN(n13618) );
  OAI21HSV0 U16488 ( .A1(n16570), .A2(n13617), .B(n13618), .ZN(n13619) );
  NAND2HSV0 U16489 ( .A1(\pe8/bq[9] ), .A2(\pe8/aot [15]), .ZN(n13620) );
  CLKNAND2HSV0 U16490 ( .A1(n13620), .A2(n13619), .ZN(n13621) );
  OAI21HSV0 U16491 ( .A1(n13619), .A2(n13620), .B(n13621), .ZN(n13622) );
  NAND2HSV0 U16492 ( .A1(\pe8/aot [8]), .A2(n25539), .ZN(n13623) );
  CLKNAND2HSV0 U16493 ( .A1(n13623), .A2(n13622), .ZN(n13624) );
  OAI21HSV0 U16494 ( .A1(n13622), .A2(n13623), .B(n13624), .ZN(n13625) );
  XOR2HSV4 U16495 ( .A1(n13616), .A2(n13625), .Z(n16571) );
  CLKNHSV0 U16496 ( .I(n15941), .ZN(n13626) );
  NAND2HSV0 U16497 ( .A1(\pe3/pvq [8]), .A2(\pe3/ctrq ), .ZN(n13627) );
  NAND2HSV2 U16498 ( .A1(n13627), .A2(\pe3/phq [8]), .ZN(n13628) );
  OAI21HSV2 U16499 ( .A1(\pe3/phq [8]), .A2(n13627), .B(n13628), .ZN(n13629)
         );
  MUX2NHSV0 U16500 ( .I0(n15941), .I1(n13626), .S(n13629), .ZN(n15213) );
  AO22HSV2 U16501 ( .A1(\pe1/aot [4]), .A2(\pe1/bq[13] ), .B1(\pe1/bq[5] ), 
        .B2(\pe1/aot [12]), .Z(n13630) );
  OAI21HSV2 U16502 ( .A1(n26858), .A2(n26439), .B(n13630), .ZN(n26440) );
  CLKNHSV0 U16503 ( .I(n20160), .ZN(n13631) );
  MUX2NHSV4 U16504 ( .I0(n20160), .I1(n13631), .S(n20161), .ZN(n20188) );
  NAND2HSV0 U16505 ( .A1(n15845), .A2(n25131), .ZN(n13632) );
  NOR2HSV2 U16506 ( .A1(n15846), .A2(n13632), .ZN(n15891) );
  INAND2HSV2 U16507 ( .A1(\pe8/ti_7t [1]), .B1(n16504), .ZN(n16414) );
  NAND2HSV0 U16508 ( .A1(\pe6/ti_1 ), .A2(\pe6/got [13]), .ZN(n13633) );
  NAND2HSV0 U16509 ( .A1(n13634), .A2(n13633), .ZN(n13635) );
  OAI21HSV2 U16510 ( .A1(n13633), .A2(n13634), .B(n13635), .ZN(n14168) );
  INOR2HSV2 U16511 ( .A1(\pe6/ti_7t [5]), .B1(n14698), .ZN(n14368) );
  AOI22HSV0 U16512 ( .A1(\pe9/bq[5] ), .A2(\pe9/aot [3]), .B1(\pe9/aot [1]), 
        .B2(\pe9/bq[7] ), .ZN(n13636) );
  IAO21HSV2 U16513 ( .A1(n28325), .A2(n28324), .B(n13636), .ZN(n28327) );
  CLKNHSV0 U16514 ( .I(n17700), .ZN(n13637) );
  MUX2NHSV1 U16515 ( .I0(n17700), .I1(n13637), .S(n13638), .ZN(n17706) );
  OA21HSV4 U16516 ( .A1(n17951), .A2(n18214), .B(n18338), .Z(n17991) );
  NAND2HSV0 U16517 ( .A1(n20987), .A2(n24634), .ZN(n13639) );
  INHSV2 U16518 ( .I(n21889), .ZN(n13640) );
  MUX2NHSV2 U16519 ( .I0(n21889), .I1(n13640), .S(n21890), .ZN(n21904) );
  XOR2HSV0 U16520 ( .A1(n15735), .A2(n15736), .Z(n13641) );
  XOR2HSV0 U16521 ( .A1(n15730), .A2(n15729), .Z(n13642) );
  XOR2HSV0 U16522 ( .A1(n13641), .A2(n13642), .Z(n13643) );
  CLKNHSV0 U16523 ( .I(n22001), .ZN(n13644) );
  MUX2NHSV0 U16524 ( .I0(n13644), .I1(n22001), .S(n15738), .ZN(n13645) );
  XOR2HSV0 U16525 ( .A1(n13643), .A2(n15739), .Z(n13646) );
  XOR2HSV0 U16526 ( .A1(n13645), .A2(n13646), .Z(n13647) );
  NAND2HSV0 U16527 ( .A1(n13996), .A2(n28653), .ZN(n13648) );
  NAND2HSV2 U16528 ( .A1(n13648), .A2(n13647), .ZN(n13649) );
  OAI21HSV2 U16529 ( .A1(n13647), .A2(n13648), .B(n13649), .ZN(n13650) );
  NAND2HSV0 U16530 ( .A1(n28671), .A2(\pe4/got [8]), .ZN(n13651) );
  NAND2HSV0 U16531 ( .A1(n13651), .A2(n13650), .ZN(n13652) );
  OAI21HSV0 U16532 ( .A1(n13650), .A2(n13651), .B(n13652), .ZN(n13653) );
  NAND2HSV0 U16533 ( .A1(n27739), .A2(\pe4/got [10]), .ZN(n13654) );
  NAND2HSV0 U16534 ( .A1(n13654), .A2(n13653), .ZN(n13655) );
  OAI21HSV2 U16535 ( .A1(n13653), .A2(n13654), .B(n13655), .ZN(n15741) );
  INHSV4 U16536 ( .I(n16744), .ZN(n13656) );
  AOI31HSV2 U16537 ( .A1(n19703), .A2(n19683), .A3(n19682), .B(n19765), .ZN(
        n13657) );
  INHSV2 U16538 ( .I(n21156), .ZN(n13659) );
  MUX2NHSV2 U16539 ( .I0(n13659), .I1(n21156), .S(n21155), .ZN(n13660) );
  CLKNHSV0 U16540 ( .I(n23559), .ZN(n13661) );
  NAND2HSV0 U16541 ( .A1(\pe7/got [3]), .A2(n24284), .ZN(n13662) );
  MUX2NHSV1 U16542 ( .I0(n13661), .I1(n23559), .S(n13662), .ZN(\pe7/poht [13])
         );
  CLKNHSV0 U16543 ( .I(\pe10/pq ), .ZN(n13663) );
  MUX2NHSV0 U16544 ( .I0(n13663), .I1(n26185), .S(n28811), .ZN(\pe10/ti_1t )
         );
  NAND2HSV0 U16545 ( .A1(n23757), .A2(n25203), .ZN(n13664) );
  CLKNAND2HSV0 U16546 ( .A1(n13664), .A2(n23774), .ZN(n13665) );
  OAI21HSV0 U16547 ( .A1(n23774), .A2(n13664), .B(n13665), .ZN(n13666) );
  NAND2HSV0 U16548 ( .A1(n26231), .A2(\pe8/got [5]), .ZN(n13667) );
  CLKNAND2HSV0 U16549 ( .A1(n13667), .A2(n13666), .ZN(n13668) );
  OAI21HSV0 U16550 ( .A1(n13666), .A2(n13667), .B(n13668), .ZN(n13669) );
  NAND2HSV0 U16551 ( .A1(\pe8/got [6]), .A2(n26229), .ZN(n13670) );
  OAI21HSV0 U16552 ( .A1(n13669), .A2(n13670), .B(n13671), .ZN(\pe8/poht [10])
         );
  CLKNHSV0 U16553 ( .I(n18629), .ZN(n13672) );
  OAI21HSV0 U16554 ( .A1(n25689), .A2(n25688), .B(n25687), .ZN(n13675) );
  MUX2NHSV1 U16555 ( .I0(n13674), .I1(n25690), .S(n13675), .ZN(n28980) );
  AOI22HSV2 U16556 ( .A1(n25517), .A2(n12260), .B1(n25520), .B2(n25521), .ZN(
        n29018) );
  OAI21HSV0 U16557 ( .A1(n26730), .A2(n16166), .B(n23442), .ZN(n13676) );
  OAI31HSV0 U16558 ( .A1(n26730), .A2(n23442), .A3(n16166), .B(n13676), .ZN(
        n13677) );
  INAND3HSV0 U16559 ( .A1(n23441), .B1(n23439), .B2(n23440), .ZN(n13678) );
  CLKNAND2HSV0 U16560 ( .A1(n13678), .A2(n13677), .ZN(n13679) );
  OAI21HSV0 U16561 ( .A1(n13677), .A2(n13678), .B(n13679), .ZN(n29035) );
  IOA21HSV4 U16562 ( .A1(n23454), .A2(n20698), .B(n20782), .ZN(n28918) );
  CLKNAND2HSV0 U16563 ( .A1(n13680), .A2(n13681), .ZN(n13682) );
  OAI21HSV0 U16564 ( .A1(n13680), .A2(n13681), .B(n13682), .ZN(\pe5/poht [5])
         );
  CLKNHSV0 U16565 ( .I(n26821), .ZN(n13683) );
  XOR2HSV0 U16566 ( .A1(n26820), .A2(n26819), .Z(n13684) );
  MUX2NHSV0 U16567 ( .I0(n13683), .I1(n26821), .S(n13684), .ZN(n13685) );
  NAND3HSV0 U16568 ( .A1(n26827), .A2(\pe1/got [1]), .A3(n26828), .ZN(n13686)
         );
  CLKNAND2HSV0 U16569 ( .A1(n13686), .A2(n13685), .ZN(n13687) );
  OAI21HSV0 U16570 ( .A1(n13685), .A2(n13686), .B(n13687), .ZN(n13688) );
  NAND2HSV0 U16571 ( .A1(n26909), .A2(\pe1/got [2]), .ZN(n13689) );
  CLKNAND2HSV0 U16572 ( .A1(n13689), .A2(n13688), .ZN(n13690) );
  OAI21HSV0 U16573 ( .A1(n13688), .A2(n13689), .B(n13690), .ZN(n13691) );
  NAND2HSV0 U16574 ( .A1(\pe1/got [3]), .A2(n28600), .ZN(n13692) );
  CLKNAND2HSV0 U16575 ( .A1(n13692), .A2(n13691), .ZN(n13693) );
  OAI21HSV0 U16576 ( .A1(n13691), .A2(n13692), .B(n13693), .ZN(\pe1/poht [13])
         );
  CLKNAND2HSV0 U16577 ( .A1(n25633), .A2(n28688), .ZN(n13694) );
  NAND2HSV0 U16578 ( .A1(n13694), .A2(n25634), .ZN(n13695) );
  OAI21HSV0 U16579 ( .A1(n25634), .A2(n13694), .B(n13695), .ZN(n29003) );
  CLKNHSV0 U16580 ( .I(n11858), .ZN(n13696) );
  OAI21HSV0 U16581 ( .A1(n27134), .A2(n13696), .B(n25629), .ZN(n13697) );
  OAI31HSV0 U16582 ( .A1(n27134), .A2(n25629), .A3(n13696), .B(n13697), .ZN(
        n29017) );
  CLKNAND2HSV0 U16583 ( .A1(n25880), .A2(n27218), .ZN(n13698) );
  NAND2HSV0 U16584 ( .A1(n13698), .A2(n23461), .ZN(n13699) );
  OAI21HSV0 U16585 ( .A1(n23461), .A2(n13698), .B(n13699), .ZN(n29048) );
  NAND2HSV2 U16586 ( .A1(n15937), .A2(\pe3/pvq [12]), .ZN(n13700) );
  NAND2HSV2 U16587 ( .A1(n13700), .A2(\pe3/phq [12]), .ZN(n13701) );
  OAI21HSV2 U16588 ( .A1(\pe3/phq [12]), .A2(n13700), .B(n13701), .ZN(n15938)
         );
  NAND2HSV0 U16589 ( .A1(n15737), .A2(\pe4/bq[12] ), .ZN(n13703) );
  NAND2HSV2 U16590 ( .A1(n13703), .A2(n13702), .ZN(n13704) );
  OAI21HSV2 U16591 ( .A1(n13702), .A2(n13703), .B(n13704), .ZN(n15459) );
  NAND2HSV0 U16592 ( .A1(\pe5/aot [7]), .A2(\pe5/bq[2] ), .ZN(n13705) );
  CLKNHSV0 U16593 ( .I(n23254), .ZN(n13706) );
  AOI22HSV0 U16594 ( .A1(n23255), .A2(n13705), .B1(n24389), .B2(n13706), .ZN(
        n23256) );
  AOI22HSV0 U16595 ( .A1(\pe7/bq[2] ), .A2(\pe7/aot [15]), .B1(\pe7/bq[1] ), 
        .B2(n14078), .ZN(n13707) );
  IAO21HSV2 U16596 ( .A1(n25303), .A2(n25302), .B(n13707), .ZN(n25304) );
  AOI22HSV0 U16597 ( .A1(\pe10/bq[3] ), .A2(\pe10/aot [6]), .B1(\pe10/bq[4] ), 
        .B2(\pe10/aot [5]), .ZN(n13708) );
  IAO21HSV0 U16598 ( .A1(n22769), .A2(n22601), .B(n13708), .ZN(n22575) );
  INOR2HSV0 U16599 ( .A1(\pe7/ti_7t [3]), .B1(n25494), .ZN(n19282) );
  INOR2HSV0 U16600 ( .A1(\pe8/ti_7t [5]), .B1(n18787), .ZN(n16508) );
  CLKNAND2HSV2 U16601 ( .A1(\pe4/pvq [1]), .A2(\pe4/phq [1]), .ZN(n13709) );
  NOR2HSV0 U16602 ( .A1(n15502), .A2(n13709), .ZN(n15341) );
  INAND2HSV2 U16603 ( .A1(n23666), .B1(\pe3/ti_7t [15]), .ZN(n23802) );
  INAND2HSV0 U16604 ( .A1(\pe2/ti_7t [3]), .B1(n21901), .ZN(n17702) );
  INAND2HSV0 U16605 ( .A1(\pe6/ti_7t [7]), .B1(n19055), .ZN(n14400) );
  INOR2HSV0 U16606 ( .A1(\pe7/ti_7t [12]), .B1(n19623), .ZN(n19696) );
  INAND2HSV0 U16607 ( .A1(\pe5/ti_7t [10]), .B1(ctro5), .ZN(n20987) );
  INAND2HSV2 U16608 ( .A1(\pe10/ti_7t [4]), .B1(n17119), .ZN(n16735) );
  NAND2HSV0 U16609 ( .A1(\pe6/bq[14] ), .A2(\pe6/aot [16]), .ZN(n13710) );
  NAND2HSV0 U16610 ( .A1(\pe6/aot [14]), .A2(\pe6/bq[16] ), .ZN(n13711) );
  NAND2HSV0 U16611 ( .A1(n13711), .A2(n13710), .ZN(n13712) );
  OAI21HSV2 U16612 ( .A1(n13710), .A2(n13711), .B(n13712), .ZN(n14141) );
  INAND2HSV2 U16613 ( .A1(\pe8/ti_7t [8]), .B1(n22138), .ZN(n18655) );
  INHSV4 U16614 ( .I(n17869), .ZN(n13713) );
  MUX2NHSV4 U16615 ( .I0(n17869), .I1(n13713), .S(n13714), .ZN(n29039) );
  INOR2HSV0 U16616 ( .A1(\pe3/ti_7t [2]), .B1(n15191), .ZN(n15096) );
  NAND2HSV0 U16617 ( .A1(n26068), .A2(\pe6/got [2]), .ZN(n13715) );
  NAND2HSV0 U16618 ( .A1(n14008), .A2(n25952), .ZN(n13717) );
  NAND2HSV0 U16619 ( .A1(n13717), .A2(n13716), .ZN(n13718) );
  OAI21HSV0 U16620 ( .A1(n25981), .A2(n25951), .B(n13719), .ZN(n13720) );
  OAI31HSV0 U16621 ( .A1(n25981), .A2(n13719), .A3(n25951), .B(n13720), .ZN(
        n25972) );
  INOR2HSV1 U16622 ( .A1(\pe4/ti_7t [4]), .B1(n15484), .ZN(n15491) );
  AND2HSV2 U16623 ( .A1(\pe5/got [15]), .A2(n14474), .Z(n14496) );
  XOR2HSV0 U16624 ( .A1(n28314), .A2(n28313), .Z(n13721) );
  NAND2HSV0 U16625 ( .A1(n28394), .A2(n28405), .ZN(n13722) );
  CLKNAND2HSV0 U16626 ( .A1(n13722), .A2(n13721), .ZN(n13723) );
  OAI21HSV0 U16627 ( .A1(n13721), .A2(n13722), .B(n13723), .ZN(n13724) );
  NAND3HSV2 U16628 ( .A1(n28403), .A2(n28369), .A3(n28373), .ZN(n13725) );
  OAI21HSV2 U16629 ( .A1(n13724), .A2(n13725), .B(n13726), .ZN(n13727) );
  NAND2HSV0 U16630 ( .A1(n28643), .A2(n28390), .ZN(n13728) );
  CLKNAND2HSV0 U16631 ( .A1(n13728), .A2(n13727), .ZN(n13729) );
  OAI21HSV0 U16632 ( .A1(n13727), .A2(n13728), .B(n13729), .ZN(\pe9/poht [11])
         );
  XOR2HSV0 U16633 ( .A1(n27733), .A2(n27732), .Z(n13730) );
  XOR2HSV0 U16634 ( .A1(n27734), .A2(n13730), .Z(n13731) );
  OAI21HSV0 U16635 ( .A1(n13731), .A2(n13732), .B(n13733), .ZN(n13734) );
  NAND2HSV0 U16636 ( .A1(n14052), .A2(n27727), .ZN(n13736) );
  CLKNAND2HSV0 U16637 ( .A1(n13736), .A2(n13735), .ZN(n13737) );
  OAI21HSV0 U16638 ( .A1(n13735), .A2(n13736), .B(n13737), .ZN(\pe2/poht [13])
         );
  NAND2HSV0 U16639 ( .A1(n28426), .A2(\pe8/got [8]), .ZN(n13738) );
  CLKNAND2HSV0 U16640 ( .A1(n13738), .A2(n23756), .ZN(n13739) );
  OAI21HSV0 U16641 ( .A1(n23756), .A2(n13738), .B(n13739), .ZN(n13740) );
  NAND2HSV0 U16642 ( .A1(n23721), .A2(n25525), .ZN(n13741) );
  CLKNAND2HSV0 U16643 ( .A1(n13741), .A2(n13740), .ZN(n13742) );
  OAI21HSV0 U16644 ( .A1(n13740), .A2(n13741), .B(n13742), .ZN(n13743) );
  NAND2HSV0 U16645 ( .A1(\pe8/got [10]), .A2(n26229), .ZN(n13744) );
  OAI21HSV0 U16646 ( .A1(n13743), .A2(n13744), .B(n13745), .ZN(\pe8/poht [6])
         );
  MUX2NHSV2 U16647 ( .I0(n16310), .I1(n13746), .S(n16309), .ZN(n29012) );
  CLKNHSV0 U16648 ( .I(n23668), .ZN(n13747) );
  AOI32HSV0 U16649 ( .A1(n24522), .A2(n23668), .A3(n26413), .B1(n13747), .B2(
        n23669), .ZN(n28979) );
  XOR2HSV0 U16650 ( .A1(n23326), .A2(n23325), .Z(n13748) );
  AOI21HSV0 U16651 ( .A1(n24893), .A2(\pe11/got [1]), .B(n13748), .ZN(n13749)
         );
  NAND2HSV0 U16652 ( .A1(n25182), .A2(\pe11/got [3]), .ZN(n13751) );
  CLKNAND2HSV0 U16653 ( .A1(n13751), .A2(n13750), .ZN(n13752) );
  OAI21HSV0 U16654 ( .A1(n13750), .A2(n13751), .B(n13752), .ZN(\pe11/poht [13]) );
  MUX2NHSV1 U16655 ( .I0(n25258), .I1(n25257), .S(n25690), .ZN(n13753) );
  XOR2HSV4 U16656 ( .A1(n25254), .A2(n25253), .Z(n13754) );
  CLKNAND2HSV0 U16657 ( .A1(n13757), .A2(n13758), .ZN(n13759) );
  CLKNHSV0 U16658 ( .I(n23843), .ZN(n13760) );
  NAND2HSV0 U16659 ( .A1(n24277), .A2(\pe7/got [6]), .ZN(n13761) );
  CLKNHSV0 U16660 ( .I(bo10[14]), .ZN(n13762) );
  MUX2NHSV0 U16661 ( .I0(n13762), .I1(n23509), .S(n23510), .ZN(n28900) );
  INAND3HSV0 U16662 ( .A1(n23463), .B1(n23465), .B2(n23464), .ZN(n13763) );
  NAND2HSV0 U16663 ( .A1(n13763), .A2(n23466), .ZN(n13764) );
  OAI21HSV0 U16664 ( .A1(n23466), .A2(n13763), .B(n13764), .ZN(n28962) );
  CLKNHSV0 U16665 ( .I(\pe9/pq ), .ZN(n13765) );
  MUX2NHSV0 U16666 ( .I0(n13765), .I1(n21334), .S(n27093), .ZN(\pe9/ti_1t ) );
  CLKNHSV0 U16667 ( .I(n27135), .ZN(n13766) );
  OAI211HSV0 U16668 ( .A1(n27134), .A2(n27133), .B(n27132), .C(n27131), .ZN(
        n13767) );
  MUX2NHSV0 U16669 ( .I0(n27135), .I1(n13766), .S(n13767), .ZN(n28983) );
  CLKNHSV0 U16670 ( .I(\pe3/pq ), .ZN(n13768) );
  CLKNHSV0 U16671 ( .I(bo2[9]), .ZN(n13769) );
  MUX2NHSV0 U16672 ( .I0(n13769), .I1(n23502), .S(n23503), .ZN(n28827) );
  CLKNHSV0 U16673 ( .I(n25680), .ZN(n13770) );
  MUX2NHSV0 U16674 ( .I0(n12282), .I1(n13770), .S(n25679), .ZN(n13771) );
  OAI21HSV0 U16675 ( .A1(n27139), .A2(n25678), .B(n13771), .ZN(n13772) );
  OAI31HSV0 U16676 ( .A1(n27139), .A2(n13771), .A3(n25678), .B(n13772), .ZN(
        pov1[12]) );
  CLKNHSV0 U16677 ( .I(bo1[12]), .ZN(n13773) );
  MUX2NHSV0 U16678 ( .I0(n13773), .I1(n27070), .S(n14024), .ZN(n28742) );
  NOR2HSV0 U16679 ( .A1(n27191), .A2(n24683), .ZN(n13774) );
  NAND2HSV0 U16680 ( .A1(n14071), .A2(n24406), .ZN(n13775) );
  NAND2HSV0 U16681 ( .A1(n13775), .A2(n13774), .ZN(n13776) );
  OAI21HSV2 U16682 ( .A1(n13774), .A2(n13775), .B(n13776), .ZN(n14849) );
  IOA22HSV0 U16683 ( .B1(n22000), .B2(n27846), .A1(n28683), .A2(\pe4/bq[3] ), 
        .ZN(n13777) );
  OAI21HSV2 U16684 ( .A1(n22001), .A2(n22960), .B(n13777), .ZN(n13778) );
  NAND2HSV0 U16685 ( .A1(\pe4/aot [3]), .A2(n26948), .ZN(n13779) );
  NAND2HSV2 U16686 ( .A1(n13779), .A2(n13778), .ZN(n13780) );
  OAI21HSV2 U16687 ( .A1(n13778), .A2(n13779), .B(n13780), .ZN(n22009) );
  CLKNHSV0 U16688 ( .I(n23560), .ZN(n13781) );
  AOI22HSV0 U16689 ( .A1(\pe8/bq[3] ), .A2(\pe8/aot [10]), .B1(\pe8/aot [11]), 
        .B2(\pe8/bq[2] ), .ZN(n13782) );
  AOI21HSV2 U16690 ( .A1(n23561), .A2(n13781), .B(n13782), .ZN(n23565) );
  AOI22HSV0 U16691 ( .A1(\pe3/bq[5] ), .A2(\pe3/aot [7]), .B1(\pe3/aot [2]), 
        .B2(\pe3/bq[10] ), .ZN(n13783) );
  IAO21HSV2 U16692 ( .A1(n26605), .A2(n26604), .B(n13783), .ZN(n26607) );
  CLKNAND2HSV2 U16693 ( .A1(n14669), .A2(n14670), .ZN(n13784) );
  NAND2HSV2 U16694 ( .A1(n22430), .A2(n20136), .ZN(n20134) );
  CLKNHSV0 U16695 ( .I(\pe4/phq [4]), .ZN(n13786) );
  MUX2NHSV1 U16696 ( .I0(\pe4/phq [4]), .I1(n13786), .S(n13787), .ZN(n15378)
         );
  XOR2HSV0 U16697 ( .A1(n20392), .A2(n20391), .Z(n13789) );
  MUX2NHSV4 U16698 ( .I0(n13788), .I1(n20393), .S(n13789), .ZN(n20452) );
  INOR2HSV0 U16699 ( .A1(\pe9/ti_7t [8]), .B1(n18219), .ZN(n18274) );
  INOR2HSV0 U16700 ( .A1(\pe5/ti_7t [9]), .B1(n14757), .ZN(n14865) );
  INOR2HSV0 U16701 ( .A1(\pe4/ti_7t [8]), .B1(n15394), .ZN(n15700) );
  NAND2HSV0 U16702 ( .A1(\pe2/bq[2] ), .A2(\pe2/aot [3]), .ZN(n13790) );
  OAI21HSV0 U16703 ( .A1(n27693), .A2(n27692), .B(n13790), .ZN(n13791) );
  OAI31HSV0 U16704 ( .A1(n27693), .A2(n13790), .A3(n27692), .B(n13791), .ZN(
        n27697) );
  NAND2HSV0 U16705 ( .A1(n25419), .A2(n14400), .ZN(n13792) );
  AOI21HSV2 U16706 ( .A1(n15242), .A2(n15096), .B(n15099), .ZN(n13793) );
  CLKNHSV0 U16707 ( .I(n23470), .ZN(n13794) );
  OAI21HSV0 U16708 ( .A1(n23460), .A2(n13794), .B(poh11[7]), .ZN(n13795) );
  OAI31HSV0 U16709 ( .A1(n23460), .A2(poh11[7]), .A3(n13794), .B(n13795), .ZN(
        po[8]) );
  NAND2HSV0 U16710 ( .A1(\pe10/got [4]), .A2(n23219), .ZN(n13797) );
  CLKNAND2HSV0 U16711 ( .A1(n13797), .A2(n13796), .ZN(n13798) );
  OAI21HSV0 U16712 ( .A1(n13796), .A2(n13797), .B(n13798), .ZN(\pe10/poht [12]) );
  AOI21HSV0 U16713 ( .A1(n23870), .A2(n18767), .B(n23869), .ZN(n13799) );
  XOR2HSV0 U16714 ( .A1(n23864), .A2(n23863), .Z(n13800) );
  XOR2HSV0 U16715 ( .A1(n23865), .A2(n13800), .Z(n13801) );
  NAND2HSV0 U16716 ( .A1(\pe8/got [5]), .A2(n23757), .ZN(n13802) );
  CLKNAND2HSV0 U16717 ( .A1(n13802), .A2(n13801), .ZN(n13803) );
  OAI21HSV0 U16718 ( .A1(n13801), .A2(n13802), .B(n13803), .ZN(n13804) );
  NAND2HSV0 U16719 ( .A1(\pe8/got [6]), .A2(n25525), .ZN(n13805) );
  NAND2HSV0 U16720 ( .A1(n13805), .A2(n13804), .ZN(n13806) );
  OAI21HSV2 U16721 ( .A1(n13804), .A2(n13805), .B(n13806), .ZN(n13807) );
  CLKNAND2HSV0 U16722 ( .A1(n13808), .A2(n13807), .ZN(n13809) );
  CLKNHSV0 U16723 ( .I(n23718), .ZN(n13811) );
  OAI21HSV0 U16724 ( .A1(n23717), .A2(n13811), .B(n23719), .ZN(n13812) );
  NAND3HSV0 U16725 ( .A1(n25371), .A2(n25369), .A3(n25370), .ZN(n13814) );
  NAND2HSV0 U16726 ( .A1(n13814), .A2(n25372), .ZN(n13815) );
  OAI21HSV0 U16727 ( .A1(n25372), .A2(n13814), .B(n13815), .ZN(pov4[15]) );
  CLKNHSV0 U16728 ( .I(n22051), .ZN(n13816) );
  NAND2HSV0 U16729 ( .A1(\pe11/got [10]), .A2(n24957), .ZN(n13818) );
  CLKNAND2HSV0 U16730 ( .A1(n13818), .A2(n13817), .ZN(n13819) );
  OAI21HSV0 U16731 ( .A1(n13817), .A2(n13818), .B(n13819), .ZN(\pe11/poht [6])
         );
  NAND2HSV2 U16732 ( .A1(n24322), .A2(\pe5/got [5]), .ZN(n13821) );
  XOR2HSV0 U16733 ( .A1(n23700), .A2(n23699), .Z(n13823) );
  NAND2HSV0 U16734 ( .A1(n28652), .A2(n28648), .ZN(n13824) );
  NAND2HSV0 U16735 ( .A1(n26760), .A2(\pe3/got [9]), .ZN(n13826) );
  CLKNAND2HSV0 U16736 ( .A1(n13826), .A2(n13825), .ZN(n13827) );
  OAI21HSV0 U16737 ( .A1(n13825), .A2(n13826), .B(n13827), .ZN(n13828) );
  NAND2HSV0 U16738 ( .A1(\pe3/got [10]), .A2(n28661), .ZN(n13829) );
  NAND2HSV0 U16739 ( .A1(n13829), .A2(n13828), .ZN(n13830) );
  OAI21HSV0 U16740 ( .A1(n13828), .A2(n13829), .B(n13830), .ZN(\pe3/poht [6])
         );
  CLKNHSV0 U16741 ( .I(\pe11/pq ), .ZN(n13831) );
  MUX2NHSV0 U16742 ( .I0(n13831), .I1(n22112), .S(n28639), .ZN(\pe11/ti_1t )
         );
  CLKNHSV0 U16743 ( .I(bo11[1]), .ZN(n13832) );
  MUX2NHSV0 U16744 ( .I0(n13832), .I1(n25413), .S(n23499), .ZN(n28727) );
  CLKNAND2HSV0 U16745 ( .A1(n26189), .A2(n26220), .ZN(n13833) );
  NAND2HSV0 U16746 ( .A1(n13833), .A2(n23484), .ZN(n13834) );
  OAI21HSV0 U16747 ( .A1(n13833), .A2(n23484), .B(n13834), .ZN(n28998) );
  CLKNHSV0 U16748 ( .I(bo10[13]), .ZN(n13835) );
  MUX2NHSV0 U16749 ( .I0(n13835), .I1(n23511), .S(n23512), .ZN(n28902) );
  INHSV2 U16750 ( .I(n25639), .ZN(n13836) );
  CLKNHSV0 U16751 ( .I(n25638), .ZN(n13837) );
  MUX2NHSV0 U16752 ( .I0(n13837), .I1(n25638), .S(n25637), .ZN(n13838) );
  MUX2NHSV1 U16753 ( .I0(n13836), .I1(n25639), .S(n13838), .ZN(n29002) );
  CLKNHSV0 U16754 ( .I(n23449), .ZN(n13839) );
  CLKNHSV0 U16755 ( .I(n23448), .ZN(n13840) );
  AO32HSV1 U16756 ( .A1(n18564), .A2(n13839), .A3(n13840), .B1(n23449), .B2(
        n23447), .Z(pov9[11]) );
  CLKNHSV0 U16757 ( .I(bo9[12]), .ZN(n13841) );
  MUX2NHSV0 U16758 ( .I0(n13841), .I1(n27101), .S(n27093), .ZN(n28778) );
  NAND2HSV0 U16759 ( .A1(n25578), .A2(n25523), .ZN(n13842) );
  NAND2HSV0 U16760 ( .A1(n13842), .A2(n22092), .ZN(n13843) );
  OAI21HSV0 U16761 ( .A1(n22092), .A2(n13842), .B(n13843), .ZN(n29009) );
  CLKNHSV0 U16762 ( .I(n14034), .ZN(n13844) );
  MUX2NHSV1 U16763 ( .I0(n13844), .I1(n14034), .S(n25650), .ZN(n13845) );
  OAI21HSV0 U16764 ( .A1(n25652), .A2(n25651), .B(n13845), .ZN(n13846) );
  OAI31HSV0 U16765 ( .A1(n25652), .A2(n13845), .A3(n25651), .B(n13846), .ZN(
        n29008) );
  CLKNHSV0 U16766 ( .I(\pe8/pq ), .ZN(n13847) );
  MUX2NHSV0 U16767 ( .I0(n13847), .I1(n25531), .S(n23545), .ZN(\pe8/ti_1t ) );
  NAND2HSV0 U16768 ( .A1(n11936), .A2(n28610), .ZN(n13848) );
  NAND2HSV0 U16769 ( .A1(n13848), .A2(n22091), .ZN(n13849) );
  OAI21HSV0 U16770 ( .A1(n22091), .A2(n13848), .B(n13849), .ZN(n28987) );
  CLKNHSV0 U16771 ( .I(n25665), .ZN(n13850) );
  NAND2HSV0 U16772 ( .A1(n28816), .A2(n28587), .ZN(n13851) );
  NAND2HSV0 U16773 ( .A1(n13851), .A2(n25664), .ZN(n13852) );
  OAI21HSV2 U16774 ( .A1(n25664), .A2(n13851), .B(n13852), .ZN(n13853) );
  MUX2NHSV1 U16775 ( .I0(n13850), .I1(n25665), .S(n13853), .ZN(\pov7[10] ) );
  CLKNHSV0 U16776 ( .I(\pe7/pq ), .ZN(n13854) );
  MUX2NHSV0 U16777 ( .I0(n13854), .I1(n19243), .S(n28876), .ZN(\pe7/ti_1t ) );
  CLKNHSV0 U16778 ( .I(bo7[8]), .ZN(n13855) );
  MUX2NHSV0 U16779 ( .I0(n13855), .I1(n23497), .S(n27082), .ZN(n28878) );
  NOR2HSV2 U16780 ( .A1(n24962), .A2(n24963), .ZN(n13856) );
  NAND2HSV0 U16781 ( .A1(n13856), .A2(n24964), .ZN(n13857) );
  OAI21HSV0 U16782 ( .A1(n13856), .A2(n24964), .B(n13857), .ZN(n29024) );
  CLKNHSV0 U16783 ( .I(\pe6/pq ), .ZN(n13858) );
  MUX2NHSV0 U16784 ( .I0(n13858), .I1(n13237), .S(n28867), .ZN(\pe6/ti_1t ) );
  CLKNHSV0 U16785 ( .I(bo6[13]), .ZN(n13859) );
  MUX2NHSV0 U16786 ( .I0(n13859), .I1(n22107), .S(n23498), .ZN(n28870) );
  MUX2HSV0 U16787 ( .I0(n25626), .I1(\pe5/pq ), .S(n27051), .Z(\pe5/ti_1t ) );
  CLKNAND2HSV0 U16788 ( .A1(n27052), .A2(bo5[9]), .ZN(n13860) );
  OAI21HSV0 U16789 ( .A1(n27049), .A2(n27052), .B(n13860), .ZN(n28713) );
  NAND2HSV0 U16790 ( .A1(n23482), .A2(n15813), .ZN(n13861) );
  NAND2HSV0 U16791 ( .A1(n13861), .A2(n23483), .ZN(n13862) );
  OAI21HSV0 U16792 ( .A1(n23483), .A2(n13861), .B(n13862), .ZN(n29034) );
  CLKNHSV0 U16793 ( .I(bo3[12]), .ZN(n13863) );
  MUX2NHSV0 U16794 ( .I0(n13863), .I1(n24535), .S(n23518), .ZN(n28840) );
  CLKNHSV0 U16795 ( .I(bo2[7]), .ZN(n13864) );
  MUX2NHSV0 U16796 ( .I0(n13864), .I1(n27461), .S(n27311), .ZN(n28830) );
  CLKNHSV0 U16797 ( .I(n23478), .ZN(n13865) );
  MUX2NHSV0 U16798 ( .I0(n13865), .I1(n23478), .S(n23479), .ZN(n29049) );
  CLKNHSV0 U16799 ( .I(bo1[3]), .ZN(n13866) );
  MUX2NHSV0 U16800 ( .I0(n13866), .I1(n27157), .S(n27062), .ZN(n28821) );
  CLKNHSV0 U16801 ( .I(\pe5/bq[10] ), .ZN(n13867) );
  OAI21HSV0 U16802 ( .A1(n14883), .A2(n13867), .B(n14781), .ZN(n14649) );
  AOI22HSV0 U16803 ( .A1(\pe1/bq[7] ), .A2(\pe1/aot [6]), .B1(\pe1/aot [3]), 
        .B2(\pe1/bq[10] ), .ZN(n13868) );
  IAO21HSV0 U16804 ( .A1(n26770), .A2(n26769), .B(n13868), .ZN(n26771) );
  NOR2HSV0 U16805 ( .A1(n24346), .A2(n21573), .ZN(n13869) );
  OAI22HSV0 U16806 ( .A1(n24389), .A2(n13869), .B1(n21560), .B2(n23233), .ZN(
        n21561) );
  AOI22HSV0 U16807 ( .A1(n27103), .A2(\pe7/aot [3]), .B1(\pe7/aot [2]), .B2(
        n27083), .ZN(n13870) );
  IAO21HSV0 U16808 ( .A1(n25277), .A2(n25276), .B(n13870), .ZN(n25282) );
  AOI22HSV0 U16809 ( .A1(\pe3/bq[7] ), .A2(\pe3/aot [5]), .B1(\pe3/aot [4]), 
        .B2(\pe3/bq[8] ), .ZN(n13871) );
  IAO21HSV0 U16810 ( .A1(n26610), .A2(n26700), .B(n13871), .ZN(n26611) );
  AOI22HSV0 U16811 ( .A1(\pe8/bq[2] ), .A2(\pe8/aot [9]), .B1(\pe8/aot [4]), 
        .B2(\pe8/bq[7] ), .ZN(n13872) );
  IAO21HSV0 U16812 ( .A1(n23727), .A2(n23726), .B(n13872), .ZN(n23728) );
  AOI22HSV0 U16813 ( .A1(\pe10/bq[4] ), .A2(\pe10/aot [3]), .B1(\pe10/bq[3] ), 
        .B2(\pe10/aot [4]), .ZN(n13875) );
  IAO21HSV0 U16814 ( .A1(n22766), .A2(n22703), .B(n13875), .ZN(n22425) );
  AOI22HSV0 U16815 ( .A1(\pe1/bq[9] ), .A2(\pe1/aot [5]), .B1(\pe1/aot [1]), 
        .B2(\pe1/bq[13] ), .ZN(n13876) );
  IAO21HSV0 U16816 ( .A1(n27021), .A2(n27020), .B(n13876), .ZN(n27023) );
  INAND2HSV0 U16817 ( .A1(\pe4/ti_7t [10]), .B1(n28812), .ZN(n15837) );
  INAND2HSV0 U16818 ( .A1(\pe3/ti_7t [9]), .B1(n16159), .ZN(n15964) );
  INOR2HSV0 U16819 ( .A1(\pe4/ti_7t [5]), .B1(n15484), .ZN(n15476) );
  INAND2HSV0 U16820 ( .A1(\pe9/ti_7t [9]), .B1(n18194), .ZN(n18276) );
  INAND2HSV0 U16821 ( .A1(\pe3/ti_7t [5]), .B1(n15238), .ZN(n15202) );
  INAND2HSV0 U16822 ( .A1(\pe1/ti_7t [13]), .B1(n22050), .ZN(n26827) );
  CLKNAND2HSV0 U16823 ( .A1(n11804), .A2(n20775), .ZN(n13877) );
  CLKNAND2HSV0 U16824 ( .A1(n23469), .A2(n13877), .ZN(n13878) );
  OAI211HSV0 U16825 ( .A1(n13877), .A2(n23469), .B(n13878), .C(n23470), .ZN(
        n13879) );
  CLKNAND2HSV0 U16826 ( .A1(n13879), .A2(poh11[5]), .ZN(n13880) );
  OAI21HSV0 U16827 ( .A1(poh11[5]), .A2(n13879), .B(n13880), .ZN(po[6]) );
  INAND2HSV0 U16828 ( .A1(\pe8/ti_7t [7]), .B1(n16504), .ZN(n18716) );
  XOR2HSV0 U16829 ( .A1(n23274), .A2(n23273), .Z(n13881) );
  CLKNAND2HSV0 U16830 ( .A1(n13882), .A2(n13881), .ZN(n13883) );
  OAI21HSV0 U16831 ( .A1(n13882), .A2(n13881), .B(n13883), .ZN(\pe5/poht [8])
         );
  OAI21HSV0 U16832 ( .A1(n23433), .A2(n27731), .B(n21714), .ZN(n13884) );
  AOI21HSV0 U16833 ( .A1(n28590), .A2(n23433), .B(n13884), .ZN(n13885) );
  CLKNAND2HSV0 U16834 ( .A1(n13886), .A2(n23435), .ZN(n13887) );
  OAI21HSV0 U16835 ( .A1(n23435), .A2(n13886), .B(n13887), .ZN(n13888) );
  OAI21HSV0 U16836 ( .A1(n13885), .A2(n23434), .B(n13888), .ZN(n13889) );
  OAI31HSV0 U16837 ( .A1(n13885), .A2(n13888), .A3(n23434), .B(n13889), .ZN(
        n28970) );
  IOA21HSV0 U16838 ( .A1(n23244), .A2(pov9[14]), .B(n23245), .ZN(
        \pe9/ti_7[14] ) );
  INOR2HSV0 U16839 ( .A1(\pe11/aot [1]), .B1(n25413), .ZN(n13890) );
  CLKNAND2HSV0 U16840 ( .A1(\pe11/got [1]), .A2(n24957), .ZN(n13891) );
  CLKNAND2HSV0 U16841 ( .A1(n13891), .A2(n13890), .ZN(n13892) );
  OAI21HSV0 U16842 ( .A1(n13890), .A2(n13891), .B(n13892), .ZN(\pe11/poht [15]) );
  CLKNAND2HSV0 U16843 ( .A1(n22328), .A2(n22329), .ZN(n13893) );
  CLKNAND2HSV0 U16844 ( .A1(n13895), .A2(n13894), .ZN(n13896) );
  OAI21HSV0 U16845 ( .A1(n13894), .A2(n13895), .B(n13896), .ZN(\pe8/poht [3])
         );
  INOR2HSV0 U16846 ( .A1(\pe7/aot [1]), .B1(n27095), .ZN(n13897) );
  CLKNAND2HSV0 U16847 ( .A1(n24277), .A2(\pe7/got [1]), .ZN(n13898) );
  CLKNAND2HSV0 U16848 ( .A1(n13898), .A2(n13897), .ZN(n13899) );
  OAI21HSV0 U16849 ( .A1(n13897), .A2(n13898), .B(n13899), .ZN(\pe7/poht [15])
         );
  XOR2HSV0 U16850 ( .A1(n25817), .A2(n25816), .Z(n13900) );
  CLKNAND2HSV0 U16851 ( .A1(n26084), .A2(\pe6/got [9]), .ZN(n13901) );
  CLKNAND2HSV0 U16852 ( .A1(n13901), .A2(n13900), .ZN(n13902) );
  OAI21HSV0 U16853 ( .A1(n13900), .A2(n13901), .B(n13902), .ZN(n13903) );
  CLKNAND2HSV0 U16854 ( .A1(\pe6/got [10]), .A2(n25784), .ZN(n13904) );
  CLKNAND2HSV0 U16855 ( .A1(n13904), .A2(n13903), .ZN(n13905) );
  OAI21HSV0 U16856 ( .A1(n13903), .A2(n13904), .B(n13905), .ZN(\pe6/poht [6])
         );
  CLKNHSV0 U16857 ( .I(n26309), .ZN(n13906) );
  MUX2NHSV0 U16858 ( .I0(n13906), .I1(n26309), .S(n23679), .ZN(n13907) );
  XOR2HSV0 U16859 ( .A1(n23680), .A2(n13907), .Z(n13908) );
  CLKNAND2HSV0 U16860 ( .A1(n24522), .A2(\pe3/got [2]), .ZN(n13909) );
  CLKNAND2HSV0 U16861 ( .A1(n13909), .A2(n13908), .ZN(n13910) );
  OAI21HSV0 U16862 ( .A1(n13908), .A2(n13909), .B(n13910), .ZN(n13911) );
  CLKNAND2HSV0 U16863 ( .A1(n26679), .A2(n26751), .ZN(n13912) );
  CLKNAND2HSV0 U16864 ( .A1(n13912), .A2(n13911), .ZN(n13913) );
  OAI21HSV0 U16865 ( .A1(n13911), .A2(n13912), .B(n13913), .ZN(\pe3/poht [13])
         );
  CLKNHSV0 U16866 ( .I(bo11[11]), .ZN(n13914) );
  MUX2NHSV0 U16867 ( .I0(n13914), .I1(n24314), .S(n27055), .ZN(n28728) );
  MUX2NHSV0 U16868 ( .I0(n13915), .I1(n22102), .S(n22103), .ZN(n13916) );
  XOR2HSV0 U16869 ( .A1(n13916), .A2(n22105), .Z(n28944) );
  NOR2HSV0 U16870 ( .A1(n23474), .A2(n23473), .ZN(n13917) );
  AOI211HSV0 U16871 ( .A1(n23474), .A2(n23473), .B(n22419), .C(n13917), .ZN(
        n13918) );
  NOR2HSV0 U16872 ( .A1(n13918), .A2(n23475), .ZN(n13919) );
  CLKNAND2HSV0 U16873 ( .A1(n13919), .A2(n23476), .ZN(n13920) );
  OAI21HSV0 U16874 ( .A1(n13919), .A2(n23476), .B(n13920), .ZN(n28982) );
  CLKNHSV0 U16875 ( .I(n25676), .ZN(n13921) );
  MUX2NHSV0 U16876 ( .I0(n13921), .I1(n25676), .S(n25677), .ZN(n13922) );
  CLKNAND2HSV0 U16877 ( .A1(n26220), .A2(n28585), .ZN(n13923) );
  CLKNAND2HSV0 U16878 ( .A1(n13923), .A2(n13922), .ZN(n13924) );
  OAI21HSV0 U16879 ( .A1(n13922), .A2(n13923), .B(n13924), .ZN(pov10[10]) );
  CLKNHSV0 U16880 ( .I(n23716), .ZN(n13925) );
  MUX2NHSV0 U16881 ( .I0(n23716), .I1(n13925), .S(n23715), .ZN(n28995) );
  CLKNHSV0 U16882 ( .I(bo10[1]), .ZN(n13926) );
  MUX2NHSV0 U16883 ( .I0(n13926), .I1(n26163), .S(n23510), .ZN(n28912) );
  CLKNHSV0 U16884 ( .I(bo9[11]), .ZN(n13927) );
  MUX2NHSV0 U16885 ( .I0(n13927), .I1(n23531), .S(n27093), .ZN(n28897) );
  CLKNHSV0 U16886 ( .I(n21320), .ZN(n13928) );
  MUX2NHSV0 U16887 ( .I0(n21320), .I1(n13928), .S(n21319), .ZN(n13929) );
  CLKNAND2HSV0 U16888 ( .A1(n28457), .A2(\pe8/got [16]), .ZN(n13930) );
  CLKNAND2HSV0 U16889 ( .A1(n13930), .A2(n13929), .ZN(n13931) );
  OAI21HSV0 U16890 ( .A1(n13929), .A2(n13930), .B(n13931), .ZN(n29005) );
  CLKNHSV0 U16891 ( .I(bo8[10]), .ZN(n13932) );
  MUX2NHSV0 U16892 ( .I0(n13932), .I1(n23723), .S(n23528), .ZN(n28887) );
  NAND3HSV0 U16893 ( .A1(n25346), .A2(n25345), .A3(n25344), .ZN(n13933) );
  XOR2HSV0 U16894 ( .A1(n25348), .A2(n13933), .Z(n28975) );
  CLKNHSV0 U16895 ( .I(bo7[5]), .ZN(n13934) );
  MUX2NHSV0 U16896 ( .I0(n13934), .I1(n27097), .S(n27099), .ZN(n28775) );
  CLKNHSV0 U16897 ( .I(n27212), .ZN(n13935) );
  CLKNHSV0 U16898 ( .I(n27210), .ZN(n13936) );
  MUX2NHSV0 U16899 ( .I0(n13936), .I1(n27210), .S(n27211), .ZN(n13937) );
  MUX2NHSV0 U16900 ( .I0(n27212), .I1(n13935), .S(n13937), .ZN(n28993) );
  CLKNAND2HSV0 U16901 ( .A1(n25849), .A2(n25647), .ZN(n13938) );
  CLKNAND2HSV0 U16902 ( .A1(n13938), .A2(n12068), .ZN(n13939) );
  OAI21HSV0 U16903 ( .A1(n25648), .A2(n13938), .B(n13939), .ZN(n28991) );
  CLKNAND2HSV0 U16904 ( .A1(n25764), .A2(n25058), .ZN(n13940) );
  CLKNAND2HSV0 U16905 ( .A1(n13940), .A2(n12297), .ZN(n13941) );
  OAI21HSV0 U16906 ( .A1(n12297), .A2(n13940), .B(n13941), .ZN(n29022) );
  CLKNAND2HSV0 U16907 ( .A1(n24305), .A2(bo6[6]), .ZN(n13942) );
  OAI21HSV0 U16908 ( .A1(n25706), .A2(n24305), .B(n13942), .ZN(n28749) );
  CLKNHSV0 U16909 ( .I(n25659), .ZN(n13943) );
  MUX2NHSV0 U16910 ( .I0(n25659), .I1(n13943), .S(n14613), .ZN(n13944) );
  CLKNAND2HSV0 U16911 ( .A1(n25656), .A2(n25657), .ZN(n13945) );
  CLKNAND2HSV0 U16912 ( .A1(n13945), .A2(n13944), .ZN(n13946) );
  OAI21HSV0 U16913 ( .A1(n13944), .A2(n13945), .B(n13946), .ZN(n29025) );
  CLKNAND2HSV0 U16914 ( .A1(n27051), .A2(bo5[7]), .ZN(n13947) );
  OAI21HSV0 U16915 ( .A1(n23504), .A2(n27051), .B(n13947), .ZN(n28863) );
  CLKNHSV0 U16916 ( .I(n27228), .ZN(n13948) );
  MUX2NHSV0 U16917 ( .I0(n27228), .I1(n13948), .S(n27229), .ZN(n29032) );
  CLKNAND2HSV0 U16918 ( .A1(n15813), .A2(n27957), .ZN(n13949) );
  CLKNAND2HSV0 U16919 ( .A1(n13949), .A2(n25663), .ZN(n13950) );
  OAI21HSV0 U16920 ( .A1(n13949), .A2(n25663), .B(n13950), .ZN(n29030) );
  CLKNAND2HSV0 U16921 ( .A1(n15176), .A2(n23480), .ZN(n13951) );
  CLKNAND2HSV0 U16922 ( .A1(n13951), .A2(n23481), .ZN(n13952) );
  OAI21HSV0 U16923 ( .A1(n23481), .A2(n13951), .B(n13952), .ZN(n29038) );
  CLKNHSV0 U16924 ( .I(bo3[11]), .ZN(n13953) );
  MUX2NHSV0 U16925 ( .I0(n13953), .I1(n24527), .S(n23518), .ZN(n28845) );
  CLKNHSV0 U16926 ( .I(\pe2/pq ), .ZN(n13954) );
  MUX2NHSV0 U16927 ( .I0(n13954), .I1(n17782), .S(n25623), .ZN(\pe2/ti_1t ) );
  CLKNHSV0 U16928 ( .I(bo2[2]), .ZN(n13955) );
  MUX2NHSV0 U16929 ( .I0(n13955), .I1(n27554), .S(n28835), .ZN(n28834) );
  CLKNHSV0 U16930 ( .I(bo1[1]), .ZN(n13956) );
  MUX2NHSV0 U16931 ( .I0(n13956), .I1(n27064), .S(n27065), .ZN(n28738) );
  BUFHSV8 U16932 ( .I(n19267), .Z(n19466) );
  INHSV4 U16933 ( .I(n19699), .ZN(n19695) );
  INHSV4 U16934 ( .I(n25494), .ZN(n25499) );
  INHSV6 U16935 ( .I(ctro10), .ZN(n16638) );
  BUFHSV6 U16936 ( .I(n16740), .Z(n16844) );
  INHSV4 U16937 ( .I(n20559), .ZN(n21785) );
  CLKNHSV6 U16938 ( .I(n20636), .ZN(n20770) );
  INHSV4 U16939 ( .I(n19141), .ZN(n19055) );
  INHSV8 U16940 ( .I(n18416), .ZN(n27093) );
  INHSV2 U16941 ( .I(n22995), .ZN(n26034) );
  INHSV4 U16942 ( .I(n26034), .ZN(n14029) );
  AND2HSV4 U16943 ( .A1(n22080), .A2(n22079), .Z(n27232) );
  INHSV4 U16944 ( .I(n27232), .ZN(n27657) );
  INHSV4 U16945 ( .I(n27232), .ZN(n27667) );
  CLKNHSV6 U16946 ( .I(n22490), .ZN(n28585) );
  INHSV4 U16947 ( .I(n22374), .ZN(n28437) );
  BUFHSV2 U16948 ( .I(n16331), .Z(n22125) );
  CLKNHSV0 U16949 ( .I(n18657), .ZN(n19830) );
  CLKNHSV6 U16950 ( .I(ctro5), .ZN(n14506) );
  BUFHSV8 U16951 ( .I(n14506), .Z(n21422) );
  INHSV4 U16952 ( .I(n23373), .ZN(n14054) );
  INHSV4 U16953 ( .I(n22373), .ZN(n28317) );
  INHSV4 U16954 ( .I(n22373), .ZN(n28231) );
  INHSV4 U16955 ( .I(n26418), .ZN(n26830) );
  INHSV4 U16956 ( .I(n15007), .ZN(n26380) );
  INHSV4 U16957 ( .I(n23459), .ZN(n28588) );
  CLKAND2HSV2 U16958 ( .A1(n17350), .A2(\pe1/got [15]), .Z(n13957) );
  BUFHSV4 U16959 ( .I(ctro4), .Z(n15534) );
  INHSV6 U16960 ( .I(\pe1/got [15]), .ZN(n26536) );
  INHSV4 U16961 ( .I(n20336), .ZN(n20157) );
  INHSV4 U16962 ( .I(n15919), .ZN(n16112) );
  INHSV2 U16963 ( .I(\pe1/got [13]), .ZN(n17364) );
  INHSV4 U16964 ( .I(n24685), .ZN(n14071) );
  INHSV2 U16965 ( .I(n18330), .ZN(n18194) );
  INHSV4 U16966 ( .I(n18628), .ZN(n18330) );
  INHSV4 U16967 ( .I(n15963), .ZN(n16163) );
  INHSV2 U16968 ( .I(n21313), .ZN(n23382) );
  INHSV2 U16969 ( .I(n21159), .ZN(n17652) );
  INHSV6 U16970 ( .I(n23508), .ZN(n21332) );
  INHSV4 U16971 ( .I(n18325), .ZN(n18462) );
  INHSV4 U16972 ( .I(n18325), .ZN(n18628) );
  INHSV4 U16973 ( .I(n19267), .ZN(n19674) );
  BUFHSV4 U16974 ( .I(\pe2/got [15]), .Z(n17862) );
  INHSV4 U16975 ( .I(n17862), .ZN(n17773) );
  INHSV4 U16976 ( .I(n17862), .ZN(n17863) );
  BUFHSV4 U16977 ( .I(n20551), .Z(n20698) );
  INHSV4 U16978 ( .I(n14559), .ZN(n14497) );
  INHSV2 U16979 ( .I(n14559), .ZN(n14482) );
  INHSV4 U16980 ( .I(n16948), .ZN(n17120) );
  INHSV4 U16981 ( .I(n21880), .ZN(n17767) );
  INHSV4 U16982 ( .I(n21164), .ZN(n21144) );
  INHSV4 U16983 ( .I(n28667), .ZN(n25523) );
  INHSV4 U16984 ( .I(n16304), .ZN(n16307) );
  INHSV4 U16985 ( .I(n16554), .ZN(n19969) );
  BUFHSV4 U16986 ( .I(n15534), .Z(n15693) );
  CLKNHSV0 U16987 ( .I(n23798), .ZN(n28606) );
  CLKNHSV0 U16988 ( .I(n23793), .ZN(n28607) );
  CLKNHSV0 U16989 ( .I(n23793), .ZN(n28604) );
  INHSV6 U16990 ( .I(n14535), .ZN(n20977) );
  INHSV8 U16991 ( .I(\pe5/bq[12] ), .ZN(n14766) );
  INHSV2 U16992 ( .I(n27190), .ZN(n14631) );
  INHSV4 U16993 ( .I(n20074), .ZN(n26096) );
  INHSV2 U16994 ( .I(\pe7/got [8]), .ZN(n19479) );
  INHSV2 U16995 ( .I(\pe7/got [6]), .ZN(n19532) );
  INHSV4 U16996 ( .I(n17038), .ZN(n16973) );
  BUFHSV4 U16997 ( .I(n16740), .Z(n16998) );
  INHSV4 U16998 ( .I(n21422), .ZN(n20870) );
  INHSV4 U16999 ( .I(n21422), .ZN(n21412) );
  INHSV2 U17000 ( .I(\pe6/got [7]), .ZN(n14418) );
  INHSV4 U17001 ( .I(n21117), .ZN(n27231) );
  INHSV2 U17002 ( .I(\pe11/bq[12] ), .ZN(n20267) );
  CLKAND2HSV2 U17003 ( .A1(n22129), .A2(n16393), .Z(n13958) );
  CLKNHSV0 U17004 ( .I(\pe5/bq[3] ), .ZN(n21572) );
  INHSV4 U17005 ( .I(\pe11/phq [2]), .ZN(n20165) );
  INHSV6 U17006 ( .I(\pe1/aot [15]), .ZN(n17374) );
  INHSV6 U17007 ( .I(n14979), .ZN(n26431) );
  INHSV4 U17008 ( .I(n16809), .ZN(n17084) );
  INHSV6 U17009 ( .I(n16312), .ZN(n16511) );
  INHSV6 U17010 ( .I(\pe8/ti_1 ), .ZN(n16312) );
  INHSV4 U17011 ( .I(n25057), .ZN(n23041) );
  INHSV4 U17012 ( .I(\pe4/got [11]), .ZN(n27871) );
  INHSV2 U17013 ( .I(\pe11/bq[10] ), .ZN(n20384) );
  INHSV4 U17014 ( .I(n15176), .ZN(n16031) );
  INHSV4 U17015 ( .I(n23477), .ZN(n28621) );
  INHSV4 U17016 ( .I(n20568), .ZN(n20506) );
  INHSV6 U17017 ( .I(n17973), .ZN(n21761) );
  INHSV6 U17018 ( .I(n17781), .ZN(n27543) );
  INHSV2 U17019 ( .I(\pe2/got [7]), .ZN(n27686) );
  INHSV4 U17020 ( .I(\pe5/got [13]), .ZN(n14544) );
  INHSV4 U17021 ( .I(n20869), .ZN(n14852) );
  INHSV4 U17022 ( .I(n14544), .ZN(n14503) );
  INHSV6 U17023 ( .I(n24128), .ZN(n14022) );
  INHSV4 U17024 ( .I(n16554), .ZN(n16504) );
  INHSV4 U17025 ( .I(n17651), .ZN(n21234) );
  INHSV4 U17026 ( .I(n17651), .ZN(n28693) );
  BUFHSV4 U17027 ( .I(n14506), .Z(n14815) );
  BUFHSV4 U17028 ( .I(n22931), .Z(n22825) );
  INHSV4 U17029 ( .I(n15393), .ZN(n26919) );
  INHSV4 U17030 ( .I(n25027), .ZN(n20227) );
  INHSV4 U17031 ( .I(n26536), .ZN(n14056) );
  INHSV4 U17032 ( .I(n26536), .ZN(n17230) );
  CLKNHSV0 U17033 ( .I(\pe2/aot [2]), .ZN(n27250) );
  INHSV4 U17034 ( .I(n20370), .ZN(n20565) );
  INHSV4 U17035 ( .I(n15189), .ZN(n16164) );
  INHSV2 U17036 ( .I(n21722), .ZN(n16015) );
  INHSV4 U17037 ( .I(\pe10/got [13]), .ZN(n16729) );
  INHSV6 U17038 ( .I(n16729), .ZN(n28479) );
  INHSV6 U17039 ( .I(n27140), .ZN(n28434) );
  INHSV2 U17040 ( .I(\pe4/got [12]), .ZN(n15614) );
  INHSV4 U17041 ( .I(n15614), .ZN(n28428) );
  INHSV4 U17042 ( .I(n22822), .ZN(n25128) );
  INHSV6 U17043 ( .I(\pe7/got [15]), .ZN(n19279) );
  BUFHSV4 U17044 ( .I(\pe7/got [15]), .Z(n19212) );
  INHSV4 U17045 ( .I(n19212), .ZN(n19512) );
  INHSV2 U17046 ( .I(n19526), .ZN(n25339) );
  CLKNHSV6 U17047 ( .I(ctro2), .ZN(n17808) );
  INHSV4 U17048 ( .I(n21901), .ZN(n21641) );
  INHSV6 U17049 ( .I(n15835), .ZN(n15813) );
  INHSV4 U17050 ( .I(n22895), .ZN(n15621) );
  INHSV4 U17051 ( .I(n25052), .ZN(n25504) );
  BUFHSV6 U17052 ( .I(n14815), .Z(n14628) );
  INHSV2 U17053 ( .I(\pe4/got [5]), .ZN(n21997) );
  CLKNHSV0 U17054 ( .I(\pe3/got [11]), .ZN(n26296) );
  INHSV4 U17055 ( .I(n15702), .ZN(n22918) );
  INHSV4 U17056 ( .I(n22137), .ZN(n18773) );
  INHSV4 U17057 ( .I(n26852), .ZN(n28435) );
  BUFHSV4 U17058 ( .I(n19267), .Z(n19765) );
  INHSV6 U17059 ( .I(n22637), .ZN(n26132) );
  INHSV4 U17060 ( .I(n23244), .ZN(n18641) );
  INHSV6 U17061 ( .I(n18855), .ZN(n14236) );
  INHSV2 U17062 ( .I(\pe5/got [2]), .ZN(n23260) );
  BUFHSV2 U17063 ( .I(n18050), .Z(n23244) );
  INHSV4 U17064 ( .I(\pe2/got [1]), .ZN(n27677) );
  INHSV4 U17065 ( .I(\pe3/got [8]), .ZN(n26601) );
  INHSV2 U17066 ( .I(\pe5/got [3]), .ZN(n24364) );
  BUFHSV2 U17067 ( .I(n15973), .Z(n15333) );
  INHSV4 U17068 ( .I(n20698), .ZN(n20637) );
  INHSV4 U17069 ( .I(n20551), .ZN(n20302) );
  INHSV4 U17070 ( .I(n16331), .ZN(n18657) );
  INHSV2 U17071 ( .I(n16166), .ZN(n15017) );
  CLKNHSV0 U17072 ( .I(\pe10/got [12]), .ZN(n23548) );
  BUFHSV4 U17073 ( .I(\pe10/got [12]), .Z(n16876) );
  BUFHSV8 U17074 ( .I(\pe9/got [1]), .Z(n28658) );
  INHSV2 U17075 ( .I(\pe9/got [1]), .ZN(n28303) );
  OR2HSV1 U17076 ( .A1(n19824), .A2(n25602), .Z(n13959) );
  INHSV4 U17077 ( .I(n21332), .ZN(n27089) );
  BUFHSV4 U17078 ( .I(n20551), .Z(n24889) );
  INHSV2 U17079 ( .I(n22125), .ZN(n18767) );
  CLKNHSV0 U17080 ( .I(n23798), .ZN(n28595) );
  CLKNHSV0 U17081 ( .I(\pe8/got [6]), .ZN(n22142) );
  BUFHSV4 U17082 ( .I(n15060), .Z(n15973) );
  INHSV2 U17083 ( .I(n18788), .ZN(n18787) );
  INHSV4 U17084 ( .I(n14911), .ZN(n21523) );
  BUFHSV4 U17085 ( .I(n23528), .Z(n23519) );
  INHSV4 U17086 ( .I(n14642), .ZN(n14630) );
  INHSV4 U17087 ( .I(n22378), .ZN(n23822) );
  INHSV4 U17088 ( .I(n14303), .ZN(n19045) );
  INHSV4 U17089 ( .I(n18927), .ZN(n18992) );
  INHSV2 U17090 ( .I(n21312), .ZN(n16172) );
  AND2HSV2 U17091 ( .A1(\pe7/got [4]), .A2(n25408), .Z(n13960) );
  NOR2HSV2 U17092 ( .A1(n14578), .A2(n14517), .ZN(n14472) );
  INHSV2 U17093 ( .I(n14472), .ZN(n14473) );
  CLKAND2HSV2 U17094 ( .A1(n22134), .A2(n23422), .Z(n13961) );
  CLKNHSV0 U17095 ( .I(n14549), .ZN(n14572) );
  INHSV4 U17096 ( .I(n21713), .ZN(n21235) );
  INHSV2 U17097 ( .I(n21007), .ZN(n17813) );
  CLKAND2HSV2 U17098 ( .A1(n14736), .A2(n14396), .Z(n13964) );
  CLKXOR2HSV4 U17099 ( .A1(n15329), .A2(n15328), .Z(n13965) );
  INHSV4 U17100 ( .I(n19160), .ZN(n19073) );
  XNOR2HSV1 U17101 ( .A1(n22874), .A2(n22873), .ZN(n13966) );
  CLKNAND2HSV2 U17102 ( .A1(n18613), .A2(\pe9/ti_7t [1]), .ZN(n17945) );
  CLKNHSV0 U17103 ( .I(n19975), .ZN(n19981) );
  NOR2HSV2 U17104 ( .A1(n14629), .A2(n14614), .ZN(n13967) );
  INHSV2 U17105 ( .I(n21977), .ZN(n22800) );
  INHSV4 U17106 ( .I(n18050), .ZN(n18650) );
  INHSV4 U17107 ( .I(n23115), .ZN(n23116) );
  CLKAND2HSV2 U17108 ( .A1(n17236), .A2(n17230), .Z(n13971) );
  INHSV6 U17109 ( .I(\pe4/bq[16] ), .ZN(n15363) );
  INHSV6 U17110 ( .I(n15416), .ZN(n15428) );
  XNOR3HSV2 U17111 ( .A1(n15445), .A2(n15444), .A3(n15443), .ZN(n13973) );
  XNOR3HSV2 U17112 ( .A1(n22678), .A2(n22677), .A3(n22676), .ZN(n13974) );
  CLKNHSV0 U17113 ( .I(\pe6/bq[8] ), .ZN(n24307) );
  CLKAND2HSV2 U17114 ( .A1(n14238), .A2(n14239), .Z(n13975) );
  INHSV2 U17115 ( .I(n23137), .ZN(n25292) );
  INHSV4 U17116 ( .I(n15140), .ZN(n23480) );
  INHSV4 U17117 ( .I(n15223), .ZN(n26255) );
  INHSV4 U17118 ( .I(n17374), .ZN(n28468) );
  AO21HSV1 U17119 ( .A1(n20292), .A2(n28918), .B(n20837), .Z(n13976) );
  INHSV4 U17120 ( .I(n21254), .ZN(n17785) );
  CLKNHSV0 U17121 ( .I(\pe7/got [7]), .ZN(n25373) );
  CLKNHSV0 U17122 ( .I(n21066), .ZN(n17830) );
  BUFHSV4 U17123 ( .I(n21066), .Z(n21260) );
  INHSV2 U17124 ( .I(n15284), .ZN(n15194) );
  INHSV6 U17125 ( .I(\pe11/ctrq ), .ZN(n20164) );
  CLKNAND2HSV2 U17126 ( .A1(n16159), .A2(\pe3/ti_7t [1]), .ZN(n13977) );
  CLKAND2HSV4 U17127 ( .A1(n15629), .A2(n15626), .Z(n13979) );
  INHSV6 U17128 ( .I(\pe4/ctrq ), .ZN(n15502) );
  INHSV4 U17129 ( .I(\pe10/ctrq ), .ZN(n16976) );
  INHSV2 U17130 ( .I(n22086), .ZN(n21154) );
  BUFHSV4 U17131 ( .I(n22086), .Z(n21150) );
  CLKNHSV0 U17132 ( .I(n15628), .ZN(n15632) );
  BUFHSV4 U17133 ( .I(\pe3/got [14]), .Z(n28930) );
  CLKNHSV0 U17134 ( .I(n18774), .ZN(n19952) );
  CLKNAND2HSV4 U17135 ( .A1(n18705), .A2(n18704), .ZN(n18774) );
  INHSV2 U17136 ( .I(\pe5/got [9]), .ZN(n24685) );
  INHSV6 U17137 ( .I(n19357), .ZN(n24271) );
  CLKNHSV0 U17138 ( .I(\pe2/got [12]), .ZN(n17792) );
  BUFHSV4 U17139 ( .I(\pe6/got [11]), .Z(n28586) );
  INHSV2 U17140 ( .I(n22994), .ZN(n14086) );
  INHSV4 U17141 ( .I(n26417), .ZN(n28425) );
  INHSV6 U17142 ( .I(n14547), .ZN(n24635) );
  CLKNHSV0 U17143 ( .I(\pe8/got [5]), .ZN(n22283) );
  CLKNHSV0 U17144 ( .I(\pe6/got [8]), .ZN(n26032) );
  CLKNHSV0 U17145 ( .I(\pe6/got [9]), .ZN(n25698) );
  INHSV4 U17146 ( .I(\pe7/bq[4] ), .ZN(n19649) );
  BUFHSV4 U17147 ( .I(n15534), .Z(n15627) );
  BUFHSV4 U17148 ( .I(n15752), .Z(n27976) );
  INHSV4 U17149 ( .I(n16998), .ZN(n20148) );
  INHSV2 U17150 ( .I(n16708), .ZN(n20142) );
  INHSV2 U17151 ( .I(n16740), .ZN(n16669) );
  INHSV2 U17152 ( .I(\pe3/bq[4] ), .ZN(n23349) );
  BUFHSV4 U17153 ( .I(n14815), .Z(n20848) );
  INHSV4 U17154 ( .I(n24313), .ZN(n28628) );
  INHSV6 U17155 ( .I(\pe3/got [13]), .ZN(n24313) );
  INHSV4 U17156 ( .I(n19972), .ZN(n16311) );
  INHSV2 U17157 ( .I(n18001), .ZN(n28669) );
  CLKNHSV6 U17158 ( .I(n18308), .ZN(n28423) );
  INHSV6 U17159 ( .I(n18691), .ZN(n22136) );
  INHSV4 U17160 ( .I(n19905), .ZN(n23653) );
  INHSV6 U17161 ( .I(\pe10/got [11]), .ZN(n22636) );
  INHSV2 U17162 ( .I(\pe4/got [8]), .ZN(n27827) );
  BUFHSV4 U17163 ( .I(n23372), .Z(n21722) );
  INHSV6 U17164 ( .I(\pe7/got [13]), .ZN(n19242) );
  INHSV4 U17165 ( .I(\pe9/got [9]), .ZN(n28067) );
  INHSV6 U17166 ( .I(n28067), .ZN(n14073) );
  INHSV6 U17167 ( .I(\pe2/got [11]), .ZN(n17781) );
  CLKNHSV0 U17168 ( .I(\pe2/got [15]), .ZN(n21225) );
  INHSV6 U17169 ( .I(n17773), .ZN(n22085) );
  INHSV6 U17170 ( .I(\pe9/got [10]), .ZN(n22116) );
  BUFHSV4 U17171 ( .I(n18325), .Z(n18219) );
  INHSV6 U17172 ( .I(n19264), .ZN(n28610) );
  OA21HSV2 U17173 ( .A1(n14698), .A2(\pe6/ti_7t [5]), .B(n25058), .Z(n13980)
         );
  INHSV4 U17174 ( .I(\pe5/got [11]), .ZN(n14535) );
  INHSV2 U17175 ( .I(\pe8/got [2]), .ZN(n28650) );
  OA21HSV2 U17176 ( .A1(n15487), .A2(\pe4/ti_7t [5]), .B(n15813), .Z(n13981)
         );
  INHSV2 U17177 ( .I(\pe6/got [2]), .ZN(n28651) );
  INHSV2 U17178 ( .I(n20215), .ZN(n20623) );
  INHSV4 U17179 ( .I(n23402), .ZN(n26240) );
  INHSV4 U17180 ( .I(\pe1/got [6]), .ZN(n27140) );
  INHSV4 U17181 ( .I(\pe10/got [4]), .ZN(n22637) );
  INHSV4 U17182 ( .I(n17773), .ZN(n17774) );
  CLKNHSV0 U17183 ( .I(n28802), .ZN(n17214) );
  AND2HSV2 U17184 ( .A1(n15491), .A2(n15813), .Z(n13982) );
  INHSV2 U17185 ( .I(\pe4/ti_7t [3]), .ZN(n15423) );
  CLKNHSV0 U17186 ( .I(\pe5/bq[1] ), .ZN(n24326) );
  INHSV4 U17187 ( .I(n17533), .ZN(n26595) );
  BUFHSV4 U17188 ( .I(n18325), .Z(n18543) );
  INHSV6 U17189 ( .I(\pe10/got [2]), .ZN(n27194) );
  CLKNHSV0 U17190 ( .I(\pe7/got [5]), .ZN(n23191) );
  INHSV4 U17191 ( .I(n21554), .ZN(n24686) );
  BUFHSV4 U17192 ( .I(n21813), .Z(n27354) );
  INHSV4 U17193 ( .I(\pe2/got [6]), .ZN(n27498) );
  INHSV2 U17194 ( .I(n27498), .ZN(n14006) );
  INHSV4 U17195 ( .I(\pe5/got [4]), .ZN(n24414) );
  INHSV2 U17196 ( .I(n24414), .ZN(n13999) );
  INHSV4 U17197 ( .I(\pe4/got [7]), .ZN(n27969) );
  INHSV2 U17198 ( .I(n27969), .ZN(n14000) );
  INHSV2 U17199 ( .I(n26416), .ZN(n27002) );
  INHSV2 U17200 ( .I(n25079), .ZN(n28001) );
  INHSV4 U17201 ( .I(n27194), .ZN(n14065) );
  INHSV4 U17202 ( .I(n27194), .ZN(n28637) );
  INHSV4 U17203 ( .I(\pe6/got [5]), .ZN(n26014) );
  INHSV4 U17204 ( .I(n24311), .ZN(n28612) );
  INHSV4 U17205 ( .I(n17359), .ZN(n28802) );
  INHSV4 U17206 ( .I(n22117), .ZN(n22826) );
  BUFHSV4 U17207 ( .I(n14303), .Z(n14698) );
  INHSV4 U17208 ( .I(n11851), .ZN(n20372) );
  INHSV2 U17209 ( .I(n14506), .ZN(n21003) );
  INHSV4 U17210 ( .I(n28929), .ZN(n26413) );
  INHSV4 U17211 ( .I(n16031), .ZN(n15242) );
  INHSV4 U17212 ( .I(n28929), .ZN(n15176) );
  INHSV4 U17213 ( .I(\pe8/got [4]), .ZN(n22230) );
  INHSV2 U17214 ( .I(n19045), .ZN(n19127) );
  INHSV4 U17215 ( .I(n19820), .ZN(n19940) );
  BUFHSV4 U17216 ( .I(n19940), .Z(n25602) );
  INHSV2 U17217 ( .I(n15900), .ZN(n21968) );
  INHSV4 U17218 ( .I(n15693), .ZN(n15531) );
  INHSV4 U17219 ( .I(n21117), .ZN(n28429) );
  INHSV4 U17220 ( .I(n18029), .ZN(n18469) );
  AO21HSV1 U17221 ( .A1(n25696), .A2(n19151), .B(n19056), .Z(n13983) );
  INHSV4 U17222 ( .I(n19695), .ZN(n19623) );
  AO21HSV1 U17223 ( .A1(n18630), .A2(n18646), .B(n23448), .Z(n13984) );
  INHSV4 U17224 ( .I(n23986), .ZN(n28624) );
  INHSV4 U17225 ( .I(\pe3/got [5]), .ZN(n23329) );
  INHSV4 U17226 ( .I(n22848), .ZN(n28591) );
  NOR2HSV2 U17227 ( .A1(n18997), .A2(n14745), .ZN(n13985) );
  CLKAND2HSV2 U17228 ( .A1(n19707), .A2(n19702), .Z(n13986) );
  BUFHSV2 U17229 ( .I(n18915), .Z(n18927) );
  CLKNHSV0 U17230 ( .I(n18558), .ZN(n18524) );
  NAND2HSV0 U17231 ( .A1(n19830), .A2(n19835), .ZN(n13987) );
  INHSV2 U17232 ( .I(n22801), .ZN(n26923) );
  INHSV4 U17233 ( .I(n19808), .ZN(n18463) );
  CLKNHSV0 U17234 ( .I(n18538), .ZN(n18539) );
  INHSV4 U17235 ( .I(n14925), .ZN(n14926) );
  BUFHSV4 U17236 ( .I(n22111), .Z(n23499) );
  BUFHSV4 U17237 ( .I(n20470), .Z(n20650) );
  INHSV4 U17238 ( .I(n17819), .ZN(n21701) );
  INHSV4 U17239 ( .I(n22069), .ZN(n25678) );
  INHSV2 U17240 ( .I(n16284), .ZN(n28422) );
  INHSV4 U17241 ( .I(n22069), .ZN(n17598) );
  INHSV2 U17242 ( .I(n23372), .ZN(n16054) );
  BUFHSV4 U17243 ( .I(n28639), .Z(n27055) );
  BUFHSV4 U17244 ( .I(n28639), .Z(n22111) );
  BUFHSV4 U17245 ( .I(n23541), .Z(n23543) );
  BUFHSV4 U17246 ( .I(n23516), .Z(n23517) );
  BUFHSV4 U17247 ( .I(n23516), .Z(n23518) );
  BUFHSV4 U17248 ( .I(n23524), .Z(n23520) );
  BUFHSV4 U17249 ( .I(n21335), .Z(n23524) );
  BUFHSV4 U17250 ( .I(n28876), .Z(n27102) );
  INHSV2 U17251 ( .I(n14972), .ZN(n22069) );
  INHSV4 U17252 ( .I(\pe9/got [2]), .ZN(n28286) );
  INHSV4 U17253 ( .I(n28286), .ZN(n28654) );
  CLKNHSV0 U17254 ( .I(n24884), .ZN(n20768) );
  INHSV6 U17255 ( .I(n25932), .ZN(n14008) );
  INHSV4 U17256 ( .I(\pe9/got [12]), .ZN(n28016) );
  OR2HSV1 U17257 ( .A1(n22913), .A2(n21968), .Z(n13991) );
  INHSV4 U17258 ( .I(n16569), .ZN(n25532) );
  INHSV6 U17259 ( .I(\pe1/ctrq ), .ZN(n24316) );
  INHSV2 U17260 ( .I(\pe3/bq[13] ), .ZN(n26246) );
  INHSV2 U17261 ( .I(\pe1/bq[5] ), .ZN(n26659) );
  CLKNHSV0 U17262 ( .I(\pe4/bq[2] ), .ZN(n27088) );
  INHSV4 U17263 ( .I(\pe4/got [10]), .ZN(n27825) );
  INHSV4 U17264 ( .I(\pe2/got [3]), .ZN(n27633) );
  INHSV6 U17265 ( .I(\pe6/got [13]), .ZN(n18855) );
  INHSV4 U17266 ( .I(\pe5/got [13]), .ZN(n20869) );
  INHSV2 U17267 ( .I(\pe7/got [12]), .ZN(n24321) );
  INHSV2 U17268 ( .I(n16312), .ZN(n25624) );
  INHSV2 U17269 ( .I(n25624), .ZN(n25531) );
  CLKNHSV0 U17270 ( .I(\pe9/aot [16]), .ZN(n23546) );
  CLKNHSV0 U17271 ( .I(n23799), .ZN(n28601) );
  CLKNHSV0 U17272 ( .I(\pe7/got [16]), .ZN(n27134) );
  INHSV4 U17273 ( .I(n14676), .ZN(n14478) );
  CLKNHSV0 U17274 ( .I(n17668), .ZN(n21702) );
  INHSV2 U17275 ( .I(n16876), .ZN(n26091) );
  INHSV4 U17276 ( .I(n23548), .ZN(n26212) );
  NOR2HSV2 U17277 ( .A1(n26091), .A2(n22419), .ZN(n17006) );
  NOR2HSV2 U17278 ( .A1(n17023), .A2(n26091), .ZN(n16782) );
  INHSV4 U17279 ( .I(n24414), .ZN(n13993) );
  INHSV4 U17280 ( .I(n27871), .ZN(n13994) );
  CLKNHSV0 U17281 ( .I(n16795), .ZN(n13995) );
  CLKNHSV0 U17282 ( .I(\pe10/got [15]), .ZN(n16795) );
  CLKNHSV0 U17283 ( .I(n16795), .ZN(n22508) );
  NAND2HSV0 U17284 ( .A1(n28480), .A2(n13996), .ZN(n27936) );
  INHSV4 U17285 ( .I(n27969), .ZN(n13996) );
  INHSV4 U17286 ( .I(\pe2/ti_1 ), .ZN(n17782) );
  INHSV2 U17287 ( .I(n20051), .ZN(n13997) );
  INHSV4 U17288 ( .I(n13997), .ZN(n13998) );
  CLKNHSV0 U17289 ( .I(n20058), .ZN(n20051) );
  NAND2HSV0 U17290 ( .A1(n24674), .A2(n24637), .ZN(n14898) );
  INHSV6 U17291 ( .I(n16393), .ZN(n20058) );
  CLKNHSV0 U17292 ( .I(n27686), .ZN(n14046) );
  INHSV2 U17293 ( .I(n16976), .ZN(n14001) );
  INHSV4 U17294 ( .I(n27498), .ZN(n14003) );
  NAND2HSV0 U17295 ( .A1(n27784), .A2(n13994), .ZN(n22824) );
  NAND2HSV0 U17296 ( .A1(n15853), .A2(n13994), .ZN(n15888) );
  CLKNHSV0 U17297 ( .I(n24316), .ZN(n14004) );
  CLKNHSV0 U17298 ( .I(n24316), .ZN(n14005) );
  NAND2HSV0 U17299 ( .A1(n23327), .A2(n11891), .ZN(n16156) );
  NAND2HSV0 U17300 ( .A1(n27106), .A2(n13993), .ZN(n24339) );
  NAND2HSV0 U17301 ( .A1(n12517), .A2(n13993), .ZN(n24449) );
  NAND2HSV0 U17302 ( .A1(n28803), .A2(n13993), .ZN(n23267) );
  NAND2HSV0 U17303 ( .A1(n28699), .A2(\pe6/got [13]), .ZN(n23053) );
  NAND2HSV0 U17304 ( .A1(n19121), .A2(n14236), .ZN(n19039) );
  CLKNHSV0 U17305 ( .I(n23339), .ZN(n26751) );
  NAND2HSV0 U17306 ( .A1(n28803), .A2(n24637), .ZN(n24427) );
  CLKNHSV0 U17307 ( .I(n17230), .ZN(n14007) );
  NAND2HSV0 U17308 ( .A1(n28803), .A2(n28647), .ZN(n24370) );
  NAND2HSV0 U17309 ( .A1(n26082), .A2(n14008), .ZN(n24007) );
  NAND2HSV0 U17310 ( .A1(n28699), .A2(\pe6/got [3]), .ZN(n21779) );
  NAND2HSV0 U17311 ( .A1(n26031), .A2(n14008), .ZN(n19170) );
  NAND2HSV0 U17312 ( .A1(n25767), .A2(n14008), .ZN(n25768) );
  NAND2HSV0 U17313 ( .A1(\pe6/bq[13] ), .A2(\pe6/aot [10]), .ZN(n25835) );
  NAND2HSV0 U17314 ( .A1(n25950), .A2(\pe6/got [4]), .ZN(n21781) );
  NAND2HSV0 U17315 ( .A1(n28699), .A2(\pe6/got [4]), .ZN(n19172) );
  INHSV6 U17316 ( .I(\pe6/got [3]), .ZN(n25932) );
  CLKNHSV0 U17317 ( .I(\pe10/bq[7] ), .ZN(n14009) );
  CLKNHSV0 U17318 ( .I(n14009), .ZN(n14010) );
  CLKNHSV0 U17319 ( .I(\pe6/bq[9] ), .ZN(n14011) );
  CLKNHSV0 U17320 ( .I(n14011), .ZN(n14012) );
  CLKNHSV0 U17321 ( .I(\pe2/bq[13] ), .ZN(n14013) );
  CLKNHSV0 U17322 ( .I(n14013), .ZN(n14014) );
  CLKNHSV0 U17323 ( .I(\pe2/bq[12] ), .ZN(n14015) );
  CLKNHSV0 U17324 ( .I(n14015), .ZN(n14016) );
  CLKNHSV0 U17325 ( .I(\pe2/bq[10] ), .ZN(n14017) );
  CLKNHSV0 U17326 ( .I(n14017), .ZN(n14018) );
  CLKNHSV0 U17327 ( .I(n14956), .ZN(n14019) );
  NAND2HSV0 U17328 ( .A1(\pe2/bq[13] ), .A2(\pe2/aot [16]), .ZN(n17724) );
  INHSV2 U17329 ( .I(n21128), .ZN(n14020) );
  CLKNHSV0 U17330 ( .I(n28537), .ZN(n28921) );
  CLKNHSV0 U17331 ( .I(n28921), .ZN(n14021) );
  INHSV4 U17332 ( .I(\pe7/got [11]), .ZN(n24128) );
  NAND2HSV0 U17333 ( .A1(\pe6/bq[16] ), .A2(\pe6/aot [10]), .ZN(n14311) );
  CLKNHSV0 U17334 ( .I(n28921), .ZN(n14023) );
  INHSV2 U17335 ( .I(n24316), .ZN(n14024) );
  CLKNHSV0 U17336 ( .I(\pe3/bq[14] ), .ZN(n14025) );
  INHSV2 U17337 ( .I(n14025), .ZN(n14026) );
  NAND2HSV2 U17338 ( .A1(\pe6/bq[12] ), .A2(\pe6/aot [14]), .ZN(n14308) );
  NAND2HSV2 U17339 ( .A1(\pe3/bq[14] ), .A2(\pe3/aot [16]), .ZN(n15161) );
  CLKNHSV0 U17340 ( .I(\pe6/bq[16] ), .ZN(n14027) );
  INHSV2 U17341 ( .I(n14027), .ZN(n14028) );
  NAND2HSV0 U17342 ( .A1(n25060), .A2(n26218), .ZN(n26219) );
  CLKNAND2HSV2 U17343 ( .A1(n22432), .A2(n26218), .ZN(n20137) );
  NAND2HSV0 U17344 ( .A1(n21632), .A2(n21696), .ZN(n21633) );
  NAND3HSV2 U17345 ( .A1(\pe2/phq [2]), .A2(\pe2/ti_1 ), .A3(\pe2/got [15]), 
        .ZN(n17626) );
  INHSV2 U17346 ( .I(\pe2/got [15]), .ZN(n17668) );
  OAI21HSV0 U17347 ( .A1(n21737), .A2(n25261), .B(n17123), .ZN(n17125) );
  NAND2HSV0 U17348 ( .A1(n28480), .A2(\pe4/got [10]), .ZN(n27779) );
  NAND2HSV0 U17349 ( .A1(\pe4/ti_7[7] ), .A2(\pe4/got [10]), .ZN(n22038) );
  NAND2HSV4 U17350 ( .A1(n19698), .A2(n23112), .ZN(n28926) );
  INHSV4 U17351 ( .I(n28687), .ZN(n14031) );
  INHSV2 U17352 ( .I(n14032), .ZN(n14033) );
  OAI21HSV2 U17353 ( .A1(n15843), .A2(n15842), .B(n15841), .ZN(n21980) );
  OAI21HSV2 U17354 ( .A1(n21993), .A2(n15842), .B(n15751), .ZN(n25666) );
  AND2HSV4 U17355 ( .A1(n16040), .A2(n23414), .Z(n16045) );
  CLKNHSV0 U17356 ( .I(n28929), .ZN(n23414) );
  INHSV4 U17357 ( .I(n16308), .ZN(n16358) );
  CLKNHSV0 U17358 ( .I(\pe6/got [14]), .ZN(n14361) );
  CLKNHSV0 U17359 ( .I(\pe2/got [7]), .ZN(n27572) );
  CLKNHSV0 U17360 ( .I(n16430), .ZN(n14034) );
  CLKNHSV0 U17361 ( .I(n16430), .ZN(n25649) );
  NAND3HSV2 U17362 ( .A1(n19569), .A2(n19565), .A3(n27133), .ZN(n19610) );
  NAND2HSV4 U17363 ( .A1(n19459), .A2(n22089), .ZN(n19565) );
  BUFHSV4 U17364 ( .I(n23513), .Z(n14035) );
  BUFHSV4 U17365 ( .I(n23536), .Z(n23513) );
  CLKNHSV0 U17366 ( .I(n20690), .ZN(n20687) );
  OAI22HSV2 U17367 ( .A1(n20611), .A2(n20556), .B1(n20690), .B2(n20372), .ZN(
        n20557) );
  INHSV2 U17368 ( .I(n28623), .ZN(n14036) );
  NAND2HSV0 U17369 ( .A1(n26229), .A2(\pe8/got [8]), .ZN(n25213) );
  NAND2HSV0 U17370 ( .A1(n26229), .A2(\pe8/got [2]), .ZN(n26237) );
  BUFHSV8 U17371 ( .I(\pe6/got [1]), .Z(n28608) );
  INHSV2 U17372 ( .I(n28523), .ZN(n14037) );
  CLKNHSV6 U17373 ( .I(n14037), .ZN(n14038) );
  NAND2HSV0 U17374 ( .A1(n25879), .A2(n26595), .ZN(n17468) );
  NAND2HSV0 U17375 ( .A1(n26030), .A2(\pe6/got [8]), .ZN(n25817) );
  NAND2HSV0 U17376 ( .A1(n28662), .A2(\pe6/got [8]), .ZN(n25739) );
  NAND2HSV0 U17377 ( .A1(n19076), .A2(\pe6/got [8]), .ZN(n18889) );
  CLKNHSV0 U17378 ( .I(n18398), .ZN(n28142) );
  INHSV4 U17379 ( .I(n28142), .ZN(n14039) );
  INHSV2 U17380 ( .I(n15108), .ZN(n14040) );
  CLKNHSV0 U17381 ( .I(n15108), .ZN(n28465) );
  INHSV4 U17382 ( .I(n15301), .ZN(n15086) );
  NAND2HSV4 U17383 ( .A1(n15085), .A2(n15084), .ZN(n29037) );
  CLKNAND2HSV4 U17384 ( .A1(n15083), .A2(n15082), .ZN(n15084) );
  NAND2HSV0 U17385 ( .A1(n15837), .A2(n28592), .ZN(n15838) );
  NAND2HSV0 U17386 ( .A1(n22043), .A2(n22042), .ZN(n28523) );
  NAND2HSV2 U17387 ( .A1(n22043), .A2(n22042), .ZN(n27907) );
  OR2HSV1 U17388 ( .A1(n18916), .A2(n19069), .Z(n18854) );
  CLKNAND2HSV4 U17389 ( .A1(n29019), .A2(n14698), .ZN(n25697) );
  CLKNAND2HSV2 U17390 ( .A1(n20369), .A2(n20368), .ZN(n14043) );
  CLKNAND2HSV2 U17391 ( .A1(n20369), .A2(n20368), .ZN(n20601) );
  INHSV2 U17392 ( .I(n28809), .ZN(n14044) );
  INHSV2 U17393 ( .I(n28809), .ZN(n21102) );
  CLKNHSV0 U17394 ( .I(\pe5/got [16]), .ZN(n27190) );
  NAND2HSV0 U17395 ( .A1(n28806), .A2(n14045), .ZN(n14692) );
  CLKNHSV0 U17396 ( .I(n23839), .ZN(n25272) );
  INHSV2 U17397 ( .I(n19794), .ZN(n18200) );
  NAND2HSV2 U17398 ( .A1(\pe7/aot [14]), .A2(\pe7/bq[16] ), .ZN(n19185) );
  BUFHSV8 U17399 ( .I(\pe7/bq[16] ), .Z(n25273) );
  CLKNHSV0 U17400 ( .I(n21817), .ZN(n21753) );
  NAND2HSV0 U17401 ( .A1(n21246), .A2(n21817), .ZN(n21283) );
  NAND2HSV0 U17402 ( .A1(n21817), .A2(n27544), .ZN(n21052) );
  CLKNHSV0 U17403 ( .I(\pe11/got [12]), .ZN(n24800) );
  INHSV4 U17404 ( .I(n24800), .ZN(n14049) );
  CLKNHSV0 U17405 ( .I(\pe7/aot [13]), .ZN(n14051) );
  INHSV4 U17406 ( .I(n14051), .ZN(n14050) );
  INHSV2 U17407 ( .I(\pe7/aot [13]), .ZN(n19247) );
  NAND2HSV0 U17408 ( .A1(n26925), .A2(n22903), .ZN(n22899) );
  INHSV4 U17409 ( .I(n26925), .ZN(n26916) );
  NAND2HSV2 U17410 ( .A1(n26925), .A2(n26924), .ZN(n22796) );
  CLKNHSV0 U17411 ( .I(n21979), .ZN(n22905) );
  INHSV4 U17412 ( .I(n16518), .ZN(n28627) );
  INHSV4 U17413 ( .I(n27633), .ZN(n14052) );
  NAND2HSV0 U17414 ( .A1(\pe6/bq[11] ), .A2(\pe6/aot [15]), .ZN(n14306) );
  BUFHSV8 U17415 ( .I(\pe6/aot [15]), .Z(n28680) );
  INHSV4 U17416 ( .I(n27677), .ZN(n14055) );
  INHSV2 U17417 ( .I(\pe2/aot [16]), .ZN(n21254) );
  CLKNHSV0 U17418 ( .I(\pe11/got [15]), .ZN(n25052) );
  INHSV4 U17419 ( .I(n21075), .ZN(n27312) );
  NAND2HSV0 U17420 ( .A1(n19900), .A2(n19825), .ZN(n19826) );
  NAND2HSV2 U17421 ( .A1(\pe9/ti_1 ), .A2(\pe9/got [16]), .ZN(n17888) );
  NOR2HSV4 U17422 ( .A1(n14480), .A2(n14481), .ZN(n14057) );
  NOR2HSV2 U17423 ( .A1(n14481), .A2(n14480), .ZN(n14786) );
  NAND2HSV4 U17424 ( .A1(n21318), .A2(n21317), .ZN(n14059) );
  INHSV4 U17425 ( .I(n23869), .ZN(n14060) );
  BUFHSV4 U17426 ( .I(n14086), .Z(n14061) );
  CLKNHSV0 U17427 ( .I(n27633), .ZN(n14062) );
  INHSV4 U17428 ( .I(n21321), .ZN(n28684) );
  INHSV2 U17429 ( .I(n28684), .ZN(n14063) );
  INHSV4 U17430 ( .I(n28684), .ZN(n14064) );
  NAND2HSV0 U17431 ( .A1(n17940), .A2(\pe9/ti_1 ), .ZN(n17900) );
  INHSV2 U17432 ( .I(n28673), .ZN(n14066) );
  INHSV8 U17433 ( .I(n28673), .ZN(n14067) );
  NAND2HSV0 U17434 ( .A1(n26030), .A2(n26065), .ZN(n25943) );
  NAND2HSV0 U17435 ( .A1(n26030), .A2(n28593), .ZN(n25871) );
  NAND2HSV0 U17436 ( .A1(n26030), .A2(n28586), .ZN(n25745) );
  NAND2HSV0 U17437 ( .A1(n26030), .A2(\pe6/got [7]), .ZN(n25780) );
  NAND2HSV0 U17438 ( .A1(n26030), .A2(\pe6/got [9]), .ZN(n26025) );
  NAND2HSV4 U17439 ( .A1(n25697), .A2(n25696), .ZN(n26030) );
  CLKNHSV0 U17440 ( .I(n23869), .ZN(n14068) );
  INHSV6 U17441 ( .I(\pe8/got [7]), .ZN(n23869) );
  NAND2HSV0 U17442 ( .A1(n28600), .A2(n27218), .ZN(n26480) );
  NAND2HSV0 U17443 ( .A1(n28600), .A2(\pe1/got [6]), .ZN(n26851) );
  NAND2HSV0 U17444 ( .A1(n28600), .A2(\pe1/got [8]), .ZN(n26886) );
  NAND2HSV0 U17445 ( .A1(n28600), .A2(\pe1/got [7]), .ZN(n26678) );
  NAND2HSV0 U17446 ( .A1(n28600), .A2(\pe1/got [11]), .ZN(n27189) );
  NAND2HSV0 U17447 ( .A1(n28600), .A2(\pe1/got [9]), .ZN(n23983) );
  CLKNHSV0 U17448 ( .I(\pe9/ti_1 ), .ZN(n21334) );
  CLKNHSV0 U17449 ( .I(n24685), .ZN(n14069) );
  INHSV4 U17450 ( .I(\pe7/aot [16]), .ZN(n14077) );
  CLKNHSV0 U17451 ( .I(\pe10/got [14]), .ZN(n26153) );
  INHSV4 U17452 ( .I(n26153), .ZN(n14070) );
  NAND2HSV0 U17453 ( .A1(\pe8/bq[7] ), .A2(\pe8/aot [11]), .ZN(n23615) );
  NAND2HSV0 U17454 ( .A1(\pe8/aot [9]), .A2(\pe8/bq[7] ), .ZN(n23727) );
  INHSV2 U17455 ( .I(\pe8/aot [15]), .ZN(n19995) );
  CLKNHSV0 U17456 ( .I(n17792), .ZN(n27544) );
  BUFHSV4 U17457 ( .I(\pe5/got [5]), .Z(n14072) );
  INHSV8 U17458 ( .I(n14217), .ZN(n28593) );
  CLKNHSV0 U17459 ( .I(n26601), .ZN(n14074) );
  INHSV8 U17460 ( .I(n26601), .ZN(n28648) );
  NAND2HSV0 U17461 ( .A1(\pe1/bq[10] ), .A2(\pe1/aot [16]), .ZN(n17149) );
  CLKNHSV0 U17462 ( .I(\pe3/bq[6] ), .ZN(n14075) );
  CLKNHSV0 U17463 ( .I(n14075), .ZN(n14076) );
  NAND2HSV2 U17464 ( .A1(n28424), .A2(\pe10/bq[12] ), .ZN(n16683) );
  NAND2HSV0 U17465 ( .A1(\pe1/aot [14]), .A2(\pe1/bq[14] ), .ZN(n17432) );
  NAND2HSV0 U17466 ( .A1(\pe2/aot [8]), .A2(\pe2/bq[15] ), .ZN(n27299) );
  INHSV2 U17467 ( .I(n11855), .ZN(n14078) );
  CLKNHSV0 U17468 ( .I(n28038), .ZN(n14079) );
  NAND2HSV0 U17469 ( .A1(\pe2/aot [14]), .A2(\pe2/bq[15] ), .ZN(n17718) );
  NAND2HSV0 U17470 ( .A1(\pe2/aot [14]), .A2(\pe2/bq[14] ), .ZN(n17681) );
  NAND2HSV2 U17471 ( .A1(n17172), .A2(\pe1/got [11]), .ZN(n17195) );
  NAND2HSV4 U17472 ( .A1(n16183), .A2(n16239), .ZN(n17172) );
  NAND2HSV4 U17473 ( .A1(\pe10/bq[16] ), .A2(\pe10/aot [16]), .ZN(n16609) );
  CLKNAND2HSV2 U17474 ( .A1(n19464), .A2(n19465), .ZN(n19515) );
  XOR4HSV2 U17475 ( .A1(n14428), .A2(n14427), .A3(n14426), .A4(n14425), .Z(
        n14429) );
  XNOR2HSV4 U17476 ( .A1(n14417), .A2(n25835), .ZN(n14426) );
  CLKNAND2HSV4 U17477 ( .A1(n14469), .A2(n20848), .ZN(n14553) );
  NOR2HSV4 U17478 ( .A1(n21870), .A2(n21869), .ZN(n23453) );
  NOR2HSV2 U17479 ( .A1(n28704), .A2(n20145), .ZN(n16622) );
  CLKNAND2HSV2 U17480 ( .A1(n19050), .A2(n19049), .ZN(n19051) );
  XNOR2HSV4 U17481 ( .A1(n18902), .A2(n18901), .ZN(n18914) );
  XNOR2HSV1 U17482 ( .A1(n18900), .A2(n18899), .ZN(n18902) );
  XNOR2HSV2 U17483 ( .A1(n20700), .A2(n20699), .ZN(n20776) );
  NAND3HSV2 U17484 ( .A1(n21842), .A2(n17635), .A3(\pe2/aot [15]), .ZN(n17636)
         );
  CLKXOR2HSV2 U17485 ( .A1(n17724), .A2(\pe2/phq [4]), .Z(n17726) );
  XOR2HSV4 U17486 ( .A1(n21127), .A2(n21126), .Z(n21136) );
  XOR2HSV4 U17487 ( .A1(n21125), .A2(n21124), .Z(n21126) );
  INHSV4 U17488 ( .I(n17131), .ZN(n17129) );
  NAND2HSV4 U17489 ( .A1(n26481), .A2(n26482), .ZN(n28600) );
  NAND2HSV4 U17490 ( .A1(n14860), .A2(n14859), .ZN(n14930) );
  NAND3HSV4 U17491 ( .A1(n18712), .A2(n18711), .A3(n18710), .ZN(n18713) );
  CLKNAND2HSV2 U17492 ( .A1(n15834), .A2(n15833), .ZN(n21973) );
  MUX2NHSV4 U17493 ( .I0(n20051), .I1(n25650), .S(n14034), .ZN(n19883) );
  NAND2HSV2 U17494 ( .A1(n14905), .A2(n14820), .ZN(n14813) );
  MUX2NHSV1 U17495 ( .I0(n19315), .I1(n28816), .S(n19312), .ZN(n19311) );
  NAND3HSV4 U17496 ( .A1(n15822), .A2(n15824), .A3(n15823), .ZN(n21745) );
  NAND3HSV3 U17497 ( .A1(n16535), .A2(n16459), .A3(n19830), .ZN(n16443) );
  NAND2HSV2 U17498 ( .A1(n20317), .A2(\pe11/got [15]), .ZN(n20195) );
  OAI21HSV2 U17499 ( .A1(pov6[11]), .A2(n18924), .B(n18923), .ZN(n18985) );
  NOR2HSV0 U17500 ( .A1(n27941), .A2(n21997), .ZN(n27966) );
  OAI21HSV4 U17501 ( .A1(n16358), .A2(n16357), .B(n28599), .ZN(n16364) );
  NAND2HSV2 U17502 ( .A1(n27106), .A2(n14069), .ZN(n24376) );
  CLKNHSV0 U17503 ( .I(n23549), .ZN(n23550) );
  CLKNAND2HSV4 U17504 ( .A1(n17687), .A2(n17686), .ZN(n17656) );
  NOR2HSV4 U17505 ( .A1(n17688), .A2(n25630), .ZN(n17701) );
  NAND2HSV2 U17506 ( .A1(n24377), .A2(n14503), .ZN(n24434) );
  INHSV4 U17507 ( .I(n20074), .ZN(n17068) );
  CLKNHSV0 U17508 ( .I(n19043), .ZN(n19046) );
  INHSV4 U17509 ( .I(n14298), .ZN(n14299) );
  AOI21HSV4 U17510 ( .A1(n18153), .A2(n18151), .B(n18150), .ZN(n18152) );
  NOR2HSV4 U17511 ( .A1(n24312), .A2(n16029), .ZN(n15035) );
  BUFHSV4 U17512 ( .I(n12295), .Z(n28189) );
  NAND2HSV4 U17513 ( .A1(n17473), .A2(n25680), .ZN(n17481) );
  NAND3HSV2 U17514 ( .A1(n14286), .A2(n14285), .A3(n14284), .ZN(n14296) );
  NAND2HSV0 U17515 ( .A1(\pe6/aot [13]), .A2(\pe6/bq[14] ), .ZN(n14082) );
  NAND2HSV0 U17516 ( .A1(\pe6/bq[13] ), .A2(\pe6/aot [14]), .ZN(n14081) );
  XOR2HSV2 U17517 ( .A1(n14082), .A2(n14081), .Z(n14085) );
  NAND2HSV0 U17518 ( .A1(\pe6/aot [11]), .A2(\pe6/bq[16] ), .ZN(n14084) );
  NAND2HSV0 U17519 ( .A1(\pe6/aot [16]), .A2(\pe6/bq[11] ), .ZN(n14083) );
  NAND2HSV0 U17520 ( .A1(\pe6/bq[15] ), .A2(\pe6/aot [12]), .ZN(n14088) );
  INHSV2 U17521 ( .I(\pe6/got [11]), .ZN(n22994) );
  BUFHSV8 U17522 ( .I(\pe6/ti_1 ), .Z(n19021) );
  CLKNAND2HSV1 U17523 ( .A1(n14086), .A2(n19021), .ZN(n14087) );
  XOR2HSV0 U17524 ( .A1(n14088), .A2(n14087), .Z(n14089) );
  XOR2HSV0 U17525 ( .A1(n14090), .A2(n14089), .Z(n14122) );
  CLKNAND2HSV2 U17526 ( .A1(\pe6/got [16]), .A2(\pe6/ti_1 ), .ZN(n14093) );
  INHSV6 U17527 ( .I(\pe6/got [16]), .ZN(n14118) );
  NOR2HSV4 U17528 ( .A1(n18955), .A2(n14118), .ZN(n14092) );
  MUX2NHSV4 U17529 ( .I0(n14093), .I1(n14092), .S(n14091), .ZN(n14115) );
  INHSV2 U17530 ( .I(\pe6/phq [1]), .ZN(n14095) );
  INHSV2 U17531 ( .I(\pe6/pvq [1]), .ZN(n14094) );
  NOR2HSV2 U17532 ( .A1(n14095), .A2(n14094), .ZN(n14097) );
  AOI21HSV4 U17533 ( .A1(n14220), .A2(\pe6/pvq [1]), .B(\pe6/phq [1]), .ZN(
        n14096) );
  AOI21HSV4 U17534 ( .A1(n21764), .A2(n14097), .B(n14096), .ZN(n14114) );
  XNOR2HSV4 U17535 ( .A1(n14115), .A2(n14114), .ZN(n28579) );
  INHSV6 U17536 ( .I(ctro6), .ZN(n18852) );
  CLKBUFHSV4 U17537 ( .I(n18852), .Z(n14303) );
  CLKNAND2HSV4 U17538 ( .A1(n28579), .A2(n14257), .ZN(n14099) );
  CLKAND2HSV2 U17539 ( .A1(n14281), .A2(\pe6/ti_7t [1]), .Z(n14152) );
  INHSV2 U17540 ( .I(n14152), .ZN(n14098) );
  CLKNAND2HSV4 U17541 ( .A1(n14099), .A2(n14098), .ZN(n14139) );
  INHSV2 U17542 ( .I(n14139), .ZN(n24963) );
  INHSV2 U17543 ( .I(n12437), .ZN(n14316) );
  INHSV2 U17544 ( .I(n14316), .ZN(n27073) );
  INHSV4 U17545 ( .I(\pe6/bq[12] ), .ZN(n18879) );
  INHSV2 U17546 ( .I(n18879), .ZN(n25701) );
  NAND2HSV2 U17547 ( .A1(n28680), .A2(n25701), .ZN(n14100) );
  XNOR2HSV4 U17548 ( .A1(n14101), .A2(n14100), .ZN(n14103) );
  CLKNHSV0 U17549 ( .I(\pe6/got [12]), .ZN(n14105) );
  INHSV1 U17550 ( .I(n14105), .ZN(n14102) );
  CLKNAND2HSV1 U17551 ( .A1(n14103), .A2(n14102), .ZN(n14107) );
  INHSV4 U17552 ( .I(n14139), .ZN(n14156) );
  INHSV2 U17553 ( .I(n14103), .ZN(n14104) );
  OAI21HSV4 U17554 ( .A1(n14156), .A2(n14105), .B(n14104), .ZN(n14106) );
  OAI21HSV4 U17555 ( .A1(n24963), .A2(n14107), .B(n14106), .ZN(n14121) );
  NAND2HSV2 U17556 ( .A1(n14110), .A2(n14109), .ZN(n14111) );
  INHSV3 U17557 ( .I(\pe6/got [15]), .ZN(n19056) );
  NOR2HSV4 U17558 ( .A1(n19056), .A2(n18955), .ZN(n14113) );
  XNOR2HSV4 U17559 ( .A1(n14145), .A2(n14144), .ZN(n14117) );
  XNOR2HSV4 U17560 ( .A1(n14115), .A2(n14114), .ZN(n14119) );
  CLKBUFHSV4 U17561 ( .I(n18852), .Z(n18915) );
  CLKBUFHSV4 U17562 ( .I(n18915), .Z(n14280) );
  INHSV2 U17563 ( .I(n14118), .ZN(n28472) );
  NAND2HSV2 U17564 ( .A1(n14280), .A2(n28472), .ZN(n14406) );
  INHSV2 U17565 ( .I(n14406), .ZN(n14396) );
  NAND2HSV4 U17566 ( .A1(n14117), .A2(n14181), .ZN(n14148) );
  CLKBUFHSV4 U17567 ( .I(n14280), .Z(n19141) );
  NAND2HSV2 U17568 ( .A1(n19045), .A2(\pe6/ti_7t [2]), .ZN(n14182) );
  INHSV2 U17569 ( .I(n14182), .ZN(n14146) );
  INHSV2 U17570 ( .I(n14146), .ZN(n14116) );
  BUFHSV2 U17571 ( .I(\pe6/got [16]), .Z(n25647) );
  BUFHSV2 U17572 ( .I(n14303), .Z(n18920) );
  XOR3HSV2 U17573 ( .A1(n14122), .A2(n14121), .A3(n14120), .Z(n14166) );
  CLKNAND2HSV1 U17574 ( .A1(\pe6/got [14]), .A2(\pe6/ti_1 ), .ZN(n14126) );
  MUX2NHSV4 U17575 ( .I0(n14126), .I1(n14125), .S(n14124), .ZN(n14133) );
  CLKNHSV0 U17576 ( .I(n14048), .ZN(n18871) );
  CLKNAND2HSV1 U17577 ( .A1(n14220), .A2(\pe6/pvq [3]), .ZN(n14127) );
  INHSV2 U17578 ( .I(\pe6/phq [3]), .ZN(n14129) );
  CLKNAND2HSV1 U17579 ( .A1(n14127), .A2(n14129), .ZN(n14132) );
  INHSV2 U17580 ( .I(\pe6/pvq [3]), .ZN(n14128) );
  NOR2HSV2 U17581 ( .A1(n14129), .A2(n14128), .ZN(n14130) );
  NAND2HSV2 U17582 ( .A1(n14130), .A2(n12437), .ZN(n14131) );
  NAND2HSV2 U17583 ( .A1(n14133), .A2(n14134), .ZN(n14138) );
  INHSV2 U17584 ( .I(n14133), .ZN(n14136) );
  CLKNAND2HSV3 U17585 ( .A1(n14136), .A2(n14135), .ZN(n14137) );
  XNOR2HSV4 U17586 ( .A1(n14142), .A2(n14141), .ZN(n27210) );
  INHSV2 U17587 ( .I(n27210), .ZN(n14140) );
  INHSV4 U17588 ( .I(n14139), .ZN(n25455) );
  NAND2HSV2 U17589 ( .A1(n14140), .A2(n25455), .ZN(n14192) );
  XNOR2HSV4 U17590 ( .A1(n14142), .A2(n14141), .ZN(n14158) );
  INHSV4 U17591 ( .I(n19056), .ZN(n18847) );
  CLKNHSV0 U17592 ( .I(n19055), .ZN(n14143) );
  OAI21HSV2 U17593 ( .A1(n14158), .A2(n18847), .B(n14143), .ZN(n14244) );
  INHSV2 U17594 ( .I(n14244), .ZN(n14189) );
  XNOR2HSV4 U17595 ( .A1(n14145), .A2(n14144), .ZN(n24964) );
  INHSV2 U17596 ( .I(n28472), .ZN(n14745) );
  INHSV2 U17597 ( .I(n14745), .ZN(n25058) );
  INHSV4 U17598 ( .I(n14148), .ZN(n14149) );
  NOR2HSV8 U17599 ( .A1(n14150), .A2(n14149), .ZN(n14157) );
  CLKNAND2HSV1 U17600 ( .A1(n14189), .A2(n27212), .ZN(n14151) );
  INHSV2 U17601 ( .I(n14151), .ZN(n14164) );
  CLKNAND2HSV1 U17602 ( .A1(n14152), .A2(n18847), .ZN(n14155) );
  CLKNAND2HSV0 U17603 ( .A1(n19160), .A2(n18847), .ZN(n14153) );
  INAND2HSV2 U17604 ( .A1(n14153), .B1(n28579), .ZN(n14154) );
  CLKNAND2HSV2 U17605 ( .A1(n14155), .A2(n14154), .ZN(n27211) );
  NAND2HSV2 U17606 ( .A1(n27210), .A2(n27211), .ZN(n14191) );
  CLKBUFHSV4 U17607 ( .I(\pe6/got [14]), .Z(n28686) );
  AND2HSV2 U17608 ( .A1(n14191), .A2(n28686), .Z(n14163) );
  NAND2HSV2 U17609 ( .A1(n27210), .A2(n14156), .ZN(n14186) );
  NAND2HSV0 U17610 ( .A1(n14186), .A2(\pe6/got [14]), .ZN(n14161) );
  BUFHSV2 U17611 ( .I(n19056), .Z(n14253) );
  AOI21HSV4 U17612 ( .A1(n14158), .A2(n14253), .B(n19055), .ZN(n14251) );
  CLKNAND2HSV3 U17613 ( .A1(n14157), .A2(n14251), .ZN(n14188) );
  CLKNHSV0 U17614 ( .I(n14187), .ZN(n14160) );
  NAND2HSV2 U17615 ( .A1(n18992), .A2(\pe6/ti_7t [3]), .ZN(n14326) );
  CLKNHSV0 U17616 ( .I(\pe6/got [14]), .ZN(n18996) );
  OR2HSV1 U17617 ( .A1(n14326), .A2(n18996), .Z(n14159) );
  OAI31HSV2 U17618 ( .A1(n14161), .A2(n14188), .A3(n14160), .B(n14159), .ZN(
        n14162) );
  AOI31HSV2 U17619 ( .A1(n14192), .A2(n14164), .A3(n14163), .B(n14162), .ZN(
        n14165) );
  XOR2HSV4 U17620 ( .A1(n14166), .A2(n14165), .Z(n14209) );
  XNOR2HSV4 U17621 ( .A1(n14168), .A2(n14167), .ZN(n14172) );
  NAND2HSV2 U17622 ( .A1(\pe6/bq[15] ), .A2(\pe6/aot [14]), .ZN(n14170) );
  INHSV2 U17623 ( .I(n14047), .ZN(n23525) );
  NAND2HSV2 U17624 ( .A1(n23525), .A2(\pe6/pvq [4]), .ZN(n14169) );
  XOR3HSV2 U17625 ( .A1(\pe6/phq [4]), .A2(n14170), .A3(n14169), .Z(n14171) );
  XNOR2HSV4 U17626 ( .A1(n14172), .A2(n14171), .ZN(n14176) );
  OAI21HSV0 U17627 ( .A1(n14303), .A2(\pe6/ti_7t [1]), .B(\pe6/got [14]), .ZN(
        n14173) );
  CLKNHSV0 U17628 ( .I(n14173), .ZN(n14174) );
  OAI21HSV2 U17629 ( .A1(n28579), .A2(n19045), .B(n14174), .ZN(n14175) );
  XNOR2HSV4 U17630 ( .A1(n14176), .A2(n14175), .ZN(n14200) );
  INHSV2 U17631 ( .I(n18927), .ZN(n19147) );
  NOR2HSV1 U17632 ( .A1(n19147), .A2(n14253), .ZN(n14177) );
  CLKAND2HSV2 U17633 ( .A1(n14178), .A2(n14177), .Z(n14180) );
  NAND2HSV2 U17634 ( .A1(n14180), .A2(n14179), .ZN(n14199) );
  NAND2HSV4 U17635 ( .A1(n13969), .A2(n24964), .ZN(n14198) );
  OR2HSV1 U17636 ( .A1(n14182), .A2(n14253), .Z(n14183) );
  NAND3HSV3 U17637 ( .A1(n14198), .A2(n14199), .A3(n14183), .ZN(n14184) );
  XNOR2HSV4 U17638 ( .A1(n14200), .A2(n14184), .ZN(n25648) );
  INHSV2 U17639 ( .I(\pe6/got [15]), .ZN(n14304) );
  INHSV2 U17640 ( .I(n14304), .ZN(n25420) );
  CLKNAND2HSV3 U17641 ( .A1(n14187), .A2(n14186), .ZN(n14250) );
  NOR2HSV4 U17642 ( .A1(n14188), .A2(n14250), .ZN(n14328) );
  INHSV4 U17643 ( .I(n14328), .ZN(n14284) );
  INHSV2 U17644 ( .I(n14284), .ZN(n14195) );
  NAND2HSV4 U17645 ( .A1(n14192), .A2(n14191), .ZN(n14247) );
  INHSV4 U17646 ( .I(n14247), .ZN(n14288) );
  NAND2HSV2 U17647 ( .A1(n14289), .A2(n14288), .ZN(n14193) );
  INHSV2 U17648 ( .I(n19151), .ZN(n19160) );
  OR2HSV4 U17649 ( .A1(n28472), .A2(n19045), .Z(n18907) );
  NAND2HSV2 U17650 ( .A1(n19055), .A2(\pe6/ti_7t [4]), .ZN(n14291) );
  INHSV2 U17651 ( .I(n14291), .ZN(n14287) );
  CLKNAND2HSV1 U17652 ( .A1(n14213), .A2(n14291), .ZN(n14203) );
  NAND3HSV2 U17653 ( .A1(n14286), .A2(n14284), .A3(n14291), .ZN(n14202) );
  OA21HSV2 U17654 ( .A1(n14285), .A2(n14287), .B(n25420), .Z(n14201) );
  NAND3HSV2 U17655 ( .A1(n14203), .A2(n14202), .A3(n14201), .ZN(n14204) );
  INHSV2 U17656 ( .I(n14208), .ZN(n14206) );
  CLKNAND2HSV2 U17657 ( .A1(n14209), .A2(n14208), .ZN(n14210) );
  INHSV2 U17658 ( .I(n14285), .ZN(n14212) );
  AOI21HSV4 U17659 ( .A1(n14214), .A2(n14259), .B(n14287), .ZN(n14270) );
  NAND2HSV0 U17660 ( .A1(\pe6/aot [14]), .A2(\pe6/bq[14] ), .ZN(n14216) );
  INHSV4 U17661 ( .I(\pe6/got [12]), .ZN(n14217) );
  NAND2HSV2 U17662 ( .A1(\pe6/got [12]), .A2(\pe6/ti_1 ), .ZN(n14218) );
  NAND2HSV2 U17663 ( .A1(n18871), .A2(\pe6/pvq [5]), .ZN(n14222) );
  NAND2HSV0 U17664 ( .A1(\pe6/aot [15]), .A2(\pe6/bq[13] ), .ZN(n14221) );
  NAND2HSV2 U17665 ( .A1(\pe6/aot [16]), .A2(\pe6/bq[12] ), .ZN(n14223) );
  XNOR2HSV1 U17666 ( .A1(n14223), .A2(\pe6/phq [5]), .ZN(n14224) );
  NAND2HSV4 U17667 ( .A1(n14226), .A2(n14225), .ZN(n14228) );
  CLKNAND2HSV3 U17668 ( .A1(n14227), .A2(n14228), .ZN(n14238) );
  CLKNHSV2 U17669 ( .I(n14227), .ZN(n14230) );
  CLKNAND2HSV2 U17670 ( .A1(n14228), .A2(n22992), .ZN(n14229) );
  NOR2HSV4 U17671 ( .A1(n14230), .A2(n14229), .ZN(n14233) );
  AOI22HSV4 U17672 ( .A1(n14361), .A2(n14238), .B1(n14233), .B2(n14231), .ZN(
        n14235) );
  INHSV1 U17673 ( .I(n14239), .ZN(n14232) );
  CLKNAND2HSV2 U17674 ( .A1(n14233), .A2(n14232), .ZN(n14234) );
  CLKNAND2HSV4 U17675 ( .A1(n14235), .A2(n14234), .ZN(n14242) );
  INHSV2 U17676 ( .I(n25455), .ZN(n14321) );
  CLKNAND2HSV2 U17677 ( .A1(n14321), .A2(n14236), .ZN(n14240) );
  INHSV2 U17678 ( .I(n14240), .ZN(n14237) );
  NAND2HSV4 U17679 ( .A1(n14242), .A2(n14237), .ZN(n14263) );
  CLKNAND2HSV3 U17680 ( .A1(n13975), .A2(n12766), .ZN(n14241) );
  OAI22HSV4 U17681 ( .A1(n14243), .A2(n14242), .B1(n14241), .B2(n14240), .ZN(
        n14265) );
  NOR2HSV0 U17682 ( .A1(n14244), .A2(n14253), .ZN(n14245) );
  CLKNAND2HSV1 U17683 ( .A1(n14245), .A2(n27212), .ZN(n14246) );
  INHSV2 U17684 ( .I(n14246), .ZN(n14249) );
  INHSV2 U17685 ( .I(n14247), .ZN(n14248) );
  NAND2HSV4 U17686 ( .A1(n14249), .A2(n14248), .ZN(n14262) );
  INHSV2 U17687 ( .I(n14250), .ZN(n14256) );
  CLKNAND2HSV1 U17688 ( .A1(n14251), .A2(n18847), .ZN(n14252) );
  NOR2HSV2 U17689 ( .A1(n27212), .A2(n14252), .ZN(n14255) );
  NOR2HSV2 U17690 ( .A1(n14326), .A2(n14253), .ZN(n14254) );
  AOI21HSV4 U17691 ( .A1(n14256), .A2(n14255), .B(n14254), .ZN(n14264) );
  CLKNHSV0 U17692 ( .I(n19138), .ZN(n14257) );
  NAND3HSV4 U17693 ( .A1(n14264), .A2(n14263), .A3(n14262), .ZN(n14266) );
  INHSV2 U17694 ( .I(n14281), .ZN(n14267) );
  NAND3HSV4 U17695 ( .A1(n14275), .A2(n14274), .A3(n13980), .ZN(n14277) );
  CLKNAND2HSV2 U17696 ( .A1(n14276), .A2(n14277), .ZN(n14338) );
  INHSV3 U17697 ( .I(n14277), .ZN(n14279) );
  CLKNAND2HSV3 U17698 ( .A1(n14279), .A2(n14278), .ZN(n14337) );
  INHSV2 U17699 ( .I(n14303), .ZN(n19142) );
  NAND2HSV2 U17700 ( .A1(n19142), .A2(\pe6/ti_7t [6]), .ZN(n14339) );
  BUFHSV2 U17701 ( .I(n14280), .Z(n19069) );
  INHSV2 U17702 ( .I(n14369), .ZN(n14281) );
  NAND2HSV2 U17703 ( .A1(n14281), .A2(n14339), .ZN(n14282) );
  CLKNAND2HSV4 U17704 ( .A1(n14283), .A2(n14282), .ZN(n14397) );
  INHSV2 U17705 ( .I(n14745), .ZN(n25419) );
  AND2HSV2 U17706 ( .A1(n19160), .A2(n25419), .Z(n14285) );
  INHSV2 U17707 ( .I(n25648), .ZN(n14295) );
  NOR2HSV0 U17708 ( .A1(n14328), .A2(n14287), .ZN(n14290) );
  CLKNAND2HSV3 U17709 ( .A1(n14289), .A2(n14288), .ZN(n14329) );
  AOI21HSV2 U17710 ( .A1(n14290), .A2(n14329), .B(n24962), .ZN(n14293) );
  NAND2HSV2 U17711 ( .A1(n25648), .A2(n14291), .ZN(n14292) );
  CLKNAND2HSV1 U17712 ( .A1(n14293), .A2(n14292), .ZN(n14294) );
  NAND2HSV2 U17713 ( .A1(n14297), .A2(n14298), .ZN(n14302) );
  INHSV2 U17714 ( .I(n14297), .ZN(n14300) );
  CLKNAND2HSV3 U17715 ( .A1(n14300), .A2(n14299), .ZN(n14301) );
  CLKNAND2HSV4 U17716 ( .A1(n14301), .A2(n14302), .ZN(n14367) );
  INHSV2 U17717 ( .I(n14368), .ZN(n14360) );
  INHSV2 U17718 ( .I(n18852), .ZN(n19151) );
  INHSV2 U17719 ( .I(\pe6/got [15]), .ZN(n19048) );
  AO21HSV1 U17720 ( .A1(n14360), .A2(n19151), .B(n19048), .Z(n14305) );
  AOI21HSV4 U17721 ( .A1(n14367), .A2(n14360), .B(n14305), .ZN(n14336) );
  CLKNAND2HSV2 U17722 ( .A1(n14391), .A2(n28686), .ZN(n14334) );
  CLKNHSV2 U17723 ( .I(n14306), .ZN(n14307) );
  XNOR2HSV4 U17724 ( .A1(n14308), .A2(n14307), .ZN(n14310) );
  CLKNAND2HSV0 U17725 ( .A1(n19021), .A2(\pe6/got [10]), .ZN(n14309) );
  XNOR2HSV4 U17726 ( .A1(n14310), .A2(n14309), .ZN(n14314) );
  NAND2HSV0 U17727 ( .A1(\pe6/aot [13]), .A2(\pe6/bq[13] ), .ZN(n18875) );
  NAND2HSV0 U17728 ( .A1(\pe6/aot [11]), .A2(\pe6/bq[15] ), .ZN(n14315) );
  XOR2HSV0 U17729 ( .A1(n18875), .A2(n14315), .Z(n14318) );
  INHSV4 U17730 ( .I(n14316), .ZN(n27072) );
  NAND2HSV2 U17731 ( .A1(n27072), .A2(\pe6/pvq [7]), .ZN(n14317) );
  XNOR2HSV1 U17732 ( .A1(n14318), .A2(n14317), .ZN(n14319) );
  XNOR2HSV4 U17733 ( .A1(n14320), .A2(n14319), .ZN(n14323) );
  CLKNAND2HSV1 U17734 ( .A1(n14321), .A2(n28586), .ZN(n14322) );
  XNOR2HSV4 U17735 ( .A1(n14323), .A2(n14322), .ZN(n14325) );
  NAND2HSV0 U17736 ( .A1(n28798), .A2(n28593), .ZN(n14324) );
  XNOR2HSV4 U17737 ( .A1(n14325), .A2(n14324), .ZN(n14332) );
  CLKNHSV1 U17738 ( .I(n14326), .ZN(n14327) );
  NOR2HSV2 U17739 ( .A1(n14328), .A2(n14327), .ZN(n14330) );
  NAND2HSV4 U17740 ( .A1(n14330), .A2(n14329), .ZN(n28793) );
  XNOR2HSV4 U17741 ( .A1(n14336), .A2(n14335), .ZN(n14736) );
  CLKNAND2HSV1 U17742 ( .A1(n14338), .A2(n14337), .ZN(n28966) );
  AOI21HSV4 U17743 ( .A1(n14340), .A2(n14339), .B(n19048), .ZN(n14366) );
  INHSV3 U17744 ( .I(n25455), .ZN(\pe6/ti_7[1] ) );
  NAND2HSV2 U17745 ( .A1(\pe6/ti_7[1] ), .A2(\pe6/got [10]), .ZN(n14355) );
  CLKNAND2HSV1 U17746 ( .A1(\pe6/aot [11]), .A2(\pe6/bq[14] ), .ZN(n23021) );
  NAND2HSV0 U17747 ( .A1(\pe6/aot [15]), .A2(\pe6/bq[10] ), .ZN(n14341) );
  NAND2HSV0 U17748 ( .A1(\pe6/aot [14]), .A2(\pe6/bq[11] ), .ZN(n14343) );
  NAND2HSV0 U17749 ( .A1(\pe6/aot [9]), .A2(\pe6/bq[16] ), .ZN(n14342) );
  XOR2HSV0 U17750 ( .A1(n14343), .A2(n14342), .Z(n14344) );
  NAND2HSV0 U17751 ( .A1(\pe6/bq[15] ), .A2(\pe6/aot [10]), .ZN(n14346) );
  NAND2HSV0 U17752 ( .A1(\pe6/aot [16]), .A2(\pe6/bq[9] ), .ZN(n14345) );
  XOR2HSV0 U17753 ( .A1(n14346), .A2(n14345), .Z(n14350) );
  NAND2HSV0 U17754 ( .A1(\pe6/bq[13] ), .A2(\pe6/aot [12]), .ZN(n14348) );
  NAND2HSV0 U17755 ( .A1(\pe6/got [9]), .A2(n19021), .ZN(n14347) );
  XOR2HSV0 U17756 ( .A1(n14348), .A2(n14347), .Z(n14349) );
  XOR2HSV0 U17757 ( .A1(n14350), .A2(n14349), .Z(n14351) );
  XNOR2HSV4 U17758 ( .A1(n14352), .A2(n14351), .ZN(n14354) );
  CLKBUFHSV4 U17759 ( .I(n28798), .Z(n18930) );
  NAND2HSV2 U17760 ( .A1(n18930), .A2(\pe6/got [11]), .ZN(n14353) );
  XOR3HSV2 U17761 ( .A1(n14355), .A2(n14354), .A3(n14353), .Z(n14357) );
  NAND2HSV0 U17762 ( .A1(n28793), .A2(n28593), .ZN(n14356) );
  XNOR2HSV1 U17763 ( .A1(n14357), .A2(n14356), .ZN(n14359) );
  NAND2HSV0 U17764 ( .A1(n14391), .A2(n14236), .ZN(n14358) );
  XNOR2HSV1 U17765 ( .A1(n14359), .A2(n14358), .ZN(n14364) );
  INHSV2 U17766 ( .I(n19151), .ZN(n14369) );
  CLKNAND2HSV1 U17767 ( .A1(n22992), .A2(n14369), .ZN(n14362) );
  OAI22HSV2 U17768 ( .A1(n14367), .A2(n14362), .B1(n14361), .B2(n14360), .ZN(
        n14363) );
  XNOR2HSV4 U17769 ( .A1(n14364), .A2(n14363), .ZN(n14365) );
  NAND2HSV2 U17770 ( .A1(n14696), .A2(n25058), .ZN(n18849) );
  INHSV4 U17771 ( .I(n14367), .ZN(n28678) );
  NAND2HSV0 U17772 ( .A1(\pe6/bq[16] ), .A2(\pe6/aot [8]), .ZN(n14371) );
  CLKNAND2HSV0 U17773 ( .A1(n19021), .A2(\pe6/got [8]), .ZN(n14370) );
  XOR2HSV0 U17774 ( .A1(n14371), .A2(n14370), .Z(n14375) );
  NAND2HSV0 U17775 ( .A1(\pe6/bq[14] ), .A2(\pe6/aot [10]), .ZN(n14373) );
  NAND2HSV0 U17776 ( .A1(\pe6/aot [14]), .A2(\pe6/bq[10] ), .ZN(n14372) );
  XOR2HSV0 U17777 ( .A1(n14373), .A2(n14372), .Z(n14374) );
  XOR2HSV0 U17778 ( .A1(n14375), .A2(n14374), .Z(n14381) );
  INHSV4 U17779 ( .I(n23525), .ZN(n27074) );
  NAND2HSV0 U17780 ( .A1(\pe6/aot [9]), .A2(\pe6/bq[15] ), .ZN(n14377) );
  NAND2HSV0 U17781 ( .A1(\pe6/aot [13]), .A2(\pe6/bq[11] ), .ZN(n14376) );
  XOR2HSV0 U17782 ( .A1(n14377), .A2(n14376), .Z(n14378) );
  XNOR2HSV4 U17783 ( .A1(n14379), .A2(n14378), .ZN(n14380) );
  XOR2HSV0 U17784 ( .A1(n14381), .A2(n14380), .Z(n14389) );
  NAND2HSV0 U17785 ( .A1(\pe6/aot [11]), .A2(\pe6/bq[13] ), .ZN(n14383) );
  NAND2HSV0 U17786 ( .A1(n28680), .A2(\pe6/bq[9] ), .ZN(n14382) );
  XOR2HSV0 U17787 ( .A1(n14383), .A2(n14382), .Z(n14387) );
  NAND2HSV0 U17788 ( .A1(\pe6/bq[12] ), .A2(\pe6/aot [12]), .ZN(n14385) );
  BUFHSV2 U17789 ( .I(\pe6/aot [16]), .Z(n28681) );
  CLKNAND2HSV1 U17790 ( .A1(n28681), .A2(\pe6/bq[8] ), .ZN(n14384) );
  XOR2HSV0 U17791 ( .A1(n14385), .A2(n14384), .Z(n14386) );
  XOR2HSV0 U17792 ( .A1(n14387), .A2(n14386), .Z(n14388) );
  INHSV2 U17793 ( .I(n28793), .ZN(n22996) );
  INHSV4 U17794 ( .I(n22996), .ZN(n19076) );
  INHSV2 U17795 ( .I(n14391), .ZN(n18968) );
  INHSV4 U17796 ( .I(n18968), .ZN(n19109) );
  XNOR2HSV4 U17797 ( .A1(n14393), .A2(n14392), .ZN(n14395) );
  XNOR2HSV4 U17798 ( .A1(n14395), .A2(n14394), .ZN(n14403) );
  INHSV2 U17799 ( .I(n14397), .ZN(n28526) );
  NOR2HSV2 U17800 ( .A1(n14736), .A2(n19045), .ZN(n14399) );
  INHSV2 U17801 ( .I(n14400), .ZN(n14738) );
  NOR2HSV1 U17802 ( .A1(n14738), .A2(n19048), .ZN(n14401) );
  XNOR2HSV4 U17803 ( .A1(n14403), .A2(n14402), .ZN(n25059) );
  CLKNAND2HSV2 U17804 ( .A1(n25059), .A2(n14267), .ZN(n14404) );
  CLKNHSV2 U17805 ( .I(n14404), .ZN(n14405) );
  CLKNAND2HSV3 U17806 ( .A1(n18849), .A2(n14405), .ZN(n14407) );
  INHSV2 U17807 ( .I(n18915), .ZN(n19138) );
  CLKBUFHSV4 U17808 ( .I(n28938), .Z(n19121) );
  INHSV2 U17809 ( .I(\pe6/ti_7t [8]), .ZN(n14697) );
  AOI21HSV2 U17810 ( .A1(n14697), .A2(n18992), .B(n19048), .ZN(n14410) );
  NAND2HSV2 U17811 ( .A1(n28681), .A2(\pe6/bq[7] ), .ZN(n14718) );
  NAND2HSV0 U17812 ( .A1(\pe6/aot [11]), .A2(n25701), .ZN(n18881) );
  XOR2HSV0 U17813 ( .A1(n14718), .A2(n18881), .Z(n14428) );
  NAND2HSV0 U17814 ( .A1(\pe6/aot [12]), .A2(\pe6/bq[11] ), .ZN(n14412) );
  NAND2HSV0 U17815 ( .A1(n28680), .A2(\pe6/bq[8] ), .ZN(n14411) );
  XOR2HSV0 U17816 ( .A1(n14412), .A2(n14411), .Z(n14416) );
  NAND2HSV0 U17817 ( .A1(\pe6/bq[15] ), .A2(\pe6/aot [8]), .ZN(n14414) );
  NAND2HSV0 U17818 ( .A1(\pe6/aot [9]), .A2(\pe6/bq[14] ), .ZN(n14413) );
  XOR2HSV0 U17819 ( .A1(n14414), .A2(n14413), .Z(n14415) );
  XNOR2HSV1 U17820 ( .A1(n14416), .A2(n14415), .ZN(n14427) );
  INHSV2 U17821 ( .I(n14316), .ZN(n23498) );
  NAND2HSV0 U17822 ( .A1(\pe6/aot [13]), .A2(\pe6/bq[10] ), .ZN(n14420) );
  NAND2HSV0 U17823 ( .A1(\pe6/got [7]), .A2(n19021), .ZN(n14419) );
  XOR2HSV0 U17824 ( .A1(n14420), .A2(n14419), .Z(n14424) );
  NAND2HSV0 U17825 ( .A1(\pe6/aot [7]), .A2(\pe6/bq[16] ), .ZN(n14422) );
  NAND2HSV0 U17826 ( .A1(\pe6/aot [14]), .A2(\pe6/bq[9] ), .ZN(n14421) );
  XOR2HSV0 U17827 ( .A1(n14422), .A2(n14421), .Z(n14423) );
  XOR2HSV0 U17828 ( .A1(n14424), .A2(n14423), .Z(n14425) );
  INHSV2 U17829 ( .I(n14433), .ZN(n21374) );
  NAND2HSV0 U17830 ( .A1(n21374), .A2(\pe5/aot [13]), .ZN(n14435) );
  NAND2HSV0 U17831 ( .A1(\pe5/aot [12]), .A2(\pe5/bq[16] ), .ZN(n14434) );
  INAND2HSV1 U17832 ( .A1(n14766), .B1(\pe5/aot [16]), .ZN(n14437) );
  INHSV2 U17833 ( .I(n14777), .ZN(n14646) );
  NAND2HSV2 U17834 ( .A1(n14646), .A2(\pe5/pvq [5]), .ZN(n14438) );
  CLKNAND2HSV1 U17835 ( .A1(\pe5/bq[13] ), .A2(\pe5/aot [14]), .ZN(n14534) );
  CLKNHSV0 U17836 ( .I(\pe5/aot [15]), .ZN(n14883) );
  INHSV2 U17837 ( .I(\pe5/bq[13] ), .ZN(n21357) );
  NAND2HSV0 U17838 ( .A1(\pe5/bq[14] ), .A2(\pe5/aot [14]), .ZN(n14439) );
  OAI21HSV2 U17839 ( .A1(n14883), .A2(n21357), .B(n14439), .ZN(n14440) );
  NAND2HSV2 U17840 ( .A1(n20870), .A2(\pe5/ti_7t [1]), .ZN(n14441) );
  INHSV4 U17841 ( .I(n14443), .ZN(n14458) );
  INHSV4 U17842 ( .I(n14444), .ZN(n14457) );
  CLKNAND2HSV3 U17843 ( .A1(n28455), .A2(n14631), .ZN(n14519) );
  INHSV4 U17844 ( .I(\pe5/pvq [2]), .ZN(n14447) );
  INHSV4 U17845 ( .I(\pe5/phq [2]), .ZN(n14446) );
  OAI21HSV4 U17846 ( .A1(n14448), .A2(n14447), .B(n14446), .ZN(n14449) );
  XNOR2HSV4 U17847 ( .A1(n14452), .A2(n14451), .ZN(n14456) );
  CLKXOR2HSV4 U17848 ( .A1(n14454), .A2(n14453), .Z(n14455) );
  XNOR2HSV4 U17849 ( .A1(n14456), .A2(n14455), .ZN(n27192) );
  CLKNAND2HSV3 U17850 ( .A1(n14458), .A2(n14457), .ZN(n14460) );
  INAND2HSV2 U17851 ( .A1(n27190), .B1(n21342), .ZN(n14459) );
  INHSV2 U17852 ( .I(n14459), .ZN(n14909) );
  INHSV4 U17853 ( .I(n21422), .ZN(n21421) );
  NAND2HSV2 U17854 ( .A1(n21421), .A2(\pe5/ti_7t [2]), .ZN(n14518) );
  INHSV4 U17855 ( .I(n14058), .ZN(n14552) );
  INHSV2 U17856 ( .I(\pe5/got [14]), .ZN(n14547) );
  XNOR2HSV4 U17857 ( .A1(n14462), .A2(n14461), .ZN(n14493) );
  NAND2HSV2 U17858 ( .A1(n21421), .A2(\pe5/ti_7t [3]), .ZN(n14578) );
  INHSV2 U17859 ( .I(\pe5/got [15]), .ZN(n14676) );
  INHSV2 U17860 ( .I(n14478), .ZN(n14517) );
  INHSV2 U17861 ( .I(\pe5/got [16]), .ZN(n14559) );
  CLKAND2HSV1 U17862 ( .A1(n14473), .A2(n14482), .Z(n14463) );
  NAND2HSV2 U17863 ( .A1(\pe5/pvq [3]), .A2(\pe5/ctrq ), .ZN(n14465) );
  NAND2HSV2 U17864 ( .A1(\pe5/ti_1 ), .A2(\pe5/got [14]), .ZN(n14464) );
  CLKNAND2HSV1 U17865 ( .A1(\pe5/aot [15]), .A2(\pe5/bq[15] ), .ZN(n14468) );
  CLKNAND2HSV2 U17866 ( .A1(\pe5/bq[15] ), .A2(\pe5/aot [15]), .ZN(n14466) );
  CLKNAND2HSV2 U17867 ( .A1(n14466), .A2(\pe5/phq [3]), .ZN(n14467) );
  NAND2HSV2 U17868 ( .A1(n25644), .A2(n13992), .ZN(n14469) );
  XNOR2HSV4 U17869 ( .A1(n14471), .A2(n14470), .ZN(n14484) );
  INAND2HSV2 U17870 ( .A1(n14474), .B1(n25644), .ZN(n14558) );
  INHSV2 U17871 ( .I(n14558), .ZN(n14576) );
  INHSV2 U17872 ( .I(n14478), .ZN(n14684) );
  NAND2HSV0 U17873 ( .A1(\pe5/got [15]), .A2(n14482), .ZN(n14483) );
  INHSV2 U17874 ( .I(n14501), .ZN(n14549) );
  NOR2HSV4 U17875 ( .A1(n14487), .A2(n14486), .ZN(n14573) );
  OAI21HSV4 U17876 ( .A1(n14491), .A2(n14490), .B(n14489), .ZN(n14492) );
  XNOR2HSV4 U17877 ( .A1(n14493), .A2(n14492), .ZN(n14620) );
  CLKNAND2HSV2 U17878 ( .A1(n14496), .A2(n14495), .ZN(n14555) );
  INHSV2 U17879 ( .I(n14497), .ZN(n14498) );
  NOR2HSV2 U17880 ( .A1(n14553), .A2(n14498), .ZN(n14499) );
  NAND3HSV3 U17881 ( .A1(n14573), .A2(n24406), .A3(n14502), .ZN(n22097) );
  NAND2HSV2 U17882 ( .A1(n22094), .A2(n22097), .ZN(n14525) );
  NAND2HSV0 U17883 ( .A1(\pe5/aot [15]), .A2(\pe5/bq[14] ), .ZN(n14504) );
  CLKNHSV0 U17884 ( .I(\pe5/aot [16]), .ZN(n23789) );
  NOR2HSV2 U17885 ( .A1(n23789), .A2(n21357), .ZN(n20953) );
  BUFHSV2 U17886 ( .I(n14506), .Z(n14757) );
  INHSV2 U17887 ( .I(n14757), .ZN(n14616) );
  INHSV2 U17888 ( .I(\pe5/got [14]), .ZN(n21411) );
  CLKNAND2HSV1 U17889 ( .A1(n14507), .A2(n14508), .ZN(n14512) );
  INHSV2 U17890 ( .I(n14508), .ZN(n14509) );
  CLKNAND2HSV3 U17891 ( .A1(n14510), .A2(n14509), .ZN(n14511) );
  NOR2HSV1 U17892 ( .A1(n14513), .A2(n14517), .ZN(n14516) );
  INHSV2 U17893 ( .I(n14514), .ZN(n14515) );
  CLKNAND2HSV1 U17894 ( .A1(n14516), .A2(n14515), .ZN(n14522) );
  OR2HSV1 U17895 ( .A1(n14518), .A2(n14517), .Z(n14521) );
  NAND3HSV2 U17896 ( .A1(n14519), .A2(n21347), .A3(n27192), .ZN(n14520) );
  NAND3HSV2 U17897 ( .A1(n14522), .A2(n14521), .A3(n14520), .ZN(n14527) );
  XNOR2HSV4 U17898 ( .A1(n14528), .A2(n14527), .ZN(n14524) );
  CLKAND2HSV2 U17899 ( .A1(n21421), .A2(\pe5/ti_7t [4]), .Z(n14523) );
  AOI21HSV4 U17900 ( .A1(n14525), .A2(n14524), .B(n14523), .ZN(n14606) );
  XOR2HSV2 U17901 ( .A1(n14528), .A2(n14527), .Z(n22099) );
  CLKNAND2HSV4 U17902 ( .A1(n14529), .A2(n22099), .ZN(n14605) );
  INHSV2 U17903 ( .I(\pe5/ti_7t [5]), .ZN(n14530) );
  NAND2HSV2 U17904 ( .A1(n14530), .A2(n21345), .ZN(n14632) );
  CLKAND2HSV2 U17905 ( .A1(n14632), .A2(n14497), .Z(n14680) );
  NAND2HSV0 U17906 ( .A1(\pe5/aot [11]), .A2(\pe5/bq[16] ), .ZN(n14532) );
  NAND2HSV0 U17907 ( .A1(\pe5/aot [12]), .A2(\pe5/bq[15] ), .ZN(n14531) );
  XOR2HSV0 U17908 ( .A1(n14532), .A2(n14531), .Z(n14533) );
  INHSV2 U17909 ( .I(n14766), .ZN(n23909) );
  NAND2HSV2 U17910 ( .A1(n14646), .A2(\pe5/pvq [6]), .ZN(n14538) );
  XOR2HSV0 U17911 ( .A1(n14538), .A2(\pe5/phq [6]), .Z(n14539) );
  INHSV2 U17912 ( .I(\pe5/got [12]), .ZN(n20979) );
  NOR2HSV2 U17913 ( .A1(n14583), .A2(n20979), .ZN(n14542) );
  XNOR2HSV4 U17914 ( .A1(n14543), .A2(n14542), .ZN(n14546) );
  XNOR2HSV4 U17915 ( .A1(n14546), .A2(n14545), .ZN(n14565) );
  NAND2HSV0 U17916 ( .A1(\pe5/got [14]), .A2(\pe5/got [16]), .ZN(n14548) );
  NOR2HSV1 U17917 ( .A1(n14549), .A2(n14548), .ZN(n14551) );
  NOR2HSV1 U17918 ( .A1(n14578), .A2(n21411), .ZN(n14550) );
  AOI31HSV2 U17919 ( .A1(n14552), .A2(n14551), .A3(n14573), .B(n14550), .ZN(
        n14563) );
  CLKNHSV2 U17920 ( .I(n14553), .ZN(n14554) );
  INHSV2 U17921 ( .I(n14554), .ZN(n14557) );
  CLKNHSV2 U17922 ( .I(n14555), .ZN(n14556) );
  NOR2HSV4 U17923 ( .A1(n14557), .A2(n14556), .ZN(n14580) );
  CLKNAND2HSV0 U17924 ( .A1(n14558), .A2(\pe5/got [14]), .ZN(n14560) );
  NOR2HSV4 U17925 ( .A1(n14057), .A2(n14559), .ZN(n14577) );
  NOR2HSV2 U17926 ( .A1(n14560), .A2(n14577), .ZN(n14561) );
  NAND2HSV2 U17927 ( .A1(n14563), .A2(n14562), .ZN(n14564) );
  XNOR2HSV4 U17928 ( .A1(n14565), .A2(n14564), .ZN(n14674) );
  NAND2HSV2 U17929 ( .A1(n14675), .A2(n14674), .ZN(n14567) );
  INHSV4 U17930 ( .I(n14675), .ZN(n14683) );
  CLKNHSV0 U17931 ( .I(n14680), .ZN(n14568) );
  NAND2HSV2 U17932 ( .A1(n14569), .A2(n14681), .ZN(n14570) );
  INHSV2 U17933 ( .I(n14577), .ZN(n25645) );
  CLKNHSV3 U17934 ( .I(n25645), .ZN(n14574) );
  INHSV2 U17935 ( .I(n14578), .ZN(n22093) );
  AOI21HSV4 U17936 ( .A1(n14579), .A2(n14580), .B(n22093), .ZN(n14581) );
  INAND2HSV2 U17937 ( .A1(n14766), .B1(\pe5/aot [14]), .ZN(n14584) );
  XNOR2HSV4 U17938 ( .A1(n14585), .A2(n14584), .ZN(n14588) );
  XOR2HSV0 U17939 ( .A1(n14586), .A2(\pe5/phq [7]), .Z(n14587) );
  XNOR2HSV4 U17940 ( .A1(n14588), .A2(n14587), .ZN(n14592) );
  NAND2HSV0 U17941 ( .A1(\pe5/aot [10]), .A2(\pe5/bq[16] ), .ZN(n14590) );
  BUFHSV2 U17942 ( .I(\pe5/ti_1 ), .Z(n25626) );
  INHSV2 U17943 ( .I(\pe5/got [10]), .ZN(n14643) );
  CLKNAND2HSV1 U17944 ( .A1(n25626), .A2(\pe5/got [10]), .ZN(n14589) );
  XOR2HSV0 U17945 ( .A1(n14590), .A2(n14589), .Z(n14591) );
  XNOR2HSV4 U17946 ( .A1(n14592), .A2(n14591), .ZN(n14599) );
  NAND2HSV2 U17947 ( .A1(\pe5/aot [16]), .A2(\pe5/bq[10] ), .ZN(n14650) );
  NAND2HSV0 U17948 ( .A1(n21374), .A2(\pe5/aot [11]), .ZN(n14593) );
  XOR2HSV0 U17949 ( .A1(n14650), .A2(n14593), .Z(n14597) );
  NAND2HSV0 U17950 ( .A1(\pe5/bq[13] ), .A2(\pe5/aot [13]), .ZN(n14595) );
  XNOR2HSV4 U17951 ( .A1(n14597), .A2(n14596), .ZN(n14598) );
  XNOR2HSV4 U17952 ( .A1(n14599), .A2(n14598), .ZN(n14601) );
  INHSV2 U17953 ( .I(\pe5/got [12]), .ZN(n21349) );
  NOR2HSV1 U17954 ( .A1(n14058), .A2(n21349), .ZN(n14600) );
  XOR3HSV2 U17955 ( .A1(n14602), .A2(n14601), .A3(n14600), .Z(n14603) );
  XNOR2HSV4 U17956 ( .A1(n14604), .A2(n14603), .ZN(n14608) );
  INHSV3 U17957 ( .I(n14608), .ZN(n14609) );
  CLKNHSV0 U17958 ( .I(\pe5/got [15]), .ZN(n14862) );
  INHSV2 U17959 ( .I(n14862), .ZN(n14820) );
  NOR2HSV2 U17960 ( .A1(n14820), .A2(n21412), .ZN(n14626) );
  INHSV2 U17961 ( .I(n14626), .ZN(n14614) );
  OAI21HSV2 U17962 ( .A1(n14815), .A2(\pe5/ti_7t [6]), .B(n14497), .ZN(n14617)
         );
  INHSV2 U17963 ( .I(n14617), .ZN(n25656) );
  NOR2HSV2 U17964 ( .A1(n25656), .A2(n14614), .ZN(n14615) );
  INHSV4 U17965 ( .I(n14620), .ZN(n14635) );
  CLKNAND2HSV1 U17966 ( .A1(n14621), .A2(n14620), .ZN(n14622) );
  CLKNAND2HSV4 U17967 ( .A1(n28990), .A2(n14628), .ZN(n14625) );
  NAND2HSV2 U17968 ( .A1(n20870), .A2(\pe5/ti_7t [5]), .ZN(n14624) );
  CLKNAND2HSV1 U17969 ( .A1(n25656), .A2(n14626), .ZN(n14627) );
  INHSV2 U17970 ( .I(n21422), .ZN(n14763) );
  INHSV1 U17971 ( .I(n21422), .ZN(n21345) );
  NOR2HSV2 U17972 ( .A1(n28664), .A2(n21345), .ZN(n14636) );
  INHSV2 U17973 ( .I(n14635), .ZN(n14638) );
  NOR2HSV2 U17974 ( .A1(n21412), .A2(n14045), .ZN(n14914) );
  INHSV2 U17975 ( .I(n14914), .ZN(n14924) );
  CLKAND2HSV1 U17976 ( .A1(n14632), .A2(n24635), .Z(n14633) );
  NAND2HSV0 U17977 ( .A1(n28664), .A2(n14909), .ZN(n14637) );
  CLKNHSV1 U17978 ( .I(n14637), .ZN(n14639) );
  CLKNAND2HSV1 U17979 ( .A1(n14639), .A2(n14638), .ZN(n14640) );
  NAND2HSV2 U17980 ( .A1(n14641), .A2(n14640), .ZN(n14673) );
  NAND2HSV0 U17981 ( .A1(n14852), .A2(n24411), .ZN(n14671) );
  CLKNAND2HSV1 U17982 ( .A1(n14894), .A2(n24636), .ZN(n14665) );
  NAND2HSV0 U17983 ( .A1(\pe5/aot [9]), .A2(\pe5/bq[16] ), .ZN(n14644) );
  XOR2HSV0 U17984 ( .A1(n14645), .A2(n14644), .Z(n14648) );
  XNOR2HSV1 U17985 ( .A1(n14648), .A2(n14647), .ZN(n14653) );
  CLKNAND2HSV1 U17986 ( .A1(n14031), .A2(\pe5/bq[9] ), .ZN(n14779) );
  NAND2HSV0 U17987 ( .A1(\pe5/aot [16]), .A2(\pe5/bq[9] ), .ZN(n14781) );
  OAI21HSV2 U17988 ( .A1(n14779), .A2(n14650), .B(n14649), .ZN(n14651) );
  NAND2HSV0 U17989 ( .A1(\pe5/bq[11] ), .A2(\pe5/aot [14]), .ZN(n24391) );
  XNOR2HSV1 U17990 ( .A1(n14651), .A2(n24391), .ZN(n14652) );
  XNOR2HSV4 U17991 ( .A1(n14653), .A2(n14652), .ZN(n14661) );
  NAND2HSV0 U17992 ( .A1(\pe5/aot [10]), .A2(\pe5/bq[15] ), .ZN(n14655) );
  NAND2HSV0 U17993 ( .A1(\pe5/aot [12]), .A2(\pe5/bq[13] ), .ZN(n14654) );
  XOR2HSV0 U17994 ( .A1(n14655), .A2(n14654), .Z(n14659) );
  NAND2HSV0 U17995 ( .A1(\pe5/aot [11]), .A2(\pe5/bq[14] ), .ZN(n14657) );
  NAND2HSV0 U17996 ( .A1(\pe5/aot [13]), .A2(n23909), .ZN(n14656) );
  XOR2HSV0 U17997 ( .A1(n14657), .A2(n14656), .Z(n14658) );
  XOR2HSV0 U17998 ( .A1(n14659), .A2(n14658), .Z(n14660) );
  XNOR2HSV4 U17999 ( .A1(n14661), .A2(n14660), .ZN(n14663) );
  INHSV1 U18000 ( .I(n14057), .ZN(n28594) );
  NAND2HSV0 U18001 ( .A1(n20977), .A2(n14552), .ZN(n14662) );
  XOR3HSV2 U18002 ( .A1(n14664), .A2(n14663), .A3(n14662), .Z(n14666) );
  CLKNAND2HSV1 U18003 ( .A1(n14665), .A2(n14666), .ZN(n14670) );
  CLKNHSV1 U18004 ( .I(n14665), .ZN(n14668) );
  CLKNHSV1 U18005 ( .I(n14666), .ZN(n14667) );
  CLKNAND2HSV1 U18006 ( .A1(n14668), .A2(n14667), .ZN(n14669) );
  CLKAND2HSV2 U18007 ( .A1(\pe5/ti_7t [6]), .A2(n20870), .Z(n14805) );
  INHSV1 U18008 ( .I(n14803), .ZN(n14678) );
  OAI21HSV2 U18009 ( .A1(n14675), .A2(n14674), .B(n20848), .ZN(n14802) );
  NOR2HSV2 U18010 ( .A1(n14802), .A2(n13992), .ZN(n14677) );
  OAI21HSV2 U18011 ( .A1(n14685), .A2(n14678), .B(n14677), .ZN(n14679) );
  INHSV2 U18012 ( .I(n14679), .ZN(n14682) );
  CLKNAND2HSV4 U18013 ( .A1(n14681), .A2(n14680), .ZN(n14807) );
  AOI22HSV2 U18014 ( .A1(n14820), .A2(n14805), .B1(n14682), .B2(n14807), .ZN(
        n14691) );
  NOR2HSV2 U18015 ( .A1(n14807), .A2(n14684), .ZN(n14689) );
  INHSV2 U18016 ( .I(n14685), .ZN(n14804) );
  MUX2NHSV1 U18017 ( .I0(n14630), .I1(n14683), .S(n14804), .ZN(n14687) );
  AOI21HSV2 U18018 ( .A1(n14685), .A2(n14684), .B(n21412), .ZN(n14686) );
  CLKNAND2HSV1 U18019 ( .A1(n14687), .A2(n14686), .ZN(n14688) );
  INHSV2 U18020 ( .I(n14688), .ZN(n14808) );
  CLKNAND2HSV1 U18021 ( .A1(n14689), .A2(n14808), .ZN(n14690) );
  INHSV2 U18022 ( .I(n14910), .ZN(n14693) );
  INHSV2 U18023 ( .I(n14693), .ZN(n14915) );
  NAND2HSV2 U18024 ( .A1(n14824), .A2(n14915), .ZN(n14695) );
  NAND3HSV2 U18025 ( .A1(n14760), .A2(n14759), .A3(n14758), .ZN(n28806) );
  CLKNAND2HSV2 U18026 ( .A1(n14693), .A2(n14692), .ZN(n14694) );
  CLKNAND2HSV2 U18027 ( .A1(n14695), .A2(n14694), .ZN(n28989) );
  NOR2HSV2 U18028 ( .A1(n14698), .A2(n14697), .ZN(n18857) );
  INHSV2 U18029 ( .I(n18857), .ZN(n18856) );
  BUFHSV2 U18030 ( .I(\pe6/got [14]), .Z(n22992) );
  INAND2HSV2 U18031 ( .A1(n22995), .B1(\pe6/got [11]), .ZN(n14733) );
  NAND2HSV0 U18032 ( .A1(n28793), .A2(\pe6/got [9]), .ZN(n14731) );
  CLKNAND2HSV1 U18033 ( .A1(n18930), .A2(\pe6/got [8]), .ZN(n14700) );
  NOR2HSV1 U18034 ( .A1(n24963), .A2(n14418), .ZN(n14699) );
  XNOR2HSV1 U18035 ( .A1(n14700), .A2(n14699), .ZN(n14728) );
  NAND2HSV0 U18036 ( .A1(\pe6/aot [7]), .A2(\pe6/bq[15] ), .ZN(n14702) );
  NAND2HSV0 U18037 ( .A1(\pe6/bq[8] ), .A2(\pe6/aot [14]), .ZN(n14701) );
  XOR2HSV0 U18038 ( .A1(n14702), .A2(n14701), .Z(n14706) );
  NAND2HSV0 U18039 ( .A1(\pe6/aot [13]), .A2(\pe6/bq[9] ), .ZN(n14704) );
  NAND2HSV0 U18040 ( .A1(\pe6/aot [9]), .A2(\pe6/bq[13] ), .ZN(n14703) );
  XOR2HSV0 U18041 ( .A1(n14704), .A2(n14703), .Z(n14705) );
  XOR2HSV0 U18042 ( .A1(n14706), .A2(n14705), .Z(n14714) );
  NAND2HSV0 U18043 ( .A1(\pe6/aot [8]), .A2(\pe6/bq[14] ), .ZN(n14708) );
  NAND2HSV0 U18044 ( .A1(\pe6/aot [11]), .A2(\pe6/bq[11] ), .ZN(n14707) );
  XOR2HSV0 U18045 ( .A1(n14708), .A2(n14707), .Z(n14712) );
  INHSV2 U18046 ( .I(\pe6/got [6]), .ZN(n25785) );
  CLKNAND2HSV0 U18047 ( .A1(n19021), .A2(\pe6/got [6]), .ZN(n14710) );
  NAND2HSV0 U18048 ( .A1(\pe6/aot [6]), .A2(\pe6/bq[16] ), .ZN(n14709) );
  XOR2HSV0 U18049 ( .A1(n14710), .A2(n14709), .Z(n14711) );
  XOR2HSV0 U18050 ( .A1(n14712), .A2(n14711), .Z(n14713) );
  XOR2HSV0 U18051 ( .A1(n14714), .A2(n14713), .Z(n14726) );
  CLKNAND2HSV1 U18052 ( .A1(n23498), .A2(\pe6/pvq [11]), .ZN(n14715) );
  XNOR2HSV1 U18053 ( .A1(n14715), .A2(\pe6/phq [11]), .ZN(n14720) );
  INHSV2 U18054 ( .I(\pe6/bq[6] ), .ZN(n25706) );
  CLKNAND2HSV0 U18055 ( .A1(n28680), .A2(\pe6/bq[6] ), .ZN(n18866) );
  CLKNHSV0 U18056 ( .I(\pe6/aot [16]), .ZN(n18934) );
  NAND2HSV0 U18057 ( .A1(n28680), .A2(\pe6/bq[7] ), .ZN(n14716) );
  OAI21HSV1 U18058 ( .A1(n18934), .A2(n25706), .B(n14716), .ZN(n14717) );
  OAI21HSV1 U18059 ( .A1(n14718), .A2(n18866), .B(n14717), .ZN(n14719) );
  XOR2HSV0 U18060 ( .A1(n14720), .A2(n14719), .Z(n14724) );
  NAND2HSV0 U18061 ( .A1(\pe6/aot [10]), .A2(\pe6/bq[12] ), .ZN(n14722) );
  NAND2HSV0 U18062 ( .A1(\pe6/bq[10] ), .A2(\pe6/aot [12]), .ZN(n14721) );
  XOR2HSV0 U18063 ( .A1(n14722), .A2(n14721), .Z(n14723) );
  XNOR2HSV1 U18064 ( .A1(n14724), .A2(n14723), .ZN(n14725) );
  XNOR2HSV1 U18065 ( .A1(n14726), .A2(n14725), .ZN(n14727) );
  XNOR2HSV1 U18066 ( .A1(n14728), .A2(n14727), .ZN(n14730) );
  CLKNAND2HSV1 U18067 ( .A1(\pe6/got [10]), .A2(n19109), .ZN(n14729) );
  XOR3HSV2 U18068 ( .A1(n14731), .A2(n14730), .A3(n14729), .Z(n14732) );
  XNOR2HSV1 U18069 ( .A1(n14733), .A2(n14732), .ZN(n14735) );
  NAND2HSV0 U18070 ( .A1(n28526), .A2(n28593), .ZN(n14734) );
  CLKXOR2HSV4 U18071 ( .A1(n14735), .A2(n14734), .Z(n14741) );
  NOR2HSV2 U18072 ( .A1(n14738), .A2(n18855), .ZN(n14739) );
  CLKNHSV0 U18073 ( .I(n28938), .ZN(n14742) );
  NOR2HSV2 U18074 ( .A1(n14742), .A2(n19142), .ZN(n14743) );
  NOR2HSV2 U18075 ( .A1(n28938), .A2(n19073), .ZN(n14744) );
  NOR2HSV1 U18076 ( .A1(n18852), .A2(\pe6/ti_7t [10]), .ZN(n18997) );
  INHSV2 U18077 ( .I(\pe11/pvq [1]), .ZN(n14746) );
  INHSV4 U18078 ( .I(n20164), .ZN(n20264) );
  INHSV2 U18079 ( .I(n20264), .ZN(n14747) );
  NAND4HSV4 U18080 ( .A1(n20264), .A2(n20272), .A3(\pe11/got [16]), .A4(
        \pe11/pvq [1]), .ZN(n14749) );
  CLKNHSV2 U18081 ( .I(\pe11/phq [1]), .ZN(n14752) );
  INHSV2 U18082 ( .I(ctro11), .ZN(n20551) );
  INHSV2 U18083 ( .I(n20551), .ZN(n20215) );
  CLKNAND2HSV2 U18084 ( .A1(n20181), .A2(n20623), .ZN(n20319) );
  NAND2HSV2 U18085 ( .A1(\pe11/ti_7t [1]), .A2(n20215), .ZN(n20320) );
  CLKNAND2HSV3 U18086 ( .A1(n20319), .A2(n20320), .ZN(n28629) );
  INHSV2 U18087 ( .I(\pe5/ti_7t [11]), .ZN(n14756) );
  NOR2HSV2 U18088 ( .A1(n14815), .A2(n14756), .ZN(n20868) );
  CLKNAND2HSV3 U18089 ( .A1(n14910), .A2(n14757), .ZN(n14819) );
  NOR2HSV4 U18090 ( .A1(n14819), .A2(n14762), .ZN(n14908) );
  INHSV2 U18091 ( .I(n14911), .ZN(n21465) );
  NAND2HSV4 U18092 ( .A1(n14825), .A2(n21465), .ZN(n14816) );
  CLKNAND2HSV1 U18093 ( .A1(\pe5/bq[13] ), .A2(\pe5/aot [11]), .ZN(n21358) );
  XOR2HSV0 U18094 ( .A1(n14765), .A2(n21358), .Z(n14770) );
  INAND2HSV0 U18095 ( .A1(n14766), .B1(\pe5/aot [12]), .ZN(n14768) );
  NAND2HSV0 U18096 ( .A1(\pe5/aot [14]), .A2(\pe5/bq[10] ), .ZN(n14767) );
  XOR2HSV0 U18097 ( .A1(n14768), .A2(n14767), .Z(n14769) );
  XOR2HSV0 U18098 ( .A1(n14770), .A2(n14769), .Z(n14795) );
  NAND2HSV0 U18099 ( .A1(n21374), .A2(\pe5/aot [9]), .ZN(n14772) );
  INHSV1 U18100 ( .I(\pe5/got [8]), .ZN(n24421) );
  INHSV2 U18101 ( .I(n24421), .ZN(n28632) );
  CLKNAND2HSV0 U18102 ( .A1(n25626), .A2(n28632), .ZN(n14771) );
  XOR2HSV0 U18103 ( .A1(n14772), .A2(n14771), .Z(n14776) );
  NAND2HSV0 U18104 ( .A1(\pe5/aot [10]), .A2(\pe5/bq[14] ), .ZN(n14774) );
  BUFHSV2 U18105 ( .I(\pe5/bq[16] ), .Z(n25349) );
  NAND2HSV0 U18106 ( .A1(\pe5/aot [8]), .A2(n25349), .ZN(n14773) );
  XOR2HSV0 U18107 ( .A1(n14774), .A2(n14773), .Z(n14775) );
  XNOR2HSV1 U18108 ( .A1(n14776), .A2(n14775), .ZN(n14785) );
  INHSV2 U18109 ( .I(n27052), .ZN(n23505) );
  CLKNAND2HSV0 U18110 ( .A1(n23505), .A2(\pe5/pvq [9]), .ZN(n14778) );
  XOR2HSV0 U18111 ( .A1(n14778), .A2(\pe5/phq [9]), .Z(n14783) );
  NAND2HSV0 U18112 ( .A1(n14031), .A2(\pe5/bq[8] ), .ZN(n14836) );
  INHSV2 U18113 ( .I(\pe5/bq[8] ), .ZN(n23923) );
  OAI21HSV0 U18114 ( .A1(n23789), .A2(n23923), .B(n14779), .ZN(n14780) );
  OAI21HSV1 U18115 ( .A1(n14836), .A2(n14781), .B(n14780), .ZN(n14782) );
  XOR2HSV0 U18116 ( .A1(n14783), .A2(n14782), .Z(n14784) );
  XNOR2HSV1 U18117 ( .A1(n14785), .A2(n14784), .ZN(n14794) );
  NAND2HSV0 U18118 ( .A1(n24406), .A2(n24637), .ZN(n14787) );
  CLKNAND2HSV0 U18119 ( .A1(n14787), .A2(n14788), .ZN(n14792) );
  CLKNHSV0 U18120 ( .I(n14788), .ZN(n14789) );
  NAND2HSV2 U18121 ( .A1(n14792), .A2(n14791), .ZN(n14793) );
  XOR3HSV2 U18122 ( .A1(n14795), .A2(n14794), .A3(n14793), .Z(n14797) );
  CLKNAND2HSV1 U18123 ( .A1(n14848), .A2(n20977), .ZN(n14796) );
  NAND2HSV0 U18124 ( .A1(n28664), .A2(n24636), .ZN(n14798) );
  XNOR2HSV4 U18125 ( .A1(n14801), .A2(n14800), .ZN(n14811) );
  AOI21HSV0 U18126 ( .A1(n14804), .A2(n14803), .B(n14802), .ZN(n14806) );
  INHSV2 U18127 ( .I(n14807), .ZN(n14809) );
  XNOR2HSV4 U18128 ( .A1(n14811), .A2(n14810), .ZN(n14812) );
  XNOR2HSV4 U18129 ( .A1(n14813), .A2(n14812), .ZN(n14863) );
  NAND3HSV3 U18130 ( .A1(n14864), .A2(n14863), .A3(n14628), .ZN(n14814) );
  INHSV4 U18131 ( .I(n14814), .ZN(n14928) );
  INHSV2 U18132 ( .I(n14865), .ZN(n14817) );
  OAI21HSV4 U18133 ( .A1(n14818), .A2(n14863), .B(n14817), .ZN(n14927) );
  NOR2HSV4 U18134 ( .A1(n14928), .A2(n14927), .ZN(n20978) );
  INHSV2 U18135 ( .I(n14819), .ZN(n14822) );
  CLKNAND2HSV1 U18136 ( .A1(n14965), .A2(n14820), .ZN(n14821) );
  IOA21HSV4 U18137 ( .A1(n14825), .A2(n14824), .B(n14823), .ZN(n14857) );
  INHSV2 U18138 ( .I(n14857), .ZN(n14856) );
  NAND2HSV2 U18139 ( .A1(n28806), .A2(n24635), .ZN(n14854) );
  NAND2HSV0 U18140 ( .A1(\pe5/bq[9] ), .A2(\pe5/aot [14]), .ZN(n14827) );
  NAND2HSV0 U18141 ( .A1(\pe5/aot [10]), .A2(\pe5/bq[13] ), .ZN(n14826) );
  XOR2HSV0 U18142 ( .A1(n14827), .A2(n14826), .Z(n14847) );
  NAND2HSV0 U18143 ( .A1(\pe5/aot [12]), .A2(\pe5/bq[11] ), .ZN(n14829) );
  BUFHSV4 U18144 ( .I(\pe5/got [7]), .Z(n28645) );
  NAND2HSV0 U18145 ( .A1(n28645), .A2(n25626), .ZN(n14828) );
  XOR2HSV0 U18146 ( .A1(n14829), .A2(n14828), .Z(n14832) );
  CLKNAND2HSV0 U18147 ( .A1(n23505), .A2(\pe5/pvq [10]), .ZN(n14830) );
  XOR2HSV0 U18148 ( .A1(n14830), .A2(\pe5/phq [10]), .Z(n14831) );
  XOR2HSV0 U18149 ( .A1(n14832), .A2(n14831), .Z(n14846) );
  CLKNAND2HSV0 U18150 ( .A1(\pe5/aot [9]), .A2(\pe5/bq[7] ), .ZN(n24651) );
  CLKNHSV0 U18151 ( .I(\pe5/aot [9]), .ZN(n21493) );
  CLKNHSV0 U18152 ( .I(\pe5/bq[14] ), .ZN(n20889) );
  CLKNHSV0 U18153 ( .I(\pe5/aot [16]), .ZN(n14833) );
  INHSV2 U18154 ( .I(n14833), .ZN(n21488) );
  CLKNAND2HSV1 U18155 ( .A1(n21488), .A2(\pe5/bq[7] ), .ZN(n14885) );
  OAI21HSV1 U18156 ( .A1(n21493), .A2(n20889), .B(n14885), .ZN(n14834) );
  OAI21HSV0 U18157 ( .A1(n24651), .A2(n14835), .B(n14834), .ZN(n14837) );
  XNOR2HSV1 U18158 ( .A1(n14837), .A2(n14836), .ZN(n14845) );
  NAND2HSV0 U18159 ( .A1(\pe5/aot [11]), .A2(n23909), .ZN(n14839) );
  BUFHSV2 U18160 ( .I(n21374), .Z(n24647) );
  NAND2HSV0 U18161 ( .A1(\pe5/aot [8]), .A2(n24647), .ZN(n14838) );
  XOR2HSV0 U18162 ( .A1(n14839), .A2(n14838), .Z(n14843) );
  NAND2HSV0 U18163 ( .A1(n25349), .A2(\pe5/aot [7]), .ZN(n14841) );
  NAND2HSV0 U18164 ( .A1(\pe5/aot [13]), .A2(\pe5/bq[10] ), .ZN(n14840) );
  XOR2HSV0 U18165 ( .A1(n14841), .A2(n14840), .Z(n14842) );
  XOR2HSV2 U18166 ( .A1(n14843), .A2(n14842), .Z(n14844) );
  XOR4HSV1 U18167 ( .A1(n14847), .A2(n14846), .A3(n14845), .A4(n14844), .Z(
        n14850) );
  INHSV2 U18168 ( .I(\pe5/got [8]), .ZN(n24683) );
  NAND2HSV0 U18169 ( .A1(n28664), .A2(n20977), .ZN(n14851) );
  XNOR2HSV4 U18170 ( .A1(n14854), .A2(n14853), .ZN(n14858) );
  CLKNHSV3 U18171 ( .I(n14858), .ZN(n14855) );
  CLKNAND2HSV3 U18172 ( .A1(n14856), .A2(n14855), .ZN(n14860) );
  CLKNAND2HSV1 U18173 ( .A1(n14858), .A2(n14857), .ZN(n14859) );
  CLKXOR2HSV4 U18174 ( .A1(n20978), .A2(n14930), .Z(n14861) );
  NAND2HSV2 U18175 ( .A1(n20987), .A2(n14045), .ZN(n20855) );
  AOI21HSV4 U18176 ( .A1(n14861), .A2(n20848), .B(n20855), .ZN(n14923) );
  NOR2HSV0 U18177 ( .A1(n14535), .A2(n14931), .ZN(n14901) );
  NAND2HSV0 U18178 ( .A1(n24340), .A2(n24406), .ZN(n14867) );
  XNOR2HSV1 U18179 ( .A1(n14867), .A2(n14866), .ZN(n14893) );
  BUFHSV4 U18180 ( .I(\pe5/got [6]), .Z(n28647) );
  NAND2HSV0 U18181 ( .A1(n25626), .A2(n28647), .ZN(n14869) );
  NAND2HSV0 U18182 ( .A1(\pe5/aot [9]), .A2(\pe5/bq[13] ), .ZN(n14868) );
  XOR2HSV0 U18183 ( .A1(n14869), .A2(n14868), .Z(n14873) );
  NAND2HSV0 U18184 ( .A1(\pe5/aot [8]), .A2(\pe5/bq[14] ), .ZN(n14871) );
  NAND2HSV0 U18185 ( .A1(\pe5/bq[8] ), .A2(\pe5/aot [14]), .ZN(n14870) );
  XOR2HSV0 U18186 ( .A1(n14871), .A2(n14870), .Z(n14872) );
  XOR2HSV0 U18187 ( .A1(n14873), .A2(n14872), .Z(n14881) );
  NAND2HSV0 U18188 ( .A1(n21374), .A2(\pe5/aot [7]), .ZN(n14875) );
  NAND2HSV0 U18189 ( .A1(\pe5/aot [6]), .A2(n25349), .ZN(n14874) );
  XOR2HSV0 U18190 ( .A1(n14875), .A2(n14874), .Z(n14879) );
  NAND2HSV0 U18191 ( .A1(\pe5/aot [11]), .A2(\pe5/bq[11] ), .ZN(n14877) );
  NAND2HSV0 U18192 ( .A1(\pe5/aot [12]), .A2(\pe5/bq[10] ), .ZN(n14876) );
  XOR2HSV0 U18193 ( .A1(n14877), .A2(n14876), .Z(n14878) );
  XOR2HSV0 U18194 ( .A1(n14879), .A2(n14878), .Z(n14880) );
  XOR2HSV0 U18195 ( .A1(n14881), .A2(n14880), .Z(n14891) );
  CLKNAND2HSV0 U18196 ( .A1(n23505), .A2(\pe5/pvq [11]), .ZN(n14882) );
  XOR2HSV0 U18197 ( .A1(n14882), .A2(\pe5/phq [11]), .Z(n14887) );
  NAND2HSV0 U18198 ( .A1(n14031), .A2(\pe5/bq[6] ), .ZN(n14954) );
  CLKNHSV0 U18199 ( .I(\pe5/bq[7] ), .ZN(n23504) );
  CLKNAND2HSV1 U18200 ( .A1(n21488), .A2(\pe5/bq[6] ), .ZN(n14955) );
  OAI21HSV0 U18201 ( .A1(n23504), .A2(n14883), .B(n14955), .ZN(n14884) );
  OAI21HSV1 U18202 ( .A1(n14954), .A2(n14885), .B(n14884), .ZN(n14886) );
  XNOR2HSV1 U18203 ( .A1(n14887), .A2(n14886), .ZN(n14889) );
  CLKNHSV0 U18204 ( .I(\pe5/aot [13]), .ZN(n14956) );
  INHSV2 U18205 ( .I(\pe5/bq[9] ), .ZN(n27049) );
  NOR2HSV2 U18206 ( .A1(n14956), .A2(n27049), .ZN(n24388) );
  INAND2HSV0 U18207 ( .A1(n14766), .B1(\pe5/aot [10]), .ZN(n14951) );
  XOR2HSV0 U18208 ( .A1(n24388), .A2(n14951), .Z(n14888) );
  XNOR2HSV1 U18209 ( .A1(n14889), .A2(n14888), .ZN(n14890) );
  XNOR2HSV1 U18210 ( .A1(n14891), .A2(n14890), .ZN(n14892) );
  XNOR2HSV1 U18211 ( .A1(n14893), .A2(n14892), .ZN(n14897) );
  CLKNHSV0 U18212 ( .I(n14894), .ZN(n14895) );
  INHSV2 U18213 ( .I(n14895), .ZN(n28614) );
  NAND2HSV0 U18214 ( .A1(n28614), .A2(n14069), .ZN(n14896) );
  XNOR2HSV1 U18215 ( .A1(n14897), .A2(n14896), .ZN(n14899) );
  INHSV2 U18216 ( .I(n14630), .ZN(n24674) );
  XNOR2HSV1 U18217 ( .A1(n14899), .A2(n14898), .ZN(n14900) );
  NOR2HSV2 U18218 ( .A1(n21325), .A2(n21349), .ZN(n14903) );
  XNOR2HSV1 U18219 ( .A1(n14904), .A2(n14903), .ZN(n14907) );
  CLKBUFHSV4 U18220 ( .I(n14905), .Z(n24378) );
  XNOR2HSV4 U18221 ( .A1(n14907), .A2(n14906), .ZN(n14920) );
  CLKNHSV0 U18222 ( .I(n14908), .ZN(n14918) );
  INHSV2 U18223 ( .I(n14909), .ZN(n14925) );
  NOR2HSV0 U18224 ( .A1(n14910), .A2(n14925), .ZN(n14912) );
  CLKNAND2HSV1 U18225 ( .A1(n14912), .A2(n21523), .ZN(n14917) );
  NAND2HSV0 U18226 ( .A1(n14965), .A2(n24635), .ZN(n14913) );
  AOI21HSV2 U18227 ( .A1(n14915), .A2(n14914), .B(n14913), .ZN(n14916) );
  XNOR2HSV4 U18228 ( .A1(n14920), .A2(n14919), .ZN(n14921) );
  XNOR2HSV4 U18229 ( .A1(n14922), .A2(n14921), .ZN(n20860) );
  NOR2HSV2 U18230 ( .A1(n14930), .A2(n14924), .ZN(n20917) );
  NAND2HSV2 U18231 ( .A1(n14930), .A2(n14926), .ZN(n14929) );
  NOR2HSV4 U18232 ( .A1(n14928), .A2(n14927), .ZN(n20983) );
  NOR2HSV2 U18233 ( .A1(n14929), .A2(n20983), .ZN(n20920) );
  CLKBUFHSV4 U18234 ( .I(n14930), .Z(n20985) );
  INHSV1 U18235 ( .I(n14931), .ZN(n21352) );
  INHSV2 U18236 ( .I(n21352), .ZN(n20931) );
  INHSV2 U18237 ( .I(\pe5/got [10]), .ZN(n21510) );
  NOR2HSV4 U18238 ( .A1(n20931), .A2(n21510), .ZN(n14962) );
  NAND2HSV0 U18239 ( .A1(n28645), .A2(n28594), .ZN(n14933) );
  CLKNAND2HSV0 U18240 ( .A1(\pe5/aot [6]), .A2(n24647), .ZN(n14935) );
  NAND2HSV0 U18241 ( .A1(\pe5/aot [8]), .A2(\pe5/bq[13] ), .ZN(n14934) );
  XOR2HSV0 U18242 ( .A1(n14935), .A2(n14934), .Z(n14939) );
  NAND2HSV0 U18243 ( .A1(\pe5/bq[7] ), .A2(\pe5/aot [14]), .ZN(n14937) );
  NAND2HSV0 U18244 ( .A1(\pe5/aot [12]), .A2(\pe5/bq[9] ), .ZN(n14936) );
  XOR2HSV0 U18245 ( .A1(n14937), .A2(n14936), .Z(n14938) );
  XOR2HSV0 U18246 ( .A1(n14939), .A2(n14938), .Z(n14947) );
  NAND2HSV0 U18247 ( .A1(\pe5/aot [11]), .A2(\pe5/bq[10] ), .ZN(n14941) );
  NAND2HSV0 U18248 ( .A1(\pe5/aot [5]), .A2(\pe5/bq[16] ), .ZN(n14940) );
  XOR2HSV0 U18249 ( .A1(n14941), .A2(n14940), .Z(n14945) );
  NAND2HSV0 U18250 ( .A1(\pe5/aot [7]), .A2(\pe5/bq[14] ), .ZN(n14943) );
  XOR2HSV0 U18251 ( .A1(n14943), .A2(n14942), .Z(n14944) );
  XOR2HSV0 U18252 ( .A1(n14945), .A2(n14944), .Z(n14946) );
  CLKBUFHSV4 U18253 ( .I(n23505), .Z(n28682) );
  CLKNAND2HSV0 U18254 ( .A1(n28682), .A2(\pe5/pvq [12]), .ZN(n14948) );
  XNOR2HSV1 U18255 ( .A1(n14948), .A2(\pe5/phq [12]), .ZN(n14953) );
  NAND2HSV0 U18256 ( .A1(\pe5/aot [9]), .A2(\pe5/bq[11] ), .ZN(n20881) );
  NAND2HSV0 U18257 ( .A1(\pe5/aot [10]), .A2(\pe5/bq[11] ), .ZN(n14949) );
  OAI21HSV0 U18258 ( .A1(n21493), .A2(n14766), .B(n14949), .ZN(n14950) );
  OAI21HSV1 U18259 ( .A1(n20881), .A2(n14951), .B(n14950), .ZN(n14952) );
  XOR2HSV0 U18260 ( .A1(n14953), .A2(n14952), .Z(n14958) );
  CLKNAND2HSV0 U18261 ( .A1(n14031), .A2(\pe5/bq[5] ), .ZN(n21470) );
  NAND2HSV0 U18262 ( .A1(n24674), .A2(n14071), .ZN(n14959) );
  XNOR2HSV1 U18263 ( .A1(n14960), .A2(n14959), .ZN(n14961) );
  XNOR2HSV4 U18264 ( .A1(n14962), .A2(n14961), .ZN(n14964) );
  INHSV2 U18265 ( .I(n21325), .ZN(n21504) );
  XOR2HSV2 U18266 ( .A1(n14964), .A2(n14963), .Z(n14970) );
  NAND2HSV1 U18267 ( .A1(n24378), .A2(n24636), .ZN(n14969) );
  CLKNHSV0 U18268 ( .I(n14965), .ZN(n14966) );
  NOR2HSV2 U18269 ( .A1(n14966), .A2(n20869), .ZN(n14967) );
  OAI21HSV4 U18270 ( .A1(n28989), .A2(n14763), .B(n14967), .ZN(n14968) );
  INHSV4 U18271 ( .I(\pe1/aot [16]), .ZN(n17373) );
  INHSV4 U18272 ( .I(\pe1/bq[15] ), .ZN(n14979) );
  INHSV2 U18273 ( .I(\pe1/bq[15] ), .ZN(n14971) );
  NOR2HSV4 U18274 ( .A1(n17373), .A2(n14971), .ZN(n14974) );
  CLKXOR2HSV4 U18275 ( .A1(n14974), .A2(n14975), .Z(n16197) );
  INHSV4 U18276 ( .I(ctro1), .ZN(n16184) );
  NOR2HSV2 U18277 ( .A1(n16185), .A2(\pe1/got [16]), .ZN(n16198) );
  INHSV3 U18278 ( .I(n16197), .ZN(n16201) );
  INHSV2 U18279 ( .I(\pe1/got [16]), .ZN(n14972) );
  NOR2HSV2 U18280 ( .A1(n16284), .A2(ctro1), .ZN(n17602) );
  INHSV4 U18281 ( .I(\pe1/bq[16] ), .ZN(n14990) );
  NOR2HSV8 U18282 ( .A1(n17373), .A2(n14990), .ZN(n29052) );
  NAND2HSV0 U18283 ( .A1(n17602), .A2(n29052), .ZN(n14973) );
  INHSV2 U18284 ( .I(n14973), .ZN(n16200) );
  BUFHSV4 U18285 ( .I(n16184), .Z(n17359) );
  IOA21HSV4 U18286 ( .A1(\pe1/ti_7t [2]), .A2(n17531), .B(n14976), .ZN(n16199)
         );
  AOI21HSV4 U18287 ( .A1(n16201), .A2(n16200), .B(n16199), .ZN(n14977) );
  IOA21HSV4 U18288 ( .A1(n16197), .A2(n16198), .B(n14977), .ZN(n26444) );
  INHSV4 U18289 ( .I(n26444), .ZN(n16211) );
  INHSV4 U18290 ( .I(n16211), .ZN(n28814) );
  INHSV4 U18291 ( .I(\pe1/got [16]), .ZN(n16284) );
  INHSV4 U18292 ( .I(n16284), .ZN(n17617) );
  CLKNAND2HSV3 U18293 ( .A1(n28814), .A2(n17617), .ZN(n15000) );
  NOR2HSV4 U18294 ( .A1(n14978), .A2(n26536), .ZN(n14981) );
  NAND2HSV2 U18295 ( .A1(n28468), .A2(n26431), .ZN(n16216) );
  CLKNHSV0 U18296 ( .I(\pe1/ti_7t [1]), .ZN(n14980) );
  NAND2HSV0 U18297 ( .A1(n14980), .A2(ctro1), .ZN(n14985) );
  NAND3HSV2 U18298 ( .A1(n14981), .A2(n16216), .A3(n14985), .ZN(n14984) );
  INHSV1 U18299 ( .I(n16216), .ZN(n14987) );
  INHSV2 U18300 ( .I(n14981), .ZN(n14982) );
  CLKNAND2HSV2 U18301 ( .A1(n14984), .A2(n14983), .ZN(n14989) );
  CLKNHSV1 U18302 ( .I(n14985), .ZN(n14986) );
  CLKAND2HSV2 U18303 ( .A1(n14987), .A2(n14986), .Z(n14988) );
  NOR2HSV4 U18304 ( .A1(n14989), .A2(n14988), .ZN(n14998) );
  CLKNHSV1 U18305 ( .I(n14990), .ZN(n14991) );
  NAND2HSV0 U18306 ( .A1(\pe1/bq[14] ), .A2(\pe1/aot [16]), .ZN(n14993) );
  CLKNHSV2 U18307 ( .I(n14992), .ZN(n14995) );
  CLKNHSV2 U18308 ( .I(n14993), .ZN(n14994) );
  NAND2HSV4 U18309 ( .A1(n14995), .A2(n14994), .ZN(n14996) );
  NAND2HSV4 U18310 ( .A1(n14997), .A2(n14996), .ZN(n16214) );
  XNOR2HSV4 U18311 ( .A1(n14998), .A2(n16214), .ZN(n15001) );
  INHSV3 U18312 ( .I(n15001), .ZN(n14999) );
  CLKNAND2HSV3 U18313 ( .A1(n15000), .A2(n14999), .ZN(n15003) );
  NOR2HSV2 U18314 ( .A1(n23345), .A2(\pe3/phq [1]), .ZN(n15005) );
  NOR2HSV4 U18315 ( .A1(n15006), .A2(n15005), .ZN(n15014) );
  NAND2HSV0 U18316 ( .A1(\pe3/ti_1 ), .A2(\pe3/got [16]), .ZN(n15010) );
  INHSV3 U18317 ( .I(\pe3/got [16]), .ZN(n16042) );
  NOR2HSV2 U18318 ( .A1(n16042), .A2(n15007), .ZN(n15009) );
  MUX2NHSV2 U18319 ( .I0(n15010), .I1(n15009), .S(n15008), .ZN(n15013) );
  INHSV2 U18320 ( .I(n15013), .ZN(n15011) );
  NAND2HSV2 U18321 ( .A1(n15014), .A2(n15013), .ZN(n15015) );
  INHSV2 U18322 ( .I(n15089), .ZN(n24312) );
  INHSV2 U18323 ( .I(n26240), .ZN(n16166) );
  INHSV2 U18324 ( .I(n15161), .ZN(n15019) );
  INHSV2 U18325 ( .I(\pe3/bq[16] ), .ZN(n15062) );
  CLKNAND2HSV1 U18326 ( .A1(n15019), .A2(n15018), .ZN(n15021) );
  CLKBUFHSV4 U18327 ( .I(\pe3/bq[16] ), .Z(n23336) );
  NAND3HSV2 U18328 ( .A1(n15161), .A2(n23336), .A3(\pe3/aot [14]), .ZN(n15020)
         );
  NAND2HSV2 U18329 ( .A1(n15021), .A2(n15020), .ZN(n15028) );
  INHSV4 U18330 ( .I(\pe3/got [14]), .ZN(n15301) );
  AOI21HSV2 U18331 ( .A1(n15044), .A2(n15086), .B(\pe3/phq [3]), .ZN(n15024)
         );
  NAND2HSV2 U18332 ( .A1(\pe3/ti_1 ), .A2(\pe3/phq [3]), .ZN(n15022) );
  NOR2HSV2 U18333 ( .A1(n15301), .A2(n15022), .ZN(n15023) );
  NOR2HSV4 U18334 ( .A1(n15024), .A2(n15023), .ZN(n15027) );
  INHSV2 U18335 ( .I(n15027), .ZN(n15025) );
  NAND2HSV2 U18336 ( .A1(n15028), .A2(n15027), .ZN(n15029) );
  NAND2HSV2 U18337 ( .A1(n21335), .A2(\pe3/pvq [3]), .ZN(n15032) );
  NAND2HSV0 U18338 ( .A1(\pe3/aot [15]), .A2(\pe3/bq[15] ), .ZN(n15031) );
  XNOR2HSV1 U18339 ( .A1(n15032), .A2(n15031), .ZN(n15033) );
  XNOR2HSV4 U18340 ( .A1(n15034), .A2(n15033), .ZN(n15093) );
  CLKNAND2HSV0 U18341 ( .A1(n15035), .A2(n15093), .ZN(n15039) );
  INHSV2 U18342 ( .I(n15035), .ZN(n15037) );
  NAND2HSV2 U18343 ( .A1(n15039), .A2(n15038), .ZN(n15055) );
  INHSV2 U18344 ( .I(\pe3/phq [2]), .ZN(n15040) );
  CLKNAND2HSV2 U18345 ( .A1(n23345), .A2(\pe3/pvq [2]), .ZN(n15042) );
  XNOR2HSV4 U18346 ( .A1(n15043), .A2(n15042), .ZN(n15051) );
  CLKBUFHSV4 U18347 ( .I(\pe3/got [15]), .Z(n15157) );
  NAND2HSV2 U18348 ( .A1(n15044), .A2(n15157), .ZN(n15048) );
  CLKNHSV1 U18349 ( .I(n15048), .ZN(n15046) );
  NAND2HSV2 U18350 ( .A1(\pe3/bq[16] ), .A2(\pe3/aot [15]), .ZN(n15047) );
  CLKNHSV1 U18351 ( .I(n15047), .ZN(n15045) );
  CLKNAND2HSV1 U18352 ( .A1(n15046), .A2(n15045), .ZN(n15050) );
  CLKNAND2HSV1 U18353 ( .A1(n15048), .A2(n15047), .ZN(n15049) );
  INHSV4 U18354 ( .I(ctro3), .ZN(n15060) );
  BUFHSV8 U18355 ( .I(n15060), .Z(n15056) );
  BUFHSV8 U18356 ( .I(n15056), .Z(n15057) );
  INHSV2 U18357 ( .I(n15191), .ZN(n15238) );
  BUFHSV8 U18358 ( .I(n15057), .Z(n15191) );
  INHSV2 U18359 ( .I(\pe3/got [16]), .ZN(n28929) );
  NAND2HSV2 U18360 ( .A1(n15057), .A2(n15176), .ZN(n15052) );
  CLKNHSV3 U18361 ( .I(n15052), .ZN(n15285) );
  CLKAND2HSV2 U18362 ( .A1(n15089), .A2(n15285), .Z(n15053) );
  CLKNAND2HSV3 U18363 ( .A1(n15054), .A2(n15097), .ZN(n28677) );
  XNOR2HSV4 U18364 ( .A1(n15055), .A2(n28677), .ZN(n15059) );
  BUFHSV2 U18365 ( .I(n15056), .Z(n23372) );
  BUFHSV2 U18366 ( .I(n23372), .Z(n23666) );
  OAI21HSV2 U18367 ( .A1(n15191), .A2(\pe3/ti_7t [3]), .B(n15176), .ZN(n15058)
         );
  AOI21HSV4 U18368 ( .A1(n15059), .A2(n23666), .B(n15058), .ZN(n15080) );
  CLKBUFHSV4 U18369 ( .I(n15060), .Z(n15963) );
  CLKNAND2HSV2 U18370 ( .A1(n15089), .A2(n15333), .ZN(n15061) );
  CLKBUFHSV4 U18371 ( .I(n15973), .Z(n15189) );
  INHSV4 U18372 ( .I(n15189), .ZN(n16159) );
  INHSV3 U18373 ( .I(n15062), .ZN(n26351) );
  NAND2HSV2 U18374 ( .A1(\pe3/aot [13]), .A2(n26351), .ZN(n15064) );
  NAND2HSV0 U18375 ( .A1(\pe3/aot [16]), .A2(\pe3/bq[13] ), .ZN(n15063) );
  CLKXOR2HSV2 U18376 ( .A1(n15064), .A2(n15063), .Z(n15071) );
  BUFHSV2 U18377 ( .I(\pe3/ctrq ), .Z(n23516) );
  NAND2HSV2 U18378 ( .A1(\pe3/aot [15]), .A2(\pe3/bq[14] ), .ZN(n15066) );
  CLKNHSV0 U18379 ( .I(\pe3/pvq [4]), .ZN(n15065) );
  NOR2HSV1 U18380 ( .A1(n15066), .A2(n15065), .ZN(n15069) );
  BUFHSV2 U18381 ( .I(\pe3/ctrq ), .Z(n23541) );
  INHSV2 U18382 ( .I(n15066), .ZN(n15067) );
  AOI21HSV2 U18383 ( .A1(n23541), .A2(\pe3/pvq [4]), .B(n15067), .ZN(n15068)
         );
  AOI21HSV2 U18384 ( .A1(n23516), .A2(n15069), .B(n15068), .ZN(n15070) );
  NOR2HSV2 U18385 ( .A1(n24313), .A2(n15162), .ZN(n15072) );
  NAND2HSV2 U18386 ( .A1(n28677), .A2(n15157), .ZN(n15075) );
  NAND2HSV2 U18387 ( .A1(n15074), .A2(n15075), .ZN(n15079) );
  INHSV2 U18388 ( .I(n15075), .ZN(n15076) );
  NAND2HSV4 U18389 ( .A1(n15077), .A2(n15076), .ZN(n15078) );
  CLKNAND2HSV3 U18390 ( .A1(n15079), .A2(n15078), .ZN(n15081) );
  CLKNAND2HSV2 U18391 ( .A1(n15080), .A2(n15081), .ZN(n15085) );
  INHSV2 U18392 ( .I(n15080), .ZN(n15083) );
  INHSV2 U18393 ( .I(n15081), .ZN(n15082) );
  NAND2HSV2 U18394 ( .A1(\pe3/ti_7t [4]), .A2(n15238), .ZN(n15146) );
  INHSV4 U18395 ( .I(n15963), .ZN(n21720) );
  INHSV2 U18396 ( .I(n15086), .ZN(n23383) );
  AO21HSV1 U18397 ( .A1(n15146), .A2(n21720), .B(n23383), .Z(n15087) );
  NOR2HSV2 U18398 ( .A1(n15088), .A2(n15087), .ZN(n15125) );
  NOR2HSV2 U18399 ( .A1(n15089), .A2(n16163), .ZN(n15091) );
  OAI21HSV2 U18400 ( .A1(n15973), .A2(\pe3/ti_7t [1]), .B(n15157), .ZN(n15090)
         );
  NOR2HSV4 U18401 ( .A1(n15091), .A2(n15090), .ZN(n15092) );
  XNOR2HSV4 U18402 ( .A1(n15093), .A2(n15092), .ZN(n25636) );
  NOR2HSV2 U18403 ( .A1(n15095), .A2(n15094), .ZN(n15099) );
  CLKNAND2HSV1 U18404 ( .A1(n15097), .A2(n15333), .ZN(n15098) );
  NOR2HSV2 U18405 ( .A1(n15099), .A2(n15098), .ZN(n15100) );
  CLKNAND2HSV2 U18406 ( .A1(n25636), .A2(n15100), .ZN(n15102) );
  NAND2HSV2 U18407 ( .A1(n21720), .A2(\pe3/ti_7t [3]), .ZN(n15101) );
  BUFHSV2 U18408 ( .I(n15160), .Z(n15272) );
  NOR2HSV3 U18409 ( .A1(n15272), .A2(n24313), .ZN(n15123) );
  NAND2HSV0 U18410 ( .A1(\pe3/got [10]), .A2(n26380), .ZN(n15104) );
  NAND2HSV0 U18411 ( .A1(\pe3/aot [11]), .A2(\pe3/bq[15] ), .ZN(n15103) );
  XOR2HSV0 U18412 ( .A1(n15104), .A2(n15103), .Z(n15117) );
  BUFHSV4 U18413 ( .I(\pe3/ctrq ), .Z(n21335) );
  CLKNAND2HSV1 U18414 ( .A1(\pe3/aot [14]), .A2(\pe3/bq[12] ), .ZN(n26243) );
  NAND2HSV0 U18415 ( .A1(\pe3/aot [12]), .A2(\pe3/bq[14] ), .ZN(n26310) );
  NAND2HSV2 U18416 ( .A1(\pe3/aot [14]), .A2(\pe3/bq[14] ), .ZN(n15135) );
  CLKNAND2HSV2 U18417 ( .A1(\pe3/aot [12]), .A2(\pe3/bq[12] ), .ZN(n16080) );
  NOR2HSV2 U18418 ( .A1(n15135), .A2(n16080), .ZN(n15105) );
  AOI21HSV2 U18419 ( .A1(n26243), .A2(n26310), .B(n15105), .ZN(n15106) );
  NAND2HSV0 U18420 ( .A1(\pe3/aot [15]), .A2(\pe3/bq[11] ), .ZN(n15109) );
  NAND2HSV0 U18421 ( .A1(\pe3/aot [13]), .A2(\pe3/bq[13] ), .ZN(n15111) );
  XOR2HSV0 U18422 ( .A1(n15112), .A2(n15111), .Z(n15113) );
  XOR2HSV0 U18423 ( .A1(n15114), .A2(n15113), .Z(n15115) );
  XOR3HSV2 U18424 ( .A1(n15117), .A2(n15116), .A3(n15115), .Z(n15121) );
  INHSV2 U18425 ( .I(n15118), .ZN(n15140) );
  INHSV4 U18426 ( .I(n23480), .ZN(n15223) );
  NAND2HSV2 U18427 ( .A1(n26255), .A2(\pe3/got [11]), .ZN(n15120) );
  INHSV4 U18428 ( .I(n28677), .ZN(n15302) );
  INHSV3 U18429 ( .I(n15302), .ZN(n15979) );
  NAND2HSV0 U18430 ( .A1(n15979), .A2(n15245), .ZN(n15119) );
  XOR3HSV2 U18431 ( .A1(n15121), .A2(n15120), .A3(n15119), .Z(n15122) );
  XNOR2HSV4 U18432 ( .A1(n15123), .A2(n15122), .ZN(n15124) );
  XNOR2HSV4 U18433 ( .A1(n15125), .A2(n15124), .ZN(n15155) );
  NAND2HSV2 U18434 ( .A1(n29037), .A2(n15242), .ZN(n15126) );
  INHSV4 U18435 ( .I(n15127), .ZN(n15178) );
  INHSV2 U18436 ( .I(\pe3/got [12]), .ZN(n26241) );
  NAND2HSV0 U18437 ( .A1(\pe3/aot [12]), .A2(n23336), .ZN(n15128) );
  XOR2HSV0 U18438 ( .A1(n15128), .A2(n15129), .Z(n15131) );
  XOR2HSV0 U18439 ( .A1(n15131), .A2(n15130), .Z(n15139) );
  INHSV1 U18440 ( .I(\pe3/aot [15]), .ZN(n16066) );
  NOR2HSV2 U18441 ( .A1(n16066), .A2(n26246), .ZN(n15133) );
  NAND2HSV0 U18442 ( .A1(n28465), .A2(\pe3/bq[12] ), .ZN(n15132) );
  XOR2HSV0 U18443 ( .A1(n15133), .A2(n15132), .Z(n15137) );
  NAND2HSV0 U18444 ( .A1(\pe3/aot [13]), .A2(\pe3/bq[15] ), .ZN(n15134) );
  XOR2HSV0 U18445 ( .A1(n15134), .A2(n15135), .Z(n15136) );
  XOR2HSV0 U18446 ( .A1(n15137), .A2(n15136), .Z(n15138) );
  NAND2HSV2 U18447 ( .A1(n23480), .A2(n28628), .ZN(n15141) );
  NOR2HSV2 U18448 ( .A1(n15302), .A2(n23383), .ZN(n15142) );
  XNOR2HSV4 U18449 ( .A1(n15143), .A2(n15142), .ZN(n15150) );
  AOI21HSV4 U18450 ( .A1(n15145), .A2(n25635), .B(n15144), .ZN(n15226) );
  NOR2HSV4 U18451 ( .A1(n15226), .A2(n16166), .ZN(n15149) );
  XNOR2HSV4 U18452 ( .A1(n15150), .A2(n15149), .ZN(n15239) );
  CLKNAND2HSV4 U18453 ( .A1(n15178), .A2(n15239), .ZN(n27117) );
  INHSV2 U18454 ( .I(\pe3/got [15]), .ZN(n23402) );
  AND2HSV2 U18455 ( .A1(n15202), .A2(n26240), .Z(n15154) );
  CLKNAND2HSV2 U18456 ( .A1(n27117), .A2(n15154), .ZN(n15152) );
  NOR2HSV1 U18457 ( .A1(n16164), .A2(n16031), .ZN(n15148) );
  NAND2HSV2 U18458 ( .A1(n15241), .A2(n15148), .ZN(n15151) );
  XNOR2HSV4 U18459 ( .A1(n15150), .A2(n15149), .ZN(n15181) );
  INHSV4 U18460 ( .I(n15181), .ZN(n15243) );
  NOR2HSV4 U18461 ( .A1(n15151), .A2(n15181), .ZN(n15205) );
  NOR2HSV2 U18462 ( .A1(n15152), .A2(n15205), .ZN(n15153) );
  INAND2HSV4 U18463 ( .A1(n15155), .B1(n15153), .ZN(n15288) );
  INHSV4 U18464 ( .I(n15288), .ZN(n15188) );
  CLKNAND2HSV2 U18465 ( .A1(n27117), .A2(n15154), .ZN(n15156) );
  OAI21HSV4 U18466 ( .A1(n15156), .A2(n15205), .B(n15155), .ZN(n15284) );
  INHSV1 U18467 ( .I(\pe3/ti_7t [4]), .ZN(n15158) );
  INHSV2 U18468 ( .I(n15157), .ZN(n16029) );
  AOI21HSV2 U18469 ( .A1(n15158), .A2(n16163), .B(n16029), .ZN(n15159) );
  OAI21HSV4 U18470 ( .A1(n14041), .A2(n16164), .B(n15159), .ZN(n15175) );
  NAND2HSV2 U18471 ( .A1(n15979), .A2(n28628), .ZN(n15173) );
  NAND2HSV0 U18472 ( .A1(\pe3/aot [14]), .A2(\pe3/bq[13] ), .ZN(n15167) );
  NAND2HSV2 U18473 ( .A1(\pe3/bq[11] ), .A2(\pe3/aot [13]), .ZN(n15304) );
  NAND2HSV2 U18474 ( .A1(\pe3/got [11]), .A2(n26380), .ZN(n15164) );
  NAND2HSV0 U18475 ( .A1(\pe3/aot [11]), .A2(n26351), .ZN(n15163) );
  NAND2HSV2 U18476 ( .A1(n21335), .A2(\pe3/pvq [6]), .ZN(n15171) );
  NAND2HSV0 U18477 ( .A1(\pe3/aot [12]), .A2(\pe3/bq[15] ), .ZN(n15169) );
  NAND2HSV0 U18478 ( .A1(\pe3/aot [15]), .A2(\pe3/bq[12] ), .ZN(n15168) );
  XOR2HSV0 U18479 ( .A1(n15169), .A2(n15168), .Z(n15170) );
  XOR3HSV2 U18480 ( .A1(\pe3/phq [6]), .A2(n15171), .A3(n15170), .Z(n15172) );
  INHSV2 U18481 ( .I(n26241), .ZN(n15245) );
  XNOR2HSV4 U18482 ( .A1(n15175), .A2(n15174), .ZN(n15186) );
  INHSV6 U18483 ( .I(n15186), .ZN(n27119) );
  NAND2HSV2 U18484 ( .A1(n15285), .A2(n14041), .ZN(n15182) );
  CLKNAND2HSV0 U18485 ( .A1(n15202), .A2(n15176), .ZN(n27115) );
  INHSV2 U18486 ( .I(n27115), .ZN(n15183) );
  CLKNAND2HSV2 U18487 ( .A1(n15182), .A2(n15183), .ZN(n15177) );
  AOI22HSV4 U18488 ( .A1(n16015), .A2(\pe3/ti_7t [6]), .B1(n27119), .B2(n15289), .ZN(n15187) );
  NOR2HSV1 U18489 ( .A1(n15182), .A2(n15181), .ZN(n27116) );
  CLKNAND2HSV1 U18490 ( .A1(n15183), .A2(n23382), .ZN(n15184) );
  NOR2HSV2 U18491 ( .A1(n27116), .A2(n15184), .ZN(n15185) );
  NAND3HSV4 U18492 ( .A1(n15186), .A2(n15185), .A3(n27117), .ZN(n15291) );
  OAI21HSV2 U18493 ( .A1(n15188), .A2(n15194), .B(n28707), .ZN(n15190) );
  NOR2HSV2 U18494 ( .A1(n21722), .A2(\pe3/ti_7t [7]), .ZN(n15286) );
  OR2HSV1 U18495 ( .A1(n15286), .A2(n16031), .Z(n15195) );
  INHSV2 U18496 ( .I(n15195), .ZN(n15192) );
  CLKAND2HSV2 U18497 ( .A1(n15288), .A2(n15284), .Z(n15197) );
  NOR2HSV2 U18498 ( .A1(n28707), .A2(n15195), .ZN(n15196) );
  NAND2HSV2 U18499 ( .A1(n15197), .A2(n15196), .ZN(n15198) );
  NAND2HSV0 U18500 ( .A1(n15241), .A2(n26413), .ZN(n15201) );
  NOR2HSV2 U18501 ( .A1(n15243), .A2(n16164), .ZN(n15200) );
  AND2HSV2 U18502 ( .A1(n15202), .A2(n28930), .Z(n15203) );
  NAND2HSV2 U18503 ( .A1(n15241), .A2(n28628), .ZN(n15231) );
  NAND2HSV0 U18504 ( .A1(n15979), .A2(\pe3/got [11]), .ZN(n15229) );
  NAND2HSV0 U18505 ( .A1(\pe3/aot [12]), .A2(\pe3/bq[13] ), .ZN(n15208) );
  NAND2HSV0 U18506 ( .A1(\pe3/bq[9] ), .A2(\pe3/aot [16]), .ZN(n15207) );
  XOR2HSV0 U18507 ( .A1(n15208), .A2(n15207), .Z(n15212) );
  NAND2HSV0 U18508 ( .A1(\pe3/bq[10] ), .A2(\pe3/aot [15]), .ZN(n15210) );
  INHSV2 U18509 ( .I(\pe3/got [9]), .ZN(n26680) );
  XOR2HSV2 U18510 ( .A1(n15210), .A2(n15209), .Z(n15211) );
  XNOR2HSV4 U18511 ( .A1(n15212), .A2(n15211), .ZN(n15214) );
  CLKNHSV2 U18512 ( .I(\pe3/aot [10]), .ZN(n15260) );
  CLKNHSV0 U18513 ( .I(\pe3/bq[15] ), .ZN(n15252) );
  NOR2HSV2 U18514 ( .A1(n15260), .A2(n15252), .ZN(n15941) );
  XNOR2HSV1 U18515 ( .A1(n15214), .A2(n15213), .ZN(n15222) );
  NAND2HSV0 U18516 ( .A1(\pe3/aot [14]), .A2(\pe3/bq[11] ), .ZN(n15216) );
  NAND2HSV0 U18517 ( .A1(n11932), .A2(\pe3/bq[12] ), .ZN(n15215) );
  XOR2HSV0 U18518 ( .A1(n15216), .A2(n15215), .Z(n15220) );
  NAND2HSV0 U18519 ( .A1(\pe3/aot [9]), .A2(n26351), .ZN(n15218) );
  NAND2HSV0 U18520 ( .A1(\pe3/aot [11]), .A2(\pe3/bq[14] ), .ZN(n15217) );
  XOR2HSV0 U18521 ( .A1(n15218), .A2(n15217), .Z(n15219) );
  XOR2HSV0 U18522 ( .A1(n15220), .A2(n15219), .Z(n15221) );
  CLKXOR2HSV2 U18523 ( .A1(n15222), .A2(n15221), .Z(n15225) );
  INHSV4 U18524 ( .I(n15223), .ZN(n26367) );
  CLKNAND2HSV1 U18525 ( .A1(n26367), .A2(\pe3/got [10]), .ZN(n15224) );
  XNOR2HSV1 U18526 ( .A1(n15225), .A2(n15224), .ZN(n15228) );
  INHSV3 U18527 ( .I(n15226), .ZN(n28920) );
  XOR3HSV2 U18528 ( .A1(n15229), .A2(n15228), .A3(n15227), .Z(n15230) );
  XNOR2HSV4 U18529 ( .A1(n15231), .A2(n15230), .ZN(n15232) );
  XNOR2HSV4 U18530 ( .A1(n15233), .A2(n15232), .ZN(n15234) );
  INHSV2 U18531 ( .I(n15236), .ZN(n15905) );
  NAND2HSV2 U18532 ( .A1(n15905), .A2(n16159), .ZN(n16021) );
  CLKNAND2HSV1 U18533 ( .A1(n16021), .A2(n15017), .ZN(n15237) );
  NOR2HSV4 U18534 ( .A1(n16023), .A2(n15237), .ZN(n15281) );
  CLKNAND2HSV3 U18535 ( .A1(n15288), .A2(n15284), .ZN(n15294) );
  INHSV4 U18536 ( .I(n15294), .ZN(n15909) );
  NAND2HSV2 U18537 ( .A1(\pe3/ti_7t [7]), .A2(n15238), .ZN(n16016) );
  INHSV2 U18538 ( .I(n16016), .ZN(n16056) );
  INHSV4 U18539 ( .I(n15241), .ZN(n15919) );
  INHSV2 U18540 ( .I(n15963), .ZN(n21313) );
  NAND2HSV0 U18541 ( .A1(\pe3/aot [14]), .A2(\pe3/bq[9] ), .ZN(n15251) );
  NAND2HSV2 U18542 ( .A1(n23345), .A2(\pe3/pvq [10]), .ZN(n15246) );
  XNOR2HSV1 U18543 ( .A1(n15246), .A2(\pe3/phq [10]), .ZN(n15250) );
  NAND2HSV0 U18544 ( .A1(\pe3/aot [11]), .A2(\pe3/bq[12] ), .ZN(n15248) );
  NAND2HSV0 U18545 ( .A1(n11932), .A2(\pe3/bq[10] ), .ZN(n15247) );
  XOR2HSV0 U18546 ( .A1(n15248), .A2(n15247), .Z(n15249) );
  XOR3HSV2 U18547 ( .A1(n15251), .A2(n15250), .A3(n15249), .Z(n15269) );
  NAND2HSV2 U18548 ( .A1(n26255), .A2(n28648), .ZN(n15268) );
  NAND2HSV0 U18549 ( .A1(\pe3/aot [7]), .A2(n26351), .ZN(n15254) );
  INHSV2 U18550 ( .I(n15252), .ZN(n26373) );
  CLKNAND2HSV0 U18551 ( .A1(\pe3/aot [8]), .A2(n26373), .ZN(n15253) );
  XOR2HSV0 U18552 ( .A1(n15254), .A2(n15253), .Z(n15259) );
  CLKNHSV0 U18553 ( .I(n14040), .ZN(n15255) );
  INHSV2 U18554 ( .I(n15255), .ZN(n26358) );
  CLKNAND2HSV1 U18555 ( .A1(n26358), .A2(\pe3/bq[7] ), .ZN(n15257) );
  NAND2HSV0 U18556 ( .A1(\pe3/got [7]), .A2(n26380), .ZN(n15256) );
  XOR2HSV0 U18557 ( .A1(n15257), .A2(n15256), .Z(n15258) );
  XOR2HSV0 U18558 ( .A1(n15259), .A2(n15258), .Z(n15266) );
  NAND2HSV0 U18559 ( .A1(\pe3/aot [9]), .A2(\pe3/bq[14] ), .ZN(n15262) );
  NAND2HSV0 U18560 ( .A1(\pe3/bq[8] ), .A2(\pe3/aot [15]), .ZN(n15261) );
  XOR2HSV0 U18561 ( .A1(n15262), .A2(n15261), .Z(n15263) );
  XOR2HSV0 U18562 ( .A1(n15264), .A2(n15263), .Z(n15265) );
  XOR2HSV0 U18563 ( .A1(n15266), .A2(n15265), .Z(n15267) );
  XOR3HSV2 U18564 ( .A1(n15269), .A2(n15268), .A3(n15267), .Z(n15271) );
  INHSV2 U18565 ( .I(n26680), .ZN(n26642) );
  NAND2HSV0 U18566 ( .A1(n15979), .A2(n26642), .ZN(n15270) );
  XNOR2HSV1 U18567 ( .A1(n15271), .A2(n15270), .ZN(n15274) );
  INHSV2 U18568 ( .I(n15272), .ZN(n26242) );
  NAND2HSV0 U18569 ( .A1(n26242), .A2(\pe3/got [10]), .ZN(n15273) );
  AOI22HSV4 U18570 ( .A1(n16159), .A2(\pe3/ti_7t [6]), .B1(n27119), .B2(n15289), .ZN(n15275) );
  CLKNAND2HSV4 U18571 ( .A1(n15275), .A2(n15291), .ZN(n23683) );
  XNOR2HSV4 U18572 ( .A1(n15277), .A2(n15276), .ZN(n15280) );
  INHSV4 U18573 ( .I(n15283), .ZN(n26625) );
  NOR2HSV2 U18574 ( .A1(n26625), .A2(n24313), .ZN(n15299) );
  INHSV1 U18575 ( .I(n15299), .ZN(n15300) );
  OR2HSV1 U18576 ( .A1(n15286), .A2(n16029), .Z(n15287) );
  AOI31HSV2 U18577 ( .A1(n13978), .A2(n23683), .A3(n15288), .B(n15287), .ZN(
        n15297) );
  CLKNHSV0 U18578 ( .I(n15291), .ZN(n15292) );
  NOR2HSV2 U18579 ( .A1(n15293), .A2(n15292), .ZN(n15295) );
  CLKNAND2HSV1 U18580 ( .A1(n15295), .A2(n15294), .ZN(n15296) );
  CLKNAND2HSV2 U18581 ( .A1(n15297), .A2(n15296), .ZN(n15298) );
  MUX2NHSV2 U18582 ( .I0(n15300), .I1(n15299), .S(n15298), .ZN(n15330) );
  INHSV2 U18583 ( .I(n15301), .ZN(n26348) );
  NAND2HSV2 U18584 ( .A1(n23683), .A2(n26348), .ZN(n15329) );
  NAND2HSV0 U18585 ( .A1(n16112), .A2(n15245), .ZN(n15327) );
  INHSV2 U18586 ( .I(n15302), .ZN(n26350) );
  NAND2HSV0 U18587 ( .A1(n26350), .A2(\pe3/got [10]), .ZN(n15325) );
  CLKNAND2HSV1 U18588 ( .A1(\pe3/bq[13] ), .A2(\pe3/aot [11]), .ZN(n15996) );
  XOR2HSV0 U18589 ( .A1(n16080), .A2(n15996), .Z(n15306) );
  BUFHSV2 U18590 ( .I(\pe3/bq[15] ), .Z(n16115) );
  NAND2HSV0 U18591 ( .A1(n16115), .A2(\pe3/aot [9]), .ZN(n15303) );
  XOR2HSV0 U18592 ( .A1(n15303), .A2(n15304), .Z(n15305) );
  XOR2HSV0 U18593 ( .A1(n15306), .A2(n15305), .Z(n15322) );
  NAND2HSV0 U18594 ( .A1(n26367), .A2(n26642), .ZN(n15321) );
  NAND2HSV0 U18595 ( .A1(\pe3/aot [14]), .A2(\pe3/bq[10] ), .ZN(n15308) );
  NAND2HSV0 U18596 ( .A1(\pe3/aot [10]), .A2(\pe3/bq[14] ), .ZN(n15307) );
  XOR2HSV0 U18597 ( .A1(n15308), .A2(n15307), .Z(n15312) );
  NAND2HSV0 U18598 ( .A1(\pe3/got [8]), .A2(n26380), .ZN(n15310) );
  NAND2HSV0 U18599 ( .A1(\pe3/aot [15]), .A2(\pe3/bq[9] ), .ZN(n15309) );
  XOR2HSV0 U18600 ( .A1(n15310), .A2(n15309), .Z(n15311) );
  XOR2HSV0 U18601 ( .A1(n15312), .A2(n15311), .Z(n15319) );
  NAND2HSV0 U18602 ( .A1(\pe3/bq[8] ), .A2(n14040), .ZN(n15314) );
  NAND2HSV0 U18603 ( .A1(\pe3/aot [8]), .A2(n23336), .ZN(n15313) );
  XOR2HSV0 U18604 ( .A1(n15314), .A2(n15313), .Z(n15317) );
  CLKNAND2HSV0 U18605 ( .A1(n21335), .A2(\pe3/pvq [9]), .ZN(n15315) );
  XOR2HSV0 U18606 ( .A1(n15315), .A2(\pe3/phq [9]), .Z(n15316) );
  XOR2HSV0 U18607 ( .A1(n15317), .A2(n15316), .Z(n15318) );
  XOR2HSV0 U18608 ( .A1(n15319), .A2(n15318), .Z(n15320) );
  XOR3HSV2 U18609 ( .A1(n15322), .A2(n15321), .A3(n15320), .Z(n15324) );
  NAND2HSV0 U18610 ( .A1(n26242), .A2(\pe3/got [11]), .ZN(n15323) );
  XOR3HSV2 U18611 ( .A1(n15325), .A2(n15324), .A3(n15323), .Z(n15326) );
  XNOR2HSV1 U18612 ( .A1(n15327), .A2(n15326), .ZN(n15328) );
  XNOR2HSV4 U18613 ( .A1(n15330), .A2(n13965), .ZN(n15961) );
  XNOR2HSV4 U18614 ( .A1(n15332), .A2(n15331), .ZN(n28611) );
  NOR2HSV2 U18615 ( .A1(n28611), .A2(n21720), .ZN(n15336) );
  CLKAND2HSV2 U18616 ( .A1(n15964), .A2(n15242), .Z(n15334) );
  OAI21HSV4 U18617 ( .A1(n15961), .A2(n15906), .B(n15334), .ZN(n15335) );
  AOI21HSV4 U18618 ( .A1(n15961), .A2(n15336), .B(n15335), .ZN(n15974) );
  XNOR2HSV4 U18619 ( .A1(n15975), .A2(n15974), .ZN(n28708) );
  INHSV6 U18620 ( .I(\pe10/aot [16]), .ZN(n16774) );
  INHSV4 U18621 ( .I(n16774), .ZN(n28424) );
  INHSV4 U18622 ( .I(\pe4/aot [16]), .ZN(n15379) );
  NOR2HSV2 U18623 ( .A1(n15363), .A2(n15379), .ZN(n15339) );
  CLKNAND2HSV0 U18624 ( .A1(\pe4/bq[16] ), .A2(\pe4/aot [16]), .ZN(n15338) );
  NAND2HSV2 U18625 ( .A1(\pe4/ti_1 ), .A2(\pe4/got [16]), .ZN(n15337) );
  MUX2NHSV4 U18626 ( .I0(n15339), .I1(n15338), .S(n15337), .ZN(n15342) );
  INHSV2 U18627 ( .I(n15502), .ZN(n15382) );
  AOI21HSV4 U18628 ( .A1(n15382), .A2(\pe4/pvq [1]), .B(\pe4/phq [1]), .ZN(
        n15340) );
  NOR2HSV4 U18629 ( .A1(n15341), .A2(n15340), .ZN(n15343) );
  NAND2HSV2 U18630 ( .A1(n15342), .A2(n15343), .ZN(n15347) );
  INHSV4 U18631 ( .I(n15342), .ZN(n15345) );
  INHSV4 U18632 ( .I(n15343), .ZN(n15344) );
  CLKNAND2HSV4 U18633 ( .A1(n15345), .A2(n15344), .ZN(n15346) );
  CLKNAND2HSV4 U18634 ( .A1(n15347), .A2(n15346), .ZN(n15416) );
  CLKNHSV3 U18635 ( .I(n15417), .ZN(n15418) );
  NOR2HSV4 U18636 ( .A1(n15428), .A2(n15418), .ZN(n15389) );
  INHSV2 U18637 ( .I(\pe4/got [15]), .ZN(n22987) );
  INHSV2 U18638 ( .I(n22987), .ZN(n15393) );
  NOR2HSV4 U18639 ( .A1(n15389), .A2(n26919), .ZN(n15362) );
  NAND2HSV2 U18640 ( .A1(\pe4/aot [14]), .A2(\pe4/bq[16] ), .ZN(n15349) );
  XNOR2HSV4 U18641 ( .A1(n15349), .A2(n15348), .ZN(n15354) );
  CLKNAND2HSV1 U18642 ( .A1(\pe4/phq [3]), .A2(\pe4/bq[14] ), .ZN(n15350) );
  NOR2HSV2 U18643 ( .A1(n15379), .A2(n15350), .ZN(n15352) );
  CLKNHSV4 U18644 ( .I(n15379), .ZN(n15737) );
  AOI21HSV2 U18645 ( .A1(n15737), .A2(\pe4/bq[14] ), .B(\pe4/phq [3]), .ZN(
        n15351) );
  NOR2HSV4 U18646 ( .A1(n15352), .A2(n15351), .ZN(n15353) );
  XNOR2HSV4 U18647 ( .A1(n15354), .A2(n15353), .ZN(n15357) );
  INHSV2 U18648 ( .I(n26958), .ZN(n15538) );
  INHSV4 U18649 ( .I(\pe4/aot [15]), .ZN(n15871) );
  NOR2HSV2 U18650 ( .A1(n15538), .A2(n15871), .ZN(n15356) );
  NAND2HSV0 U18651 ( .A1(\pe4/got [14]), .A2(\pe4/ti_1 ), .ZN(n15355) );
  XOR2HSV0 U18652 ( .A1(n15356), .A2(n15355), .Z(n15358) );
  CLKNAND2HSV2 U18653 ( .A1(n15357), .A2(n15358), .ZN(n15415) );
  INHSV4 U18654 ( .I(n15357), .ZN(n15360) );
  INHSV2 U18655 ( .I(n15358), .ZN(n15359) );
  CLKNAND2HSV4 U18656 ( .A1(n15360), .A2(n15359), .ZN(n15414) );
  CLKNAND2HSV3 U18657 ( .A1(n15415), .A2(n15414), .ZN(n15361) );
  XNOR2HSV4 U18658 ( .A1(n15361), .A2(n15362), .ZN(n15408) );
  INHSV3 U18659 ( .I(n15408), .ZN(n15376) );
  XNOR2HSV4 U18660 ( .A1(n15365), .A2(n15364), .ZN(n15369) );
  CLKNAND2HSV1 U18661 ( .A1(\pe4/got [15]), .A2(\pe4/ti_1 ), .ZN(n15367) );
  XOR2HSV2 U18662 ( .A1(n15367), .A2(n15366), .Z(n15368) );
  XNOR2HSV4 U18663 ( .A1(n15369), .A2(n15368), .ZN(n15372) );
  INHSV2 U18664 ( .I(\pe4/got [16]), .ZN(n22895) );
  CLKNHSV0 U18665 ( .I(ctro4), .ZN(n15370) );
  INAND2HSV2 U18666 ( .A1(n22895), .B1(n15370), .ZN(n21976) );
  NOR2HSV2 U18667 ( .A1(n15416), .A2(n21976), .ZN(n15371) );
  AOI22HSV4 U18668 ( .A1(ctro4), .A2(\pe4/ti_7t [2]), .B1(n15372), .B2(n15371), 
        .ZN(n15398) );
  INHSV4 U18669 ( .I(n15372), .ZN(n23483) );
  CLKBUFHSV4 U18670 ( .I(n15534), .Z(n15702) );
  INHSV2 U18671 ( .I(n15627), .ZN(n15394) );
  CLKNAND2HSV3 U18672 ( .A1(n15428), .A2(n15621), .ZN(n15395) );
  NAND3HSV4 U18673 ( .A1(n23483), .A2(n15394), .A3(n15395), .ZN(n15373) );
  NAND2HSV4 U18674 ( .A1(n15398), .A2(n15373), .ZN(n15413) );
  CLKAND2HSV2 U18675 ( .A1(n15413), .A2(n15531), .Z(n15375) );
  NOR2HSV2 U18676 ( .A1(n15394), .A2(\pe4/ti_7t [3]), .ZN(n15497) );
  NOR2HSV2 U18677 ( .A1(n15497), .A2(n22895), .ZN(n15406) );
  INHSV2 U18678 ( .I(n15406), .ZN(n15374) );
  INHSV2 U18679 ( .I(n15627), .ZN(n15487) );
  CLKBUFHSV4 U18680 ( .I(\pe4/ti_1 ), .Z(n27128) );
  CLKNAND2HSV1 U18681 ( .A1(\pe4/got [13]), .A2(n27128), .ZN(n15377) );
  XNOR2HSV1 U18682 ( .A1(n15378), .A2(n15377), .ZN(n15392) );
  INHSV2 U18683 ( .I(\pe4/bq[14] ), .ZN(n15507) );
  NOR2HSV2 U18684 ( .A1(n15507), .A2(n15871), .ZN(n15381) );
  INHSV4 U18685 ( .I(\pe4/bq[13] ), .ZN(n15596) );
  INHSV2 U18686 ( .I(n15596), .ZN(n15643) );
  INAND2HSV2 U18687 ( .A1(n15379), .B1(n15643), .ZN(n15380) );
  XNOR2HSV4 U18688 ( .A1(n15381), .A2(n15380), .ZN(n15386) );
  NAND2HSV2 U18689 ( .A1(n15382), .A2(\pe4/pvq [4]), .ZN(n15384) );
  NAND2HSV2 U18690 ( .A1(\pe4/aot [13]), .A2(\pe4/bq[16] ), .ZN(n15383) );
  XNOR2HSV4 U18691 ( .A1(n15386), .A2(n15385), .ZN(n15391) );
  INHSV2 U18692 ( .I(\pe4/ti_7t [1]), .ZN(n15419) );
  INAND2HSV4 U18693 ( .A1(n15419), .B1(n15418), .ZN(n15514) );
  INHSV2 U18694 ( .I(\pe4/got [14]), .ZN(n22880) );
  AOI21HSV0 U18695 ( .A1(n15514), .A2(n15534), .B(n22880), .ZN(n15387) );
  INHSV2 U18696 ( .I(n15387), .ZN(n15388) );
  NOR2HSV4 U18697 ( .A1(n15389), .A2(n15388), .ZN(n15390) );
  XOR3HSV2 U18698 ( .A1(n15392), .A2(n15391), .A3(n15390), .Z(n15399) );
  CLKNAND2HSV0 U18699 ( .A1(n15395), .A2(\pe4/got [15]), .ZN(n15396) );
  OAI22HSV2 U18700 ( .A1(n15398), .A2(n15748), .B1(n15397), .B2(n15396), .ZN(
        n15400) );
  INHSV2 U18701 ( .I(n15399), .ZN(n15402) );
  INHSV2 U18702 ( .I(n15400), .ZN(n15401) );
  CLKNAND2HSV1 U18703 ( .A1(n15404), .A2(n15403), .ZN(n15410) );
  CLKNHSV0 U18704 ( .I(n15413), .ZN(n25108) );
  CLKAND2HSV1 U18705 ( .A1(n15406), .A2(n15487), .Z(n15407) );
  OAI21HSV2 U18706 ( .A1(n15408), .A2(n25108), .B(n15407), .ZN(n15482) );
  NOR2HSV2 U18707 ( .A1(n15483), .A2(n15482), .ZN(n15409) );
  INHSV2 U18708 ( .I(n15702), .ZN(n15484) );
  AOI21HSV2 U18709 ( .A1(n15410), .A2(n15409), .B(n15491), .ZN(n15411) );
  INHSV2 U18710 ( .I(n28923), .ZN(n15724) );
  INHSV2 U18711 ( .I(\pe4/got [14]), .ZN(n24311) );
  NOR2HSV4 U18712 ( .A1(n15724), .A2(n24311), .ZN(n15450) );
  INHSV4 U18713 ( .I(n15413), .ZN(n15453) );
  INHSV4 U18714 ( .I(n15453), .ZN(n15469) );
  INHSV2 U18715 ( .I(\pe4/got [16]), .ZN(n15835) );
  CLKNAND2HSV4 U18716 ( .A1(n15469), .A2(n15813), .ZN(n15457) );
  INHSV4 U18717 ( .I(n15417), .ZN(n15535) );
  CLKBUFHSV4 U18718 ( .I(n15535), .Z(n21979) );
  AOI21HSV2 U18719 ( .A1(n15419), .A2(n15418), .B(n22987), .ZN(n15420) );
  XNOR2HSV4 U18720 ( .A1(n15422), .A2(n15421), .ZN(n15455) );
  XNOR2HSV4 U18721 ( .A1(n15457), .A2(n15455), .ZN(n29033) );
  NOR2HSV2 U18722 ( .A1(n29033), .A2(n15535), .ZN(n15426) );
  CLKNAND2HSV0 U18723 ( .A1(n15535), .A2(n15423), .ZN(n15424) );
  BUFHSV2 U18724 ( .I(\pe4/got [13]), .Z(n28463) );
  CLKNAND2HSV1 U18725 ( .A1(n15424), .A2(n28463), .ZN(n15425) );
  NOR2HSV2 U18726 ( .A1(n15426), .A2(n15425), .ZN(n15427) );
  INHSV2 U18727 ( .I(n15427), .ZN(n15447) );
  INHSV3 U18728 ( .I(n15453), .ZN(n15854) );
  NAND2HSV2 U18729 ( .A1(n15854), .A2(n25128), .ZN(n15430) );
  CLKNAND2HSV3 U18730 ( .A1(n15428), .A2(n22918), .ZN(n15515) );
  NAND2HSV4 U18731 ( .A1(n15515), .A2(n15514), .ZN(n23482) );
  NAND2HSV0 U18732 ( .A1(n23482), .A2(n13994), .ZN(n15429) );
  XNOR2HSV4 U18733 ( .A1(n15430), .A2(n15429), .ZN(n15446) );
  INHSV2 U18734 ( .I(n15596), .ZN(n26961) );
  NAND2HSV0 U18735 ( .A1(\pe4/aot [13]), .A2(n26961), .ZN(n15432) );
  INHSV4 U18736 ( .I(n15363), .ZN(n22834) );
  NAND2HSV0 U18737 ( .A1(\pe4/aot [10]), .A2(n22834), .ZN(n15431) );
  XOR2HSV0 U18738 ( .A1(n15432), .A2(n15431), .Z(n15445) );
  NAND2HSV0 U18739 ( .A1(\pe4/got [10]), .A2(\pe4/ti_1 ), .ZN(n15434) );
  NAND2HSV0 U18740 ( .A1(n15737), .A2(\pe4/bq[10] ), .ZN(n15433) );
  XOR2HSV0 U18741 ( .A1(n15434), .A2(n15433), .Z(n15436) );
  INHSV4 U18742 ( .I(n15502), .ZN(n23508) );
  INHSV2 U18743 ( .I(n21332), .ZN(n27105) );
  XNOR2HSV1 U18744 ( .A1(n15436), .A2(n15435), .ZN(n15444) );
  NAND2HSV0 U18745 ( .A1(\pe4/aot [11]), .A2(n26958), .ZN(n15438) );
  NAND2HSV0 U18746 ( .A1(\pe4/aot [14]), .A2(\pe4/bq[12] ), .ZN(n15437) );
  XOR2HSV0 U18747 ( .A1(n15438), .A2(n15437), .Z(n15442) );
  BUFHSV2 U18748 ( .I(\pe4/aot [15]), .Z(n15784) );
  NAND2HSV0 U18749 ( .A1(n15784), .A2(\pe4/bq[11] ), .ZN(n15440) );
  NAND2HSV0 U18750 ( .A1(\pe4/aot [12]), .A2(\pe4/bq[14] ), .ZN(n15439) );
  XOR2HSV0 U18751 ( .A1(n15440), .A2(n15439), .Z(n15441) );
  XOR2HSV0 U18752 ( .A1(n15442), .A2(n15441), .Z(n15443) );
  XNOR2HSV4 U18753 ( .A1(n15450), .A2(n15449), .ZN(n15477) );
  NAND2HSV2 U18754 ( .A1(n28974), .A2(n15813), .ZN(n15566) );
  CLKNHSV0 U18755 ( .I(n15621), .ZN(n15451) );
  NOR2HSV0 U18756 ( .A1(n15534), .A2(n15451), .ZN(n15452) );
  INHSV2 U18757 ( .I(n15453), .ZN(n15640) );
  NOR2HSV2 U18758 ( .A1(n15497), .A2(n26919), .ZN(n15454) );
  CLKNAND2HSV4 U18759 ( .A1(n15499), .A2(n15454), .ZN(n15472) );
  INHSV2 U18760 ( .I(n15455), .ZN(n15456) );
  INHSV4 U18761 ( .I(n15500), .ZN(n15474) );
  INHSV2 U18762 ( .I(n21332), .ZN(n21759) );
  NAND2HSV2 U18763 ( .A1(n21759), .A2(\pe4/pvq [5]), .ZN(n15458) );
  XNOR2HSV4 U18764 ( .A1(n15459), .A2(n15458), .ZN(n15466) );
  NAND2HSV0 U18765 ( .A1(n26958), .A2(\pe4/aot [13]), .ZN(n15461) );
  NAND2HSV0 U18766 ( .A1(\pe4/bq[14] ), .A2(\pe4/aot [14]), .ZN(n15460) );
  INAND2HSV4 U18767 ( .A1(n15596), .B1(\pe4/aot [15]), .ZN(n15599) );
  NAND2HSV2 U18768 ( .A1(\pe4/aot [12]), .A2(\pe4/bq[16] ), .ZN(n15462) );
  XOR2HSV2 U18769 ( .A1(n15599), .A2(n15462), .Z(n15463) );
  CLKXOR2HSV4 U18770 ( .A1(n15466), .A2(n15465), .Z(n15468) );
  BUFHSV2 U18771 ( .I(\pe4/got [13]), .Z(n25131) );
  CLKXOR2HSV4 U18772 ( .A1(n15468), .A2(n15467), .Z(n15471) );
  CLKNAND2HSV3 U18773 ( .A1(n15469), .A2(n25134), .ZN(n15470) );
  XNOR2HSV4 U18774 ( .A1(n15471), .A2(n15470), .ZN(n15473) );
  OAI21HSV4 U18775 ( .A1(n15472), .A2(n15474), .B(n15473), .ZN(n15478) );
  INHSV2 U18776 ( .I(n21976), .ZN(n15839) );
  INHSV2 U18777 ( .I(n15476), .ZN(n15475) );
  INHSV2 U18778 ( .I(\pe4/got [15]), .ZN(n15748) );
  BUFHSV2 U18779 ( .I(n15535), .Z(n15900) );
  CLKNAND2HSV2 U18780 ( .A1(n15479), .A2(n15478), .ZN(n27229) );
  INAND2HSV2 U18781 ( .A1(n15835), .B1(n15487), .ZN(n15480) );
  NOR2HSV2 U18782 ( .A1(n15492), .A2(n15485), .ZN(n15486) );
  INHSV2 U18783 ( .I(n15496), .ZN(n15494) );
  NAND2HSV2 U18784 ( .A1(n15494), .A2(n15495), .ZN(n15530) );
  NOR2HSV0 U18785 ( .A1(n15497), .A2(n22880), .ZN(n15498) );
  NAND3HSV2 U18786 ( .A1(n15500), .A2(n15499), .A3(n15498), .ZN(n15521) );
  NAND2HSV0 U18787 ( .A1(n15640), .A2(n25131), .ZN(n15501) );
  INHSV1 U18788 ( .I(n15501), .ZN(n15520) );
  CLKNHSV0 U18789 ( .I(\pe4/aot [14]), .ZN(n22115) );
  XNOR2HSV4 U18790 ( .A1(n15504), .A2(n15503), .ZN(n15513) );
  NAND2HSV0 U18791 ( .A1(n26958), .A2(\pe4/aot [12]), .ZN(n15506) );
  CLKNAND2HSV1 U18792 ( .A1(\pe4/got [11]), .A2(n27128), .ZN(n15505) );
  XOR2HSV2 U18793 ( .A1(n15506), .A2(n15505), .Z(n15511) );
  INHSV2 U18794 ( .I(\pe4/aot [13]), .ZN(n22000) );
  NOR2HSV2 U18795 ( .A1(n22000), .A2(n15507), .ZN(n15509) );
  NAND2HSV0 U18796 ( .A1(\pe4/aot [11]), .A2(\pe4/bq[16] ), .ZN(n15508) );
  XOR2HSV0 U18797 ( .A1(n15509), .A2(n15508), .Z(n15510) );
  XOR2HSV0 U18798 ( .A1(n15511), .A2(n15510), .Z(n15512) );
  XNOR2HSV4 U18799 ( .A1(n15513), .A2(n15512), .ZN(n15517) );
  NAND2HSV4 U18800 ( .A1(n15515), .A2(n15514), .ZN(n28653) );
  NAND2HSV0 U18801 ( .A1(n28653), .A2(n28428), .ZN(n15516) );
  XNOR2HSV4 U18802 ( .A1(n15517), .A2(n15516), .ZN(n15519) );
  AOI21HSV2 U18803 ( .A1(n15854), .A2(n25131), .B(n15519), .ZN(n15518) );
  CLKNAND2HSV2 U18804 ( .A1(n28923), .A2(\pe4/got [15]), .ZN(n15523) );
  NAND2HSV2 U18805 ( .A1(n15522), .A2(n15523), .ZN(n15527) );
  INHSV2 U18806 ( .I(n15522), .ZN(n15525) );
  INHSV2 U18807 ( .I(n15523), .ZN(n15524) );
  CLKNAND2HSV3 U18808 ( .A1(n15527), .A2(n15526), .ZN(n15528) );
  MUX2NHSV4 U18809 ( .I0(n15530), .I1(n15529), .S(n15528), .ZN(n15570) );
  CLKNAND2HSV4 U18810 ( .A1(n15570), .A2(n15531), .ZN(n15580) );
  NAND2HSV2 U18811 ( .A1(\pe4/ti_7t [6]), .A2(n15702), .ZN(n15579) );
  NAND2HSV2 U18812 ( .A1(n15580), .A2(n15579), .ZN(n22931) );
  NOR2HSV4 U18813 ( .A1(n15532), .A2(n21979), .ZN(n15622) );
  INHSV2 U18814 ( .I(n28933), .ZN(n15533) );
  CLKNAND2HSV3 U18815 ( .A1(n15622), .A2(n15533), .ZN(n15686) );
  CLKAND2HSV2 U18816 ( .A1(n15638), .A2(n15813), .Z(n15681) );
  NAND3HSV4 U18817 ( .A1(n15685), .A2(n15686), .A3(n15681), .ZN(n15628) );
  BUFHSV2 U18818 ( .I(n15535), .Z(n15752) );
  BUFHSV2 U18819 ( .I(n15752), .Z(n28812) );
  INHSV2 U18820 ( .I(\pe4/got [12]), .ZN(n22822) );
  NOR2HSV2 U18821 ( .A1(n15723), .A2(n22822), .ZN(n15561) );
  CLKNAND2HSV1 U18822 ( .A1(n28653), .A2(\pe4/got [10]), .ZN(n15536) );
  CLKNHSV0 U18823 ( .I(\pe4/aot [10]), .ZN(n15597) );
  NOR2HSV1 U18824 ( .A1(n15597), .A2(n15538), .ZN(n15540) );
  NAND2HSV0 U18825 ( .A1(\pe4/bq[9] ), .A2(n28683), .ZN(n15539) );
  XOR2HSV0 U18826 ( .A1(n15540), .A2(n15539), .Z(n15544) );
  INHSV2 U18827 ( .I(\pe4/got [9]), .ZN(n27826) );
  CLKNAND2HSV0 U18828 ( .A1(\pe4/got [9]), .A2(\pe4/ti_1 ), .ZN(n15542) );
  NAND2HSV0 U18829 ( .A1(\pe4/bq[11] ), .A2(\pe4/aot [14]), .ZN(n15541) );
  XOR2HSV0 U18830 ( .A1(n15542), .A2(n15541), .Z(n15543) );
  XOR2HSV0 U18831 ( .A1(n15544), .A2(n15543), .Z(n15549) );
  INHSV2 U18832 ( .I(n21332), .ZN(n27129) );
  NAND2HSV2 U18833 ( .A1(n27129), .A2(\pe4/pvq [8]), .ZN(n15545) );
  XNOR2HSV1 U18834 ( .A1(n15545), .A2(\pe4/phq [8]), .ZN(n15547) );
  NAND2HSV0 U18835 ( .A1(\pe4/aot [12]), .A2(n26961), .ZN(n15546) );
  XNOR2HSV1 U18836 ( .A1(n15547), .A2(n15546), .ZN(n15548) );
  XNOR2HSV1 U18837 ( .A1(n15549), .A2(n15548), .ZN(n15557) );
  NAND2HSV0 U18838 ( .A1(\pe4/aot [9]), .A2(n22834), .ZN(n15551) );
  NAND2HSV0 U18839 ( .A1(n15784), .A2(\pe4/bq[10] ), .ZN(n15550) );
  XOR2HSV0 U18840 ( .A1(n15551), .A2(n15550), .Z(n15555) );
  BUFHSV4 U18841 ( .I(\pe4/bq[14] ), .Z(n27060) );
  NAND2HSV0 U18842 ( .A1(\pe4/aot [11]), .A2(n27060), .ZN(n15553) );
  NAND2HSV0 U18843 ( .A1(\pe4/aot [13]), .A2(\pe4/bq[12] ), .ZN(n15552) );
  XOR2HSV0 U18844 ( .A1(n15553), .A2(n15552), .Z(n15554) );
  XOR2HSV0 U18845 ( .A1(n15555), .A2(n15554), .Z(n15556) );
  XNOR2HSV1 U18846 ( .A1(n15557), .A2(n15556), .ZN(n15558) );
  XNOR2HSV4 U18847 ( .A1(n15561), .A2(n15560), .ZN(n15563) );
  BUFHSV4 U18848 ( .I(n28923), .Z(n22827) );
  NAND2HSV0 U18849 ( .A1(n22827), .A2(n25131), .ZN(n15562) );
  XNOR2HSV4 U18850 ( .A1(n15563), .A2(n15562), .ZN(n15569) );
  NAND2HSV2 U18851 ( .A1(n28696), .A2(n25134), .ZN(n15568) );
  XNOR2HSV4 U18852 ( .A1(n15569), .A2(n15568), .ZN(n15573) );
  CLKNHSV0 U18853 ( .I(\pe4/ti_7t [6]), .ZN(n15571) );
  AO21HSV1 U18854 ( .A1(n15571), .A2(n15752), .B(n15748), .Z(n15572) );
  AOI21HSV4 U18855 ( .A1(n23985), .A2(n22918), .B(n15572), .ZN(n15574) );
  INHSV4 U18856 ( .I(n15573), .ZN(n15576) );
  INHSV3 U18857 ( .I(n15574), .ZN(n15575) );
  CLKNAND2HSV8 U18858 ( .A1(n15578), .A2(n15577), .ZN(n15688) );
  NOR2HSV2 U18859 ( .A1(n15723), .A2(n27825), .ZN(n15611) );
  NAND2HSV0 U18860 ( .A1(n15854), .A2(\pe4/got [9]), .ZN(n15582) );
  CLKNHSV0 U18861 ( .I(n28653), .ZN(n22932) );
  NOR2HSV2 U18862 ( .A1(n22932), .A2(n27827), .ZN(n15581) );
  XNOR2HSV1 U18863 ( .A1(n15582), .A2(n15581), .ZN(n15609) );
  NAND2HSV0 U18864 ( .A1(\pe4/aot [9]), .A2(n27060), .ZN(n15584) );
  NAND2HSV0 U18865 ( .A1(\pe4/aot [11]), .A2(\pe4/bq[12] ), .ZN(n15583) );
  XOR2HSV0 U18866 ( .A1(n15584), .A2(n15583), .Z(n15588) );
  BUFHSV2 U18867 ( .I(n22834), .Z(n26948) );
  NAND2HSV0 U18868 ( .A1(\pe4/aot [7]), .A2(n26948), .ZN(n15586) );
  NAND2HSV0 U18869 ( .A1(\pe4/aot [13]), .A2(\pe4/bq[10] ), .ZN(n15585) );
  XOR2HSV0 U18870 ( .A1(n15586), .A2(n15585), .Z(n15587) );
  XOR2HSV0 U18871 ( .A1(n15588), .A2(n15587), .Z(n15595) );
  NAND2HSV0 U18872 ( .A1(\pe4/bq[9] ), .A2(\pe4/aot [14]), .ZN(n15590) );
  NAND2HSV0 U18873 ( .A1(n15737), .A2(\pe4/bq[7] ), .ZN(n15589) );
  XOR2HSV0 U18874 ( .A1(n15590), .A2(n15589), .Z(n15593) );
  INHSV2 U18875 ( .I(n21332), .ZN(n28924) );
  CLKNAND2HSV1 U18876 ( .A1(n28924), .A2(\pe4/pvq [10]), .ZN(n15591) );
  XOR2HSV0 U18877 ( .A1(n15591), .A2(\pe4/phq [10]), .Z(n15592) );
  XOR2HSV0 U18878 ( .A1(n15593), .A2(n15592), .Z(n15594) );
  XOR2HSV0 U18879 ( .A1(n15595), .A2(n15594), .Z(n15607) );
  CLKNAND2HSV0 U18880 ( .A1(\pe4/aot [10]), .A2(\pe4/bq[8] ), .ZN(n22838) );
  NAND2HSV0 U18881 ( .A1(n15784), .A2(\pe4/bq[8] ), .ZN(n15787) );
  OAI21HSV0 U18882 ( .A1(n15597), .A2(n15596), .B(n15787), .ZN(n15598) );
  OAI21HSV1 U18883 ( .A1(n15599), .A2(n22838), .B(n15598), .ZN(n15601) );
  NAND2HSV0 U18884 ( .A1(\pe4/got [7]), .A2(n27128), .ZN(n15600) );
  XNOR2HSV1 U18885 ( .A1(n15601), .A2(n15600), .ZN(n15605) );
  NAND2HSV0 U18886 ( .A1(\pe4/aot [12]), .A2(\pe4/bq[11] ), .ZN(n15603) );
  NAND2HSV0 U18887 ( .A1(\pe4/aot [8]), .A2(n26958), .ZN(n15602) );
  XOR2HSV0 U18888 ( .A1(n15603), .A2(n15602), .Z(n15604) );
  XNOR2HSV1 U18889 ( .A1(n15605), .A2(n15604), .ZN(n15606) );
  XNOR2HSV1 U18890 ( .A1(n15607), .A2(n15606), .ZN(n15608) );
  XNOR2HSV1 U18891 ( .A1(n15609), .A2(n15608), .ZN(n15610) );
  XNOR2HSV4 U18892 ( .A1(n15611), .A2(n15610), .ZN(n15613) );
  NAND2HSV0 U18893 ( .A1(n22827), .A2(n13994), .ZN(n15612) );
  XNOR2HSV4 U18894 ( .A1(n15613), .A2(n15612), .ZN(n15616) );
  CLKNAND2HSV1 U18895 ( .A1(n28696), .A2(n28428), .ZN(n15615) );
  XNOR2HSV4 U18896 ( .A1(n15616), .A2(n15615), .ZN(n15617) );
  XNOR2HSV4 U18897 ( .A1(n15618), .A2(n15617), .ZN(n15625) );
  CLKNAND2HSV0 U18898 ( .A1(n15638), .A2(n28612), .ZN(n15619) );
  AOI31HSV2 U18899 ( .A1(n15620), .A2(n15853), .A3(n15839), .B(n15619), .ZN(
        n15623) );
  CLKNAND2HSV4 U18900 ( .A1(n28933), .A2(n15621), .ZN(n15711) );
  CLKNAND2HSV3 U18901 ( .A1(n15711), .A2(n15622), .ZN(n15849) );
  CLKNAND2HSV1 U18902 ( .A1(n15623), .A2(n15849), .ZN(n15624) );
  XNOR2HSV4 U18903 ( .A1(n15625), .A2(n15624), .ZN(n15629) );
  INHSV2 U18904 ( .I(n15748), .ZN(n28592) );
  OAI21HSV2 U18905 ( .A1(n15417), .A2(\pe4/ti_7t [8]), .B(n28592), .ZN(n15630)
         );
  INHSV1 U18906 ( .I(n15630), .ZN(n15626) );
  OAI21HSV4 U18907 ( .A1(n29031), .A2(n15627), .B(n13979), .ZN(n15822) );
  NOR2HSV1 U18908 ( .A1(n15698), .A2(n27976), .ZN(n15636) );
  INHSV2 U18909 ( .I(n15629), .ZN(n15635) );
  CLKNHSV0 U18910 ( .I(n15688), .ZN(n15631) );
  AOI31HSV2 U18911 ( .A1(n15632), .A2(n15631), .A3(n15417), .B(n15630), .ZN(
        n15633) );
  INHSV2 U18912 ( .I(n15633), .ZN(n15634) );
  NAND2HSV4 U18913 ( .A1(n15635), .A2(n15634), .ZN(n15823) );
  NAND2HSV2 U18914 ( .A1(n15837), .A2(n15813), .ZN(n15696) );
  NOR2HSV2 U18915 ( .A1(n15697), .A2(n15696), .ZN(n15699) );
  INHSV1 U18916 ( .I(n15638), .ZN(n15847) );
  NOR2HSV2 U18917 ( .A1(n15847), .A2(n26919), .ZN(n15639) );
  CLKAND2HSV4 U18918 ( .A1(n15849), .A2(n15639), .Z(n15676) );
  CLKNAND2HSV2 U18919 ( .A1(n15676), .A2(n15852), .ZN(n15674) );
  CLKNAND2HSV0 U18920 ( .A1(n15640), .A2(\pe4/got [10]), .ZN(n15642) );
  NAND2HSV0 U18921 ( .A1(n23482), .A2(\pe4/got [9]), .ZN(n15641) );
  XNOR2HSV1 U18922 ( .A1(n15642), .A2(n15641), .ZN(n15664) );
  CLKNAND2HSV0 U18923 ( .A1(n15784), .A2(\pe4/bq[9] ), .ZN(n15645) );
  NAND2HSV0 U18924 ( .A1(\pe4/aot [11]), .A2(n15643), .ZN(n15644) );
  XOR2HSV0 U18925 ( .A1(n15645), .A2(n15644), .Z(n15649) );
  BUFHSV2 U18926 ( .I(\pe4/bq[15] ), .Z(n22943) );
  NAND2HSV0 U18927 ( .A1(n22943), .A2(\pe4/aot [9]), .ZN(n15647) );
  NAND2HSV0 U18928 ( .A1(\pe4/got [8]), .A2(n27128), .ZN(n15646) );
  XOR2HSV0 U18929 ( .A1(n15647), .A2(n15646), .Z(n15648) );
  XOR2HSV0 U18930 ( .A1(n15649), .A2(n15648), .Z(n15656) );
  NAND2HSV0 U18931 ( .A1(n15737), .A2(\pe4/bq[8] ), .ZN(n15651) );
  NAND2HSV0 U18932 ( .A1(\pe4/aot [12]), .A2(\pe4/bq[12] ), .ZN(n15650) );
  XOR2HSV0 U18933 ( .A1(n15651), .A2(n15650), .Z(n15654) );
  CLKNAND2HSV0 U18934 ( .A1(n21759), .A2(\pe4/pvq [9]), .ZN(n15652) );
  XOR2HSV0 U18935 ( .A1(n15652), .A2(\pe4/phq [9]), .Z(n15653) );
  XOR2HSV0 U18936 ( .A1(n15654), .A2(n15653), .Z(n15655) );
  XOR2HSV0 U18937 ( .A1(n15656), .A2(n15655), .Z(n15662) );
  INHSV2 U18938 ( .I(\pe4/bq[11] ), .ZN(n26968) );
  NOR2HSV2 U18939 ( .A1(n22000), .A2(n26968), .ZN(n15874) );
  NAND2HSV0 U18940 ( .A1(\pe4/bq[10] ), .A2(\pe4/aot [14]), .ZN(n22957) );
  XOR2HSV0 U18941 ( .A1(n15874), .A2(n22957), .Z(n15660) );
  NAND2HSV0 U18942 ( .A1(\pe4/aot [8]), .A2(n26948), .ZN(n15658) );
  NAND2HSV0 U18943 ( .A1(\pe4/aot [10]), .A2(n27060), .ZN(n15657) );
  XOR2HSV0 U18944 ( .A1(n15658), .A2(n15657), .Z(n15659) );
  XOR2HSV0 U18945 ( .A1(n15660), .A2(n15659), .Z(n15661) );
  XNOR2HSV1 U18946 ( .A1(n15662), .A2(n15661), .ZN(n15663) );
  XNOR2HSV1 U18947 ( .A1(n15664), .A2(n15663), .ZN(n15667) );
  NOR2HSV2 U18948 ( .A1(n15723), .A2(n27871), .ZN(n15666) );
  CLKNAND2HSV1 U18949 ( .A1(n22827), .A2(n28428), .ZN(n15665) );
  CLKNAND2HSV1 U18950 ( .A1(n15668), .A2(n15669), .ZN(n15673) );
  INHSV2 U18951 ( .I(n15669), .ZN(n15670) );
  CLKNAND2HSV3 U18952 ( .A1(n15673), .A2(n15672), .ZN(n15675) );
  CLKNAND2HSV2 U18953 ( .A1(n15680), .A2(n29031), .ZN(n15695) );
  CLKNHSV0 U18954 ( .I(n15686), .ZN(n15683) );
  CLKNAND2HSV1 U18955 ( .A1(n15685), .A2(n15681), .ZN(n15682) );
  NOR2HSV2 U18956 ( .A1(n15683), .A2(n15682), .ZN(n15684) );
  CLKAND2HSV2 U18957 ( .A1(n15688), .A2(n15684), .Z(n15691) );
  NAND2HSV2 U18958 ( .A1(n15686), .A2(n15685), .ZN(n15687) );
  OAI21HSV2 U18959 ( .A1(n15689), .A2(n15688), .B(n15370), .ZN(n15690) );
  NOR2HSV2 U18960 ( .A1(n15691), .A2(n15690), .ZN(n15692) );
  AOI22HSV4 U18961 ( .A1(\pe4/ti_7t [9]), .A2(n15693), .B1(n15692), .B2(n25663), .ZN(n15694) );
  CLKNAND2HSV4 U18962 ( .A1(n15695), .A2(n15694), .ZN(n15747) );
  INHSV3 U18963 ( .I(n15747), .ZN(n15821) );
  INHSV4 U18964 ( .I(n15821), .ZN(n27784) );
  INHSV6 U18965 ( .I(n21992), .ZN(n15844) );
  AOI21HSV4 U18966 ( .A1(n15844), .A2(n15697), .B(n15696), .ZN(n15751) );
  INHSV2 U18967 ( .I(n15698), .ZN(n15824) );
  INHSV2 U18968 ( .I(n15700), .ZN(n23058) );
  NAND2HSV2 U18969 ( .A1(n23058), .A2(n27976), .ZN(n15845) );
  NAND2HSV2 U18970 ( .A1(n15845), .A2(n28612), .ZN(n15701) );
  NOR2HSV4 U18971 ( .A1(n15846), .A2(n15701), .ZN(n15746) );
  NOR2HSV0 U18972 ( .A1(n15702), .A2(n22822), .ZN(n15703) );
  AND2HSV2 U18973 ( .A1(n28933), .A2(n15703), .Z(n15718) );
  INHSV2 U18974 ( .I(n15704), .ZN(n15712) );
  INHSV4 U18975 ( .I(n15712), .ZN(n15758) );
  CLKNAND2HSV1 U18976 ( .A1(n15718), .A2(n15758), .ZN(n15706) );
  NOR2HSV2 U18977 ( .A1(n15706), .A2(n15705), .ZN(n15710) );
  INHSV2 U18978 ( .I(\pe4/got [13]), .ZN(n26932) );
  NOR2HSV1 U18979 ( .A1(n15847), .A2(n26932), .ZN(n15713) );
  CLKNHSV0 U18980 ( .I(n15713), .ZN(n15707) );
  OR2HSV1 U18981 ( .A1(n15707), .A2(n21968), .Z(n15708) );
  NOR2HSV2 U18982 ( .A1(n15710), .A2(n15709), .ZN(n15722) );
  CLKNAND2HSV1 U18983 ( .A1(n12265), .A2(n15758), .ZN(n15716) );
  CLKNHSV2 U18984 ( .I(n15711), .ZN(n15759) );
  CLKNAND2HSV3 U18985 ( .A1(n15759), .A2(n15712), .ZN(n15717) );
  CLKAND2HSV2 U18986 ( .A1(n15714), .A2(n15713), .Z(n15715) );
  NAND3HSV2 U18987 ( .A1(n15716), .A2(n15717), .A3(n15715), .ZN(n15721) );
  INHSV2 U18988 ( .I(n15717), .ZN(n15719) );
  NAND2HSV2 U18989 ( .A1(n15719), .A2(n15718), .ZN(n15720) );
  NAND3HSV4 U18990 ( .A1(n15722), .A2(n15721), .A3(n15720), .ZN(n15744) );
  BUFHSV2 U18991 ( .I(n15723), .Z(n26981) );
  INHSV2 U18992 ( .I(n26981), .ZN(n28951) );
  NAND2HSV0 U18993 ( .A1(n28951), .A2(\pe4/got [9]), .ZN(n15742) );
  INHSV2 U18994 ( .I(n15724), .ZN(n27739) );
  BUFHSV2 U18995 ( .I(n15854), .Z(n28671) );
  NAND2HSV0 U18996 ( .A1(\pe4/aot [10]), .A2(\pe4/bq[12] ), .ZN(n15726) );
  NAND2HSV0 U18997 ( .A1(\pe4/aot [11]), .A2(\pe4/bq[11] ), .ZN(n15725) );
  XOR2HSV0 U18998 ( .A1(n15726), .A2(n15725), .Z(n15730) );
  INHSV2 U18999 ( .I(\pe4/got [6]), .ZN(n27905) );
  NAND2HSV0 U19000 ( .A1(\pe4/got [6]), .A2(n27128), .ZN(n15728) );
  NAND2HSV0 U19001 ( .A1(\pe4/aot [8]), .A2(n27060), .ZN(n15727) );
  XOR2HSV0 U19002 ( .A1(n15728), .A2(n15727), .Z(n15729) );
  NAND2HSV0 U19003 ( .A1(\pe4/aot [6]), .A2(n22834), .ZN(n15732) );
  NAND2HSV0 U19004 ( .A1(\pe4/aot [12]), .A2(\pe4/bq[10] ), .ZN(n15731) );
  XOR2HSV0 U19005 ( .A1(n15732), .A2(n15731), .Z(n15736) );
  NAND2HSV0 U19006 ( .A1(\pe4/bq[8] ), .A2(\pe4/aot [14]), .ZN(n15734) );
  NAND2HSV0 U19007 ( .A1(n22943), .A2(\pe4/aot [7]), .ZN(n15733) );
  XOR2HSV0 U19008 ( .A1(n15734), .A2(n15733), .Z(n15735) );
  BUFHSV2 U19009 ( .I(\pe4/bq[13] ), .Z(n23076) );
  BUFHSV2 U19010 ( .I(n15737), .Z(n28683) );
  NAND2HSV2 U19011 ( .A1(n28683), .A2(\pe4/bq[6] ), .ZN(n22001) );
  NAND2HSV0 U19012 ( .A1(\pe4/aot [13]), .A2(\pe4/bq[9] ), .ZN(n15738) );
  BUFHSV4 U19013 ( .I(n28696), .Z(n27830) );
  NAND2HSV0 U19014 ( .A1(n27830), .A2(n13994), .ZN(n15740) );
  XOR3HSV2 U19015 ( .A1(n15742), .A2(n15741), .A3(n15740), .Z(n15743) );
  XNOR2HSV4 U19016 ( .A1(n15744), .A2(n15743), .ZN(n15745) );
  XNOR2HSV4 U19017 ( .A1(n15746), .A2(n15745), .ZN(n15750) );
  INAND2HSV2 U19018 ( .A1(n15748), .B1(n15747), .ZN(n15749) );
  INHSV2 U19019 ( .I(n15370), .ZN(n22801) );
  NAND2HSV2 U19020 ( .A1(n15752), .A2(\pe4/ti_7t [11]), .ZN(n22042) );
  INHSV2 U19021 ( .I(n15834), .ZN(n15832) );
  CLKNAND2HSV1 U19022 ( .A1(n21994), .A2(n25128), .ZN(n15754) );
  CLKNHSV0 U19023 ( .I(n15754), .ZN(n15755) );
  XNOR2HSV4 U19024 ( .A1(n15759), .A2(n15758), .ZN(n28957) );
  MUX2HSV2 U19025 ( .I0(\pe4/ti_7t [7]), .I1(n28957), .S(n15531), .Z(
        \pe4/ti_7[7] ) );
  NAND2HSV0 U19026 ( .A1(\pe4/ti_7[7] ), .A2(n13994), .ZN(n15804) );
  NAND2HSV2 U19027 ( .A1(n22825), .A2(\pe4/got [10]), .ZN(n15802) );
  NAND2HSV0 U19028 ( .A1(n28951), .A2(n13996), .ZN(n15800) );
  CLKNAND2HSV0 U19029 ( .A1(n22827), .A2(\pe4/got [8]), .ZN(n15797) );
  INHSV2 U19030 ( .I(\pe4/got [6]), .ZN(n22117) );
  CLKNAND2HSV0 U19031 ( .A1(n28671), .A2(n22826), .ZN(n15761) );
  NAND2HSV0 U19032 ( .A1(n23482), .A2(\pe4/got [5]), .ZN(n15760) );
  XNOR2HSV1 U19033 ( .A1(n15761), .A2(n15760), .ZN(n15795) );
  NAND2HSV0 U19034 ( .A1(\pe4/aot [6]), .A2(n27060), .ZN(n15763) );
  NAND2HSV0 U19035 ( .A1(\pe4/aot [4]), .A2(n22834), .ZN(n15762) );
  XOR2HSV0 U19036 ( .A1(n15763), .A2(n15762), .Z(n15768) );
  CLKNHSV0 U19037 ( .I(\pe4/ti_1 ), .ZN(n15764) );
  NAND2HSV0 U19038 ( .A1(\pe4/got [4]), .A2(n27128), .ZN(n15766) );
  NAND2HSV0 U19039 ( .A1(\pe4/aot [8]), .A2(\pe4/bq[12] ), .ZN(n15765) );
  XOR2HSV0 U19040 ( .A1(n15766), .A2(n15765), .Z(n15767) );
  XOR2HSV0 U19041 ( .A1(n15768), .A2(n15767), .Z(n15776) );
  NAND2HSV0 U19042 ( .A1(\pe4/aot [11]), .A2(\pe4/bq[9] ), .ZN(n15770) );
  NAND2HSV0 U19043 ( .A1(\pe4/aot [10]), .A2(\pe4/bq[10] ), .ZN(n15769) );
  XOR2HSV0 U19044 ( .A1(n15770), .A2(n15769), .Z(n15774) );
  NAND2HSV0 U19045 ( .A1(\pe4/aot [14]), .A2(\pe4/bq[6] ), .ZN(n15772) );
  NAND2HSV0 U19046 ( .A1(\pe4/aot [13]), .A2(\pe4/bq[7] ), .ZN(n15771) );
  XOR2HSV0 U19047 ( .A1(n15772), .A2(n15771), .Z(n15773) );
  XOR2HSV0 U19048 ( .A1(n15774), .A2(n15773), .Z(n15775) );
  XOR2HSV0 U19049 ( .A1(n15776), .A2(n15775), .Z(n15793) );
  NAND2HSV0 U19050 ( .A1(\pe4/aot [9]), .A2(\pe4/bq[11] ), .ZN(n15778) );
  NAND2HSV0 U19051 ( .A1(n28683), .A2(\pe4/bq[4] ), .ZN(n15777) );
  XOR2HSV0 U19052 ( .A1(n15778), .A2(n15777), .Z(n15782) );
  NAND2HSV0 U19053 ( .A1(n22943), .A2(\pe4/aot [5]), .ZN(n15780) );
  NAND2HSV0 U19054 ( .A1(\pe4/aot [7]), .A2(n23076), .ZN(n15779) );
  XOR2HSV0 U19055 ( .A1(n15780), .A2(n15779), .Z(n15781) );
  XOR2HSV0 U19056 ( .A1(n15782), .A2(n15781), .Z(n15791) );
  CLKNAND2HSV0 U19057 ( .A1(n27066), .A2(\pe4/pvq [13]), .ZN(n15783) );
  XOR2HSV0 U19058 ( .A1(n15783), .A2(\pe4/phq [13]), .Z(n15789) );
  NAND2HSV0 U19059 ( .A1(\pe4/aot [12]), .A2(\pe4/bq[5] ), .ZN(n26939) );
  CLKNHSV0 U19060 ( .I(\pe4/bq[8] ), .ZN(n27100) );
  CLKNHSV0 U19061 ( .I(\pe4/aot [12]), .ZN(n15785) );
  CLKNAND2HSV0 U19062 ( .A1(n15784), .A2(\pe4/bq[5] ), .ZN(n26942) );
  OAI21HSV0 U19063 ( .A1(n27100), .A2(n15785), .B(n26942), .ZN(n15786) );
  OAI21HSV0 U19064 ( .A1(n26939), .A2(n15787), .B(n15786), .ZN(n15788) );
  XOR2HSV0 U19065 ( .A1(n15789), .A2(n15788), .Z(n15790) );
  XNOR2HSV1 U19066 ( .A1(n15791), .A2(n15790), .ZN(n15792) );
  XNOR2HSV1 U19067 ( .A1(n15793), .A2(n15792), .ZN(n15794) );
  XOR2HSV0 U19068 ( .A1(n15795), .A2(n15794), .Z(n15796) );
  XOR2HSV0 U19069 ( .A1(n15797), .A2(n15796), .Z(n15799) );
  NAND2HSV0 U19070 ( .A1(n27830), .A2(\pe4/got [9]), .ZN(n15798) );
  XOR3HSV2 U19071 ( .A1(n15800), .A2(n15799), .A3(n15798), .Z(n15801) );
  XNOR2HSV1 U19072 ( .A1(n15802), .A2(n15801), .ZN(n15803) );
  XNOR2HSV1 U19073 ( .A1(n15804), .A2(n15803), .ZN(n15807) );
  INHSV1 U19074 ( .I(n15807), .ZN(n15805) );
  CLKNAND2HSV2 U19075 ( .A1(n15806), .A2(n15805), .ZN(n15810) );
  CLKNAND2HSV1 U19076 ( .A1(n15808), .A2(n15807), .ZN(n15809) );
  INHSV2 U19077 ( .I(n15844), .ZN(n15811) );
  CLKAND2HSV2 U19078 ( .A1(n15693), .A2(\pe4/ti_7t [10]), .Z(n15814) );
  INHSV2 U19079 ( .I(n15814), .ZN(n15812) );
  NAND2HSV2 U19080 ( .A1(n15811), .A2(n15812), .ZN(n15820) );
  AND2HSV2 U19081 ( .A1(n15822), .A2(n15824), .Z(n15818) );
  CLKAND2HSV1 U19082 ( .A1(n15823), .A2(n15812), .Z(n15817) );
  NOR2HSV1 U19083 ( .A1(n15752), .A2(n15451), .ZN(n15815) );
  NOR2HSV2 U19084 ( .A1(n15815), .A2(n15814), .ZN(n15816) );
  AOI21HSV2 U19085 ( .A1(n15818), .A2(n15817), .B(n15816), .ZN(n15819) );
  CLKNAND2HSV1 U19086 ( .A1(n15820), .A2(n15819), .ZN(n15829) );
  NOR2HSV2 U19087 ( .A1(n15821), .A2(n15451), .ZN(n21744) );
  CLKNHSV0 U19088 ( .I(n15822), .ZN(n15826) );
  NAND3HSV2 U19089 ( .A1(n15824), .A2(n15823), .A3(n26923), .ZN(n15825) );
  NOR2HSV2 U19090 ( .A1(n15826), .A2(n15825), .ZN(n15827) );
  INAND2HSV2 U19091 ( .A1(n21744), .B1(n15827), .ZN(n15828) );
  INHSV2 U19092 ( .I(n15833), .ZN(n15831) );
  INHSV2 U19093 ( .I(n15836), .ZN(n15843) );
  CLKNHSV1 U19094 ( .I(n21745), .ZN(n15840) );
  AOI31HSV2 U19095 ( .A1(n15840), .A2(n27784), .A3(n15839), .B(n15838), .ZN(
        n15841) );
  INAND2HSV2 U19096 ( .A1(n24311), .B1(n15844), .ZN(n15892) );
  NOR2HSV0 U19097 ( .A1(n15847), .A2(n22822), .ZN(n15848) );
  CLKNAND2HSV0 U19098 ( .A1(n15849), .A2(n15848), .ZN(n15850) );
  INHSV1 U19099 ( .I(n15850), .ZN(n15851) );
  CLKNAND2HSV1 U19100 ( .A1(n12273), .A2(n15851), .ZN(n15890) );
  NOR2HSV1 U19101 ( .A1(n26981), .A2(n27827), .ZN(n15886) );
  NAND2HSV0 U19102 ( .A1(n22827), .A2(\pe4/got [9]), .ZN(n15883) );
  NAND2HSV0 U19103 ( .A1(n15640), .A2(n14000), .ZN(n15856) );
  NAND2HSV0 U19104 ( .A1(n23482), .A2(n22826), .ZN(n15855) );
  XNOR2HSV1 U19105 ( .A1(n15856), .A2(n15855), .ZN(n15881) );
  NAND2HSV0 U19106 ( .A1(\pe4/aot [5]), .A2(n26948), .ZN(n15858) );
  NAND2HSV0 U19107 ( .A1(\pe4/got [5]), .A2(n27128), .ZN(n15857) );
  XOR2HSV0 U19108 ( .A1(n15858), .A2(n15857), .Z(n15862) );
  NAND2HSV0 U19109 ( .A1(\pe4/aot [6]), .A2(n26958), .ZN(n15860) );
  NAND2HSV0 U19110 ( .A1(\pe4/aot [7]), .A2(n27060), .ZN(n15859) );
  XOR2HSV0 U19111 ( .A1(n15860), .A2(n15859), .Z(n15861) );
  XOR2HSV0 U19112 ( .A1(n15862), .A2(n15861), .Z(n15870) );
  NAND2HSV0 U19113 ( .A1(\pe4/aot [8]), .A2(n26961), .ZN(n15864) );
  NAND2HSV0 U19114 ( .A1(\pe4/bq[7] ), .A2(\pe4/aot [14]), .ZN(n15863) );
  XOR2HSV0 U19115 ( .A1(n15864), .A2(n15863), .Z(n15868) );
  NAND2HSV0 U19116 ( .A1(\pe4/aot [9]), .A2(\pe4/bq[12] ), .ZN(n15866) );
  NAND2HSV0 U19117 ( .A1(\pe4/aot [12]), .A2(\pe4/bq[9] ), .ZN(n15865) );
  XOR2HSV0 U19118 ( .A1(n15866), .A2(n15865), .Z(n15867) );
  XOR2HSV0 U19119 ( .A1(n15868), .A2(n15867), .Z(n15869) );
  XOR2HSV0 U19120 ( .A1(n15870), .A2(n15869), .Z(n15879) );
  CLKNHSV0 U19121 ( .I(\pe4/bq[6] ), .ZN(n27846) );
  BUFHSV2 U19122 ( .I(n15871), .Z(n26940) );
  NAND2HSV0 U19123 ( .A1(n28683), .A2(\pe4/bq[5] ), .ZN(n22829) );
  CLKNHSV0 U19124 ( .I(n22838), .ZN(n15873) );
  AOI22HSV0 U19125 ( .A1(\pe4/aot [13]), .A2(\pe4/bq[8] ), .B1(\pe4/bq[11] ), 
        .B2(\pe4/aot [10]), .ZN(n15872) );
  AOI21HSV1 U19126 ( .A1(n15874), .A2(n15873), .B(n15872), .ZN(n15875) );
  NAND2HSV0 U19127 ( .A1(\pe4/aot [11]), .A2(\pe4/bq[10] ), .ZN(n27832) );
  XOR2HSV0 U19128 ( .A1(n15875), .A2(n27832), .Z(n15876) );
  XNOR2HSV1 U19129 ( .A1(n15877), .A2(n15876), .ZN(n15878) );
  XNOR2HSV1 U19130 ( .A1(n15879), .A2(n15878), .ZN(n15880) );
  XOR2HSV0 U19131 ( .A1(n15881), .A2(n15880), .Z(n15882) );
  XOR2HSV0 U19132 ( .A1(n15883), .A2(n15882), .Z(n15885) );
  NAND2HSV0 U19133 ( .A1(n28696), .A2(\pe4/got [10]), .ZN(n15884) );
  XOR3HSV2 U19134 ( .A1(n15886), .A2(n15885), .A3(n15884), .Z(n15887) );
  XNOR2HSV1 U19135 ( .A1(n15888), .A2(n15887), .ZN(n15889) );
  NAND2HSV2 U19136 ( .A1(n15892), .A2(n15893), .ZN(n15897) );
  CLKNHSV1 U19137 ( .I(n15892), .ZN(n15895) );
  INHSV2 U19138 ( .I(n15893), .ZN(n15894) );
  CLKNAND2HSV1 U19139 ( .A1(n21980), .A2(n21981), .ZN(n15899) );
  CLKNAND2HSV3 U19140 ( .A1(n21983), .A2(n21984), .ZN(n15898) );
  NOR2HSV2 U19141 ( .A1(n21977), .A2(n15900), .ZN(n15903) );
  NOR2HSV2 U19142 ( .A1(n15370), .A2(\pe4/ti_7t [12]), .ZN(n22881) );
  INHSV2 U19143 ( .I(n22881), .ZN(n15901) );
  NAND2HSV2 U19144 ( .A1(n15901), .A2(\pe4/got [16]), .ZN(n15902) );
  AOI21HSV4 U19145 ( .A1(n15903), .A2(n14080), .B(n15902), .ZN(n21967) );
  NAND2HSV4 U19146 ( .A1(n15904), .A2(n21977), .ZN(n21988) );
  CLKNAND2HSV3 U19147 ( .A1(n21967), .A2(n21988), .ZN(n21974) );
  NAND2HSV0 U19148 ( .A1(n23683), .A2(\pe3/got [11]), .ZN(n15912) );
  NOR2HSV0 U19149 ( .A1(n26241), .A2(n21720), .ZN(n15911) );
  CLKNHSV0 U19150 ( .I(n15911), .ZN(n15907) );
  NOR2HSV0 U19151 ( .A1(n15912), .A2(n15907), .ZN(n15918) );
  XNOR2HSV4 U19152 ( .A1(n15909), .A2(n15908), .ZN(n28613) );
  NOR2HSV0 U19153 ( .A1(n16016), .A2(n26241), .ZN(n15914) );
  CLKNHSV0 U19154 ( .I(n15914), .ZN(n15910) );
  CLKNAND2HSV0 U19155 ( .A1(n15912), .A2(n15910), .ZN(n15916) );
  NOR2HSV0 U19156 ( .A1(n15914), .A2(n15911), .ZN(n15913) );
  MUX2NHSV1 U19157 ( .I0(n15914), .I1(n15913), .S(n15912), .ZN(n15915) );
  OAI21HSV2 U19158 ( .A1(n28613), .A2(n15916), .B(n15915), .ZN(n15917) );
  AOI21HSV2 U19159 ( .A1(n15918), .A2(n28613), .B(n15917), .ZN(n15958) );
  INHSV2 U19160 ( .I(\pe3/got [10]), .ZN(n26645) );
  NOR2HSV2 U19161 ( .A1(n26714), .A2(n26645), .ZN(n15956) );
  NAND2HSV0 U19162 ( .A1(n15240), .A2(n26642), .ZN(n15954) );
  NAND2HSV0 U19163 ( .A1(n26367), .A2(\pe3/got [6]), .ZN(n15950) );
  CLKNAND2HSV0 U19164 ( .A1(n26350), .A2(\pe3/got [7]), .ZN(n15949) );
  NAND2HSV0 U19165 ( .A1(\pe3/aot [9]), .A2(\pe3/bq[12] ), .ZN(n15921) );
  NAND2HSV0 U19166 ( .A1(\pe3/aot [7]), .A2(\pe3/bq[14] ), .ZN(n15920) );
  XOR2HSV0 U19167 ( .A1(n15921), .A2(n15920), .Z(n15925) );
  NAND2HSV0 U19168 ( .A1(\pe3/aot [5]), .A2(n26351), .ZN(n15923) );
  NAND2HSV0 U19169 ( .A1(\pe3/bq[5] ), .A2(n14040), .ZN(n15922) );
  XOR2HSV0 U19170 ( .A1(n15923), .A2(n15922), .Z(n15924) );
  XOR2HSV0 U19171 ( .A1(n15925), .A2(n15924), .Z(n15933) );
  NAND2HSV0 U19172 ( .A1(n11932), .A2(\pe3/bq[8] ), .ZN(n15927) );
  NAND2HSV0 U19173 ( .A1(\pe3/aot [14]), .A2(\pe3/bq[7] ), .ZN(n15926) );
  XOR2HSV0 U19174 ( .A1(n15927), .A2(n15926), .Z(n15931) );
  NAND2HSV0 U19175 ( .A1(\pe3/aot [12]), .A2(\pe3/bq[9] ), .ZN(n15929) );
  NAND2HSV0 U19176 ( .A1(\pe3/aot [8]), .A2(\pe3/bq[13] ), .ZN(n15928) );
  XOR2HSV0 U19177 ( .A1(n15929), .A2(n15928), .Z(n15930) );
  XOR2HSV0 U19178 ( .A1(n15931), .A2(n15930), .Z(n15932) );
  XOR2HSV0 U19179 ( .A1(n15933), .A2(n15932), .Z(n15947) );
  INHSV2 U19180 ( .I(n23329), .ZN(n26603) );
  NAND2HSV0 U19181 ( .A1(n26603), .A2(n26380), .ZN(n15935) );
  NAND2HSV0 U19182 ( .A1(\pe3/aot [15]), .A2(\pe3/bq[6] ), .ZN(n15934) );
  XOR2HSV0 U19183 ( .A1(n15935), .A2(n15934), .Z(n15939) );
  CLKNHSV0 U19184 ( .I(n15936), .ZN(n15937) );
  XNOR2HSV1 U19185 ( .A1(n15939), .A2(n15938), .ZN(n15945) );
  CLKNHSV0 U19186 ( .I(\pe3/aot [6]), .ZN(n24581) );
  INHSV2 U19187 ( .I(\pe3/bq[11] ), .ZN(n24527) );
  NOR2HSV1 U19188 ( .A1(n24581), .A2(n24527), .ZN(n26370) );
  AOI22HSV0 U19189 ( .A1(\pe3/aot [10]), .A2(\pe3/bq[11] ), .B1(n26373), .B2(
        \pe3/aot [6]), .ZN(n15940) );
  AOI21HSV1 U19190 ( .A1(n26370), .A2(n15941), .B(n15940), .ZN(n15943) );
  NAND2HSV0 U19191 ( .A1(\pe3/aot [11]), .A2(\pe3/bq[10] ), .ZN(n15942) );
  XOR2HSV0 U19192 ( .A1(n15943), .A2(n15942), .Z(n15944) );
  XNOR2HSV1 U19193 ( .A1(n15945), .A2(n15944), .ZN(n15946) );
  XNOR2HSV1 U19194 ( .A1(n15947), .A2(n15946), .ZN(n15948) );
  XOR3HSV2 U19195 ( .A1(n15950), .A2(n15949), .A3(n15948), .Z(n15952) );
  NAND2HSV0 U19196 ( .A1(n28920), .A2(n28648), .ZN(n15951) );
  XNOR2HSV1 U19197 ( .A1(n15952), .A2(n15951), .ZN(n15953) );
  XNOR2HSV1 U19198 ( .A1(n15954), .A2(n15953), .ZN(n15955) );
  XOR2HSV0 U19199 ( .A1(n15956), .A2(n15955), .Z(n15957) );
  XOR2HSV0 U19200 ( .A1(n15958), .A2(n15957), .Z(n15959) );
  NAND2HSV2 U19201 ( .A1(n16021), .A2(n26413), .ZN(n15960) );
  NOR2HSV4 U19202 ( .A1(n14053), .A2(n28931), .ZN(n15966) );
  CLKNAND2HSV1 U19203 ( .A1(n15964), .A2(n26348), .ZN(n15965) );
  NOR2HSV4 U19204 ( .A1(n15966), .A2(n15965), .ZN(n15969) );
  INHSV2 U19205 ( .I(n15973), .ZN(n23667) );
  INHSV2 U19206 ( .I(n23667), .ZN(n23664) );
  NAND2HSV2 U19207 ( .A1(n28931), .A2(\pe3/ti_7t [10]), .ZN(n16107) );
  INHSV2 U19208 ( .I(n16107), .ZN(n15976) );
  NOR2HSV2 U19209 ( .A1(n16163), .A2(n23402), .ZN(n23396) );
  XNOR2HSV4 U19210 ( .A1(n15978), .A2(n15977), .ZN(n16160) );
  NAND2HSV2 U19211 ( .A1(n28432), .A2(\pe3/got [11]), .ZN(n16014) );
  NAND2HSV0 U19212 ( .A1(n28707), .A2(n11891), .ZN(n16013) );
  CLKNAND2HSV1 U19213 ( .A1(n16112), .A2(\pe3/got [10]), .ZN(n16011) );
  NAND2HSV0 U19214 ( .A1(n26367), .A2(\pe3/got [7]), .ZN(n16007) );
  CLKNAND2HSV0 U19215 ( .A1(n15979), .A2(n28648), .ZN(n16006) );
  NAND2HSV0 U19216 ( .A1(\pe3/aot [14]), .A2(\pe3/bq[8] ), .ZN(n15981) );
  NAND2HSV0 U19217 ( .A1(\pe3/bq[7] ), .A2(\pe3/aot [15]), .ZN(n15980) );
  XOR2HSV0 U19218 ( .A1(n15981), .A2(n15980), .Z(n15985) );
  NAND2HSV0 U19219 ( .A1(\pe3/aot [8]), .A2(\pe3/bq[14] ), .ZN(n15983) );
  NAND2HSV0 U19220 ( .A1(\pe3/aot [6]), .A2(n23336), .ZN(n15982) );
  XOR2HSV0 U19221 ( .A1(n15983), .A2(n15982), .Z(n15984) );
  XOR2HSV0 U19222 ( .A1(n15985), .A2(n15984), .Z(n15993) );
  NAND2HSV0 U19223 ( .A1(\pe3/aot [7]), .A2(n16115), .ZN(n15987) );
  NAND2HSV0 U19224 ( .A1(\pe3/aot [10]), .A2(\pe3/bq[12] ), .ZN(n15986) );
  XOR2HSV0 U19225 ( .A1(n15987), .A2(n15986), .Z(n15991) );
  NAND2HSV0 U19226 ( .A1(n11932), .A2(\pe3/bq[9] ), .ZN(n15989) );
  NAND2HSV0 U19227 ( .A1(\pe3/aot [12]), .A2(\pe3/bq[10] ), .ZN(n15988) );
  XOR2HSV0 U19228 ( .A1(n15989), .A2(n15988), .Z(n15990) );
  XOR2HSV0 U19229 ( .A1(n15991), .A2(n15990), .Z(n15992) );
  XOR2HSV0 U19230 ( .A1(n15993), .A2(n15992), .Z(n16004) );
  CLKNAND2HSV0 U19231 ( .A1(\pe3/aot [9]), .A2(\pe3/bq[11] ), .ZN(n16135) );
  CLKNHSV0 U19232 ( .I(\pe3/aot [9]), .ZN(n26701) );
  NAND2HSV0 U19233 ( .A1(\pe3/aot [11]), .A2(\pe3/bq[11] ), .ZN(n15994) );
  OAI21HSV0 U19234 ( .A1(n26701), .A2(n26246), .B(n15994), .ZN(n15995) );
  OAI21HSV0 U19235 ( .A1(n16135), .A2(n15996), .B(n15995), .ZN(n15997) );
  XOR2HSV0 U19236 ( .A1(n15998), .A2(n15997), .Z(n16002) );
  NAND2HSV0 U19237 ( .A1(\pe3/bq[6] ), .A2(n14040), .ZN(n16000) );
  NAND2HSV0 U19238 ( .A1(n26380), .A2(\pe3/got [6]), .ZN(n15999) );
  XOR2HSV0 U19239 ( .A1(n16000), .A2(n15999), .Z(n16001) );
  XNOR2HSV1 U19240 ( .A1(n16002), .A2(n16001), .ZN(n16003) );
  XNOR2HSV1 U19241 ( .A1(n16004), .A2(n16003), .ZN(n16005) );
  XOR3HSV2 U19242 ( .A1(n16007), .A2(n16006), .A3(n16005), .Z(n16009) );
  NAND2HSV0 U19243 ( .A1(n28920), .A2(n26642), .ZN(n16008) );
  XNOR2HSV1 U19244 ( .A1(n16009), .A2(n16008), .ZN(n16010) );
  XOR2HSV0 U19245 ( .A1(n16011), .A2(n16010), .Z(n16012) );
  AOI21HSV2 U19246 ( .A1(n16016), .A2(n16015), .B(n24313), .ZN(n16017) );
  OAI21HSV2 U19247 ( .A1(n16018), .A2(n16056), .B(n16017), .ZN(n16019) );
  NAND2HSV0 U19248 ( .A1(n16021), .A2(n28930), .ZN(n16022) );
  NOR2HSV2 U19249 ( .A1(n16022), .A2(n16023), .ZN(n16024) );
  INHSV2 U19250 ( .I(n16024), .ZN(n16025) );
  CLKNAND2HSV3 U19251 ( .A1(n16026), .A2(n16025), .ZN(n16027) );
  CLKNAND2HSV4 U19252 ( .A1(n16027), .A2(n16028), .ZN(n25353) );
  INHSV2 U19253 ( .I(n26413), .ZN(n21719) );
  NOR2HSV2 U19254 ( .A1(n25353), .A2(n21719), .ZN(n16035) );
  NOR2HSV2 U19255 ( .A1(n16054), .A2(n16029), .ZN(n16030) );
  CLKNAND2HSV1 U19256 ( .A1(n25353), .A2(n16031), .ZN(n16032) );
  CLKNAND2HSV2 U19257 ( .A1(n16033), .A2(n16032), .ZN(n16034) );
  INHSV2 U19258 ( .I(n16106), .ZN(n16037) );
  INHSV4 U19259 ( .I(n25353), .ZN(n16052) );
  INHSV2 U19260 ( .I(n16052), .ZN(n16036) );
  NAND3HSV2 U19261 ( .A1(n16050), .A2(n23414), .A3(n16049), .ZN(n16047) );
  AND2HSV2 U19262 ( .A1(n25353), .A2(n23414), .Z(n16038) );
  CLKNAND2HSV2 U19263 ( .A1(n14054), .A2(n15017), .ZN(n16039) );
  CLKNAND2HSV3 U19264 ( .A1(n16039), .A2(n23666), .ZN(n16051) );
  INHSV2 U19265 ( .I(n16051), .ZN(n16040) );
  CLKNHSV1 U19266 ( .I(\pe3/ti_7t [11]), .ZN(n16041) );
  NOR2HSV2 U19267 ( .A1(n16042), .A2(n16041), .ZN(n16043) );
  CLKAND2HSV1 U19268 ( .A1(n16054), .A2(n16043), .Z(n16044) );
  XNOR2HSV4 U19269 ( .A1(n16048), .A2(n16160), .ZN(n21312) );
  NAND2HSV2 U19270 ( .A1(n16054), .A2(\pe3/ti_7t [9]), .ZN(n16157) );
  INHSV2 U19271 ( .I(n16157), .ZN(n23374) );
  AOI21HSV1 U19272 ( .A1(n16157), .A2(n16015), .B(n26241), .ZN(n16055) );
  OAI21HSV2 U19273 ( .A1(n14054), .A2(n23374), .B(n16055), .ZN(n16105) );
  CLKNAND2HSV1 U19274 ( .A1(n28613), .A2(n23382), .ZN(n16057) );
  CLKNAND2HSV0 U19275 ( .A1(n23328), .A2(\pe3/got [10]), .ZN(n16101) );
  NAND2HSV0 U19276 ( .A1(n16112), .A2(\pe3/got [7]), .ZN(n16096) );
  NAND2HSV0 U19277 ( .A1(n26603), .A2(n26350), .ZN(n16094) );
  NAND2HSV0 U19278 ( .A1(n26242), .A2(\pe3/got [6]), .ZN(n16093) );
  NAND2HSV0 U19279 ( .A1(\pe3/aot [14]), .A2(\pe3/bq[5] ), .ZN(n16059) );
  NAND2HSV0 U19280 ( .A1(\pe3/aot [8]), .A2(\pe3/bq[11] ), .ZN(n16058) );
  XOR2HSV0 U19281 ( .A1(n16059), .A2(n16058), .Z(n16063) );
  NAND2HSV0 U19282 ( .A1(\pe3/aot [11]), .A2(\pe3/bq[8] ), .ZN(n16061) );
  NAND2HSV0 U19283 ( .A1(n11932), .A2(\pe3/bq[6] ), .ZN(n16060) );
  XOR2HSV0 U19284 ( .A1(n16061), .A2(n16060), .Z(n16062) );
  XOR2HSV0 U19285 ( .A1(n16063), .A2(n16062), .Z(n16071) );
  NAND2HSV0 U19286 ( .A1(n23543), .A2(\pe3/pvq [14]), .ZN(n16064) );
  XNOR2HSV1 U19287 ( .A1(n16064), .A2(\pe3/phq [14]), .ZN(n16069) );
  CLKNAND2HSV0 U19288 ( .A1(\pe3/aot [15]), .A2(\pe3/bq[3] ), .ZN(n23348) );
  CLKNAND2HSV0 U19289 ( .A1(n14040), .A2(\pe3/bq[4] ), .ZN(n16137) );
  NAND2HSV0 U19290 ( .A1(n14040), .A2(\pe3/bq[3] ), .ZN(n16065) );
  OAI21HSV0 U19291 ( .A1(n16066), .A2(n23349), .B(n16065), .ZN(n16067) );
  OAI21HSV1 U19292 ( .A1(n23348), .A2(n16137), .B(n16067), .ZN(n16068) );
  XOR2HSV0 U19293 ( .A1(n16069), .A2(n16068), .Z(n16070) );
  XNOR2HSV1 U19294 ( .A1(n16071), .A2(n16070), .ZN(n16073) );
  NAND2HSV0 U19295 ( .A1(n26367), .A2(\pe3/got [4]), .ZN(n16072) );
  XOR2HSV0 U19296 ( .A1(n16073), .A2(n16072), .Z(n16091) );
  NAND2HSV0 U19297 ( .A1(\pe3/aot [10]), .A2(\pe3/bq[9] ), .ZN(n16075) );
  NAND2HSV0 U19298 ( .A1(\pe3/aot [5]), .A2(\pe3/bq[14] ), .ZN(n16074) );
  XOR2HSV0 U19299 ( .A1(n16075), .A2(n16074), .Z(n16079) );
  NAND2HSV0 U19300 ( .A1(\pe3/aot [9]), .A2(\pe3/bq[10] ), .ZN(n16077) );
  NAND2HSV0 U19301 ( .A1(\pe3/aot [6]), .A2(\pe3/bq[13] ), .ZN(n16076) );
  XOR2HSV0 U19302 ( .A1(n16077), .A2(n16076), .Z(n16078) );
  XOR2HSV0 U19303 ( .A1(n16079), .A2(n16078), .Z(n16089) );
  NAND2HSV0 U19304 ( .A1(\pe3/aot [4]), .A2(n26373), .ZN(n16087) );
  NAND2HSV0 U19305 ( .A1(\pe3/bq[7] ), .A2(\pe3/aot [7]), .ZN(n24524) );
  NOR2HSV0 U19306 ( .A1(n16080), .A2(n24524), .ZN(n16082) );
  AOI22HSV0 U19307 ( .A1(\pe3/aot [12]), .A2(\pe3/bq[7] ), .B1(\pe3/bq[12] ), 
        .B2(\pe3/aot [7]), .ZN(n16081) );
  NOR2HSV2 U19308 ( .A1(n16082), .A2(n16081), .ZN(n16086) );
  NAND2HSV0 U19309 ( .A1(\pe3/aot [3]), .A2(n26351), .ZN(n16084) );
  INHSV2 U19310 ( .I(\pe3/got [3]), .ZN(n23339) );
  NAND2HSV0 U19311 ( .A1(\pe3/got [3]), .A2(n15044), .ZN(n16083) );
  XOR2HSV0 U19312 ( .A1(n16084), .A2(n16083), .Z(n16085) );
  XOR3HSV2 U19313 ( .A1(n16087), .A2(n16086), .A3(n16085), .Z(n16088) );
  XOR2HSV0 U19314 ( .A1(n16089), .A2(n16088), .Z(n16090) );
  XNOR2HSV1 U19315 ( .A1(n16091), .A2(n16090), .ZN(n16092) );
  XOR3HSV1 U19316 ( .A1(n16094), .A2(n16093), .A3(n16092), .Z(n16095) );
  XNOR2HSV1 U19317 ( .A1(n16096), .A2(n16095), .ZN(n16099) );
  CLKBUFHSV4 U19318 ( .I(n23683), .Z(n26682) );
  NOR2HSV0 U19319 ( .A1(n26714), .A2(n26601), .ZN(n16097) );
  XNOR2HSV1 U19320 ( .A1(n16101), .A2(n16100), .ZN(n16102) );
  XNOR2HSV1 U19321 ( .A1(n16103), .A2(n16102), .ZN(n16104) );
  CLKNAND2HSV2 U19322 ( .A1(n16106), .A2(n23664), .ZN(n16108) );
  MUX2NHSV2 U19323 ( .I0(n16109), .I1(n16172), .S(n16167), .ZN(n16162) );
  CLKNAND2HSV0 U19324 ( .A1(n28432), .A2(n26642), .ZN(n16150) );
  NAND2HSV0 U19325 ( .A1(n16112), .A2(n28648), .ZN(n16148) );
  NAND2HSV0 U19326 ( .A1(n26350), .A2(\pe3/got [6]), .ZN(n16146) );
  NAND2HSV0 U19327 ( .A1(n28920), .A2(\pe3/got [7]), .ZN(n16145) );
  NAND2HSV0 U19328 ( .A1(n11932), .A2(\pe3/bq[7] ), .ZN(n16114) );
  NAND2HSV0 U19329 ( .A1(\pe3/bq[5] ), .A2(\pe3/aot [15]), .ZN(n16113) );
  XOR2HSV0 U19330 ( .A1(n16114), .A2(n16113), .Z(n16119) );
  NAND2HSV0 U19331 ( .A1(\pe3/aot [12]), .A2(\pe3/bq[8] ), .ZN(n16117) );
  NAND2HSV0 U19332 ( .A1(\pe3/aot [5]), .A2(n16115), .ZN(n16116) );
  XOR2HSV0 U19333 ( .A1(n16117), .A2(n16116), .Z(n16118) );
  XOR2HSV0 U19334 ( .A1(n16119), .A2(n16118), .Z(n16126) );
  NAND2HSV0 U19335 ( .A1(\pe3/aot [10]), .A2(\pe3/bq[10] ), .ZN(n16121) );
  NAND2HSV0 U19336 ( .A1(\pe3/aot [14]), .A2(\pe3/bq[6] ), .ZN(n16120) );
  XOR2HSV0 U19337 ( .A1(n16121), .A2(n16120), .Z(n16124) );
  NAND2HSV0 U19338 ( .A1(n23516), .A2(\pe3/pvq [13]), .ZN(n16122) );
  XOR2HSV0 U19339 ( .A1(n16122), .A2(\pe3/phq [13]), .Z(n16123) );
  XOR2HSV0 U19340 ( .A1(n16124), .A2(n16123), .Z(n16125) );
  XOR2HSV0 U19341 ( .A1(n16126), .A2(n16125), .Z(n16128) );
  NAND2HSV0 U19342 ( .A1(n26603), .A2(n26367), .ZN(n16127) );
  XNOR2HSV1 U19343 ( .A1(n16128), .A2(n16127), .ZN(n16143) );
  NAND2HSV0 U19344 ( .A1(\pe3/aot [7]), .A2(\pe3/bq[13] ), .ZN(n16130) );
  NAND2HSV0 U19345 ( .A1(\pe3/aot [6]), .A2(\pe3/bq[14] ), .ZN(n16129) );
  XOR2HSV0 U19346 ( .A1(n16130), .A2(n16129), .Z(n16134) );
  NAND2HSV0 U19347 ( .A1(\pe3/aot [4]), .A2(n23336), .ZN(n16132) );
  NAND2HSV0 U19348 ( .A1(\pe3/aot [8]), .A2(\pe3/bq[12] ), .ZN(n16131) );
  XOR2HSV0 U19349 ( .A1(n16132), .A2(n16131), .Z(n16133) );
  XOR2HSV0 U19350 ( .A1(n16134), .A2(n16133), .Z(n16141) );
  NAND2HSV0 U19351 ( .A1(\pe3/bq[9] ), .A2(\pe3/aot [11]), .ZN(n26684) );
  XOR2HSV0 U19352 ( .A1(n16135), .A2(n26684), .Z(n16139) );
  NAND2HSV0 U19353 ( .A1(\pe3/got [4]), .A2(n26380), .ZN(n16136) );
  XOR2HSV0 U19354 ( .A1(n16137), .A2(n16136), .Z(n16138) );
  XOR2HSV0 U19355 ( .A1(n16139), .A2(n16138), .Z(n16140) );
  XOR2HSV0 U19356 ( .A1(n16141), .A2(n16140), .Z(n16142) );
  XNOR2HSV1 U19357 ( .A1(n16143), .A2(n16142), .ZN(n16144) );
  XOR3HSV1 U19358 ( .A1(n16146), .A2(n16145), .A3(n16144), .Z(n16147) );
  XNOR2HSV1 U19359 ( .A1(n16148), .A2(n16147), .ZN(n16149) );
  XOR2HSV2 U19360 ( .A1(n16150), .A2(n16149), .Z(n16152) );
  NAND2HSV0 U19361 ( .A1(n26682), .A2(\pe3/got [10]), .ZN(n16151) );
  XNOR2HSV4 U19362 ( .A1(n16152), .A2(n16151), .ZN(n16154) );
  XOR2HSV2 U19363 ( .A1(n16154), .A2(n16153), .Z(n16155) );
  AOI21HSV2 U19364 ( .A1(n16157), .A2(n16015), .B(n24313), .ZN(n16158) );
  INHSV4 U19365 ( .I(n26291), .ZN(n24516) );
  CLKNAND2HSV2 U19366 ( .A1(n16160), .A2(n23664), .ZN(n21730) );
  NOR2HSV2 U19367 ( .A1(n16160), .A2(n16163), .ZN(n16169) );
  NOR2HSV1 U19368 ( .A1(n24516), .A2(n16169), .ZN(n21727) );
  NAND2HSV4 U19369 ( .A1(n21732), .A2(n16161), .ZN(n23439) );
  CLKNAND2HSV3 U19370 ( .A1(n16162), .A2(n23439), .ZN(n23419) );
  INHSV2 U19371 ( .I(\pe3/ti_7t [13]), .ZN(n21724) );
  AOI21HSV2 U19372 ( .A1(n21724), .A2(n16163), .B(n21719), .ZN(n16179) );
  INHSV2 U19373 ( .I(n16179), .ZN(n23441) );
  OR2HSV1 U19374 ( .A1(n23441), .A2(n16164), .Z(n16165) );
  INHSV2 U19375 ( .I(n21730), .ZN(n16168) );
  CLKNAND2HSV0 U19376 ( .A1(n26291), .A2(n16169), .ZN(n23395) );
  XNOR2HSV4 U19377 ( .A1(n16174), .A2(n16173), .ZN(n23442) );
  NAND2HSV2 U19378 ( .A1(n28931), .A2(\pe3/ti_7t [14]), .ZN(n16178) );
  NAND2HSV2 U19379 ( .A1(n16175), .A2(n21722), .ZN(n16177) );
  INHSV2 U19380 ( .I(n23442), .ZN(n16176) );
  NOR2HSV4 U19381 ( .A1(n16177), .A2(n16176), .ZN(n23416) );
  AND2HSV2 U19382 ( .A1(n16179), .A2(n16178), .Z(n16180) );
  NAND3HSV4 U19383 ( .A1(n23440), .A2(n23439), .A3(n16180), .ZN(n23415) );
  OAI21HSV4 U19384 ( .A1(n23417), .A2(n23416), .B(n23415), .ZN(n16181) );
  OAI21HSV4 U19385 ( .A1(n23419), .A2(n23420), .B(n16181), .ZN(n28801) );
  INHSV2 U19386 ( .I(ctro1), .ZN(n17296) );
  INHSV2 U19387 ( .I(n17359), .ZN(n16182) );
  NAND2HSV2 U19388 ( .A1(n16182), .A2(\pe1/ti_7t [6]), .ZN(n17170) );
  CLKNHSV0 U19389 ( .I(n17170), .ZN(n16256) );
  CLKBUFHSV4 U19390 ( .I(n16184), .Z(n17615) );
  CLKNAND2HSV3 U19391 ( .A1(n29050), .A2(n17478), .ZN(n16183) );
  INHSV2 U19392 ( .I(n17615), .ZN(n16240) );
  NAND2HSV2 U19393 ( .A1(n16240), .A2(\pe1/ti_7t [3]), .ZN(n16239) );
  NAND2HSV3 U19394 ( .A1(n17172), .A2(\pe1/got [14]), .ZN(n16208) );
  CLKNAND2HSV2 U19395 ( .A1(n29052), .A2(n16184), .ZN(n17155) );
  CLKNAND2HSV1 U19396 ( .A1(n17155), .A2(n17154), .ZN(n16245) );
  INHSV3 U19397 ( .I(\pe1/got [12]), .ZN(n26417) );
  CLKNAND2HSV1 U19398 ( .A1(n16245), .A2(n28425), .ZN(n16189) );
  INHSV2 U19399 ( .I(\pe1/aot [12]), .ZN(n26555) );
  INHSV2 U19400 ( .I(n26431), .ZN(n17317) );
  NOR2HSV2 U19401 ( .A1(n26555), .A2(n17317), .ZN(n16187) );
  NAND2HSV0 U19402 ( .A1(\pe1/aot [14]), .A2(\pe1/bq[13] ), .ZN(n16186) );
  XOR2HSV0 U19403 ( .A1(n16187), .A2(n16186), .Z(n16188) );
  XNOR2HSV1 U19404 ( .A1(n16189), .A2(n16188), .ZN(n16196) );
  BUFHSV4 U19405 ( .I(\pe1/bq[16] ), .Z(n26436) );
  NAND2HSV0 U19406 ( .A1(\pe1/aot [11]), .A2(n26436), .ZN(n16191) );
  NAND2HSV0 U19407 ( .A1(\pe1/aot [13]), .A2(\pe1/bq[14] ), .ZN(n16190) );
  XOR2HSV0 U19408 ( .A1(n16191), .A2(n16190), .Z(n16194) );
  INHSV2 U19409 ( .I(\pe1/bq[11] ), .ZN(n17142) );
  NAND2HSV2 U19410 ( .A1(\pe1/bq[11] ), .A2(n28468), .ZN(n16273) );
  NAND2HSV0 U19411 ( .A1(\pe1/aot [16]), .A2(\pe1/bq[12] ), .ZN(n16272) );
  INHSV4 U19412 ( .I(\pe1/bq[12] ), .ZN(n27070) );
  OAI22HSV0 U19413 ( .A1(n27070), .A2(n17374), .B1(n17373), .B2(n17142), .ZN(
        n16192) );
  OAI21HSV1 U19414 ( .A1(n16273), .A2(n16272), .B(n16192), .ZN(n16193) );
  XNOR2HSV1 U19415 ( .A1(n16194), .A2(n16193), .ZN(n16195) );
  XNOR2HSV1 U19416 ( .A1(n16196), .A2(n16195), .ZN(n16206) );
  INHSV2 U19417 ( .I(n16197), .ZN(n25627) );
  INHSV2 U19418 ( .I(n16198), .ZN(n17605) );
  OAI21HSV4 U19419 ( .A1(n25627), .A2(n17605), .B(n16202), .ZN(n17139) );
  BUFHSV3 U19420 ( .I(n17139), .Z(n26562) );
  CLKNAND2HSV2 U19421 ( .A1(n26562), .A2(\pe1/got [13]), .ZN(n16203) );
  CLKNHSV2 U19422 ( .I(n16203), .ZN(n16204) );
  CLKNAND2HSV2 U19423 ( .A1(n16206), .A2(n16204), .ZN(n16205) );
  INHSV2 U19424 ( .I(n17615), .ZN(n16230) );
  CLKNAND2HSV2 U19425 ( .A1(n12023), .A2(n17230), .ZN(n16215) );
  CLKNAND2HSV1 U19426 ( .A1(n16215), .A2(n16216), .ZN(n16209) );
  XNOR2HSV4 U19427 ( .A1(n16209), .A2(n16214), .ZN(n16210) );
  NOR2HSV4 U19428 ( .A1(n16210), .A2(n16240), .ZN(n16212) );
  NAND2HSV2 U19429 ( .A1(n16212), .A2(n16211), .ZN(n16232) );
  CLKNHSV0 U19430 ( .I(\pe1/ti_7t [3]), .ZN(n16213) );
  AOI21HSV2 U19431 ( .A1(n16213), .A2(n16185), .B(n17598), .ZN(n16231) );
  CLKNAND2HSV0 U19432 ( .A1(n26444), .A2(n17296), .ZN(n16218) );
  XOR3HSV2 U19433 ( .A1(n16216), .A2(n16215), .A3(n16214), .Z(n16217) );
  NOR2HSV2 U19434 ( .A1(n16218), .A2(n16217), .ZN(n16233) );
  NOR2HSV4 U19435 ( .A1(n23478), .A2(n16230), .ZN(n16229) );
  NAND2HSV0 U19436 ( .A1(\pe1/bq[13] ), .A2(\pe1/aot [16]), .ZN(n16221) );
  NAND2HSV0 U19437 ( .A1(\pe1/bq[14] ), .A2(\pe1/aot [15]), .ZN(n16220) );
  XOR2HSV0 U19438 ( .A1(n16221), .A2(n16220), .Z(n16224) );
  CLKNAND2HSV2 U19439 ( .A1(\pe1/aot [13]), .A2(\pe1/bq[16] ), .ZN(n17304) );
  XOR2HSV2 U19440 ( .A1(n16222), .A2(n17304), .Z(n16223) );
  CLKXOR2HSV4 U19441 ( .A1(n16224), .A2(n16223), .Z(n16226) );
  NAND2HSV2 U19442 ( .A1(n28622), .A2(\pe1/got [14]), .ZN(n16225) );
  XNOR2HSV4 U19443 ( .A1(n16226), .A2(n16225), .ZN(n16228) );
  CLKNAND2HSV3 U19444 ( .A1(n17139), .A2(n14056), .ZN(n16227) );
  XNOR2HSV4 U19445 ( .A1(n16228), .A2(n16227), .ZN(n23479) );
  AOI22HSV4 U19446 ( .A1(n16230), .A2(\pe1/ti_7t [4]), .B1(n16229), .B2(n23479), .ZN(n16237) );
  INHSV2 U19447 ( .I(n23479), .ZN(n16236) );
  NAND3HSV2 U19448 ( .A1(n16232), .A2(n16231), .A3(n17296), .ZN(n16234) );
  NOR2HSV2 U19449 ( .A1(n16234), .A2(n16233), .ZN(n16235) );
  CLKNAND2HSV2 U19450 ( .A1(n16281), .A2(n14056), .ZN(n16238) );
  BUFHSV2 U19451 ( .I(n17296), .Z(n17478) );
  INHSV2 U19452 ( .I(n17478), .ZN(n17235) );
  NOR2HSV4 U19453 ( .A1(n25653), .A2(n17235), .ZN(n16286) );
  CLKNHSV0 U19454 ( .I(n16239), .ZN(n16242) );
  AOI21HSV0 U19455 ( .A1(n16240), .A2(n16239), .B(n26536), .ZN(n16241) );
  OAI21HSV2 U19456 ( .A1(n29050), .A2(n16242), .B(n16241), .ZN(n16253) );
  NAND2HSV0 U19457 ( .A1(\pe1/aot [12]), .A2(n26436), .ZN(n16243) );
  NOR2HSV2 U19458 ( .A1(n26555), .A2(n27070), .ZN(n17188) );
  AOI22HSV0 U19459 ( .A1(n16272), .A2(n16243), .B1(n12023), .B2(n17188), .ZN(
        n16244) );
  XOR2HSV0 U19460 ( .A1(n16244), .A2(n17432), .Z(n16252) );
  NAND2HSV0 U19461 ( .A1(\pe1/bq[15] ), .A2(\pe1/aot [13]), .ZN(n16247) );
  NAND2HSV0 U19462 ( .A1(n28468), .A2(\pe1/bq[13] ), .ZN(n16246) );
  XOR2HSV0 U19463 ( .A1(n16247), .A2(n16246), .Z(n16248) );
  XNOR2HSV1 U19464 ( .A1(n16249), .A2(n16248), .ZN(n16251) );
  CLKNAND2HSV1 U19465 ( .A1(n17139), .A2(\pe1/got [14]), .ZN(n16250) );
  CLKNAND2HSV2 U19466 ( .A1(n16281), .A2(n17617), .ZN(n16257) );
  XNOR2HSV4 U19467 ( .A1(n16258), .A2(n16257), .ZN(pov1[5]) );
  INHSV1 U19468 ( .I(pov1[5]), .ZN(n16255) );
  NAND2HSV0 U19469 ( .A1(n17170), .A2(n17617), .ZN(n16254) );
  OAI22HSV2 U19470 ( .A1(n16256), .A2(n16286), .B1(n16255), .B2(n16254), .ZN(
        n16259) );
  XNOR2HSV4 U19471 ( .A1(n16258), .A2(n16257), .ZN(n17215) );
  INHSV2 U19472 ( .I(n16260), .ZN(n28418) );
  INHSV2 U19473 ( .I(n16185), .ZN(n17543) );
  CLKNHSV0 U19474 ( .I(\pe1/ti_7t [5]), .ZN(n16261) );
  AOI21HSV2 U19475 ( .A1(n16261), .A2(n16240), .B(n26536), .ZN(n16262) );
  OAI21HSV4 U19476 ( .A1(pov1[5]), .A2(n16182), .B(n16262), .ZN(n16290) );
  NAND2HSV0 U19477 ( .A1(n17172), .A2(\pe1/got [13]), .ZN(n16280) );
  NAND2HSV2 U19478 ( .A1(n28425), .A2(n28814), .ZN(n16270) );
  NAND2HSV0 U19479 ( .A1(\pe1/aot [12]), .A2(\pe1/bq[14] ), .ZN(n16264) );
  CLKBUFHSV4 U19480 ( .I(\pe1/bq[15] ), .Z(n26548) );
  NAND2HSV0 U19481 ( .A1(\pe1/aot [11]), .A2(n26548), .ZN(n16263) );
  XOR2HSV0 U19482 ( .A1(n16264), .A2(n16263), .Z(n16268) );
  NAND2HSV0 U19483 ( .A1(\pe1/aot [13]), .A2(\pe1/bq[13] ), .ZN(n16266) );
  NAND2HSV0 U19484 ( .A1(\pe1/aot [10]), .A2(n26436), .ZN(n16265) );
  XOR2HSV0 U19485 ( .A1(n16266), .A2(n16265), .Z(n16267) );
  XOR2HSV0 U19486 ( .A1(n16268), .A2(n16267), .Z(n16269) );
  CLKXOR2HSV2 U19487 ( .A1(n16270), .A2(n16269), .Z(n16278) );
  NAND2HSV0 U19488 ( .A1(\pe1/aot [14]), .A2(\pe1/bq[10] ), .ZN(n17174) );
  CLKNHSV0 U19489 ( .I(\pe1/aot [14]), .ZN(n17555) );
  OAI21HSV2 U19490 ( .A1(n27070), .A2(n17555), .B(n17149), .ZN(n16271) );
  OAI21HSV1 U19491 ( .A1(n17174), .A2(n16272), .B(n16271), .ZN(n16274) );
  XNOR2HSV1 U19492 ( .A1(n16274), .A2(n16273), .ZN(n16276) );
  NAND2HSV0 U19493 ( .A1(n28622), .A2(\pe1/got [11]), .ZN(n16275) );
  XOR2HSV0 U19494 ( .A1(n16276), .A2(n16275), .Z(n16277) );
  XNOR2HSV4 U19495 ( .A1(n16280), .A2(n16279), .ZN(n16283) );
  BUFHSV8 U19496 ( .I(n16281), .Z(n17265) );
  CLKNAND2HSV1 U19497 ( .A1(n17265), .A2(\pe1/got [14]), .ZN(n16282) );
  CLKXOR2HSV4 U19498 ( .A1(n16283), .A2(n16282), .Z(n16289) );
  XNOR2HSV4 U19499 ( .A1(n16290), .A2(n16289), .ZN(n16285) );
  INHSV2 U19500 ( .I(n28422), .ZN(n17287) );
  NAND2HSV4 U19501 ( .A1(n17225), .A2(n17223), .ZN(n17286) );
  NOR2HSV2 U19502 ( .A1(n16288), .A2(n17199), .ZN(n17222) );
  OAI21HSV4 U19503 ( .A1(n17222), .A2(n17598), .B(n16285), .ZN(n17279) );
  NAND2HSV2 U19504 ( .A1(n17286), .A2(n17279), .ZN(n16291) );
  INHSV4 U19505 ( .I(n16291), .ZN(pov1[7]) );
  NAND3HSV2 U19506 ( .A1(n16292), .A2(n16464), .A3(\pe8/aot [16]), .ZN(n16293)
         );
  NAND2HSV4 U19507 ( .A1(n16293), .A2(n16294), .ZN(n16309) );
  XNOR2HSV4 U19508 ( .A1(n16309), .A2(n16310), .ZN(n16343) );
  INHSV4 U19509 ( .I(ctro8), .ZN(n19902) );
  INHSV2 U19510 ( .I(n19902), .ZN(n16304) );
  INHSV4 U19511 ( .I(ctro8), .ZN(n16331) );
  CLKNHSV2 U19512 ( .I(n16331), .ZN(n18788) );
  NAND2HSV2 U19513 ( .A1(n18788), .A2(\pe8/ti_7t [1]), .ZN(n16295) );
  CLKNAND2HSV4 U19514 ( .A1(n16296), .A2(n16295), .ZN(n16557) );
  NAND2HSV2 U19515 ( .A1(\pe8/bq[14] ), .A2(\pe8/aot [16]), .ZN(n16297) );
  NAND2HSV2 U19516 ( .A1(\pe8/ctrq ), .A2(\pe8/pvq [3]), .ZN(n16299) );
  NAND2HSV0 U19517 ( .A1(\pe8/aot [14]), .A2(n16464), .ZN(n16303) );
  NAND2HSV0 U19518 ( .A1(\pe8/aot [15]), .A2(n16400), .ZN(n16302) );
  XNOR2HSV4 U19519 ( .A1(n16306), .A2(n16305), .ZN(n21328) );
  INHSV3 U19520 ( .I(n16304), .ZN(n22129) );
  INHSV2 U19521 ( .I(n18766), .ZN(n18784) );
  INHSV2 U19522 ( .I(\pe8/got [16]), .ZN(n19972) );
  CLKBUFHSV4 U19523 ( .I(n16331), .Z(n16554) );
  NOR2HSV4 U19524 ( .A1(n16312), .A2(n20058), .ZN(n16316) );
  INHSV2 U19525 ( .I(\pe8/phq [2]), .ZN(n16314) );
  XNOR2HSV4 U19526 ( .A1(n16316), .A2(n16315), .ZN(n16319) );
  NAND2HSV2 U19527 ( .A1(\pe8/aot [16]), .A2(n16400), .ZN(n16318) );
  NAND2HSV2 U19528 ( .A1(\pe8/aot [15]), .A2(n28663), .ZN(n16317) );
  CLKXOR2HSV2 U19529 ( .A1(n16318), .A2(n16317), .Z(n16320) );
  NAND2HSV2 U19530 ( .A1(n16319), .A2(n16320), .ZN(n16324) );
  INHSV3 U19531 ( .I(n16319), .ZN(n16322) );
  INHSV2 U19532 ( .I(n16320), .ZN(n16321) );
  NAND2HSV4 U19533 ( .A1(n16322), .A2(n16321), .ZN(n16323) );
  CLKNAND2HSV4 U19534 ( .A1(n16323), .A2(n16324), .ZN(n27226) );
  CLKAND2HSV2 U19535 ( .A1(n19969), .A2(\pe8/ti_7t [2]), .Z(n16325) );
  AOI21HSV4 U19536 ( .A1(n16326), .A2(n27226), .B(n16325), .ZN(n16330) );
  INHSV2 U19537 ( .I(n29012), .ZN(n16327) );
  BUFHSV4 U19538 ( .I(n19902), .Z(n18783) );
  INAND2HSV4 U19539 ( .A1(n19972), .B1(n18783), .ZN(n16353) );
  CLKNAND2HSV4 U19540 ( .A1(n16381), .A2(n16311), .ZN(n16394) );
  INHSV2 U19541 ( .I(n16394), .ZN(n16354) );
  CLKNAND2HSV1 U19542 ( .A1(n16354), .A2(n18787), .ZN(n16339) );
  NAND2HSV2 U19543 ( .A1(n16394), .A2(n18787), .ZN(n16332) );
  INHSV2 U19544 ( .I(n16332), .ZN(n16337) );
  INHSV2 U19545 ( .I(n28646), .ZN(n20049) );
  NAND2HSV2 U19546 ( .A1(n16343), .A2(n20049), .ZN(n16333) );
  AOI21HSV4 U19547 ( .A1(n16334), .A2(n16333), .B(n16304), .ZN(n16335) );
  OAI21HSV4 U19548 ( .A1(n16336), .A2(n21328), .B(n16335), .ZN(n16360) );
  BUFHSV4 U19549 ( .I(\pe8/got [16]), .Z(n19835) );
  INHSV2 U19550 ( .I(n19902), .ZN(n19986) );
  NOR2HSV2 U19551 ( .A1(n19835), .A2(n19986), .ZN(n19822) );
  AOI21HSV4 U19552 ( .A1(n16337), .A2(n16360), .B(n19822), .ZN(n16338) );
  OAI21HSV4 U19553 ( .A1(n16358), .A2(n16339), .B(n16338), .ZN(n16352) );
  NAND2HSV2 U19554 ( .A1(n16400), .A2(\pe8/aot [14]), .ZN(n16342) );
  NAND2HSV2 U19555 ( .A1(n16464), .A2(\pe8/aot [13]), .ZN(n16341) );
  CLKBUFHSV4 U19556 ( .I(\pe8/bq[14] ), .Z(n23627) );
  NOR2HSV4 U19557 ( .A1(n16343), .A2(n19986), .ZN(n16416) );
  INHSV2 U19558 ( .I(\pe8/got [14]), .ZN(n19987) );
  INHSV2 U19559 ( .I(n19987), .ZN(n16418) );
  CLKNAND2HSV1 U19560 ( .A1(n16414), .A2(n16418), .ZN(n16344) );
  NOR2HSV4 U19561 ( .A1(n16416), .A2(n16344), .ZN(n16345) );
  INHSV2 U19562 ( .I(n28646), .ZN(n28625) );
  NAND2HSV2 U19563 ( .A1(n16381), .A2(n28625), .ZN(n16347) );
  NAND2HSV2 U19564 ( .A1(n16346), .A2(n16347), .ZN(n16351) );
  INHSV2 U19565 ( .I(n16347), .ZN(n16348) );
  CLKNAND2HSV4 U19566 ( .A1(n16351), .A2(n16350), .ZN(n22092) );
  NAND2HSV4 U19567 ( .A1(n16352), .A2(n22092), .ZN(n16455) );
  NAND2HSV2 U19568 ( .A1(n16504), .A2(\pe8/ti_7t [4]), .ZN(n16452) );
  CLKNAND2HSV4 U19569 ( .A1(n16455), .A2(n16452), .ZN(n16423) );
  NOR2HSV4 U19570 ( .A1(n22092), .A2(n16353), .ZN(n16356) );
  INHSV2 U19571 ( .I(n16394), .ZN(n21330) );
  INHSV4 U19572 ( .I(n16360), .ZN(n16397) );
  INAND2HSV4 U19573 ( .A1(n16354), .B1(n16397), .ZN(n16463) );
  CLKNAND2HSV3 U19574 ( .A1(n16462), .A2(n16463), .ZN(n16355) );
  CLKNHSV6 U19575 ( .I(n16454), .ZN(n16424) );
  NOR2HSV4 U19576 ( .A1(n16423), .A2(n16424), .ZN(n16535) );
  NAND2HSV2 U19577 ( .A1(n19969), .A2(\pe8/ti_7t [3]), .ZN(n16392) );
  CLKNAND2HSV1 U19578 ( .A1(n21330), .A2(n16392), .ZN(n16357) );
  INHSV2 U19579 ( .I(\pe8/got [14]), .ZN(n18760) );
  INHSV2 U19580 ( .I(n18760), .ZN(n28599) );
  NAND2HSV0 U19581 ( .A1(n16394), .A2(n16392), .ZN(n16359) );
  CLKNHSV1 U19582 ( .I(n16359), .ZN(n16361) );
  NAND2HSV2 U19583 ( .A1(n16361), .A2(n16360), .ZN(n16362) );
  INHSV2 U19584 ( .I(n16362), .ZN(n16363) );
  NAND2HSV0 U19585 ( .A1(\pe8/aot [14]), .A2(\pe8/bq[13] ), .ZN(n16365) );
  XNOR2HSV4 U19586 ( .A1(n16367), .A2(\pe8/phq [6]), .ZN(n16369) );
  CLKNAND2HSV0 U19587 ( .A1(n23627), .A2(\pe8/aot [13]), .ZN(n16368) );
  XNOR2HSV4 U19588 ( .A1(n16369), .A2(n16368), .ZN(n16377) );
  NAND2HSV0 U19589 ( .A1(n16400), .A2(\pe8/aot [12]), .ZN(n16371) );
  NAND2HSV0 U19590 ( .A1(\pe8/aot [16]), .A2(\pe8/bq[11] ), .ZN(n16370) );
  XOR2HSV0 U19591 ( .A1(n16371), .A2(n16370), .Z(n16375) );
  NAND2HSV0 U19592 ( .A1(\pe8/aot [11]), .A2(n16464), .ZN(n16373) );
  XOR2HSV0 U19593 ( .A1(n16373), .A2(n16372), .Z(n16374) );
  XOR2HSV0 U19594 ( .A1(n16375), .A2(n16374), .Z(n16376) );
  XOR3HSV2 U19595 ( .A1(n16378), .A2(n16377), .A3(n16376), .Z(n16380) );
  NAND2HSV0 U19596 ( .A1(n16557), .A2(\pe8/got [12]), .ZN(n16379) );
  XNOR2HSV4 U19597 ( .A1(n16380), .A2(n16379), .ZN(n16383) );
  INHSV2 U19598 ( .I(n16381), .ZN(n16530) );
  XNOR2HSV4 U19599 ( .A1(n16383), .A2(n16382), .ZN(n16384) );
  INHSV3 U19600 ( .I(n19883), .ZN(n16429) );
  INHSV3 U19601 ( .I(n28646), .ZN(n16393) );
  CLKNAND2HSV0 U19602 ( .A1(n21328), .A2(n13958), .ZN(n16387) );
  CLKNAND2HSV1 U19603 ( .A1(n28796), .A2(n13958), .ZN(n16386) );
  CLKNAND2HSV1 U19604 ( .A1(n16387), .A2(n16386), .ZN(n16389) );
  CLKNAND2HSV1 U19605 ( .A1(n16389), .A2(n16388), .ZN(n16390) );
  INHSV2 U19606 ( .I(n16390), .ZN(n16391) );
  NAND2HSV2 U19607 ( .A1(n16391), .A2(n21330), .ZN(n16399) );
  INHSV2 U19608 ( .I(n16392), .ZN(n16460) );
  NAND2HSV0 U19609 ( .A1(n16394), .A2(n13998), .ZN(n16395) );
  INHSV2 U19610 ( .I(n16395), .ZN(n16396) );
  AOI22HSV4 U19611 ( .A1(n18784), .A2(n16460), .B1(n16397), .B2(n16396), .ZN(
        n16398) );
  NAND2HSV0 U19612 ( .A1(\pe8/aot [12]), .A2(n16464), .ZN(n16402) );
  NAND2HSV2 U19613 ( .A1(\pe8/aot [13]), .A2(n16400), .ZN(n16401) );
  XOR2HSV2 U19614 ( .A1(n16402), .A2(n16401), .Z(n16406) );
  NAND2HSV0 U19615 ( .A1(\pe8/aot [14]), .A2(\pe8/bq[14] ), .ZN(n16403) );
  XOR2HSV2 U19616 ( .A1(n16406), .A2(n16405), .Z(n16413) );
  NAND2HSV0 U19617 ( .A1(\pe8/bq[13] ), .A2(\pe8/aot [15]), .ZN(n16408) );
  XOR2HSV0 U19618 ( .A1(n16408), .A2(n16407), .Z(n16411) );
  XOR2HSV2 U19619 ( .A1(n16411), .A2(n16410), .Z(n16412) );
  CLKNAND2HSV0 U19620 ( .A1(n16414), .A2(\pe8/got [13]), .ZN(n16415) );
  NOR2HSV2 U19621 ( .A1(n16416), .A2(n16415), .ZN(n16417) );
  OAI21HSV2 U19622 ( .A1(n22128), .A2(\pe8/ti_7t [5]), .B(n25523), .ZN(n16441)
         );
  CLKNAND2HSV2 U19623 ( .A1(n16421), .A2(n19830), .ZN(n16422) );
  NOR2HSV4 U19624 ( .A1(n25652), .A2(n16422), .ZN(n16427) );
  NOR2HSV4 U19625 ( .A1(n16423), .A2(n16424), .ZN(n16496) );
  INHSV4 U19626 ( .I(n16496), .ZN(n16445) );
  INHSV2 U19627 ( .I(n25651), .ZN(n16426) );
  CLKNAND2HSV4 U19628 ( .A1(n16427), .A2(n16426), .ZN(n19884) );
  INHSV4 U19629 ( .I(n19884), .ZN(n16428) );
  CLKNAND2HSV3 U19630 ( .A1(n16429), .A2(n16428), .ZN(n16500) );
  CLKNAND2HSV2 U19631 ( .A1(n16430), .A2(n22125), .ZN(n16433) );
  NAND2HSV2 U19632 ( .A1(n19986), .A2(\pe8/ti_7t [6]), .ZN(n16446) );
  NAND2HSV0 U19633 ( .A1(n18787), .A2(n28625), .ZN(n16431) );
  CLKAND2HSV1 U19634 ( .A1(n16446), .A2(n16431), .Z(n16432) );
  NAND2HSV2 U19635 ( .A1(n16433), .A2(n16432), .ZN(n16434) );
  INHSV2 U19636 ( .I(n16434), .ZN(n16439) );
  NAND2HSV0 U19637 ( .A1(n16446), .A2(n28695), .ZN(n16435) );
  NOR2HSV2 U19638 ( .A1(n16535), .A2(n16435), .ZN(n16436) );
  INHSV2 U19639 ( .I(n16436), .ZN(n16437) );
  NOR2HSV2 U19640 ( .A1(n16437), .A2(n25649), .ZN(n16438) );
  CLKNHSV0 U19641 ( .I(n16446), .ZN(n16440) );
  NOR2HSV2 U19642 ( .A1(n16441), .A2(n16440), .ZN(n16442) );
  NAND3HSV2 U19643 ( .A1(n16443), .A2(n16442), .A3(n16444), .ZN(n16449) );
  INHSV4 U19644 ( .I(n16445), .ZN(n25582) );
  CLKAND2HSV4 U19645 ( .A1(n25582), .A2(n16446), .Z(n16447) );
  NAND3HSV4 U19646 ( .A1(n16450), .A2(n16449), .A3(n16448), .ZN(n19885) );
  NAND2HSV0 U19647 ( .A1(n16500), .A2(n19885), .ZN(n16451) );
  INHSV2 U19648 ( .I(n16451), .ZN(n16499) );
  CLKNHSV2 U19649 ( .I(n16459), .ZN(n16457) );
  OR2HSV1 U19650 ( .A1(n16452), .A2(n19972), .Z(n16453) );
  OAI211HSV2 U19651 ( .A1(n16455), .A2(n19972), .B(n16454), .C(n16453), .ZN(
        n16458) );
  NOR2HSV4 U19652 ( .A1(n28984), .A2(n16508), .ZN(n16507) );
  INHSV2 U19653 ( .I(n20049), .ZN(n18766) );
  NOR2HSV4 U19654 ( .A1(n16507), .A2(n18766), .ZN(n16497) );
  INHSV2 U19655 ( .I(n16460), .ZN(n16461) );
  NAND2HSV2 U19656 ( .A1(n28799), .A2(n22136), .ZN(n16490) );
  NAND2HSV0 U19657 ( .A1(\pe8/aot [10]), .A2(n16464), .ZN(n16466) );
  NAND2HSV0 U19658 ( .A1(\pe8/bq[11] ), .A2(\pe8/aot [15]), .ZN(n16465) );
  XOR2HSV2 U19659 ( .A1(n16466), .A2(n16465), .Z(n16470) );
  INHSV2 U19660 ( .I(\pe8/phq [7]), .ZN(n16467) );
  XNOR2HSV4 U19661 ( .A1(n16470), .A2(n16469), .ZN(n16474) );
  CLKNAND2HSV2 U19662 ( .A1(n25624), .A2(\pe8/got [10]), .ZN(n16472) );
  INHSV4 U19663 ( .I(n28623), .ZN(n23528) );
  CLKNAND2HSV2 U19664 ( .A1(n23528), .A2(\pe8/pvq [7]), .ZN(n16471) );
  XOR2HSV2 U19665 ( .A1(n16472), .A2(n16471), .Z(n16473) );
  XNOR2HSV4 U19666 ( .A1(n16474), .A2(n16473), .ZN(n16481) );
  CLKNAND2HSV1 U19667 ( .A1(\pe8/aot [14]), .A2(\pe8/bq[12] ), .ZN(n18810) );
  NAND2HSV0 U19668 ( .A1(\pe8/aot [13]), .A2(\pe8/bq[13] ), .ZN(n16475) );
  XOR2HSV0 U19669 ( .A1(n18810), .A2(n16475), .Z(n16479) );
  INHSV1 U19670 ( .I(\pe8/bq[15] ), .ZN(n16569) );
  INHSV2 U19671 ( .I(n16569), .ZN(n18720) );
  NAND2HSV0 U19672 ( .A1(\pe8/aot [11]), .A2(n18720), .ZN(n16477) );
  NAND2HSV0 U19673 ( .A1(\pe8/aot [12]), .A2(\pe8/bq[14] ), .ZN(n16476) );
  XOR2HSV0 U19674 ( .A1(n16477), .A2(n16476), .Z(n16478) );
  XOR2HSV2 U19675 ( .A1(n16479), .A2(n16478), .Z(n16480) );
  XNOR2HSV4 U19676 ( .A1(n16481), .A2(n16480), .ZN(n16483) );
  INHSV2 U19677 ( .I(\pe8/got [11]), .ZN(n19905) );
  NAND2HSV0 U19678 ( .A1(n23653), .A2(n28796), .ZN(n16482) );
  XOR2HSV2 U19679 ( .A1(n16483), .A2(n16482), .Z(n16484) );
  NAND2HSV2 U19680 ( .A1(n28788), .A2(\pe8/got [12]), .ZN(n16485) );
  NAND2HSV2 U19681 ( .A1(n16484), .A2(n16485), .ZN(n16489) );
  INHSV2 U19682 ( .I(n16484), .ZN(n16487) );
  INHSV2 U19683 ( .I(n16485), .ZN(n16486) );
  CLKNAND2HSV2 U19684 ( .A1(n16487), .A2(n16486), .ZN(n16488) );
  NAND2HSV2 U19685 ( .A1(n16490), .A2(n16491), .ZN(n16495) );
  INHSV2 U19686 ( .I(n16490), .ZN(n16493) );
  INHSV2 U19687 ( .I(n16491), .ZN(n16492) );
  CLKNAND2HSV2 U19688 ( .A1(n16493), .A2(n16492), .ZN(n16494) );
  NOR2HSV4 U19689 ( .A1(n16496), .A2(n18760), .ZN(n16582) );
  XNOR2HSV4 U19690 ( .A1(n16583), .A2(n16582), .ZN(n16606) );
  XOR2HSV4 U19691 ( .A1(n16497), .A2(n16606), .Z(n16501) );
  INHSV2 U19692 ( .I(n16501), .ZN(n16498) );
  NAND2HSV4 U19693 ( .A1(n16500), .A2(n19885), .ZN(n19931) );
  NAND2HSV2 U19694 ( .A1(n19931), .A2(n16501), .ZN(n16502) );
  NAND2HSV2 U19695 ( .A1(n18716), .A2(n16311), .ZN(n16505) );
  AOI21HSV4 U19696 ( .A1(n16506), .A2(n16307), .B(n16505), .ZN(n16550) );
  INHSV2 U19697 ( .I(n16550), .ZN(n16548) );
  CLKNAND2HSV2 U19698 ( .A1(n19931), .A2(n28625), .ZN(n16546) );
  INHSV2 U19699 ( .I(n16507), .ZN(n16510) );
  INHSV2 U19700 ( .I(n16508), .ZN(n16556) );
  AOI21HSV1 U19701 ( .A1(n16556), .A2(n18773), .B(n19987), .ZN(n16509) );
  NAND2HSV2 U19702 ( .A1(n16510), .A2(n16509), .ZN(n16544) );
  INHSV2 U19703 ( .I(\pe8/got [9]), .ZN(n19993) );
  INHSV2 U19704 ( .I(n19993), .ZN(n23721) );
  CLKNAND2HSV1 U19705 ( .A1(n23721), .A2(n25624), .ZN(n16513) );
  NAND2HSV0 U19706 ( .A1(\pe8/aot [10]), .A2(n18720), .ZN(n16512) );
  XOR2HSV0 U19707 ( .A1(n16513), .A2(n16512), .Z(n16517) );
  NAND2HSV0 U19708 ( .A1(\pe8/aot [12]), .A2(\pe8/bq[13] ), .ZN(n16515) );
  INHSV2 U19709 ( .I(n28813), .ZN(n25539) );
  NAND2HSV0 U19710 ( .A1(\pe8/aot [9]), .A2(n25539), .ZN(n16514) );
  XOR2HSV0 U19711 ( .A1(n16515), .A2(n16514), .Z(n16516) );
  XOR2HSV0 U19712 ( .A1(n16517), .A2(n16516), .Z(n16529) );
  INHSV2 U19713 ( .I(\pe8/got [10]), .ZN(n19841) );
  NOR2HSV3 U19714 ( .A1(n16385), .A2(n19841), .ZN(n16528) );
  NAND2HSV0 U19715 ( .A1(\pe8/aot [14]), .A2(\pe8/bq[11] ), .ZN(n16520) );
  CLKNHSV0 U19716 ( .I(\pe8/aot [16]), .ZN(n16518) );
  NAND2HSV0 U19717 ( .A1(n28627), .A2(\pe8/bq[9] ), .ZN(n16519) );
  XOR2HSV0 U19718 ( .A1(n16520), .A2(n16519), .Z(n16524) );
  NAND2HSV0 U19719 ( .A1(\pe8/bq[12] ), .A2(\pe8/aot [13]), .ZN(n16522) );
  NAND2HSV0 U19720 ( .A1(\pe8/bq[10] ), .A2(\pe8/aot [15]), .ZN(n16521) );
  XOR2HSV0 U19721 ( .A1(n16522), .A2(n16521), .Z(n16523) );
  XOR2HSV0 U19722 ( .A1(n16524), .A2(n16523), .Z(n16526) );
  XNOR2HSV4 U19723 ( .A1(n16526), .A2(n16525), .ZN(n16527) );
  XOR3HSV2 U19724 ( .A1(n16529), .A2(n16528), .A3(n16527), .Z(n16532) );
  INHSV2 U19725 ( .I(n16530), .ZN(n20009) );
  CLKNAND2HSV1 U19726 ( .A1(n20009), .A2(n28618), .ZN(n16531) );
  CLKXOR2HSV2 U19727 ( .A1(n16532), .A2(n16531), .Z(n16534) );
  CLKNAND2HSV1 U19728 ( .A1(n28799), .A2(\pe8/got [12]), .ZN(n16533) );
  CLKXOR2HSV2 U19729 ( .A1(n16534), .A2(n16533), .Z(n16538) );
  CLKNHSV1 U19730 ( .I(\pe8/got [13]), .ZN(n16536) );
  NOR2HSV4 U19731 ( .A1(n18823), .A2(n16536), .ZN(n16539) );
  INHSV2 U19732 ( .I(n16539), .ZN(n16537) );
  NAND2HSV2 U19733 ( .A1(n16538), .A2(n16537), .ZN(n16542) );
  INHSV2 U19734 ( .I(n16538), .ZN(n16540) );
  CLKNAND2HSV1 U19735 ( .A1(n16540), .A2(n16539), .ZN(n16541) );
  NAND2HSV2 U19736 ( .A1(n16542), .A2(n16541), .ZN(n16543) );
  XNOR2HSV4 U19737 ( .A1(n16544), .A2(n16543), .ZN(n16545) );
  XNOR2HSV4 U19738 ( .A1(n16546), .A2(n16545), .ZN(n16549) );
  INHSV3 U19739 ( .I(n16549), .ZN(n16547) );
  CLKNAND2HSV3 U19740 ( .A1(n16548), .A2(n16547), .ZN(n16553) );
  NAND2HSV2 U19741 ( .A1(n16550), .A2(n16549), .ZN(n16551) );
  INHSV2 U19742 ( .I(n18706), .ZN(n28815) );
  CLKNAND2HSV2 U19743 ( .A1(n16551), .A2(n22137), .ZN(n16552) );
  BUFHSV2 U19744 ( .I(n16554), .Z(n22128) );
  NAND2HSV2 U19745 ( .A1(n18655), .A2(n19835), .ZN(n16555) );
  INHSV2 U19746 ( .I(\pe8/got [13]), .ZN(n18691) );
  NAND2HSV0 U19747 ( .A1(n28796), .A2(n23721), .ZN(n16573) );
  NAND2HSV2 U19748 ( .A1(n20009), .A2(\pe8/got [10]), .ZN(n16572) );
  NAND2HSV0 U19749 ( .A1(\pe8/aot [10]), .A2(\pe8/bq[14] ), .ZN(n16559) );
  NAND2HSV0 U19750 ( .A1(\pe8/aot [14]), .A2(\pe8/bq[10] ), .ZN(n16558) );
  XOR2HSV0 U19751 ( .A1(n16559), .A2(n16558), .Z(n16563) );
  NAND2HSV0 U19752 ( .A1(\pe8/aot [13]), .A2(\pe8/bq[11] ), .ZN(n16561) );
  INHSV2 U19753 ( .I(\pe8/got [8]), .ZN(n28655) );
  INHSV2 U19754 ( .I(n28655), .ZN(n23605) );
  NAND2HSV0 U19755 ( .A1(n23605), .A2(n25624), .ZN(n16560) );
  XOR2HSV0 U19756 ( .A1(n16561), .A2(n16560), .Z(n16562) );
  NAND2HSV0 U19757 ( .A1(\pe8/aot [11]), .A2(\pe8/bq[13] ), .ZN(n16565) );
  NAND2HSV0 U19758 ( .A1(n28627), .A2(\pe8/bq[8] ), .ZN(n16564) );
  XOR2HSV0 U19759 ( .A1(n16565), .A2(n16564), .Z(n16568) );
  NAND2HSV2 U19760 ( .A1(n23528), .A2(\pe8/pvq [9]), .ZN(n16566) );
  XOR2HSV0 U19761 ( .A1(n16566), .A2(\pe8/phq [9]), .Z(n16567) );
  NAND2HSV0 U19762 ( .A1(\pe8/aot [9]), .A2(n25532), .ZN(n16570) );
  XOR3HSV2 U19763 ( .A1(n16573), .A2(n16572), .A3(n16571), .Z(n16575) );
  INHSV2 U19764 ( .I(n28799), .ZN(n18820) );
  INHSV2 U19765 ( .I(n18820), .ZN(n18746) );
  CLKNAND2HSV1 U19766 ( .A1(n18746), .A2(n23653), .ZN(n16574) );
  XOR2HSV0 U19767 ( .A1(n16575), .A2(n16574), .Z(n16577) );
  INAND2HSV2 U19768 ( .A1(n18823), .B1(\pe8/got [12]), .ZN(n16576) );
  XOR2HSV2 U19769 ( .A1(n16577), .A2(n16576), .Z(n16578) );
  XNOR2HSV4 U19770 ( .A1(n16579), .A2(n16578), .ZN(n16581) );
  INHSV2 U19771 ( .I(\pe8/got [14]), .ZN(n19820) );
  NAND2HSV2 U19772 ( .A1(n19931), .A2(n19940), .ZN(n16580) );
  XNOR2HSV4 U19773 ( .A1(n16581), .A2(n16580), .ZN(n16602) );
  INHSV2 U19774 ( .I(n16602), .ZN(n16600) );
  XNOR2HSV4 U19775 ( .A1(n16583), .A2(n16582), .ZN(n16587) );
  OAI21HSV1 U19776 ( .A1(n16587), .A2(n25523), .B(n22125), .ZN(n16584) );
  NOR2HSV1 U19777 ( .A1(n16607), .A2(n16584), .ZN(n16585) );
  OAI21HSV0 U19778 ( .A1(n19931), .A2(n16606), .B(n16585), .ZN(n16586) );
  CLKNHSV0 U19779 ( .I(n16586), .ZN(n16598) );
  INHSV2 U19780 ( .I(n16587), .ZN(n16590) );
  CLKAND2HSV1 U19781 ( .A1(n16590), .A2(n25523), .Z(n16588) );
  CLKNAND2HSV0 U19782 ( .A1(n16588), .A2(n18690), .ZN(n16589) );
  OAI21HSV2 U19783 ( .A1(n19931), .A2(n16590), .B(n16589), .ZN(n16595) );
  NOR2HSV1 U19784 ( .A1(n16590), .A2(n25523), .ZN(n16591) );
  NOR2HSV1 U19785 ( .A1(n16591), .A2(n18657), .ZN(n16592) );
  CLKNAND2HSV1 U19786 ( .A1(n16592), .A2(n16607), .ZN(n16594) );
  AND2HSV2 U19787 ( .A1(n18716), .A2(n13998), .Z(n16593) );
  OAI21HSV2 U19788 ( .A1(n16595), .A2(n16594), .B(n16593), .ZN(n16596) );
  CLKNAND2HSV4 U19789 ( .A1(n16604), .A2(n16603), .ZN(n18709) );
  XNOR2HSV4 U19790 ( .A1(n16605), .A2(n18709), .ZN(n29006) );
  CLKNHSV2 U19791 ( .I(n27074), .ZN(n28867) );
  XNOR2HSV4 U19792 ( .A1(n16610), .A2(n16609), .ZN(n16624) );
  XNOR2HSV4 U19793 ( .A1(n16624), .A2(n16623), .ZN(n28704) );
  CLKBUFHSV4 U19794 ( .I(n16638), .Z(n16749) );
  INHSV2 U19795 ( .I(\pe10/got [16]), .ZN(n16948) );
  INHSV2 U19796 ( .I(n16948), .ZN(n17112) );
  INHSV2 U19797 ( .I(n16739), .ZN(n28810) );
  NAND2HSV2 U19798 ( .A1(n16749), .A2(n28810), .ZN(n16886) );
  INHSV4 U19799 ( .I(n16886), .ZN(n25255) );
  INHSV2 U19800 ( .I(n25255), .ZN(n20145) );
  CLKNAND2HSV3 U19801 ( .A1(\pe10/ti_1 ), .A2(\pe10/got [15]), .ZN(n16612) );
  INHSV4 U19802 ( .I(n16774), .ZN(n16658) );
  NAND2HSV2 U19803 ( .A1(n16658), .A2(\pe10/bq[15] ), .ZN(n16611) );
  XOR3HSV2 U19804 ( .A1(\pe10/phq [2]), .A2(n16612), .A3(n16611), .Z(n16616)
         );
  NAND2HSV2 U19805 ( .A1(\pe10/pvq [2]), .A2(n14001), .ZN(n16615) );
  INHSV4 U19806 ( .I(\pe10/bq[16] ), .ZN(n16809) );
  OAI21HSV2 U19807 ( .A1(n16615), .A2(n16614), .B(n16613), .ZN(n16617) );
  INHSV2 U19808 ( .I(n16616), .ZN(n16619) );
  INHSV2 U19809 ( .I(n16617), .ZN(n16618) );
  INHSV2 U19810 ( .I(\pe10/got [16]), .ZN(n16739) );
  NOR2HSV1 U19811 ( .A1(n16666), .A2(n16739), .ZN(n16621) );
  AOI21HSV2 U19812 ( .A1(n16622), .A2(n23484), .B(n16621), .ZN(n16627) );
  XNOR2HSV4 U19813 ( .A1(n16624), .A2(n16623), .ZN(n16670) );
  NOR2HSV4 U19814 ( .A1(n23484), .A2(n16625), .ZN(n16668) );
  INHSV2 U19815 ( .I(n16668), .ZN(n16626) );
  CLKNAND2HSV3 U19816 ( .A1(n16627), .A2(n16626), .ZN(n16646) );
  INHSV4 U19817 ( .I(n16646), .ZN(n22104) );
  INHSV2 U19818 ( .I(n16638), .ZN(n20149) );
  CLKNAND2HSV1 U19819 ( .A1(\pe10/ti_7t [1]), .A2(n20149), .ZN(n16641) );
  INHSV2 U19820 ( .I(n16641), .ZN(n16663) );
  BUFHSV4 U19821 ( .I(n16638), .Z(n16995) );
  INHSV2 U19822 ( .I(n16995), .ZN(n16956) );
  INHSV2 U19823 ( .I(\pe10/got [15]), .ZN(n25256) );
  NAND2HSV2 U19824 ( .A1(n16658), .A2(\pe10/bq[14] ), .ZN(n26165) );
  NAND2HSV0 U19825 ( .A1(\pe10/aot [15]), .A2(\pe10/bq[15] ), .ZN(n16628) );
  CLKNAND2HSV1 U19826 ( .A1(n16628), .A2(\pe10/phq [3]), .ZN(n16631) );
  INHSV2 U19827 ( .I(\pe10/phq [3]), .ZN(n16629) );
  NAND3HSV2 U19828 ( .A1(n16629), .A2(\pe10/aot [15]), .A3(\pe10/bq[15] ), 
        .ZN(n16630) );
  CLKNAND2HSV2 U19829 ( .A1(n16631), .A2(n16630), .ZN(n16637) );
  CLKNAND2HSV2 U19830 ( .A1(\pe10/ti_1 ), .A2(\pe10/got [14]), .ZN(n16632) );
  NOR2HSV4 U19831 ( .A1(n16635), .A2(n16634), .ZN(n16633) );
  CLKBUFHSV4 U19832 ( .I(n16638), .Z(n16740) );
  INHSV1 U19833 ( .I(n16740), .ZN(n25259) );
  NOR2HSV1 U19834 ( .A1(n16795), .A2(n25259), .ZN(n20128) );
  AOI22HSV2 U19835 ( .A1(n16670), .A2(n20128), .B1(n16643), .B2(n22418), .ZN(
        n16639) );
  AOI21HSV2 U19836 ( .A1(n22508), .A2(n16816), .B(n22102), .ZN(n16645) );
  CLKBUFHSV4 U19837 ( .I(n16998), .Z(n17117) );
  OAI21HSV2 U19838 ( .A1(n16643), .A2(n16642), .B(n17117), .ZN(n16644) );
  NOR2HSV2 U19839 ( .A1(n16645), .A2(n16644), .ZN(n16647) );
  INHSV2 U19840 ( .I(n16638), .ZN(n16708) );
  NAND2HSV2 U19841 ( .A1(n16708), .A2(\pe10/ti_7t [3]), .ZN(n16679) );
  BUFHSV4 U19842 ( .I(\pe10/ti_1 ), .Z(n16761) );
  XNOR2HSV4 U19843 ( .A1(n16650), .A2(n16649), .ZN(n16653) );
  NAND2HSV0 U19844 ( .A1(\pe10/bq[14] ), .A2(\pe10/aot [15]), .ZN(n16651) );
  NAND2HSV2 U19845 ( .A1(n16653), .A2(n16654), .ZN(n16657) );
  INHSV3 U19846 ( .I(n16653), .ZN(n16656) );
  NAND2HSV2 U19847 ( .A1(n16658), .A2(\pe10/bq[13] ), .ZN(n16659) );
  XNOR2HSV4 U19848 ( .A1(n16659), .A2(\pe10/phq [4]), .ZN(n16660) );
  CLKBUFHSV4 U19849 ( .I(\pe10/bq[15] ), .Z(n16897) );
  XNOR2HSV4 U19850 ( .A1(n16662), .A2(n16661), .ZN(n16665) );
  INHSV2 U19851 ( .I(\pe10/got [14]), .ZN(n26156) );
  NOR2HSV2 U19852 ( .A1(n26156), .A2(n25259), .ZN(n16755) );
  XNOR2HSV4 U19853 ( .A1(n16665), .A2(n16664), .ZN(n16675) );
  INHSV3 U19854 ( .I(n16675), .ZN(n16674) );
  INHSV2 U19855 ( .I(n16666), .ZN(n16667) );
  NOR2HSV2 U19856 ( .A1(n16670), .A2(n16669), .ZN(n16672) );
  INHSV2 U19857 ( .I(n16948), .ZN(n16892) );
  AND2HSV2 U19858 ( .A1(n16749), .A2(n16739), .Z(n16671) );
  CLKNAND2HSV3 U19859 ( .A1(n16674), .A2(n16673), .ZN(n16677) );
  NAND2HSV4 U19860 ( .A1(n16677), .A2(n16676), .ZN(n16753) );
  INHSV2 U19861 ( .I(n16749), .ZN(n17119) );
  NAND2HSV2 U19862 ( .A1(n16735), .A2(n16892), .ZN(n23475) );
  INHSV2 U19863 ( .I(n23475), .ZN(n16678) );
  CLKNAND2HSV2 U19864 ( .A1(n14002), .A2(\pe10/pvq [5]), .ZN(n16684) );
  XNOR2HSV4 U19865 ( .A1(n16684), .A2(n16683), .ZN(n16685) );
  XNOR2HSV4 U19866 ( .A1(n16686), .A2(n16685), .ZN(n16692) );
  XNOR2HSV4 U19867 ( .A1(n16689), .A2(\pe10/phq [5]), .ZN(n16690) );
  XNOR2HSV4 U19868 ( .A1(n16692), .A2(n16691), .ZN(n16697) );
  CLKNHSV0 U19869 ( .I(\pe10/ti_7t [1]), .ZN(n16693) );
  AOI21HSV2 U19870 ( .A1(n16693), .A2(n25259), .B(n16729), .ZN(n16694) );
  OAI21HSV0 U19871 ( .A1(n28704), .A2(n16956), .B(n16694), .ZN(n16695) );
  INHSV2 U19872 ( .I(n16695), .ZN(n16696) );
  XNOR2HSV4 U19873 ( .A1(n16697), .A2(n16696), .ZN(n16699) );
  CLKNAND2HSV2 U19874 ( .A1(n16781), .A2(n14070), .ZN(n16700) );
  NAND2HSV2 U19875 ( .A1(n16699), .A2(n16698), .ZN(n16703) );
  INHSV2 U19876 ( .I(n16699), .ZN(n16701) );
  INHSV3 U19877 ( .I(n16704), .ZN(n16707) );
  INHSV3 U19878 ( .I(n16705), .ZN(n16706) );
  NOR2HSV2 U19879 ( .A1(n23475), .A2(n20148), .ZN(n16709) );
  NAND2HSV2 U19880 ( .A1(n17119), .A2(\pe10/ti_7t [5]), .ZN(n16796) );
  CLKNAND2HSV3 U19881 ( .A1(n16797), .A2(n16796), .ZN(n16711) );
  INHSV2 U19882 ( .I(n16761), .ZN(n26185) );
  NOR2HSV2 U19883 ( .A1(n22636), .A2(n26185), .ZN(n16714) );
  NAND2HSV0 U19884 ( .A1(n28424), .A2(\pe10/bq[11] ), .ZN(n16713) );
  XOR2HSV0 U19885 ( .A1(n16714), .A2(n16713), .Z(n16718) );
  NAND2HSV0 U19886 ( .A1(\pe10/bq[13] ), .A2(\pe10/aot [14]), .ZN(n16716) );
  INHSV2 U19887 ( .I(\pe10/aot [11]), .ZN(n24463) );
  CLKNAND2HSV1 U19888 ( .A1(\pe10/aot [11]), .A2(n17084), .ZN(n16715) );
  XOR2HSV0 U19889 ( .A1(n16716), .A2(n16715), .Z(n16717) );
  XNOR2HSV4 U19890 ( .A1(n16899), .A2(\pe10/phq [6]), .ZN(n16720) );
  BUFHSV8 U19891 ( .I(n14002), .Z(n23536) );
  NAND2HSV2 U19892 ( .A1(n23536), .A2(\pe10/pvq [6]), .ZN(n16719) );
  XNOR2HSV4 U19893 ( .A1(n16720), .A2(n16719), .ZN(n16724) );
  NAND2HSV0 U19894 ( .A1(\pe10/aot [13]), .A2(\pe10/bq[14] ), .ZN(n16722) );
  NAND2HSV0 U19895 ( .A1(\pe10/aot [12]), .A2(\pe10/bq[15] ), .ZN(n16721) );
  XOR2HSV0 U19896 ( .A1(n16722), .A2(n16721), .Z(n16723) );
  XNOR2HSV4 U19897 ( .A1(n16724), .A2(n16723), .ZN(n16725) );
  XNOR2HSV4 U19898 ( .A1(n16726), .A2(n16725), .ZN(n16728) );
  NAND2HSV2 U19899 ( .A1(n16816), .A2(n16876), .ZN(n16727) );
  XNOR2HSV4 U19900 ( .A1(n16728), .A2(n16727), .ZN(n16731) );
  NAND2HSV2 U19901 ( .A1(n16850), .A2(n28479), .ZN(n16730) );
  XNOR2HSV4 U19902 ( .A1(n16731), .A2(n16730), .ZN(n16733) );
  NAND2HSV2 U19903 ( .A1(n16848), .A2(n14070), .ZN(n16732) );
  XNOR2HSV4 U19904 ( .A1(n16733), .A2(n16732), .ZN(n16743) );
  INHSV3 U19905 ( .I(n16753), .ZN(n23473) );
  CLKNAND2HSV1 U19906 ( .A1(n16757), .A2(n25255), .ZN(n16738) );
  CLKNHSV0 U19907 ( .I(n16735), .ZN(n16736) );
  NOR2HSV0 U19908 ( .A1(n16736), .A2(n16795), .ZN(n16737) );
  INHSV2 U19909 ( .I(n16739), .ZN(n26220) );
  INHSV2 U19910 ( .I(n16803), .ZN(n16745) );
  INHSV2 U19911 ( .I(\pe10/ti_7t [6]), .ZN(n16750) );
  INHSV2 U19912 ( .I(n16749), .ZN(n16843) );
  NAND2HSV2 U19913 ( .A1(n16750), .A2(n16843), .ZN(n16804) );
  NAND2HSV2 U19914 ( .A1(n16804), .A2(n17120), .ZN(n16751) );
  AOI21HSV4 U19915 ( .A1(n16752), .A2(n20142), .B(n16751), .ZN(n16802) );
  NAND2HSV2 U19916 ( .A1(\pe10/ti_7t [4]), .A2(n16843), .ZN(n16846) );
  INHSV2 U19917 ( .I(n16846), .ZN(n16808) );
  CLKNHSV2 U19918 ( .I(n16757), .ZN(n16758) );
  NOR2HSV4 U19919 ( .A1(n16758), .A2(n17065), .ZN(n16785) );
  CLKNHSV0 U19920 ( .I(n22636), .ZN(n16759) );
  INHSV2 U19921 ( .I(\pe10/got [10]), .ZN(n16760) );
  INHSV4 U19922 ( .I(n16760), .ZN(n28644) );
  NAND2HSV0 U19923 ( .A1(n28644), .A2(n16761), .ZN(n16763) );
  NAND2HSV0 U19924 ( .A1(\pe10/aot [15]), .A2(\pe10/bq[11] ), .ZN(n16762) );
  XOR2HSV0 U19925 ( .A1(n16763), .A2(n16762), .Z(n16767) );
  NAND2HSV0 U19926 ( .A1(\pe10/aot [12]), .A2(\pe10/bq[14] ), .ZN(n16765) );
  NAND2HSV0 U19927 ( .A1(\pe10/aot [10]), .A2(n17084), .ZN(n16764) );
  XNOR2HSV4 U19928 ( .A1(n16769), .A2(n16768), .ZN(n16780) );
  NAND2HSV2 U19929 ( .A1(n23536), .A2(\pe10/pvq [7]), .ZN(n16770) );
  CLKXOR2HSV2 U19930 ( .A1(n16770), .A2(\pe10/phq [7]), .Z(n16773) );
  CLKNHSV0 U19931 ( .I(\pe10/bq[12] ), .ZN(n23535) );
  NOR2HSV2 U19932 ( .A1(n24463), .A2(n23535), .ZN(n16901) );
  AOI22HSV0 U19933 ( .A1(\pe10/bq[12] ), .A2(\pe10/aot [14]), .B1(n16897), 
        .B2(\pe10/aot [11]), .ZN(n16771) );
  XNOR2HSV4 U19934 ( .A1(n16773), .A2(n16772), .ZN(n16778) );
  NAND2HSV0 U19935 ( .A1(\pe10/aot [13]), .A2(\pe10/bq[13] ), .ZN(n16776) );
  INHSV2 U19936 ( .I(n16774), .ZN(n20083) );
  NAND2HSV0 U19937 ( .A1(n20083), .A2(\pe10/bq[10] ), .ZN(n16775) );
  XOR2HSV0 U19938 ( .A1(n16776), .A2(n16775), .Z(n16777) );
  XNOR2HSV4 U19939 ( .A1(n16778), .A2(n16777), .ZN(n16779) );
  XNOR2HSV4 U19940 ( .A1(n16780), .A2(n16779), .ZN(n16783) );
  CLKNHSV2 U19941 ( .I(n16781), .ZN(n17023) );
  CLKNAND2HSV2 U19942 ( .A1(n16785), .A2(n16784), .ZN(n16787) );
  MUX2NHSV2 U19943 ( .I0(n16789), .I1(n16788), .S(n16790), .ZN(n16794) );
  NOR2HSV1 U19944 ( .A1(n16846), .A2(n26156), .ZN(n16792) );
  OAI21HSV0 U19945 ( .A1(n16808), .A2(n17117), .B(n14070), .ZN(n16791) );
  MUX2NHSV2 U19946 ( .I0(n16792), .I1(n16791), .S(n16790), .ZN(n16793) );
  XNOR2HSV4 U19947 ( .A1(n16800), .A2(n16799), .ZN(n16801) );
  XNOR2HSV4 U19948 ( .A1(n16802), .A2(n16801), .ZN(n23462) );
  CLKNAND2HSV3 U19949 ( .A1(n23462), .A2(n16844), .ZN(n16896) );
  CLKAND2HSV2 U19950 ( .A1(n16669), .A2(\pe10/ti_7t [7]), .Z(n16887) );
  INHSV2 U19951 ( .I(n16887), .ZN(n16845) );
  CLKNHSV1 U19952 ( .I(n16804), .ZN(n16805) );
  CLKNHSV0 U19953 ( .I(\pe10/got [15]), .ZN(n25261) );
  INHSV2 U19954 ( .I(n16995), .ZN(n22442) );
  INHSV2 U19955 ( .I(\pe10/got [13]), .ZN(n17065) );
  AOI21HSV2 U19956 ( .A1(n16846), .A2(n22442), .B(n17065), .ZN(n16807) );
  NAND2HSV0 U19957 ( .A1(\pe10/aot [12]), .A2(\pe10/bq[13] ), .ZN(n16811) );
  NAND2HSV0 U19958 ( .A1(\pe10/aot [9]), .A2(n17084), .ZN(n16810) );
  XOR2HSV0 U19959 ( .A1(n16811), .A2(n16810), .Z(n16815) );
  BUFHSV2 U19960 ( .I(\pe10/ti_1 ), .Z(n22458) );
  NAND2HSV0 U19961 ( .A1(n22458), .A2(\pe10/got [9]), .ZN(n16813) );
  NAND2HSV0 U19962 ( .A1(\pe10/aot [10]), .A2(n16897), .ZN(n16812) );
  XOR2HSV0 U19963 ( .A1(n16813), .A2(n16812), .Z(n16814) );
  XOR2HSV0 U19964 ( .A1(n16815), .A2(n16814), .Z(n16830) );
  NAND2HSV2 U19965 ( .A1(n16816), .A2(n28644), .ZN(n16829) );
  CLKNHSV0 U19966 ( .I(\pe10/aot [15]), .ZN(n17038) );
  INHSV2 U19967 ( .I(\pe10/bq[10] ), .ZN(n22722) );
  CLKNAND2HSV1 U19968 ( .A1(n16973), .A2(\pe10/bq[10] ), .ZN(n16818) );
  NAND2HSV0 U19969 ( .A1(\pe10/aot [13]), .A2(\pe10/bq[12] ), .ZN(n16817) );
  XOR2HSV0 U19970 ( .A1(n16818), .A2(n16817), .Z(n16822) );
  INHSV2 U19971 ( .I(\pe10/bq[9] ), .ZN(n20081) );
  INHSV2 U19972 ( .I(n20081), .ZN(n23515) );
  CLKNAND2HSV1 U19973 ( .A1(n20083), .A2(n23515), .ZN(n16820) );
  NAND2HSV0 U19974 ( .A1(\pe10/aot [11]), .A2(\pe10/bq[14] ), .ZN(n16819) );
  XOR2HSV0 U19975 ( .A1(n16820), .A2(n16819), .Z(n16821) );
  XOR2HSV0 U19976 ( .A1(n16822), .A2(n16821), .Z(n16827) );
  BUFHSV8 U19977 ( .I(n14002), .Z(n28811) );
  NAND2HSV2 U19978 ( .A1(n14002), .A2(\pe10/pvq [8]), .ZN(n16823) );
  XNOR2HSV1 U19979 ( .A1(n16823), .A2(\pe10/phq [8]), .ZN(n16825) );
  NAND2HSV0 U19980 ( .A1(\pe10/bq[11] ), .A2(\pe10/aot [14]), .ZN(n16824) );
  XNOR2HSV1 U19981 ( .A1(n16825), .A2(n16824), .ZN(n16826) );
  NAND2HSV0 U19982 ( .A1(n28630), .A2(n16759), .ZN(n16831) );
  XNOR2HSV1 U19983 ( .A1(n16832), .A2(n16831), .ZN(n16834) );
  XNOR2HSV4 U19984 ( .A1(n16834), .A2(n16833), .ZN(n16835) );
  XOR2HSV4 U19985 ( .A1(n16836), .A2(n16835), .Z(n16839) );
  XNOR2HSV4 U19986 ( .A1(n16841), .A2(n16840), .ZN(n16891) );
  CLKAND2HSV2 U19987 ( .A1(n17002), .A2(n28810), .Z(n16884) );
  CLKNAND2HSV4 U19988 ( .A1(n23462), .A2(n16844), .ZN(n16888) );
  INHSV2 U19989 ( .I(\pe10/got [14]), .ZN(n20065) );
  NAND2HSV4 U19990 ( .A1(n16847), .A2(n16846), .ZN(n28794) );
  INHSV2 U19991 ( .I(n28679), .ZN(n16849) );
  INHSV4 U19992 ( .I(n16849), .ZN(n23474) );
  NAND2HSV0 U19993 ( .A1(n23474), .A2(n16759), .ZN(n16875) );
  INHSV2 U19994 ( .I(n16907), .ZN(n26189) );
  NAND2HSV0 U19995 ( .A1(n26189), .A2(\pe10/got [9]), .ZN(n16873) );
  NAND2HSV2 U19996 ( .A1(n16850), .A2(n28644), .ZN(n16872) );
  NAND2HSV0 U19997 ( .A1(\pe10/aot [13]), .A2(\pe10/bq[11] ), .ZN(n16852) );
  XOR2HSV0 U19998 ( .A1(n16852), .A2(n16851), .Z(n16856) );
  BUFHSV4 U19999 ( .I(\pe10/got [8]), .Z(n28642) );
  CLKNAND2HSV1 U20000 ( .A1(n22458), .A2(n28642), .ZN(n16854) );
  NAND2HSV0 U20001 ( .A1(\pe10/aot [10]), .A2(\pe10/bq[14] ), .ZN(n16853) );
  XOR2HSV0 U20002 ( .A1(n16854), .A2(n16853), .Z(n16855) );
  XOR2HSV0 U20003 ( .A1(n16856), .A2(n16855), .Z(n16863) );
  NAND2HSV0 U20004 ( .A1(\pe10/aot [12]), .A2(\pe10/bq[12] ), .ZN(n16858) );
  NAND2HSV0 U20005 ( .A1(n16973), .A2(\pe10/bq[9] ), .ZN(n16857) );
  XOR2HSV0 U20006 ( .A1(n16858), .A2(n16857), .Z(n16861) );
  NAND2HSV2 U20007 ( .A1(n28811), .A2(\pe10/pvq [9]), .ZN(n16859) );
  XOR2HSV0 U20008 ( .A1(n16859), .A2(\pe10/phq [9]), .Z(n16860) );
  XOR2HSV0 U20009 ( .A1(n16861), .A2(n16860), .Z(n16862) );
  XOR2HSV0 U20010 ( .A1(n16863), .A2(n16862), .Z(n16870) );
  NAND2HSV0 U20011 ( .A1(\pe10/aot [9]), .A2(\pe10/bq[15] ), .ZN(n16865) );
  NAND2HSV0 U20012 ( .A1(\pe10/aot [11]), .A2(\pe10/bq[13] ), .ZN(n16864) );
  XOR2HSV0 U20013 ( .A1(n16865), .A2(n16864), .Z(n16868) );
  CLKNAND2HSV1 U20014 ( .A1(n20083), .A2(\pe10/bq[8] ), .ZN(n22444) );
  NAND2HSV0 U20015 ( .A1(\pe10/bq[10] ), .A2(\pe10/aot [14]), .ZN(n16866) );
  XOR2HSV0 U20016 ( .A1(n22444), .A2(n16866), .Z(n16867) );
  XOR2HSV0 U20017 ( .A1(n16868), .A2(n16867), .Z(n16869) );
  XNOR2HSV1 U20018 ( .A1(n16870), .A2(n16869), .ZN(n16871) );
  XOR3HSV2 U20019 ( .A1(n16873), .A2(n16872), .A3(n16871), .Z(n16874) );
  NAND2HSV0 U20020 ( .A1(n28794), .A2(n16876), .ZN(n16878) );
  CLKNHSV2 U20021 ( .I(n16880), .ZN(n28582) );
  CLKNAND2HSV1 U20022 ( .A1(n28479), .A2(n28582), .ZN(n16881) );
  INHSV2 U20023 ( .I(n16999), .ZN(n28694) );
  NOR2HSV2 U20024 ( .A1(n16891), .A2(n16886), .ZN(n16890) );
  INHSV2 U20025 ( .I(n16887), .ZN(n16895) );
  CLKNAND2HSV1 U20026 ( .A1(n17002), .A2(n22508), .ZN(n16889) );
  INHSV2 U20027 ( .I(n16891), .ZN(n16954) );
  NOR2HSV2 U20028 ( .A1(n16954), .A2(n16708), .ZN(n16894) );
  INHSV4 U20029 ( .I(n16942), .ZN(n25676) );
  CLKNAND2HSV2 U20030 ( .A1(n28694), .A2(n25676), .ZN(n16939) );
  NAND2HSV4 U20031 ( .A1(n16896), .A2(n16895), .ZN(n26094) );
  NAND2HSV0 U20032 ( .A1(n26094), .A2(n14070), .ZN(n16935) );
  OR2HSV1 U20033 ( .A1(n16998), .A2(n16750), .Z(n17019) );
  NAND2HSV2 U20034 ( .A1(n17020), .A2(n17019), .ZN(n16960) );
  NAND2HSV2 U20035 ( .A1(n16960), .A2(n28479), .ZN(n16933) );
  NAND2HSV0 U20036 ( .A1(n28794), .A2(n16759), .ZN(n16929) );
  NAND2HSV0 U20037 ( .A1(\pe10/aot [8]), .A2(n16897), .ZN(n16906) );
  CLKNHSV0 U20038 ( .I(n16973), .ZN(n16898) );
  INHSV2 U20039 ( .I(\pe10/bq[8] ), .ZN(n26101) );
  NOR2HSV1 U20040 ( .A1(n16898), .A2(n26101), .ZN(n16900) );
  CLKNAND2HSV0 U20041 ( .A1(\pe10/aot [11]), .A2(\pe10/bq[8] ), .ZN(n20077) );
  OAI22HSV2 U20042 ( .A1(n16901), .A2(n16900), .B1(n16899), .B2(n20077), .ZN(
        n16905) );
  NAND2HSV0 U20043 ( .A1(\pe10/bq[9] ), .A2(\pe10/aot [14]), .ZN(n16903) );
  NAND2HSV0 U20044 ( .A1(\pe10/aot [12]), .A2(\pe10/bq[11] ), .ZN(n16902) );
  XOR2HSV0 U20045 ( .A1(n16903), .A2(n16902), .Z(n16904) );
  XOR3HSV2 U20046 ( .A1(n16906), .A2(n16905), .A3(n16904), .Z(n16923) );
  INHSV2 U20047 ( .I(n16907), .ZN(n28666) );
  CLKNAND2HSV1 U20048 ( .A1(n28666), .A2(n28642), .ZN(n16922) );
  NAND2HSV0 U20049 ( .A1(\pe10/aot [9]), .A2(\pe10/bq[14] ), .ZN(n16908) );
  XOR2HSV0 U20050 ( .A1(n16909), .A2(n16908), .Z(n16913) );
  NAND2HSV0 U20051 ( .A1(\pe10/aot [10]), .A2(\pe10/bq[13] ), .ZN(n16911) );
  NAND2HSV0 U20052 ( .A1(\pe10/bq[7] ), .A2(n20083), .ZN(n16910) );
  XOR2HSV0 U20053 ( .A1(n16911), .A2(n16910), .Z(n16912) );
  XOR2HSV0 U20054 ( .A1(n16913), .A2(n16912), .Z(n16920) );
  NAND2HSV0 U20055 ( .A1(\pe10/aot [13]), .A2(\pe10/bq[10] ), .ZN(n16915) );
  NAND2HSV0 U20056 ( .A1(n22458), .A2(\pe10/got [7]), .ZN(n16914) );
  XOR2HSV0 U20057 ( .A1(n16915), .A2(n16914), .Z(n16918) );
  NAND2HSV2 U20058 ( .A1(n23513), .A2(\pe10/pvq [10]), .ZN(n16916) );
  XOR2HSV0 U20059 ( .A1(n16916), .A2(\pe10/phq [10]), .Z(n16917) );
  XOR2HSV0 U20060 ( .A1(n16918), .A2(n16917), .Z(n16919) );
  XOR2HSV0 U20061 ( .A1(n16920), .A2(n16919), .Z(n16921) );
  XOR3HSV2 U20062 ( .A1(n16923), .A2(n16922), .A3(n16921), .Z(n16925) );
  CLKNAND2HSV0 U20063 ( .A1(n28630), .A2(\pe10/got [9]), .ZN(n16924) );
  XNOR2HSV1 U20064 ( .A1(n16925), .A2(n16924), .ZN(n16927) );
  NAND2HSV0 U20065 ( .A1(n28679), .A2(n28644), .ZN(n16926) );
  XNOR2HSV1 U20066 ( .A1(n16927), .A2(n16926), .ZN(n16928) );
  CLKBUFHSV4 U20067 ( .I(n28582), .Z(n26131) );
  NAND2HSV0 U20068 ( .A1(n28582), .A2(n16876), .ZN(n16930) );
  XOR2HSV0 U20069 ( .A1(n16931), .A2(n16930), .Z(n16932) );
  XOR2HSV0 U20070 ( .A1(n16933), .A2(n16932), .Z(n16934) );
  INHSV2 U20071 ( .I(n16936), .ZN(n16938) );
  NAND3HSV3 U20072 ( .A1(n16939), .A2(n16937), .A3(n16938), .ZN(n16941) );
  NAND2HSV2 U20073 ( .A1(n17119), .A2(\pe10/ti_7t [10]), .ZN(n16940) );
  CLKNAND2HSV4 U20074 ( .A1(n16941), .A2(n16940), .ZN(n16953) );
  NAND2HSV2 U20075 ( .A1(n16942), .A2(n25688), .ZN(n16943) );
  CLKAND2HSV2 U20076 ( .A1(n16943), .A2(n16844), .Z(n16945) );
  INHSV2 U20077 ( .I(n25677), .ZN(n16944) );
  CLKNAND2HSV2 U20078 ( .A1(n16945), .A2(n16944), .ZN(n16947) );
  NOR2HSV2 U20079 ( .A1(n16999), .A2(n25676), .ZN(n16946) );
  CLKAND2HSV2 U20080 ( .A1(n25676), .A2(n17120), .Z(n16949) );
  NAND2HSV0 U20081 ( .A1(n16999), .A2(n16949), .ZN(n16950) );
  INHSV4 U20082 ( .I(n16951), .ZN(n16952) );
  NOR2HSV8 U20083 ( .A1(n16953), .A2(n16952), .ZN(n21737) );
  INHSV4 U20084 ( .I(n21737), .ZN(n20125) );
  INHSV2 U20085 ( .I(n26220), .ZN(n25688) );
  NAND2HSV2 U20086 ( .A1(n16956), .A2(\pe10/ti_7t [8]), .ZN(n20072) );
  INHSV2 U20087 ( .I(n20072), .ZN(n17067) );
  INHSV2 U20088 ( .I(n17067), .ZN(n16957) );
  CLKNAND2HSV3 U20089 ( .A1(n28431), .A2(n16957), .ZN(n16959) );
  AOI21HSV2 U20090 ( .A1(n22442), .A2(n20072), .B(n20065), .ZN(n16958) );
  NAND2HSV0 U20091 ( .A1(n28794), .A2(n28644), .ZN(n16983) );
  NAND2HSV0 U20092 ( .A1(\pe10/aot [9]), .A2(\pe10/bq[13] ), .ZN(n16962) );
  NAND2HSV0 U20093 ( .A1(\pe10/aot [12]), .A2(\pe10/bq[10] ), .ZN(n16961) );
  XOR2HSV0 U20094 ( .A1(n16962), .A2(n16961), .Z(n16966) );
  NAND2HSV0 U20095 ( .A1(\pe10/aot [8]), .A2(\pe10/bq[14] ), .ZN(n16964) );
  NAND2HSV0 U20096 ( .A1(\pe10/aot [7]), .A2(\pe10/bq[15] ), .ZN(n16963) );
  XOR2HSV0 U20097 ( .A1(n16964), .A2(n16963), .Z(n16965) );
  NAND2HSV0 U20098 ( .A1(\pe10/aot [10]), .A2(\pe10/bq[12] ), .ZN(n16968) );
  NAND2HSV0 U20099 ( .A1(\pe10/bq[6] ), .A2(n28424), .ZN(n16967) );
  XOR2HSV0 U20100 ( .A1(n16968), .A2(n16967), .Z(n16972) );
  NAND2HSV0 U20101 ( .A1(\pe10/aot [6]), .A2(n17084), .ZN(n16970) );
  NAND2HSV0 U20102 ( .A1(n22458), .A2(\pe10/got [6]), .ZN(n16969) );
  XOR2HSV0 U20103 ( .A1(n16970), .A2(n16969), .Z(n16971) );
  NAND2HSV0 U20104 ( .A1(\pe10/bq[8] ), .A2(\pe10/aot [14]), .ZN(n16975) );
  NAND2HSV0 U20105 ( .A1(n16973), .A2(\pe10/bq[7] ), .ZN(n16974) );
  XOR2HSV0 U20106 ( .A1(n16975), .A2(n16974), .Z(n16979) );
  BUFHSV2 U20107 ( .I(n14001), .Z(n23544) );
  CLKNAND2HSV1 U20108 ( .A1(n23544), .A2(\pe10/pvq [11]), .ZN(n16977) );
  XNOR2HSV1 U20109 ( .A1(n16977), .A2(\pe10/phq [11]), .ZN(n16978) );
  XNOR2HSV1 U20110 ( .A1(n16979), .A2(n16978), .ZN(n16981) );
  NAND2HSV0 U20111 ( .A1(\pe10/aot [11]), .A2(\pe10/bq[11] ), .ZN(n25217) );
  NAND2HSV0 U20112 ( .A1(\pe10/bq[9] ), .A2(\pe10/aot [13]), .ZN(n26098) );
  XOR2HSV0 U20113 ( .A1(n25217), .A2(n26098), .Z(n16980) );
  NOR2HSV2 U20114 ( .A1(n26200), .A2(n22636), .ZN(n16984) );
  XNOR2HSV4 U20115 ( .A1(n16986), .A2(n16985), .ZN(n16990) );
  NAND2HSV2 U20116 ( .A1(n17119), .A2(\pe10/ti_7t [9]), .ZN(n17000) );
  CLKNHSV0 U20117 ( .I(n17000), .ZN(n16988) );
  AOI21HSV2 U20118 ( .A1(n17000), .A2(n20148), .B(n25261), .ZN(n16987) );
  OAI21HSV2 U20119 ( .A1(n16999), .A2(n16988), .B(n16987), .ZN(n16989) );
  XNOR2HSV4 U20120 ( .A1(n16990), .A2(n16989), .ZN(n21736) );
  NOR2HSV2 U20121 ( .A1(n21736), .A2(n20148), .ZN(n16991) );
  INHSV2 U20122 ( .I(\pe10/ti_7t [11]), .ZN(n16992) );
  NAND2HSV2 U20123 ( .A1(n16992), .A2(n20149), .ZN(n17113) );
  INHSV2 U20124 ( .I(n17113), .ZN(n20066) );
  NOR2HSV2 U20125 ( .A1(n20066), .A2(n25256), .ZN(n16993) );
  INHSV2 U20126 ( .I(n21736), .ZN(n16994) );
  INHSV2 U20127 ( .I(n16995), .ZN(n22419) );
  INHSV2 U20128 ( .I(n22419), .ZN(n22418) );
  NAND2HSV4 U20129 ( .A1(n16996), .A2(n16997), .ZN(n20070) );
  BUFHSV4 U20130 ( .I(n21737), .Z(n28674) );
  CLKNAND2HSV1 U20131 ( .A1(n21741), .A2(\pe10/got [13]), .ZN(n17058) );
  NAND2HSV0 U20132 ( .A1(n17003), .A2(n16844), .ZN(n17005) );
  NAND3HSV0 U20133 ( .A1(n22419), .A2(\pe10/ti_7t [8]), .A3(n26212), .ZN(
        n17001) );
  CLKNAND2HSV0 U20134 ( .A1(n17007), .A2(n17001), .ZN(n17004) );
  NAND2HSV2 U20135 ( .A1(n17007), .A2(n17006), .ZN(n17008) );
  NOR2HSV4 U20136 ( .A1(n17010), .A2(n17009), .ZN(n17056) );
  NAND2HSV0 U20137 ( .A1(n28794), .A2(n28642), .ZN(n17016) );
  NAND2HSV0 U20138 ( .A1(n23474), .A2(\pe10/got [7]), .ZN(n17014) );
  CLKNAND2HSV0 U20139 ( .A1(n22458), .A2(n26132), .ZN(n17012) );
  NAND2HSV0 U20140 ( .A1(\pe10/bq[6] ), .A2(\pe10/aot [14]), .ZN(n17011) );
  XOR2HSV0 U20141 ( .A1(n17012), .A2(n17011), .Z(n17013) );
  XNOR2HSV1 U20142 ( .A1(n17014), .A2(n17013), .ZN(n17015) );
  XNOR2HSV1 U20143 ( .A1(n17016), .A2(n17015), .ZN(n17018) );
  NAND2HSV0 U20144 ( .A1(n26131), .A2(\pe10/got [9]), .ZN(n17017) );
  XNOR2HSV1 U20145 ( .A1(n17018), .A2(n17017), .ZN(n17022) );
  NAND2HSV2 U20146 ( .A1(n17020), .A2(n17019), .ZN(n20074) );
  INHSV2 U20147 ( .I(\pe10/got [10]), .ZN(n26092) );
  OAI21HSV2 U20148 ( .A1(n26092), .A2(n26096), .B(n17022), .ZN(n17021) );
  OAI31HSV2 U20149 ( .A1(n17022), .A2(n26096), .A3(n26092), .B(n17021), .ZN(
        n17054) );
  INHSV2 U20150 ( .I(\pe10/got [5]), .ZN(n26095) );
  NOR2HSV2 U20151 ( .A1(n16907), .A2(n26095), .ZN(n17052) );
  NAND2HSV2 U20152 ( .A1(n28630), .A2(\pe10/got [6]), .ZN(n17051) );
  NAND2HSV0 U20153 ( .A1(\pe10/aot [7]), .A2(\pe10/bq[13] ), .ZN(n17025) );
  NAND2HSV0 U20154 ( .A1(\pe10/aot [6]), .A2(\pe10/bq[14] ), .ZN(n17024) );
  XOR2HSV0 U20155 ( .A1(n17025), .A2(n17024), .Z(n17029) );
  NAND2HSV0 U20156 ( .A1(n28424), .A2(\pe10/bq[4] ), .ZN(n17027) );
  NAND2HSV0 U20157 ( .A1(\pe10/aot [9]), .A2(\pe10/bq[11] ), .ZN(n17026) );
  XOR2HSV0 U20158 ( .A1(n17027), .A2(n17026), .Z(n17028) );
  XOR2HSV0 U20159 ( .A1(n17029), .A2(n17028), .Z(n17037) );
  NAND2HSV0 U20160 ( .A1(\pe10/aot [10]), .A2(\pe10/bq[10] ), .ZN(n17031) );
  NAND2HSV0 U20161 ( .A1(\pe10/aot [11]), .A2(\pe10/bq[9] ), .ZN(n17030) );
  XOR2HSV0 U20162 ( .A1(n17031), .A2(n17030), .Z(n17035) );
  NAND2HSV0 U20163 ( .A1(\pe10/aot [12]), .A2(\pe10/bq[8] ), .ZN(n17033) );
  NAND2HSV0 U20164 ( .A1(\pe10/aot [5]), .A2(\pe10/bq[15] ), .ZN(n17032) );
  XOR2HSV0 U20165 ( .A1(n17033), .A2(n17032), .Z(n17034) );
  XOR2HSV0 U20166 ( .A1(n17035), .A2(n17034), .Z(n17036) );
  XOR2HSV0 U20167 ( .A1(n17037), .A2(n17036), .Z(n17049) );
  NAND2HSV0 U20168 ( .A1(\pe10/aot [8]), .A2(\pe10/bq[12] ), .ZN(n17040) );
  NAND2HSV0 U20169 ( .A1(n16973), .A2(\pe10/bq[5] ), .ZN(n17039) );
  XOR2HSV0 U20170 ( .A1(n17040), .A2(n17039), .Z(n17043) );
  CLKNAND2HSV1 U20171 ( .A1(n23544), .A2(\pe10/pvq [13]), .ZN(n17041) );
  XNOR2HSV1 U20172 ( .A1(n17041), .A2(\pe10/phq [13]), .ZN(n17042) );
  XNOR2HSV1 U20173 ( .A1(n17043), .A2(n17042), .ZN(n17047) );
  NAND2HSV0 U20174 ( .A1(\pe10/aot [13]), .A2(\pe10/bq[7] ), .ZN(n17045) );
  NAND2HSV0 U20175 ( .A1(\pe10/aot [4]), .A2(\pe10/bq[16] ), .ZN(n17044) );
  XOR2HSV0 U20176 ( .A1(n17045), .A2(n17044), .Z(n17046) );
  XNOR2HSV1 U20177 ( .A1(n17047), .A2(n17046), .ZN(n17048) );
  XNOR2HSV1 U20178 ( .A1(n17049), .A2(n17048), .ZN(n17050) );
  XOR3HSV2 U20179 ( .A1(n17052), .A2(n17051), .A3(n17050), .Z(n17053) );
  XOR2HSV0 U20180 ( .A1(n17054), .A2(n17053), .Z(n17055) );
  XOR2HSV2 U20181 ( .A1(n17058), .A2(n17057), .Z(n17059) );
  XNOR2HSV4 U20182 ( .A1(n17060), .A2(n17059), .ZN(n17064) );
  BUFHSV2 U20183 ( .I(n13995), .Z(n26218) );
  AOI21HSV2 U20184 ( .A1(n16669), .A2(n20072), .B(n17065), .ZN(n17066) );
  NOR2HSV2 U20185 ( .A1(n17068), .A2(n22636), .ZN(n17105) );
  NAND2HSV0 U20186 ( .A1(n28794), .A2(\pe10/got [9]), .ZN(n17101) );
  NAND2HSV0 U20187 ( .A1(\pe10/aot [7]), .A2(\pe10/bq[14] ), .ZN(n17070) );
  NAND2HSV0 U20188 ( .A1(\pe10/aot [12]), .A2(\pe10/bq[9] ), .ZN(n17069) );
  XOR2HSV0 U20189 ( .A1(n17070), .A2(n17069), .Z(n17074) );
  NAND2HSV0 U20190 ( .A1(n22458), .A2(\pe10/got [5]), .ZN(n17072) );
  NAND2HSV0 U20191 ( .A1(\pe10/aot [6]), .A2(n16897), .ZN(n17071) );
  XOR2HSV0 U20192 ( .A1(n17072), .A2(n17071), .Z(n17073) );
  XOR2HSV0 U20193 ( .A1(n17074), .A2(n17073), .Z(n17081) );
  NAND2HSV0 U20194 ( .A1(n28424), .A2(\pe10/bq[5] ), .ZN(n17076) );
  NAND2HSV0 U20195 ( .A1(\pe10/bq[7] ), .A2(\pe10/aot [14]), .ZN(n17075) );
  XOR2HSV0 U20196 ( .A1(n17076), .A2(n17075), .Z(n17079) );
  CLKNAND2HSV0 U20197 ( .A1(n16973), .A2(\pe10/bq[6] ), .ZN(n26166) );
  NAND2HSV0 U20198 ( .A1(\pe10/aot [9]), .A2(\pe10/bq[12] ), .ZN(n17077) );
  XOR2HSV0 U20199 ( .A1(n26166), .A2(n17077), .Z(n17078) );
  XOR2HSV0 U20200 ( .A1(n17079), .A2(n17078), .Z(n17080) );
  XOR2HSV0 U20201 ( .A1(n17081), .A2(n17080), .Z(n17097) );
  CLKNAND2HSV1 U20202 ( .A1(n16850), .A2(\pe10/got [7]), .ZN(n17096) );
  NAND2HSV0 U20203 ( .A1(\pe10/aot [13]), .A2(\pe10/bq[8] ), .ZN(n17083) );
  NAND2HSV0 U20204 ( .A1(\pe10/aot [8]), .A2(\pe10/bq[13] ), .ZN(n17082) );
  XOR2HSV0 U20205 ( .A1(n17083), .A2(n17082), .Z(n17088) );
  NAND2HSV0 U20206 ( .A1(\pe10/aot [5]), .A2(n17084), .ZN(n17086) );
  NAND2HSV0 U20207 ( .A1(\pe10/aot [10]), .A2(\pe10/bq[11] ), .ZN(n17085) );
  XOR2HSV0 U20208 ( .A1(n17086), .A2(n17085), .Z(n17087) );
  XOR2HSV0 U20209 ( .A1(n17088), .A2(n17087), .Z(n17092) );
  CLKNAND2HSV1 U20210 ( .A1(n23544), .A2(\pe10/pvq [12]), .ZN(n17089) );
  XNOR2HSV1 U20211 ( .A1(n17089), .A2(\pe10/phq [12]), .ZN(n17090) );
  NAND2HSV0 U20212 ( .A1(\pe10/aot [11]), .A2(\pe10/bq[10] ), .ZN(n20080) );
  XNOR2HSV1 U20213 ( .A1(n17090), .A2(n20080), .ZN(n17091) );
  XNOR2HSV1 U20214 ( .A1(n17092), .A2(n17091), .ZN(n17094) );
  NAND2HSV0 U20215 ( .A1(n26189), .A2(\pe10/got [6]), .ZN(n17093) );
  XOR2HSV0 U20216 ( .A1(n17094), .A2(n17093), .Z(n17095) );
  XOR3HSV2 U20217 ( .A1(n17097), .A2(n17096), .A3(n17095), .Z(n17099) );
  NAND2HSV0 U20218 ( .A1(n23474), .A2(n28642), .ZN(n17098) );
  XNOR2HSV1 U20219 ( .A1(n17099), .A2(n17098), .ZN(n17100) );
  XNOR2HSV1 U20220 ( .A1(n17101), .A2(n17100), .ZN(n17103) );
  NAND2HSV0 U20221 ( .A1(n26131), .A2(n28644), .ZN(n17102) );
  XNOR2HSV1 U20222 ( .A1(n17103), .A2(n17102), .ZN(n17104) );
  NAND2HSV0 U20223 ( .A1(n26094), .A2(n26212), .ZN(n17106) );
  XOR2HSV2 U20224 ( .A1(n17107), .A2(n17106), .Z(n17108) );
  AOI21HSV0 U20225 ( .A1(n20125), .A2(n26218), .B(n17110), .ZN(n17116) );
  NOR2HSV2 U20226 ( .A1(n21737), .A2(n25256), .ZN(n17111) );
  CLKNAND2HSV0 U20227 ( .A1(n17113), .A2(n17112), .ZN(n17122) );
  NOR2HSV0 U20228 ( .A1(n17122), .A2(n22442), .ZN(n17114) );
  CLKNAND2HSV2 U20229 ( .A1(n17124), .A2(n17114), .ZN(n17115) );
  NOR2HSV3 U20230 ( .A1(n17116), .A2(n17115), .ZN(n17118) );
  XNOR2HSV4 U20231 ( .A1(n20125), .A2(n21736), .ZN(n20132) );
  CLKNAND2HSV1 U20232 ( .A1(n17119), .A2(\pe10/ti_7t [12]), .ZN(n22691) );
  INHSV2 U20233 ( .I(n22691), .ZN(n22694) );
  CLKNAND2HSV1 U20234 ( .A1(n22694), .A2(n17120), .ZN(n17121) );
  INHSV3 U20235 ( .I(n17132), .ZN(n17128) );
  INHSV2 U20236 ( .I(n17122), .ZN(n20133) );
  CLKNAND2HSV3 U20237 ( .A1(n20130), .A2(n20133), .ZN(n23715) );
  CLKNAND2HSV1 U20238 ( .A1(n22432), .A2(n25255), .ZN(n17126) );
  INHSV2 U20239 ( .I(n17126), .ZN(n17127) );
  NAND2HSV4 U20240 ( .A1(n23715), .A2(n17127), .ZN(n17130) );
  NAND3HSV4 U20241 ( .A1(n17129), .A2(n17128), .A3(n17130), .ZN(n17135) );
  OAI21HSV4 U20242 ( .A1(n17133), .A2(n17132), .B(n17131), .ZN(n17134) );
  CLKNAND2HSV3 U20243 ( .A1(n17521), .A2(n14056), .ZN(n17167) );
  NAND2HSV2 U20244 ( .A1(n16230), .A2(\pe1/ti_7t [5]), .ZN(n17136) );
  INHSV2 U20245 ( .I(n17136), .ZN(n17216) );
  INHSV2 U20246 ( .I(\pe1/got [14]), .ZN(n17533) );
  AOI21HSV2 U20247 ( .A1(n16182), .A2(n17136), .B(n17533), .ZN(n17137) );
  OAI21HSV2 U20248 ( .A1(n17215), .A2(n17216), .B(n17137), .ZN(n17165) );
  INHSV2 U20249 ( .I(n17172), .ZN(n17301) );
  INHSV2 U20250 ( .I(n17301), .ZN(n17138) );
  NAND2HSV2 U20251 ( .A1(n17138), .A2(\pe1/got [12]), .ZN(n17161) );
  NAND2HSV0 U20252 ( .A1(n17139), .A2(\pe1/got [11]), .ZN(n17147) );
  NAND2HSV0 U20253 ( .A1(n26431), .A2(\pe1/aot [10]), .ZN(n17141) );
  NAND2HSV0 U20254 ( .A1(\pe1/aot [11]), .A2(\pe1/bq[14] ), .ZN(n17140) );
  XOR2HSV0 U20255 ( .A1(n17141), .A2(n17140), .Z(n17145) );
  CLKNAND2HSV0 U20256 ( .A1(\pe1/aot [12]), .A2(\pe1/bq[13] ), .ZN(n26439) );
  NAND2HSV0 U20257 ( .A1(\pe1/aot [14]), .A2(\pe1/bq[11] ), .ZN(n17143) );
  XOR2HSV0 U20258 ( .A1(n26439), .A2(n17143), .Z(n17144) );
  XOR2HSV0 U20259 ( .A1(n17145), .A2(n17144), .Z(n17146) );
  XOR2HSV0 U20260 ( .A1(n17147), .A2(n17146), .Z(n17159) );
  NAND2HSV0 U20261 ( .A1(\pe1/aot [9]), .A2(\pe1/bq[12] ), .ZN(n17445) );
  CLKNHSV0 U20262 ( .I(\pe1/aot [13]), .ZN(n17494) );
  INHSV2 U20263 ( .I(\pe1/aot [9]), .ZN(n27158) );
  OAI22HSV0 U20264 ( .A1(n17494), .A2(n27070), .B1(n27158), .B2(n17302), .ZN(
        n17148) );
  OAI21HSV1 U20265 ( .A1(n17304), .A2(n17445), .B(n17148), .ZN(n17153) );
  CLKNAND2HSV1 U20266 ( .A1(\pe1/aot [15]), .A2(\pe1/bq[9] ), .ZN(n17173) );
  NOR2HSV0 U20267 ( .A1(n17149), .A2(n17173), .ZN(n17151) );
  AOI22HSV0 U20268 ( .A1(\pe1/aot [15]), .A2(\pe1/bq[10] ), .B1(\pe1/aot [16]), 
        .B2(\pe1/bq[9] ), .ZN(n17150) );
  NOR2HSV1 U20269 ( .A1(n17151), .A2(n17150), .ZN(n17152) );
  XOR2HSV0 U20270 ( .A1(n17153), .A2(n17152), .Z(n17157) );
  BUFHSV2 U20271 ( .I(\pe1/got [10]), .Z(n27184) );
  NAND2HSV0 U20272 ( .A1(n26426), .A2(n27184), .ZN(n17156) );
  XOR2HSV0 U20273 ( .A1(n17157), .A2(n17156), .Z(n17158) );
  XNOR2HSV1 U20274 ( .A1(n17159), .A2(n17158), .ZN(n17160) );
  NAND2HSV0 U20275 ( .A1(n17265), .A2(\pe1/got [13]), .ZN(n17162) );
  XNOR2HSV4 U20276 ( .A1(n17165), .A2(n17164), .ZN(n17166) );
  XNOR2HSV4 U20277 ( .A1(n17167), .A2(n17166), .ZN(n23461) );
  XNOR2HSV4 U20278 ( .A1(pov1[7]), .A2(n23461), .ZN(n17168) );
  OA21HSV2 U20279 ( .A1(n17296), .A2(\pe1/ti_7t [8]), .B(n17617), .Z(n17239)
         );
  CLKNAND2HSV3 U20280 ( .A1(n17240), .A2(n17239), .ZN(n17169) );
  CLKNHSV3 U20281 ( .I(n17169), .ZN(n17351) );
  NAND2HSV2 U20282 ( .A1(n17171), .A2(n17170), .ZN(n17209) );
  NAND2HSV0 U20283 ( .A1(n26426), .A2(\pe1/got [9]), .ZN(n17177) );
  INHSV2 U20284 ( .I(n17173), .ZN(n17175) );
  XOR2HSV0 U20285 ( .A1(n17175), .A2(n17174), .Z(n17176) );
  XNOR2HSV1 U20286 ( .A1(n17177), .A2(n17176), .ZN(n17179) );
  NAND2HSV0 U20287 ( .A1(\pe1/aot [8]), .A2(n26436), .ZN(n17181) );
  NAND2HSV0 U20288 ( .A1(\pe1/aot [11]), .A2(\pe1/bq[13] ), .ZN(n17180) );
  XOR2HSV0 U20289 ( .A1(n17181), .A2(n17180), .Z(n17185) );
  NAND2HSV2 U20290 ( .A1(\pe1/aot [9]), .A2(n26548), .ZN(n17183) );
  NAND2HSV0 U20291 ( .A1(\pe1/aot [13]), .A2(\pe1/bq[11] ), .ZN(n17182) );
  XOR2HSV0 U20292 ( .A1(n17183), .A2(n17182), .Z(n17184) );
  XOR2HSV0 U20293 ( .A1(n17185), .A2(n17184), .Z(n17191) );
  NAND2HSV0 U20294 ( .A1(\pe1/aot [10]), .A2(\pe1/bq[14] ), .ZN(n17187) );
  NAND2HSV0 U20295 ( .A1(\pe1/aot [16]), .A2(\pe1/bq[8] ), .ZN(n17186) );
  XOR2HSV0 U20296 ( .A1(n17187), .A2(n17186), .Z(n17189) );
  XNOR2HSV1 U20297 ( .A1(n17189), .A2(n17188), .ZN(n17190) );
  XNOR2HSV1 U20298 ( .A1(n17191), .A2(n17190), .ZN(n17192) );
  XNOR2HSV1 U20299 ( .A1(n17195), .A2(n17194), .ZN(n17197) );
  NAND2HSV2 U20300 ( .A1(n17265), .A2(\pe1/got [12]), .ZN(n17196) );
  XNOR2HSV4 U20301 ( .A1(n17197), .A2(n17196), .ZN(n17205) );
  NAND2HSV2 U20302 ( .A1(n17205), .A2(\pe1/got [14]), .ZN(n17198) );
  INHSV2 U20303 ( .I(n17198), .ZN(n17204) );
  NAND2HSV2 U20304 ( .A1(n17204), .A2(n17199), .ZN(n17202) );
  NOR2HSV0 U20305 ( .A1(n17205), .A2(\pe1/got [14]), .ZN(n17200) );
  CLKNHSV0 U20306 ( .I(n17200), .ZN(n17201) );
  CLKNAND2HSV1 U20307 ( .A1(n17202), .A2(n17201), .ZN(n17203) );
  AOI21HSV2 U20308 ( .A1(n17209), .A2(n17204), .B(n17203), .ZN(n17213) );
  INHSV2 U20309 ( .I(n17205), .ZN(n17206) );
  INHSV2 U20310 ( .I(n17209), .ZN(n17210) );
  NAND2HSV2 U20311 ( .A1(n17211), .A2(n17210), .ZN(n17212) );
  CLKNAND2HSV3 U20312 ( .A1(n17213), .A2(n17212), .ZN(n17220) );
  CLKNAND2HSV2 U20313 ( .A1(n17215), .A2(n17214), .ZN(n21755) );
  INHSV2 U20314 ( .I(n17216), .ZN(n21754) );
  NAND2HSV4 U20315 ( .A1(n21755), .A2(n21754), .ZN(n17554) );
  NAND2HSV0 U20316 ( .A1(n17554), .A2(\pe1/got [13]), .ZN(n17217) );
  INHSV2 U20317 ( .I(n17217), .ZN(n17219) );
  XNOR2HSV4 U20318 ( .A1(n17220), .A2(n17219), .ZN(n17236) );
  NOR2HSV2 U20319 ( .A1(n17236), .A2(n17230), .ZN(n17218) );
  NOR2HSV4 U20320 ( .A1(n17218), .A2(n28802), .ZN(n17350) );
  INHSV3 U20321 ( .I(n17350), .ZN(n17229) );
  XNOR2HSV4 U20322 ( .A1(n17220), .A2(n17219), .ZN(n21749) );
  INHSV4 U20323 ( .I(n21749), .ZN(n17237) );
  INHSV2 U20324 ( .I(n28802), .ZN(n17601) );
  INAND2HSV0 U20325 ( .A1(n17287), .B1(n17601), .ZN(n17221) );
  CLKNAND2HSV1 U20326 ( .A1(n17235), .A2(\pe1/ti_7t [7]), .ZN(n17224) );
  OAI21HSV1 U20327 ( .A1(n16285), .A2(n16182), .B(n17224), .ZN(n17227) );
  NAND3HSV2 U20328 ( .A1(n17225), .A2(n17224), .A3(n17223), .ZN(n17226) );
  OAI21HSV2 U20329 ( .A1(n17228), .A2(n17227), .B(n17226), .ZN(n17553) );
  AND2HSV4 U20330 ( .A1(n17237), .A2(n17553), .Z(n17348) );
  NOR2HSV4 U20331 ( .A1(n17229), .A2(n17348), .ZN(n17231) );
  NAND3HSV2 U20332 ( .A1(n17286), .A2(n17279), .A3(n17543), .ZN(n17273) );
  NAND2HSV2 U20333 ( .A1(n17235), .A2(\pe1/ti_7t [7]), .ZN(n17272) );
  NAND2HSV2 U20334 ( .A1(n17273), .A2(n17272), .ZN(n26541) );
  NAND3HSV4 U20335 ( .A1(n17351), .A2(n17231), .A3(n17347), .ZN(n17407) );
  CLKNHSV0 U20336 ( .I(n17407), .ZN(n17295) );
  CLKNHSV0 U20337 ( .I(n17272), .ZN(n17233) );
  OA21HSV2 U20338 ( .A1(n17233), .A2(n17601), .B(n14056), .Z(n17232) );
  OAI21HSV4 U20339 ( .A1(pov1[7]), .A2(n17233), .B(n17232), .ZN(n21750) );
  INHSV2 U20340 ( .I(n17234), .ZN(n17343) );
  AOI21HSV2 U20341 ( .A1(n17236), .A2(n14007), .B(n17235), .ZN(n17340) );
  CLKNAND2HSV2 U20342 ( .A1(n17343), .A2(n17340), .ZN(n17238) );
  NAND2HSV2 U20343 ( .A1(n17273), .A2(n17272), .ZN(n25880) );
  NOR2HSV2 U20344 ( .A1(n17237), .A2(n25880), .ZN(n17341) );
  CLKNHSV2 U20345 ( .I(n17239), .ZN(n17241) );
  CLKNAND2HSV1 U20346 ( .A1(n28418), .A2(\pe1/got [13]), .ZN(n17271) );
  CLKNAND2HSV0 U20347 ( .A1(n17554), .A2(\pe1/got [12]), .ZN(n17269) );
  INHSV2 U20348 ( .I(n17301), .ZN(n28481) );
  CLKNAND2HSV1 U20349 ( .A1(n28481), .A2(n27184), .ZN(n17264) );
  NAND2HSV0 U20350 ( .A1(n26426), .A2(\pe1/got [8]), .ZN(n17245) );
  NAND2HSV0 U20351 ( .A1(\pe1/aot [8]), .A2(\pe1/bq[15] ), .ZN(n17243) );
  NAND2HSV0 U20352 ( .A1(\pe1/aot [12]), .A2(\pe1/bq[11] ), .ZN(n17242) );
  XOR2HSV0 U20353 ( .A1(n17243), .A2(n17242), .Z(n17244) );
  XNOR2HSV1 U20354 ( .A1(n17245), .A2(n17244), .ZN(n17247) );
  NAND2HSV0 U20355 ( .A1(n26562), .A2(\pe1/got [9]), .ZN(n17246) );
  XOR2HSV0 U20356 ( .A1(n17247), .A2(n17246), .Z(n17262) );
  NAND2HSV0 U20357 ( .A1(\pe1/aot [11]), .A2(\pe1/bq[12] ), .ZN(n17249) );
  NAND2HSV0 U20358 ( .A1(\pe1/aot [13]), .A2(\pe1/bq[10] ), .ZN(n17248) );
  XOR2HSV0 U20359 ( .A1(n17249), .A2(n17248), .Z(n17253) );
  NAND2HSV0 U20360 ( .A1(\pe1/aot [10]), .A2(\pe1/bq[13] ), .ZN(n17251) );
  NAND2HSV0 U20361 ( .A1(\pe1/aot [9]), .A2(\pe1/bq[14] ), .ZN(n17250) );
  XOR2HSV0 U20362 ( .A1(n17251), .A2(n17250), .Z(n17252) );
  XOR2HSV0 U20363 ( .A1(n17253), .A2(n17252), .Z(n17260) );
  NAND2HSV0 U20364 ( .A1(\pe1/aot [14]), .A2(\pe1/bq[9] ), .ZN(n17255) );
  NAND2HSV0 U20365 ( .A1(\pe1/aot [15]), .A2(\pe1/bq[8] ), .ZN(n17254) );
  XOR2HSV0 U20366 ( .A1(n17255), .A2(n17254), .Z(n17258) );
  INHSV2 U20367 ( .I(\pe1/aot [7]), .ZN(n26764) );
  INHSV2 U20368 ( .I(\pe1/bq[7] ), .ZN(n27071) );
  NOR2HSV2 U20369 ( .A1(n26764), .A2(n27071), .ZN(n27025) );
  AOI22HSV0 U20370 ( .A1(\pe1/bq[7] ), .A2(\pe1/aot [16]), .B1(n26436), .B2(
        \pe1/aot [7]), .ZN(n17256) );
  AOI21HSV0 U20371 ( .A1(n27025), .A2(n12023), .B(n17256), .ZN(n17257) );
  XNOR2HSV1 U20372 ( .A1(n17258), .A2(n17257), .ZN(n17259) );
  XNOR2HSV1 U20373 ( .A1(n17260), .A2(n17259), .ZN(n17261) );
  XNOR2HSV1 U20374 ( .A1(n17262), .A2(n17261), .ZN(n17263) );
  XNOR2HSV1 U20375 ( .A1(n17264), .A2(n17263), .ZN(n17267) );
  INHSV2 U20376 ( .I(n17265), .ZN(n21327) );
  INHSV2 U20377 ( .I(n21327), .ZN(n17580) );
  NAND2HSV0 U20378 ( .A1(n17580), .A2(\pe1/got [11]), .ZN(n17266) );
  XNOR2HSV1 U20379 ( .A1(n17267), .A2(n17266), .ZN(n17268) );
  XNOR2HSV1 U20380 ( .A1(n17269), .A2(n17268), .ZN(n17270) );
  XNOR2HSV4 U20381 ( .A1(n17271), .A2(n17270), .ZN(n17274) );
  CLKNHSV2 U20382 ( .I(n17274), .ZN(n17278) );
  NAND2HSV2 U20383 ( .A1(n17273), .A2(n17272), .ZN(n17275) );
  CLKNAND2HSV2 U20384 ( .A1(n17275), .A2(n26595), .ZN(n17277) );
  BUFHSV2 U20385 ( .I(n17279), .Z(n17290) );
  INHSV2 U20386 ( .I(n17290), .ZN(n17281) );
  CLKNAND2HSV0 U20387 ( .A1(n17286), .A2(n17602), .ZN(n17280) );
  NOR2HSV4 U20388 ( .A1(n17281), .A2(n17280), .ZN(n17284) );
  INHSV2 U20389 ( .I(n23461), .ZN(n17283) );
  CLKAND2HSV2 U20390 ( .A1(n16185), .A2(\pe1/ti_7t [8]), .Z(n17282) );
  AOI21HSV4 U20391 ( .A1(n17284), .A2(n17283), .B(n17282), .ZN(n17299) );
  CLKNAND2HSV1 U20392 ( .A1(n23461), .A2(n17601), .ZN(n17285) );
  INHSV2 U20393 ( .I(n17285), .ZN(n17292) );
  CLKNHSV0 U20394 ( .I(n17286), .ZN(n17288) );
  NOR2HSV2 U20395 ( .A1(n17288), .A2(n17287), .ZN(n17289) );
  NAND2HSV2 U20396 ( .A1(n17290), .A2(n17289), .ZN(n17291) );
  CLKNHSV2 U20397 ( .I(n17363), .ZN(n17294) );
  OAI21HSV2 U20398 ( .A1(n17295), .A2(n17294), .B(n12729), .ZN(n17418) );
  NAND3HSV2 U20399 ( .A1(n17419), .A2(n17418), .A3(n17359), .ZN(n17545) );
  INHSV2 U20400 ( .I(n17296), .ZN(n17531) );
  INHSV2 U20401 ( .I(\pe1/ti_7t [10]), .ZN(n17427) );
  AOI21HSV2 U20402 ( .A1(n17531), .A2(n17427), .B(n17598), .ZN(n17546) );
  CLKNAND2HSV2 U20403 ( .A1(n17545), .A2(n17546), .ZN(n17297) );
  INHSV2 U20404 ( .I(n17297), .ZN(n17361) );
  NAND2HSV2 U20405 ( .A1(n17299), .A2(n17298), .ZN(n17402) );
  CLKNAND2HSV1 U20406 ( .A1(n17402), .A2(n26595), .ZN(n17339) );
  INHSV1 U20407 ( .I(n17553), .ZN(n17300) );
  CLKNAND2HSV1 U20408 ( .A1(n17300), .A2(\pe1/got [13]), .ZN(n17337) );
  CLKNAND2HSV1 U20409 ( .A1(n28418), .A2(\pe1/got [12]), .ZN(n17335) );
  NAND2HSV0 U20410 ( .A1(n17554), .A2(\pe1/got [11]), .ZN(n17333) );
  INHSV2 U20411 ( .I(n17301), .ZN(n27005) );
  CLKNAND2HSV1 U20412 ( .A1(n27005), .A2(\pe1/got [9]), .ZN(n17329) );
  NAND2HSV0 U20413 ( .A1(\pe1/aot [6]), .A2(\pe1/bq[9] ), .ZN(n26485) );
  CLKNHSV0 U20414 ( .I(\pe1/aot [6]), .ZN(n26653) );
  NAND2HSV0 U20415 ( .A1(\pe1/bq[9] ), .A2(\pe1/aot [13]), .ZN(n17369) );
  OAI21HSV0 U20416 ( .A1(n26653), .A2(n17302), .B(n17369), .ZN(n17303) );
  OAI21HSV0 U20417 ( .A1(n26485), .A2(n17304), .B(n17303), .ZN(n17306) );
  NAND2HSV0 U20418 ( .A1(\pe1/aot [14]), .A2(\pe1/bq[8] ), .ZN(n17305) );
  XNOR2HSV1 U20419 ( .A1(n17306), .A2(n17305), .ZN(n17308) );
  NAND2HSV0 U20420 ( .A1(n28622), .A2(\pe1/got [7]), .ZN(n17307) );
  XOR2HSV0 U20421 ( .A1(n17308), .A2(n17307), .Z(n17310) );
  NAND2HSV0 U20422 ( .A1(n28814), .A2(\pe1/got [8]), .ZN(n17309) );
  XNOR2HSV1 U20423 ( .A1(n17310), .A2(n17309), .ZN(n17327) );
  NAND2HSV0 U20424 ( .A1(n28468), .A2(\pe1/bq[7] ), .ZN(n17312) );
  NAND2HSV0 U20425 ( .A1(\pe1/bq[6] ), .A2(\pe1/aot [16]), .ZN(n17311) );
  XOR2HSV0 U20426 ( .A1(n17312), .A2(n17311), .Z(n17316) );
  NAND2HSV0 U20427 ( .A1(\pe1/aot [10]), .A2(\pe1/bq[12] ), .ZN(n17314) );
  NAND2HSV0 U20428 ( .A1(\pe1/aot [8]), .A2(\pe1/bq[14] ), .ZN(n17313) );
  XOR2HSV0 U20429 ( .A1(n17314), .A2(n17313), .Z(n17315) );
  XOR2HSV0 U20430 ( .A1(n17316), .A2(n17315), .Z(n17325) );
  NOR2HSV0 U20431 ( .A1(n26764), .A2(n17317), .ZN(n17319) );
  NAND2HSV0 U20432 ( .A1(\pe1/aot [12]), .A2(\pe1/bq[10] ), .ZN(n17318) );
  XOR2HSV0 U20433 ( .A1(n17319), .A2(n17318), .Z(n17323) );
  NAND2HSV0 U20434 ( .A1(\pe1/aot [9]), .A2(\pe1/bq[13] ), .ZN(n17321) );
  NAND2HSV0 U20435 ( .A1(\pe1/aot [11]), .A2(\pe1/bq[11] ), .ZN(n17320) );
  XOR2HSV0 U20436 ( .A1(n17321), .A2(n17320), .Z(n17322) );
  XOR2HSV0 U20437 ( .A1(n17323), .A2(n17322), .Z(n17324) );
  XOR2HSV0 U20438 ( .A1(n17325), .A2(n17324), .Z(n17326) );
  XOR2HSV0 U20439 ( .A1(n17327), .A2(n17326), .Z(n17328) );
  XNOR2HSV1 U20440 ( .A1(n17329), .A2(n17328), .ZN(n17331) );
  CLKNAND2HSV0 U20441 ( .A1(n17580), .A2(n27184), .ZN(n17330) );
  XNOR2HSV1 U20442 ( .A1(n17331), .A2(n17330), .ZN(n17332) );
  XNOR2HSV1 U20443 ( .A1(n17333), .A2(n17332), .ZN(n17334) );
  XNOR2HSV1 U20444 ( .A1(n17335), .A2(n17334), .ZN(n17336) );
  XNOR2HSV1 U20445 ( .A1(n17337), .A2(n17336), .ZN(n17338) );
  XNOR2HSV4 U20446 ( .A1(n17339), .A2(n17338), .ZN(n17355) );
  INHSV2 U20447 ( .I(n17403), .ZN(n21752) );
  CLKNAND2HSV0 U20448 ( .A1(n17340), .A2(n17230), .ZN(n17342) );
  CLKNAND2HSV1 U20449 ( .A1(n17344), .A2(n17343), .ZN(n17345) );
  NOR2HSV4 U20450 ( .A1(n21752), .A2(n17345), .ZN(n17357) );
  INHSV2 U20451 ( .I(n17357), .ZN(n17354) );
  NAND2HSV2 U20452 ( .A1(n17531), .A2(\pe1/ti_7t [9]), .ZN(n17346) );
  INHSV2 U20453 ( .I(n17346), .ZN(n17405) );
  CLKNHSV2 U20454 ( .I(n17347), .ZN(n17349) );
  INHSV3 U20455 ( .I(n17358), .ZN(n17353) );
  NAND3HSV4 U20456 ( .A1(n17355), .A2(n17354), .A3(n17353), .ZN(n17422) );
  INHSV2 U20457 ( .I(n17355), .ZN(n17356) );
  OAI21HSV4 U20458 ( .A1(n17358), .A2(n17357), .B(n17356), .ZN(n17421) );
  CLKNAND2HSV4 U20459 ( .A1(n17422), .A2(n17421), .ZN(n17544) );
  INHSV4 U20460 ( .I(n17544), .ZN(n22082) );
  NOR2HSV2 U20461 ( .A1(n17543), .A2(\pe1/ti_7t [11]), .ZN(n17549) );
  NOR2HSV0 U20462 ( .A1(n17549), .A2(n14007), .ZN(n17360) );
  INHSV2 U20463 ( .I(n17601), .ZN(n22050) );
  NOR2HSV2 U20464 ( .A1(n22082), .A2(n22050), .ZN(n17362) );
  INHSV4 U20465 ( .I(n17361), .ZN(n22083) );
  NAND2HSV4 U20466 ( .A1(n17362), .A2(n22083), .ZN(n17536) );
  INHSV2 U20467 ( .I(n17536), .ZN(n17412) );
  NAND2HSV0 U20468 ( .A1(n26541), .A2(\pe1/got [11]), .ZN(n17401) );
  CLKNAND2HSV0 U20469 ( .A1(n27005), .A2(\pe1/got [7]), .ZN(n17394) );
  NAND2HSV0 U20470 ( .A1(n28434), .A2(n26444), .ZN(n17392) );
  NAND2HSV0 U20471 ( .A1(\pe1/aot [5]), .A2(n26431), .ZN(n17366) );
  NAND2HSV0 U20472 ( .A1(\pe1/aot [10]), .A2(\pe1/bq[10] ), .ZN(n17365) );
  XOR2HSV0 U20473 ( .A1(n17366), .A2(n17365), .Z(n17371) );
  NAND2HSV0 U20474 ( .A1(\pe1/bq[7] ), .A2(\pe1/aot [11]), .ZN(n17556) );
  NAND2HSV0 U20475 ( .A1(\pe1/aot [11]), .A2(\pe1/bq[9] ), .ZN(n17367) );
  OAI21HSV0 U20476 ( .A1(n17494), .A2(n27071), .B(n17367), .ZN(n17368) );
  OAI21HSV0 U20477 ( .A1(n17556), .A2(n17369), .B(n17368), .ZN(n17370) );
  XNOR2HSV1 U20478 ( .A1(n17371), .A2(n17370), .ZN(n17377) );
  CLKNHSV0 U20479 ( .I(\pe1/aot [16]), .ZN(n17372) );
  INHSV2 U20480 ( .I(n17372), .ZN(n28485) );
  NAND2HSV0 U20481 ( .A1(n28485), .A2(\pe1/bq[4] ), .ZN(n26420) );
  NAND2HSV0 U20482 ( .A1(n28468), .A2(\pe1/bq[5] ), .ZN(n26542) );
  NOR2HSV0 U20483 ( .A1(n26659), .A2(n17373), .ZN(n17446) );
  INHSV2 U20484 ( .I(\pe1/bq[4] ), .ZN(n27141) );
  NOR2HSV0 U20485 ( .A1(n27141), .A2(n17374), .ZN(n17501) );
  AOI22HSV1 U20486 ( .A1(n26420), .A2(n26542), .B1(n17446), .B2(n17501), .ZN(
        n17375) );
  NAND2HSV0 U20487 ( .A1(\pe1/aot [14]), .A2(\pe1/bq[6] ), .ZN(n17496) );
  XOR2HSV0 U20488 ( .A1(n17375), .A2(n17496), .Z(n17376) );
  XNOR2HSV1 U20489 ( .A1(n17377), .A2(n17376), .ZN(n17391) );
  NAND2HSV0 U20490 ( .A1(n26426), .A2(\pe1/got [5]), .ZN(n17381) );
  NAND2HSV0 U20491 ( .A1(\pe1/aot [7]), .A2(\pe1/bq[13] ), .ZN(n17379) );
  BUFHSV2 U20492 ( .I(n26436), .Z(n27067) );
  NAND2HSV0 U20493 ( .A1(\pe1/aot [4]), .A2(n27067), .ZN(n17378) );
  XOR2HSV0 U20494 ( .A1(n17379), .A2(n17378), .Z(n17380) );
  XNOR2HSV1 U20495 ( .A1(n17381), .A2(n17380), .ZN(n17389) );
  NAND2HSV0 U20496 ( .A1(\pe1/aot [12]), .A2(\pe1/bq[8] ), .ZN(n17383) );
  NAND2HSV0 U20497 ( .A1(\pe1/aot [8]), .A2(\pe1/bq[12] ), .ZN(n17382) );
  XOR2HSV0 U20498 ( .A1(n17383), .A2(n17382), .Z(n17387) );
  NAND2HSV0 U20499 ( .A1(\pe1/aot [9]), .A2(\pe1/bq[11] ), .ZN(n17385) );
  NAND2HSV0 U20500 ( .A1(\pe1/aot [6]), .A2(\pe1/bq[14] ), .ZN(n17384) );
  XOR2HSV0 U20501 ( .A1(n17385), .A2(n17384), .Z(n17386) );
  XOR2HSV0 U20502 ( .A1(n17387), .A2(n17386), .Z(n17388) );
  XOR2HSV0 U20503 ( .A1(n17389), .A2(n17388), .Z(n17390) );
  XOR3HSV2 U20504 ( .A1(n17392), .A2(n17391), .A3(n17390), .Z(n17393) );
  XNOR2HSV1 U20505 ( .A1(n17394), .A2(n17393), .ZN(n17396) );
  NAND2HSV0 U20506 ( .A1(n17580), .A2(\pe1/got [8]), .ZN(n17395) );
  XNOR2HSV1 U20507 ( .A1(n17396), .A2(n17395), .ZN(n17399) );
  NAND2HSV0 U20508 ( .A1(n11886), .A2(\pe1/got [9]), .ZN(n17398) );
  INHSV2 U20509 ( .I(\pe1/got [10]), .ZN(n26539) );
  INHSV2 U20510 ( .I(n26539), .ZN(n28615) );
  CLKNAND2HSV0 U20511 ( .A1(n28615), .A2(n28418), .ZN(n17397) );
  XOR3HSV2 U20512 ( .A1(n17399), .A2(n17398), .A3(n17397), .Z(n17400) );
  NAND3HSV2 U20513 ( .A1(n17404), .A2(n17403), .A3(n17617), .ZN(n17408) );
  CLKNAND2HSV0 U20514 ( .A1(n17405), .A2(n28422), .ZN(n17406) );
  CLKNAND2HSV1 U20515 ( .A1(n17531), .A2(\pe1/ti_7t [10]), .ZN(n17532) );
  CLKNHSV0 U20516 ( .I(n17532), .ZN(n17410) );
  AOI21HSV1 U20517 ( .A1(n28802), .A2(n17532), .B(n17533), .ZN(n17409) );
  OAI21HSV4 U20518 ( .A1(n17413), .A2(n17412), .B(n17411), .ZN(n17416) );
  CLKNAND2HSV4 U20519 ( .A1(n17416), .A2(n17415), .ZN(n27223) );
  INHSV3 U20520 ( .I(n17479), .ZN(n17417) );
  NAND2HSV2 U20521 ( .A1(n17419), .A2(n17418), .ZN(n17423) );
  CLKNHSV0 U20522 ( .I(n17423), .ZN(n17420) );
  CLKNAND2HSV0 U20523 ( .A1(n17544), .A2(n17420), .ZN(n17426) );
  NAND3HSV2 U20524 ( .A1(n17423), .A2(n17422), .A3(n17421), .ZN(n17424) );
  CLKNAND2HSV1 U20525 ( .A1(n17424), .A2(n17617), .ZN(n17425) );
  INHSV4 U20526 ( .I(n17425), .ZN(n17473) );
  BUFHSV2 U20527 ( .I(n17531), .Z(n22074) );
  AOI21HSV0 U20528 ( .A1(n22074), .A2(n17427), .B(n14007), .ZN(n17428) );
  OAI21HSV2 U20529 ( .A1(n28968), .A2(n22074), .B(n17428), .ZN(n17429) );
  INHSV4 U20530 ( .I(n17429), .ZN(n25680) );
  NAND2HSV0 U20531 ( .A1(n25880), .A2(n28425), .ZN(n17464) );
  NAND2HSV0 U20532 ( .A1(n28481), .A2(\pe1/got [8]), .ZN(n17457) );
  NAND2HSV0 U20533 ( .A1(n26562), .A2(\pe1/got [7]), .ZN(n17455) );
  NAND2HSV0 U20534 ( .A1(\pe1/aot [13]), .A2(\pe1/bq[8] ), .ZN(n17431) );
  NAND2HSV0 U20535 ( .A1(n28468), .A2(\pe1/bq[6] ), .ZN(n17430) );
  XOR2HSV0 U20536 ( .A1(n17431), .A2(n17430), .Z(n17436) );
  CLKNHSV0 U20537 ( .I(n17432), .ZN(n17434) );
  AOI22HSV0 U20538 ( .A1(\pe1/aot [14]), .A2(\pe1/bq[7] ), .B1(\pe1/bq[14] ), 
        .B2(\pe1/aot [7]), .ZN(n17433) );
  AOI21HSV2 U20539 ( .A1(n27025), .A2(n17434), .B(n17433), .ZN(n17435) );
  XNOR2HSV1 U20540 ( .A1(n17436), .A2(n17435), .ZN(n17438) );
  NAND2HSV0 U20541 ( .A1(n28622), .A2(n28434), .ZN(n17437) );
  XNOR2HSV1 U20542 ( .A1(n17438), .A2(n17437), .ZN(n17454) );
  NAND2HSV0 U20543 ( .A1(\pe1/aot [12]), .A2(\pe1/bq[9] ), .ZN(n17440) );
  NAND2HSV0 U20544 ( .A1(\pe1/aot [11]), .A2(\pe1/bq[10] ), .ZN(n17439) );
  XOR2HSV0 U20545 ( .A1(n17440), .A2(n17439), .Z(n17444) );
  NAND2HSV0 U20546 ( .A1(\pe1/aot [6]), .A2(n26548), .ZN(n17442) );
  NAND2HSV0 U20547 ( .A1(\pe1/aot [8]), .A2(\pe1/bq[13] ), .ZN(n17441) );
  XOR2HSV0 U20548 ( .A1(n17442), .A2(n17441), .Z(n17443) );
  XOR2HSV0 U20549 ( .A1(n17444), .A2(n17443), .Z(n17452) );
  XOR2HSV0 U20550 ( .A1(n17446), .A2(n17445), .Z(n17450) );
  NAND2HSV0 U20551 ( .A1(\pe1/bq[11] ), .A2(\pe1/aot [10]), .ZN(n17448) );
  NAND2HSV0 U20552 ( .A1(\pe1/aot [5]), .A2(n26436), .ZN(n17447) );
  XOR2HSV0 U20553 ( .A1(n17448), .A2(n17447), .Z(n17449) );
  XOR2HSV0 U20554 ( .A1(n17450), .A2(n17449), .Z(n17451) );
  XOR2HSV0 U20555 ( .A1(n17452), .A2(n17451), .Z(n17453) );
  XOR3HSV2 U20556 ( .A1(n17455), .A2(n17454), .A3(n17453), .Z(n17456) );
  XNOR2HSV1 U20557 ( .A1(n17457), .A2(n17456), .ZN(n17459) );
  NAND2HSV0 U20558 ( .A1(n17580), .A2(\pe1/got [9]), .ZN(n17458) );
  XNOR2HSV1 U20559 ( .A1(n17459), .A2(n17458), .ZN(n17462) );
  CLKNAND2HSV1 U20560 ( .A1(n11886), .A2(n28615), .ZN(n17461) );
  CLKBUFHSV4 U20561 ( .I(n28418), .Z(n27166) );
  NAND2HSV0 U20562 ( .A1(n27166), .A2(\pe1/got [11]), .ZN(n17460) );
  XOR3HSV2 U20563 ( .A1(n17462), .A2(n17461), .A3(n17460), .Z(n17463) );
  NAND2HSV0 U20564 ( .A1(n25901), .A2(\pe1/got [13]), .ZN(n17465) );
  XNOR2HSV4 U20565 ( .A1(n17468), .A2(n17467), .ZN(n25679) );
  NOR2HSV4 U20566 ( .A1(n25679), .A2(n22074), .ZN(n22071) );
  NAND3HSV2 U20567 ( .A1(n17472), .A2(n17471), .A3(n22071), .ZN(n17469) );
  NAND2HSV2 U20568 ( .A1(n22050), .A2(\pe1/ti_7t [12]), .ZN(n17480) );
  CLKNAND2HSV1 U20569 ( .A1(n17469), .A2(n17480), .ZN(n17470) );
  INHSV2 U20570 ( .I(n17470), .ZN(n17477) );
  CLKNAND2HSV3 U20571 ( .A1(n17472), .A2(n17471), .ZN(n17482) );
  CLKAND2HSV2 U20572 ( .A1(n25679), .A2(n17543), .Z(n17474) );
  NAND3HSV4 U20573 ( .A1(n17482), .A2(n17481), .A3(n17474), .ZN(n22068) );
  INHSV2 U20574 ( .I(n22071), .ZN(n17483) );
  NOR2HSV2 U20575 ( .A1(n17481), .A2(n17483), .ZN(n17475) );
  INHSV2 U20576 ( .I(n17475), .ZN(n17476) );
  NAND3HSV4 U20577 ( .A1(n17477), .A2(n22068), .A3(n17476), .ZN(n22052) );
  CLKBUFHSV4 U20578 ( .I(n22052), .Z(n17542) );
  INHSV4 U20579 ( .I(n17542), .ZN(n22058) );
  NOR2HSV4 U20580 ( .A1(n22075), .A2(n22058), .ZN(n22047) );
  CLKNAND2HSV3 U20581 ( .A1(n17479), .A2(n17478), .ZN(n22056) );
  BUFHSV4 U20582 ( .I(n22052), .Z(n26537) );
  NOR2HSV4 U20583 ( .A1(n22056), .A2(n26537), .ZN(n26825) );
  CLKNAND2HSV1 U20584 ( .A1(n26827), .A2(n17617), .ZN(n22054) );
  CLKNHSV1 U20585 ( .I(n17480), .ZN(n27219) );
  NOR2HSV1 U20586 ( .A1(n17483), .A2(n14007), .ZN(n17484) );
  AOI22HSV2 U20587 ( .A1(n14056), .A2(n27219), .B1(n22072), .B2(n17484), .ZN(
        n17485) );
  OAI21HSV2 U20588 ( .A1(n22068), .A2(n14007), .B(n17485), .ZN(n17541) );
  INAND2HSV1 U20589 ( .A1(n26417), .B1(n12274), .ZN(n17530) );
  CLKNAND2HSV0 U20590 ( .A1(n25880), .A2(n28615), .ZN(n17526) );
  NAND2HSV0 U20591 ( .A1(n28481), .A2(n28434), .ZN(n17518) );
  NAND2HSV0 U20592 ( .A1(n26562), .A2(\pe1/got [5]), .ZN(n17516) );
  NOR2HSV0 U20593 ( .A1(n26764), .A2(n27070), .ZN(n17487) );
  NAND2HSV0 U20594 ( .A1(\pe1/aot [3]), .A2(n26436), .ZN(n17486) );
  XOR2HSV0 U20595 ( .A1(n17487), .A2(n17486), .Z(n17491) );
  NAND2HSV0 U20596 ( .A1(\pe1/aot [10]), .A2(\pe1/bq[9] ), .ZN(n17489) );
  NAND2HSV0 U20597 ( .A1(\pe1/aot [6]), .A2(\pe1/bq[13] ), .ZN(n17488) );
  XOR2HSV0 U20598 ( .A1(n17489), .A2(n17488), .Z(n17490) );
  XOR2HSV0 U20599 ( .A1(n17491), .A2(n17490), .Z(n17500) );
  NAND2HSV0 U20600 ( .A1(\pe1/aot [5]), .A2(\pe1/bq[14] ), .ZN(n17493) );
  NAND2HSV0 U20601 ( .A1(\pe1/bq[3] ), .A2(n28485), .ZN(n17492) );
  XOR2HSV0 U20602 ( .A1(n17493), .A2(n17492), .Z(n17498) );
  NAND2HSV0 U20603 ( .A1(\pe1/aot [13]), .A2(\pe1/bq[5] ), .ZN(n17557) );
  CLKNHSV0 U20604 ( .I(\pe1/bq[6] ), .ZN(n26763) );
  OAI22HSV0 U20605 ( .A1(n17494), .A2(n26763), .B1(n17555), .B2(n26659), .ZN(
        n17495) );
  OAI21HSV0 U20606 ( .A1(n17496), .A2(n17557), .B(n17495), .ZN(n17497) );
  XNOR2HSV1 U20607 ( .A1(n17498), .A2(n17497), .ZN(n17499) );
  XNOR2HSV1 U20608 ( .A1(n17500), .A2(n17499), .ZN(n17515) );
  INHSV2 U20609 ( .I(\pe1/got [4]), .ZN(n26852) );
  NAND2HSV0 U20610 ( .A1(n28622), .A2(n28435), .ZN(n17505) );
  CLKNHSV0 U20611 ( .I(n17501), .ZN(n17503) );
  NAND2HSV0 U20612 ( .A1(\pe1/aot [12]), .A2(\pe1/bq[7] ), .ZN(n17502) );
  XOR2HSV0 U20613 ( .A1(n17503), .A2(n17502), .Z(n17504) );
  XNOR2HSV1 U20614 ( .A1(n17505), .A2(n17504), .ZN(n17513) );
  NAND2HSV0 U20615 ( .A1(\pe1/aot [4]), .A2(n26548), .ZN(n17507) );
  NAND2HSV0 U20616 ( .A1(\pe1/aot [11]), .A2(\pe1/bq[8] ), .ZN(n17506) );
  XOR2HSV0 U20617 ( .A1(n17507), .A2(n17506), .Z(n17511) );
  NAND2HSV0 U20618 ( .A1(\pe1/aot [8]), .A2(\pe1/bq[11] ), .ZN(n17509) );
  NAND2HSV0 U20619 ( .A1(\pe1/aot [9]), .A2(\pe1/bq[10] ), .ZN(n17508) );
  XOR2HSV0 U20620 ( .A1(n17509), .A2(n17508), .Z(n17510) );
  XOR2HSV0 U20621 ( .A1(n17511), .A2(n17510), .Z(n17512) );
  XOR2HSV0 U20622 ( .A1(n17513), .A2(n17512), .Z(n17514) );
  XOR3HSV2 U20623 ( .A1(n17516), .A2(n17515), .A3(n17514), .Z(n17517) );
  XNOR2HSV1 U20624 ( .A1(n17518), .A2(n17517), .ZN(n17520) );
  NAND2HSV0 U20625 ( .A1(n17580), .A2(\pe1/got [7]), .ZN(n17519) );
  XNOR2HSV1 U20626 ( .A1(n17520), .A2(n17519), .ZN(n17524) );
  NAND2HSV0 U20627 ( .A1(n11886), .A2(\pe1/got [8]), .ZN(n17523) );
  NAND2HSV0 U20628 ( .A1(n17521), .A2(\pe1/got [9]), .ZN(n17522) );
  XOR3HSV2 U20629 ( .A1(n17524), .A2(n17523), .A3(n17522), .Z(n17525) );
  XNOR2HSV1 U20630 ( .A1(n17526), .A2(n17525), .ZN(n17528) );
  NAND2HSV0 U20631 ( .A1(n25901), .A2(\pe1/got [11]), .ZN(n17527) );
  XNOR2HSV1 U20632 ( .A1(n17528), .A2(n17527), .ZN(n17529) );
  XNOR2HSV1 U20633 ( .A1(n17530), .A2(n17529), .ZN(n17539) );
  NOR2HSV0 U20634 ( .A1(n17549), .A2(n17533), .ZN(n17535) );
  NAND3HSV2 U20635 ( .A1(n17536), .A2(n17535), .A3(n17534), .ZN(n17537) );
  XOR3HSV2 U20636 ( .A1(n17539), .A2(n17538), .A3(n17537), .Z(n17540) );
  XNOR2HSV4 U20637 ( .A1(n17541), .A2(n17540), .ZN(n22051) );
  CLKNAND2HSV1 U20638 ( .A1(n22082), .A2(n17543), .ZN(n17552) );
  CLKAND2HSV2 U20639 ( .A1(n17544), .A2(n17543), .Z(n17550) );
  CLKNHSV0 U20640 ( .I(n17545), .ZN(n17548) );
  INAND2HSV0 U20641 ( .A1(n17549), .B1(n17546), .ZN(n17547) );
  OAI22HSV2 U20642 ( .A1(n17550), .A2(n17549), .B1(n17548), .B2(n17547), .ZN(
        n17551) );
  OAI21HSV2 U20643 ( .A1(n17552), .A2(n22083), .B(n17551), .ZN(n23456) );
  NOR2HSV2 U20644 ( .A1(n23456), .A2(n17364), .ZN(n17597) );
  NAND2HSV0 U20645 ( .A1(n12274), .A2(\pe1/got [11]), .ZN(n17594) );
  CLKNHSV1 U20646 ( .I(n17553), .ZN(n28609) );
  CLKNAND2HSV1 U20647 ( .A1(n28609), .A2(\pe1/got [9]), .ZN(n17590) );
  NAND2HSV0 U20648 ( .A1(n11886), .A2(\pe1/got [7]), .ZN(n17586) );
  NOR2HSV0 U20649 ( .A1(n17555), .A2(n27141), .ZN(n26556) );
  NAND2HSV0 U20650 ( .A1(\pe1/bq[13] ), .A2(\pe1/aot [5]), .ZN(n27021) );
  NAND2HSV0 U20651 ( .A1(\pe1/got [4]), .A2(n26444), .ZN(n17558) );
  XOR2HSV0 U20652 ( .A1(n17559), .A2(n17558), .Z(n17584) );
  NAND2HSV0 U20653 ( .A1(n27005), .A2(\pe1/got [5]), .ZN(n17583) );
  NAND2HSV0 U20654 ( .A1(\pe1/aot [4]), .A2(\pe1/bq[14] ), .ZN(n17561) );
  NAND2HSV0 U20655 ( .A1(\pe1/aot [3]), .A2(n26431), .ZN(n17560) );
  XOR2HSV0 U20656 ( .A1(n17561), .A2(n17560), .Z(n17565) );
  NAND2HSV0 U20657 ( .A1(\pe1/aot [2]), .A2(n27067), .ZN(n17563) );
  NAND2HSV0 U20658 ( .A1(\pe1/aot [7]), .A2(\pe1/bq[11] ), .ZN(n17562) );
  XOR2HSV0 U20659 ( .A1(n17563), .A2(n17562), .Z(n17564) );
  XOR2HSV0 U20660 ( .A1(n17565), .A2(n17564), .Z(n17572) );
  NAND2HSV0 U20661 ( .A1(\pe1/aot [10]), .A2(\pe1/bq[8] ), .ZN(n17567) );
  NAND2HSV0 U20662 ( .A1(\pe1/aot [6]), .A2(\pe1/bq[12] ), .ZN(n17566) );
  XOR2HSV0 U20663 ( .A1(n17567), .A2(n17566), .Z(n17570) );
  NAND2HSV0 U20664 ( .A1(n28468), .A2(\pe1/bq[3] ), .ZN(n26421) );
  NAND2HSV0 U20665 ( .A1(\pe1/aot [12]), .A2(\pe1/bq[6] ), .ZN(n17568) );
  XOR2HSV0 U20666 ( .A1(n26421), .A2(n17568), .Z(n17569) );
  XOR2HSV0 U20667 ( .A1(n17570), .A2(n17569), .Z(n17571) );
  XOR2HSV0 U20668 ( .A1(n17572), .A2(n17571), .Z(n17579) );
  NAND2HSV0 U20669 ( .A1(\pe1/aot [8]), .A2(\pe1/bq[10] ), .ZN(n17574) );
  INHSV2 U20670 ( .I(\pe1/bq[2] ), .ZN(n26652) );
  NAND2HSV0 U20671 ( .A1(n28485), .A2(\pe1/bq[2] ), .ZN(n17573) );
  XOR2HSV0 U20672 ( .A1(n17574), .A2(n17573), .Z(n17575) );
  NAND2HSV0 U20673 ( .A1(\pe1/aot [9]), .A2(\pe1/bq[9] ), .ZN(n26487) );
  XNOR2HSV1 U20674 ( .A1(n17575), .A2(n26487), .ZN(n17577) );
  NAND2HSV0 U20675 ( .A1(n26426), .A2(\pe1/got [3]), .ZN(n17576) );
  XNOR2HSV1 U20676 ( .A1(n17577), .A2(n17576), .ZN(n17578) );
  XNOR2HSV1 U20677 ( .A1(n17579), .A2(n17578), .ZN(n17582) );
  CLKNAND2HSV0 U20678 ( .A1(n17580), .A2(n28434), .ZN(n17581) );
  XOR4HSV1 U20679 ( .A1(n17584), .A2(n17583), .A3(n17582), .A4(n17581), .Z(
        n17585) );
  XNOR2HSV1 U20680 ( .A1(n17586), .A2(n17585), .ZN(n17588) );
  NAND2HSV0 U20681 ( .A1(n27166), .A2(\pe1/got [8]), .ZN(n17587) );
  XNOR2HSV1 U20682 ( .A1(n17588), .A2(n17587), .ZN(n17589) );
  XNOR2HSV1 U20683 ( .A1(n17590), .A2(n17589), .ZN(n17592) );
  CLKNAND2HSV0 U20684 ( .A1(n25901), .A2(n28615), .ZN(n17591) );
  XNOR2HSV1 U20685 ( .A1(n17592), .A2(n17591), .ZN(n17593) );
  XNOR2HSV1 U20686 ( .A1(n17594), .A2(n17593), .ZN(n17595) );
  CLKXOR2HSV4 U20687 ( .A1(n17597), .A2(n17596), .Z(n17600) );
  XNOR2HSV4 U20688 ( .A1(n17599), .A2(n17600), .ZN(n23431) );
  INHSV2 U20689 ( .I(n23431), .ZN(n17622) );
  NOR2HSV2 U20690 ( .A1(n17622), .A2(n17598), .ZN(n17614) );
  OR2HSV1 U20691 ( .A1(n17616), .A2(n22051), .Z(n17613) );
  INHSV2 U20692 ( .I(n26825), .ZN(n17610) );
  NAND2HSV0 U20693 ( .A1(n27223), .A2(n17602), .ZN(n17603) );
  CLKNHSV1 U20694 ( .I(n17603), .ZN(n17604) );
  BUFHSV4 U20695 ( .I(n22052), .Z(n28460) );
  NOR2HSV2 U20696 ( .A1(n27223), .A2(n17605), .ZN(n26822) );
  CLKNHSV0 U20697 ( .I(n26827), .ZN(n17606) );
  OR2HSV1 U20698 ( .A1(n17606), .A2(n14007), .Z(n17607) );
  NOR2HSV2 U20699 ( .A1(n26822), .A2(n17607), .ZN(n17608) );
  CLKAND2HSV2 U20700 ( .A1(n26824), .A2(n17608), .Z(n17609) );
  CLKNAND2HSV4 U20701 ( .A1(n17610), .A2(n17609), .ZN(n23432) );
  INOR2HSV1 U20702 ( .A1(\pe1/ti_7t [15]), .B1(n17615), .ZN(n25875) );
  NOR2HSV4 U20703 ( .A1(n25874), .A2(n25875), .ZN(n26481) );
  NOR2HSV2 U20704 ( .A1(n17616), .A2(n17287), .ZN(n17620) );
  INAND2HSV2 U20705 ( .A1(n17617), .B1(n23431), .ZN(n17618) );
  NAND3HSV3 U20706 ( .A1(n17618), .A2(n17214), .A3(n23432), .ZN(n17619) );
  AOI21HSV4 U20707 ( .A1(n13962), .A2(n17620), .B(n17619), .ZN(n17621) );
  INHSV2 U20708 ( .I(\pe2/phq [2]), .ZN(n17623) );
  CLKNAND2HSV2 U20709 ( .A1(n17782), .A2(n17623), .ZN(n17625) );
  CLKNAND2HSV2 U20710 ( .A1(n17668), .A2(n17623), .ZN(n17624) );
  NAND3HSV4 U20711 ( .A1(n17625), .A2(n17626), .A3(n17624), .ZN(n17628) );
  CLKBUFHSV4 U20712 ( .I(\pe2/ctrq ), .Z(n17831) );
  NAND2HSV2 U20713 ( .A1(n17831), .A2(\pe2/pvq [2]), .ZN(n17629) );
  INHSV2 U20714 ( .I(n17629), .ZN(n17627) );
  CLKNAND2HSV2 U20715 ( .A1(n17630), .A2(n17629), .ZN(n17631) );
  NAND2HSV4 U20716 ( .A1(n17632), .A2(n17631), .ZN(n17655) );
  CLKNHSV0 U20717 ( .I(n17635), .ZN(n17634) );
  INHSV6 U20718 ( .I(\pe2/bq[16] ), .ZN(n27322) );
  NAND2HSV0 U20719 ( .A1(\pe2/aot [15]), .A2(n21842), .ZN(n17633) );
  CLKNAND2HSV1 U20720 ( .A1(n17634), .A2(n17633), .ZN(n17637) );
  XNOR2HSV4 U20721 ( .A1(n17655), .A2(n17654), .ZN(n17646) );
  CLKNAND2HSV2 U20722 ( .A1(\pe2/bq[16] ), .A2(\pe2/aot [16]), .ZN(n17638) );
  IOA21HSV4 U20723 ( .A1(\pe2/pvq [1]), .A2(\pe2/ctrq ), .B(n17638), .ZN(
        n17639) );
  CLKAND2HSV2 U20724 ( .A1(\pe2/phq [1]), .A2(\pe2/got [16]), .Z(n17641) );
  INHSV4 U20725 ( .I(n17782), .ZN(n17752) );
  AOI21HSV2 U20726 ( .A1(\pe2/ti_1 ), .A2(\pe2/got [16]), .B(\pe2/phq [1]), 
        .ZN(n17640) );
  AOI21HSV4 U20727 ( .A1(n17641), .A2(n17752), .B(n17640), .ZN(n17649) );
  CLKNAND2HSV0 U20728 ( .A1(n17649), .A2(n17650), .ZN(n17643) );
  INHSV2 U20729 ( .I(n17649), .ZN(n17647) );
  CLKNAND2HSV1 U20730 ( .A1(n17648), .A2(n17647), .ZN(n17642) );
  CLKBUFHSV4 U20731 ( .I(n17808), .Z(n21011) );
  INHSV2 U20732 ( .I(n21011), .ZN(n17714) );
  INHSV2 U20733 ( .I(\pe2/got [16]), .ZN(n17651) );
  INHSV2 U20734 ( .I(n21234), .ZN(n21168) );
  NOR2HSV4 U20735 ( .A1(n17714), .A2(n21168), .ZN(n21696) );
  INHSV2 U20736 ( .I(n17644), .ZN(n17645) );
  NAND2HSV4 U20737 ( .A1(n17646), .A2(n17645), .ZN(n17687) );
  BUFHSV2 U20738 ( .I(n17808), .Z(n17819) );
  INHSV2 U20739 ( .I(n17819), .ZN(n28932) );
  NAND2HSV2 U20740 ( .A1(n28932), .A2(\pe2/ti_7t [2]), .ZN(n17686) );
  NAND2HSV2 U20741 ( .A1(n17650), .A2(n17649), .ZN(n17672) );
  CLKNAND2HSV2 U20742 ( .A1(n17671), .A2(n17672), .ZN(n17699) );
  CLKNAND2HSV1 U20743 ( .A1(n17699), .A2(n28693), .ZN(n17653) );
  INHSV2 U20744 ( .I(n21011), .ZN(n21159) );
  CLKNAND2HSV2 U20745 ( .A1(n17653), .A2(n17652), .ZN(n17688) );
  XNOR2HSV4 U20746 ( .A1(n17655), .A2(n17654), .ZN(n25630) );
  OAI21HSV4 U20747 ( .A1(n17656), .A2(n17701), .B(n21234), .ZN(n17749) );
  CLKNAND2HSV1 U20748 ( .A1(\pe2/ctrq ), .A2(\pe2/pvq [3]), .ZN(n17658) );
  XNOR2HSV4 U20749 ( .A1(n17658), .A2(n17657), .ZN(n17661) );
  CLKXOR2HSV4 U20750 ( .A1(n17659), .A2(\pe2/phq [3]), .Z(n17660) );
  XNOR2HSV4 U20751 ( .A1(n17661), .A2(n17660), .ZN(n17664) );
  INAND2HSV2 U20752 ( .A1(n27322), .B1(\pe2/aot [14]), .ZN(n17663) );
  NAND2HSV0 U20753 ( .A1(\pe2/aot [15]), .A2(\pe2/bq[15] ), .ZN(n17662) );
  INHSV3 U20754 ( .I(n21011), .ZN(n21901) );
  INHSV2 U20755 ( .I(\pe2/ti_7t [1]), .ZN(n17673) );
  CLKBUFHSV4 U20756 ( .I(n17808), .Z(n21813) );
  CLKNHSV0 U20757 ( .I(n21813), .ZN(n21289) );
  AOI21HSV2 U20758 ( .A1(n17673), .A2(n21289), .B(n21225), .ZN(n17665) );
  OAI21HSV2 U20759 ( .A1(n17666), .A2(n21901), .B(n17665), .ZN(n17667) );
  XNOR2HSV4 U20760 ( .A1(n17700), .A2(n17667), .ZN(n17748) );
  CLKXOR2HSV4 U20761 ( .A1(n17749), .A2(n17748), .Z(n17670) );
  NAND2HSV2 U20762 ( .A1(n17702), .A2(n21702), .ZN(n17669) );
  AOI21HSV4 U20763 ( .A1(n17670), .A2(n17652), .B(n17669), .ZN(n17692) );
  NAND2HSV2 U20764 ( .A1(n17672), .A2(n17671), .ZN(n28454) );
  NOR2HSV2 U20765 ( .A1(n21813), .A2(n17673), .ZN(n17698) );
  INHSV2 U20766 ( .I(n17698), .ZN(n17715) );
  CLKBUFHSV4 U20767 ( .I(n17831), .Z(n21253) );
  NAND2HSV0 U20768 ( .A1(\pe2/aot [15]), .A2(\pe2/bq[13] ), .ZN(n17675) );
  NAND2HSV0 U20769 ( .A1(\pe2/bq[12] ), .A2(\pe2/aot [16]), .ZN(n17674) );
  XNOR2HSV1 U20770 ( .A1(n17675), .A2(n17674), .ZN(n17676) );
  CLKNAND2HSV1 U20771 ( .A1(n17752), .A2(\pe2/got [12]), .ZN(n17679) );
  NAND2HSV0 U20772 ( .A1(\pe2/aot [13]), .A2(\pe2/bq[15] ), .ZN(n17678) );
  XOR2HSV0 U20773 ( .A1(n17679), .A2(n17678), .Z(n17683) );
  INAND2HSV2 U20774 ( .A1(n27322), .B1(\pe2/aot [12]), .ZN(n17680) );
  XNOR2HSV4 U20775 ( .A1(n17681), .A2(n17680), .ZN(n17682) );
  XNOR2HSV4 U20776 ( .A1(n17683), .A2(n17682), .ZN(n17684) );
  XNOR2HSV4 U20777 ( .A1(n17685), .A2(n17684), .ZN(n17690) );
  NOR2HSV4 U20778 ( .A1(n17688), .A2(n25630), .ZN(n17707) );
  NOR2HSV4 U20779 ( .A1(n17708), .A2(n17707), .ZN(n21066) );
  INHSV2 U20780 ( .I(\pe2/got [14]), .ZN(n21164) );
  XNOR3HSV2 U20781 ( .A1(n17691), .A2(n17690), .A3(n17689), .ZN(n17693) );
  INHSV2 U20782 ( .I(n17693), .ZN(n17694) );
  CLKAND2HSV2 U20783 ( .A1(n28932), .A2(\pe2/ti_7t [5]), .Z(n17742) );
  INHSV2 U20784 ( .I(n17742), .ZN(n17696) );
  CLKNAND2HSV3 U20785 ( .A1(n17697), .A2(n17696), .ZN(n17745) );
  CLKNHSV0 U20786 ( .I(n17708), .ZN(n17705) );
  NOR2HSV2 U20787 ( .A1(n17699), .A2(n17698), .ZN(n17713) );
  NOR2HSV1 U20788 ( .A1(n17701), .A2(n21235), .ZN(n17704) );
  CLKNAND2HSV1 U20789 ( .A1(n17702), .A2(n28693), .ZN(n17703) );
  AOI31HSV2 U20790 ( .A1(n17705), .A2(n17706), .A3(n17704), .B(n17703), .ZN(
        n17711) );
  NOR2HSV4 U20791 ( .A1(n17708), .A2(n17707), .ZN(n17737) );
  INHSV2 U20792 ( .I(n17737), .ZN(n17712) );
  CLKNAND2HSV3 U20793 ( .A1(n17710), .A2(n17711), .ZN(n17747) );
  INHSV2 U20794 ( .I(n21702), .ZN(n17736) );
  INHSV2 U20795 ( .I(n17713), .ZN(n17717) );
  AOI21HSV1 U20796 ( .A1(n17715), .A2(n17714), .B(n21164), .ZN(n17716) );
  CLKNAND2HSV1 U20797 ( .A1(n17717), .A2(n17716), .ZN(n17729) );
  NAND2HSV2 U20798 ( .A1(\pe2/got [13]), .A2(\pe2/ti_1 ), .ZN(n17720) );
  XNOR2HSV4 U20799 ( .A1(n17721), .A2(n17720), .ZN(n17722) );
  XNOR2HSV4 U20800 ( .A1(n17723), .A2(n17722), .ZN(n17728) );
  INAND2HSV2 U20801 ( .A1(n27322), .B1(\pe2/aot [13]), .ZN(n17725) );
  XNOR2HSV4 U20802 ( .A1(n17726), .A2(n17725), .ZN(n17727) );
  XNOR2HSV4 U20803 ( .A1(n17728), .A2(n17727), .ZN(n17730) );
  CLKNAND2HSV1 U20804 ( .A1(n17729), .A2(n17730), .ZN(n17733) );
  CLKNAND2HSV3 U20805 ( .A1(n17735), .A2(n17734), .ZN(n17741) );
  NOR2HSV2 U20806 ( .A1(n17737), .A2(n17736), .ZN(n17739) );
  CLKNAND2HSV1 U20807 ( .A1(n17739), .A2(n17738), .ZN(n17740) );
  XNOR2HSV4 U20808 ( .A1(n17747), .A2(n17746), .ZN(n29043) );
  AOI21HSV2 U20809 ( .A1(n27354), .A2(n21116), .B(n17742), .ZN(n17743) );
  OAI21HSV4 U20810 ( .A1(n29043), .A2(n21289), .B(n17743), .ZN(n17744) );
  CLKAND2HSV2 U20811 ( .A1(n21235), .A2(\pe2/ti_7t [3]), .Z(n17798) );
  AOI21HSV2 U20812 ( .A1(n29044), .A2(n17829), .B(n17798), .ZN(n21118) );
  INHSV2 U20813 ( .I(\pe2/got [13]), .ZN(n21305) );
  NOR2HSV2 U20814 ( .A1(n21118), .A2(n21305), .ZN(n17766) );
  CLKNAND2HSV1 U20815 ( .A1(n21065), .A2(n27543), .ZN(n17763) );
  CLKBUFHSV4 U20816 ( .I(\pe2/ctrq ), .Z(n22114) );
  NAND2HSV0 U20817 ( .A1(\pe2/bq[11] ), .A2(\pe2/aot [15]), .ZN(n27255) );
  NAND2HSV0 U20818 ( .A1(\pe2/aot [11]), .A2(\pe2/bq[15] ), .ZN(n17750) );
  CLKNHSV0 U20819 ( .I(n27255), .ZN(n17751) );
  CLKNAND2HSV1 U20820 ( .A1(\pe2/got [10]), .A2(n17752), .ZN(n17754) );
  NAND2HSV0 U20821 ( .A1(\pe2/aot [14]), .A2(\pe2/bq[12] ), .ZN(n17753) );
  XOR2HSV0 U20822 ( .A1(n17754), .A2(n17753), .Z(n17758) );
  NAND2HSV0 U20823 ( .A1(\pe2/aot [13]), .A2(\pe2/bq[13] ), .ZN(n17756) );
  NAND2HSV0 U20824 ( .A1(\pe2/aot [12]), .A2(\pe2/bq[14] ), .ZN(n17755) );
  XOR2HSV0 U20825 ( .A1(n17756), .A2(n17755), .Z(n17757) );
  XOR2HSV0 U20826 ( .A1(n17758), .A2(n17757), .Z(n17759) );
  XOR3HSV2 U20827 ( .A1(n17761), .A2(n17760), .A3(n17759), .Z(n17762) );
  INHSV2 U20828 ( .I(\pe2/got [12]), .ZN(n21645) );
  NOR2HSV1 U20829 ( .A1(n21066), .A2(n21645), .ZN(n17764) );
  NAND2HSV2 U20830 ( .A1(n28932), .A2(\pe2/ti_7t [4]), .ZN(n17826) );
  INHSV2 U20831 ( .I(n17826), .ZN(n17772) );
  INHSV2 U20832 ( .I(\pe2/got [14]), .ZN(n21880) );
  OAI21HSV2 U20833 ( .A1(n17772), .A2(n21641), .B(n17767), .ZN(n17768) );
  INHSV2 U20834 ( .I(n17768), .ZN(n17769) );
  OAI21HSV4 U20835 ( .A1(n29043), .A2(n17772), .B(n17769), .ZN(n17815) );
  NOR2HSV2 U20836 ( .A1(n21260), .A2(n21305), .ZN(n17796) );
  INAND2HSV2 U20837 ( .A1(n27322), .B1(\pe2/aot [11]), .ZN(n17780) );
  NAND2HSV0 U20838 ( .A1(\pe2/aot [13]), .A2(\pe2/bq[14] ), .ZN(n17776) );
  NAND2HSV0 U20839 ( .A1(\pe2/aot [12]), .A2(\pe2/bq[15] ), .ZN(n17775) );
  CLKXOR2HSV4 U20840 ( .A1(n17776), .A2(n17775), .Z(n17779) );
  NAND2HSV0 U20841 ( .A1(n22114), .A2(\pe2/pvq [6]), .ZN(n17777) );
  XNOR2HSV1 U20842 ( .A1(n17777), .A2(\pe2/phq [6]), .ZN(n17778) );
  XOR3HSV2 U20843 ( .A1(n17780), .A2(n17779), .A3(n17778), .Z(n17791) );
  INHSV2 U20844 ( .I(n17782), .ZN(n21269) );
  NAND2HSV2 U20845 ( .A1(\pe2/got [11]), .A2(n21269), .ZN(n17784) );
  NAND2HSV0 U20846 ( .A1(\pe2/aot [14]), .A2(\pe2/bq[13] ), .ZN(n17783) );
  XOR2HSV0 U20847 ( .A1(n17784), .A2(n17783), .Z(n17789) );
  NAND2HSV0 U20848 ( .A1(\pe2/aot [15]), .A2(\pe2/bq[12] ), .ZN(n17787) );
  XOR2HSV2 U20849 ( .A1(n17789), .A2(n17788), .Z(n17790) );
  XNOR2HSV4 U20850 ( .A1(n17791), .A2(n17790), .ZN(n17794) );
  NAND2HSV0 U20851 ( .A1(n21065), .A2(\pe2/got [12]), .ZN(n17793) );
  XNOR2HSV4 U20852 ( .A1(n17794), .A2(n17793), .ZN(n17795) );
  XNOR2HSV4 U20853 ( .A1(n17796), .A2(n17795), .ZN(n17803) );
  INAND2HSV2 U20854 ( .A1(n21164), .B1(n17829), .ZN(n17797) );
  CLKNAND2HSV1 U20855 ( .A1(n17798), .A2(n21144), .ZN(n17799) );
  CLKNHSV2 U20856 ( .I(n17801), .ZN(n17802) );
  XNOR2HSV4 U20857 ( .A1(n17803), .A2(n17802), .ZN(n17806) );
  OAI21HSV4 U20858 ( .A1(n17807), .A2(n17806), .B(n17805), .ZN(n17861) );
  INHSV2 U20859 ( .I(n21009), .ZN(n17814) );
  XNOR2HSV4 U20860 ( .A1(n17807), .A2(n17806), .ZN(n21022) );
  CLKNAND2HSV1 U20861 ( .A1(n28809), .A2(n21813), .ZN(n17811) );
  BUFHSV2 U20862 ( .I(n17808), .Z(n21713) );
  CLKNHSV1 U20863 ( .I(n17864), .ZN(n17809) );
  INHSV2 U20864 ( .I(n21234), .ZN(n21116) );
  NOR2HSV2 U20865 ( .A1(n17809), .A2(n21116), .ZN(n17810) );
  OAI21HSV4 U20866 ( .A1(n21022), .A2(n17811), .B(n17810), .ZN(n21007) );
  NAND2HSV2 U20867 ( .A1(n21701), .A2(\pe2/ti_7t [7]), .ZN(n21008) );
  NOR2HSV2 U20868 ( .A1(n21008), .A2(n21116), .ZN(n17812) );
  AOI31HSV2 U20869 ( .A1(n21005), .A2(n17814), .A3(n17813), .B(n17812), .ZN(
        n17825) );
  XNOR2HSV4 U20870 ( .A1(n17816), .A2(n17815), .ZN(n21012) );
  MUX2HSV2 U20871 ( .I0(n17862), .I1(n27121), .S(n21012), .Z(n17817) );
  CLKNAND2HSV1 U20872 ( .A1(n17817), .A2(n21234), .ZN(n17821) );
  CLKBUFHSV4 U20873 ( .I(n17818), .Z(n21018) );
  INHSV4 U20874 ( .I(n14044), .ZN(n27485) );
  OAI21HSV2 U20875 ( .A1(n21018), .A2(n27485), .B(n17819), .ZN(n17820) );
  NOR2HSV2 U20876 ( .A1(n17821), .A2(n17820), .ZN(n17823) );
  NOR2HSV4 U20877 ( .A1(n21009), .A2(n21007), .ZN(n27123) );
  INHSV2 U20878 ( .I(n27123), .ZN(n17822) );
  NAND2HSV2 U20879 ( .A1(n17823), .A2(n17822), .ZN(n17824) );
  INHSV2 U20880 ( .I(\pe2/got [13]), .ZN(n21117) );
  AND2HSV2 U20881 ( .A1(n21701), .A2(\pe2/ti_7t [3]), .Z(n17828) );
  AOI21HSV2 U20882 ( .A1(n29044), .A2(n17829), .B(n17828), .ZN(n21278) );
  NOR2HSV2 U20883 ( .A1(n21278), .A2(n21645), .ZN(n17852) );
  NAND2HSV0 U20884 ( .A1(n21065), .A2(\pe2/got [10]), .ZN(n17851) );
  AND2HSV4 U20885 ( .A1(n17830), .A2(\pe2/got [11]), .Z(n17850) );
  CLKNAND2HSV0 U20886 ( .A1(n17831), .A2(\pe2/pvq [8]), .ZN(n17832) );
  XNOR2HSV1 U20887 ( .A1(n17832), .A2(\pe2/phq [8]), .ZN(n17833) );
  INHSV2 U20888 ( .I(\pe2/bq[9] ), .ZN(n23502) );
  NOR2HSV2 U20889 ( .A1(n21254), .A2(n23502), .ZN(n21130) );
  XNOR2HSV1 U20890 ( .A1(n17833), .A2(n21130), .ZN(n17848) );
  NAND2HSV0 U20891 ( .A1(\pe2/aot [13]), .A2(\pe2/bq[12] ), .ZN(n17835) );
  NAND2HSV0 U20892 ( .A1(\pe2/aot [12]), .A2(\pe2/bq[13] ), .ZN(n17834) );
  XOR2HSV0 U20893 ( .A1(n17835), .A2(n17834), .Z(n17839) );
  NAND2HSV0 U20894 ( .A1(\pe2/aot [11]), .A2(n27312), .ZN(n17837) );
  INHSV2 U20895 ( .I(\pe2/got [9]), .ZN(n21103) );
  INHSV2 U20896 ( .I(n21103), .ZN(n21246) );
  CLKNAND2HSV0 U20897 ( .A1(n21246), .A2(n21269), .ZN(n17836) );
  XOR2HSV0 U20898 ( .A1(n17837), .A2(n17836), .Z(n17838) );
  XNOR2HSV1 U20899 ( .A1(n17839), .A2(n17838), .ZN(n17847) );
  NAND2HSV0 U20900 ( .A1(\pe2/aot [15]), .A2(\pe2/bq[10] ), .ZN(n17841) );
  NAND2HSV0 U20901 ( .A1(\pe2/aot [10]), .A2(\pe2/bq[15] ), .ZN(n17840) );
  XOR2HSV0 U20902 ( .A1(n17841), .A2(n17840), .Z(n17845) );
  INAND2HSV2 U20903 ( .A1(n27322), .B1(\pe2/aot [9]), .ZN(n17843) );
  NAND2HSV0 U20904 ( .A1(\pe2/aot [14]), .A2(\pe2/bq[11] ), .ZN(n17842) );
  XOR2HSV0 U20905 ( .A1(n17843), .A2(n17842), .Z(n17844) );
  XOR2HSV0 U20906 ( .A1(n17845), .A2(n17844), .Z(n17846) );
  XOR3HSV2 U20907 ( .A1(n17848), .A2(n17847), .A3(n17846), .Z(n17849) );
  NAND2HSV2 U20908 ( .A1(n17855), .A2(\pe2/got [14]), .ZN(n17856) );
  CLKNAND2HSV2 U20909 ( .A1(n17859), .A2(n17858), .ZN(n17860) );
  CLKNAND2HSV3 U20910 ( .A1(n17860), .A2(n28693), .ZN(n21021) );
  XNOR2HSV4 U20911 ( .A1(n17861), .A2(n21021), .ZN(n17866) );
  INHSV4 U20912 ( .I(n17863), .ZN(n28421) );
  NAND2HSV2 U20913 ( .A1(n17864), .A2(n28421), .ZN(n17865) );
  AOI21HSV4 U20914 ( .A1(n17866), .A2(n17829), .B(n17865), .ZN(n17867) );
  XNOR2HSV4 U20915 ( .A1(n17868), .A2(n17867), .ZN(n17869) );
  NAND2HSV0 U20916 ( .A1(\pe9/aot [15]), .A2(\pe9/bq[13] ), .ZN(n17871) );
  BUFHSV4 U20917 ( .I(\pe9/bq[16] ), .Z(n28044) );
  NAND2HSV0 U20918 ( .A1(\pe9/aot [12]), .A2(n28044), .ZN(n17870) );
  XOR2HSV0 U20919 ( .A1(n17871), .A2(n17870), .Z(n17875) );
  INHSV4 U20920 ( .I(\pe9/bq[15] ), .ZN(n17973) );
  NAND2HSV0 U20921 ( .A1(\pe9/aot [13]), .A2(\pe9/bq[15] ), .ZN(n17873) );
  NAND2HSV0 U20922 ( .A1(\pe9/aot [14]), .A2(\pe9/bq[14] ), .ZN(n17872) );
  XOR2HSV0 U20923 ( .A1(n17873), .A2(n17872), .Z(n17874) );
  NOR2HSV1 U20924 ( .A1(n28016), .A2(n21334), .ZN(n17877) );
  XOR2HSV0 U20925 ( .A1(n17877), .A2(n17876), .Z(n17879) );
  INHSV2 U20926 ( .I(n18167), .ZN(n21760) );
  NAND2HSV2 U20927 ( .A1(n21760), .A2(\pe9/pvq [5]), .ZN(n17878) );
  INHSV2 U20928 ( .I(n17884), .ZN(n17883) );
  INHSV2 U20929 ( .I(\pe9/phq [1]), .ZN(n17882) );
  CLKNAND2HSV3 U20930 ( .A1(n17883), .A2(n17882), .ZN(n17894) );
  CLKNAND2HSV1 U20931 ( .A1(n17894), .A2(n17891), .ZN(n17890) );
  INHSV2 U20932 ( .I(n17888), .ZN(n17886) );
  NAND2HSV2 U20933 ( .A1(\pe9/pvq [1]), .A2(\pe9/ctrq ), .ZN(n17887) );
  INHSV2 U20934 ( .I(n17887), .ZN(n17885) );
  CLKNAND2HSV3 U20935 ( .A1(n17886), .A2(n17885), .ZN(n17893) );
  NAND4HSV4 U20936 ( .A1(n17894), .A2(n17893), .A3(n17892), .A4(n17891), .ZN(
        n17915) );
  NAND2HSV2 U20937 ( .A1(n17916), .A2(n17915), .ZN(n28691) );
  CLKBUFHSV4 U20938 ( .I(n17998), .Z(n18050) );
  CLKNAND2HSV2 U20939 ( .A1(n28691), .A2(n18454), .ZN(n17895) );
  INHSV2 U20940 ( .I(n18050), .ZN(n18613) );
  NAND2HSV4 U20941 ( .A1(n17895), .A2(n17945), .ZN(n18141) );
  INHSV4 U20942 ( .I(n18141), .ZN(n17962) );
  INHSV4 U20943 ( .I(n17962), .ZN(n18286) );
  BUFHSV2 U20944 ( .I(\pe9/got [13]), .Z(n18029) );
  NAND2HSV2 U20945 ( .A1(n18286), .A2(n18029), .ZN(n17919) );
  XNOR2HSV1 U20946 ( .A1(n17920), .A2(n17919), .ZN(n17918) );
  BUFHSV2 U20947 ( .I(\pe9/got [14]), .Z(n18078) );
  CLKNAND2HSV2 U20948 ( .A1(\pe9/pvq [2]), .A2(\pe9/ctrq ), .ZN(n17897) );
  NAND2HSV0 U20949 ( .A1(\pe9/bq[16] ), .A2(\pe9/aot [15]), .ZN(n17898) );
  XNOR2HSV4 U20950 ( .A1(n17899), .A2(n17898), .ZN(n17905) );
  NAND2HSV0 U20951 ( .A1(\pe9/bq[15] ), .A2(\pe9/aot [16]), .ZN(n17901) );
  INHSV1 U20952 ( .I(n17900), .ZN(n17902) );
  CLKNAND2HSV1 U20953 ( .A1(n17902), .A2(n17901), .ZN(n17903) );
  NAND2HSV2 U20954 ( .A1(n17904), .A2(n17903), .ZN(n17906) );
  NAND2HSV2 U20955 ( .A1(n17905), .A2(n17906), .ZN(n17910) );
  INHSV3 U20956 ( .I(n17905), .ZN(n17908) );
  INHSV2 U20957 ( .I(n17906), .ZN(n17907) );
  INHSV1 U20958 ( .I(n17998), .ZN(n18623) );
  INHSV2 U20959 ( .I(\pe9/got [16]), .ZN(n17988) );
  NOR2HSV4 U20960 ( .A1(n18623), .A2(n17988), .ZN(n18558) );
  CLKNAND2HSV1 U20961 ( .A1(n28691), .A2(n18558), .ZN(n17911) );
  INHSV2 U20962 ( .I(n17911), .ZN(n17913) );
  CLKAND2HSV2 U20963 ( .A1(n18628), .A2(\pe9/ti_7t [2]), .Z(n17912) );
  INHSV2 U20964 ( .I(\pe9/got [16]), .ZN(n18001) );
  INHSV2 U20965 ( .I(n18001), .ZN(n28081) );
  AOI21HSV2 U20966 ( .A1(n17946), .A2(n28081), .B(n18462), .ZN(n17917) );
  NAND2HSV2 U20967 ( .A1(n18021), .A2(n18022), .ZN(n28110) );
  CLKNAND2HSV2 U20968 ( .A1(n17918), .A2(n17921), .ZN(n17925) );
  CLKXOR2HSV4 U20969 ( .A1(n17920), .A2(n17919), .Z(n17923) );
  INHSV2 U20970 ( .I(n17921), .ZN(n17922) );
  CLKNAND2HSV2 U20971 ( .A1(n18021), .A2(n18022), .ZN(n18252) );
  INHSV2 U20972 ( .I(n18001), .ZN(n25633) );
  NAND2HSV4 U20973 ( .A1(n18252), .A2(n25633), .ZN(n18076) );
  CLKBUFHSV4 U20974 ( .I(n17998), .Z(n18325) );
  NAND2HSV2 U20975 ( .A1(n18551), .A2(\pe9/ti_7t [3]), .ZN(n18142) );
  INHSV4 U20976 ( .I(n18142), .ZN(n18147) );
  NOR2HSV2 U20977 ( .A1(n18076), .A2(n18147), .ZN(n17948) );
  NAND2HSV2 U20978 ( .A1(\pe9/ctrq ), .A2(\pe9/pvq [3]), .ZN(n17927) );
  INHSV2 U20979 ( .I(n17927), .ZN(n17926) );
  NAND3HSV2 U20980 ( .A1(n17927), .A2(\pe9/aot [15]), .A3(\pe9/bq[15] ), .ZN(
        n17928) );
  CLKNAND2HSV2 U20981 ( .A1(n17928), .A2(n17929), .ZN(n17936) );
  INHSV3 U20982 ( .I(n17936), .ZN(n17934) );
  INHSV2 U20983 ( .I(\pe9/phq [3]), .ZN(n17930) );
  CLKNAND2HSV3 U20984 ( .A1(n17932), .A2(n17931), .ZN(n17935) );
  INHSV2 U20985 ( .I(n17935), .ZN(n17933) );
  CLKNAND2HSV3 U20986 ( .A1(n17934), .A2(n17933), .ZN(n17938) );
  CLKNAND2HSV2 U20987 ( .A1(n17936), .A2(n17935), .ZN(n17937) );
  CLKNAND2HSV4 U20988 ( .A1(n17938), .A2(n17937), .ZN(n17942) );
  INHSV4 U20989 ( .I(n17940), .ZN(n17950) );
  AOI21HSV4 U20990 ( .A1(n17951), .A2(n17950), .B(n18641), .ZN(n17944) );
  XNOR2HSV4 U20991 ( .A1(n17942), .A2(n17941), .ZN(n17954) );
  NAND2HSV2 U20992 ( .A1(n17962), .A2(n17954), .ZN(n17943) );
  CLKNAND2HSV3 U20993 ( .A1(n17944), .A2(n17943), .ZN(n18073) );
  NOR2HSV2 U20994 ( .A1(n17954), .A2(n25638), .ZN(n18072) );
  NOR2HSV2 U20995 ( .A1(n18073), .A2(n18072), .ZN(n17947) );
  INHSV2 U20996 ( .I(n17947), .ZN(n18025) );
  CLKNAND2HSV2 U20997 ( .A1(n17948), .A2(n18025), .ZN(n17949) );
  INHSV2 U20998 ( .I(n17950), .ZN(n18398) );
  CLKNAND2HSV2 U20999 ( .A1(n17949), .A2(n18398), .ZN(n17959) );
  INHSV2 U21000 ( .I(n17950), .ZN(n18214) );
  INHSV2 U21001 ( .I(n18462), .ZN(n18338) );
  INHSV2 U21002 ( .I(n17954), .ZN(n25637) );
  INHSV2 U21003 ( .I(n17952), .ZN(n18077) );
  INHSV3 U21004 ( .I(n25638), .ZN(n17953) );
  CLKNAND2HSV3 U21005 ( .A1(n17954), .A2(n17953), .ZN(n17989) );
  INHSV2 U21006 ( .I(n17989), .ZN(n18075) );
  INHSV2 U21007 ( .I(n18075), .ZN(n17955) );
  AOI21HSV0 U21008 ( .A1(n18252), .A2(n28669), .B(n18147), .ZN(n17956) );
  CLKNAND2HSV1 U21009 ( .A1(n18027), .A2(n17956), .ZN(n17957) );
  INHSV2 U21010 ( .I(n17957), .ZN(n17958) );
  NOR2HSV4 U21011 ( .A1(n17959), .A2(n17958), .ZN(n17961) );
  NOR2HSV2 U21012 ( .A1(n18104), .A2(n18524), .ZN(n18000) );
  NAND2HSV0 U21013 ( .A1(\pe9/bq[14] ), .A2(\pe9/aot [15]), .ZN(n17963) );
  NAND2HSV0 U21014 ( .A1(n17963), .A2(n18302), .ZN(n17967) );
  CLKNHSV0 U21015 ( .I(n17963), .ZN(n17965) );
  CLKNHSV0 U21016 ( .I(n18302), .ZN(n17964) );
  CLKNAND2HSV1 U21017 ( .A1(n17965), .A2(n17964), .ZN(n17966) );
  CLKNAND2HSV2 U21018 ( .A1(n17967), .A2(n17966), .ZN(n17972) );
  CLKAND2HSV2 U21019 ( .A1(\pe9/pvq [4]), .A2(\pe9/phq [4]), .Z(n17970) );
  CLKNAND2HSV2 U21020 ( .A1(n27092), .A2(\pe9/pvq [4]), .ZN(n17969) );
  INHSV2 U21021 ( .I(\pe9/phq [4]), .ZN(n17968) );
  AOI22HSV4 U21022 ( .A1(n27092), .A2(n17970), .B1(n17969), .B2(n17968), .ZN(
        n17971) );
  XNOR2HSV4 U21023 ( .A1(n17972), .A2(n17971), .ZN(n17974) );
  INHSV3 U21024 ( .I(n17974), .ZN(n17977) );
  CLKNAND2HSV3 U21025 ( .A1(n17977), .A2(n17976), .ZN(n17978) );
  INHSV2 U21026 ( .I(n17980), .ZN(n17982) );
  INHSV2 U21027 ( .I(\pe9/got [14]), .ZN(n18552) );
  INHSV2 U21028 ( .I(n18552), .ZN(n18005) );
  CLKNAND2HSV1 U21029 ( .A1(n18141), .A2(n18078), .ZN(n17981) );
  INHSV2 U21030 ( .I(\pe9/got [15]), .ZN(n18647) );
  INHSV2 U21031 ( .I(n18647), .ZN(n23718) );
  INHSV2 U21032 ( .I(n23718), .ZN(n18530) );
  CLKNAND2HSV1 U21033 ( .A1(n17984), .A2(n17983), .ZN(n17987) );
  INHSV3 U21034 ( .I(n17984), .ZN(n17985) );
  INHSV2 U21035 ( .I(n17988), .ZN(n18326) );
  INHSV2 U21036 ( .I(n18326), .ZN(n18629) );
  NOR3HSV2 U21037 ( .A1(n18073), .A2(n18072), .A3(n18629), .ZN(n17996) );
  INHSV2 U21038 ( .I(n17990), .ZN(n17993) );
  NAND3HSV3 U21039 ( .A1(n17993), .A2(n17991), .A3(n17992), .ZN(n17994) );
  INHSV2 U21040 ( .I(n18147), .ZN(n18028) );
  OAI22HSV2 U21041 ( .A1(n17994), .A2(n18252), .B1(n18629), .B2(n18028), .ZN(
        n17995) );
  CLKBUFHSV4 U21042 ( .I(n17998), .Z(n18468) );
  INHSV2 U21043 ( .I(n18468), .ZN(n18551) );
  INHSV2 U21044 ( .I(n18551), .ZN(n18454) );
  CLKNAND2HSV4 U21045 ( .A1(n28961), .A2(n18219), .ZN(n19769) );
  CLKNAND2HSV0 U21046 ( .A1(n18646), .A2(\pe9/ti_7t [4]), .ZN(n17999) );
  NAND2HSV2 U21047 ( .A1(n19769), .A2(n17999), .ZN(n18231) );
  NAND2HSV2 U21048 ( .A1(n18000), .A2(n18231), .ZN(n18185) );
  NAND2HSV2 U21049 ( .A1(n18628), .A2(\pe9/ti_7t [4]), .ZN(n19768) );
  NOR2HSV2 U21050 ( .A1(n18623), .A2(n28669), .ZN(n18529) );
  INHSV2 U21051 ( .I(n18529), .ZN(n18278) );
  NOR2HSV4 U21052 ( .A1(n18002), .A2(n18278), .ZN(n18182) );
  INHSV2 U21053 ( .I(\pe9/ti_7t [5]), .ZN(n18105) );
  NAND2HSV2 U21054 ( .A1(n18105), .A2(n18613), .ZN(n18180) );
  CLKNAND2HSV0 U21055 ( .A1(n18180), .A2(n18398), .ZN(n18003) );
  NAND3HSV4 U21056 ( .A1(n18004), .A2(n18184), .A3(n18185), .ZN(n18041) );
  INHSV3 U21057 ( .I(n18041), .ZN(n18039) );
  INHSV2 U21058 ( .I(n18035), .ZN(n18033) );
  NAND2HSV0 U21059 ( .A1(\pe9/aot [13]), .A2(\pe9/bq[13] ), .ZN(n18007) );
  NAND2HSV0 U21060 ( .A1(\pe9/aot [16]), .A2(\pe9/bq[10] ), .ZN(n18006) );
  XOR2HSV0 U21061 ( .A1(n18007), .A2(n18006), .Z(n18009) );
  INHSV2 U21062 ( .I(\pe9/ctrq ), .ZN(n18416) );
  INHSV2 U21063 ( .I(n18416), .ZN(n27078) );
  NAND2HSV2 U21064 ( .A1(n27078), .A2(\pe9/pvq [7]), .ZN(n18008) );
  NAND2HSV0 U21065 ( .A1(\pe9/aot [11]), .A2(\pe9/bq[15] ), .ZN(n18117) );
  NAND2HSV0 U21066 ( .A1(\pe9/aot [10]), .A2(n28044), .ZN(n18010) );
  XOR2HSV0 U21067 ( .A1(n18117), .A2(n18010), .Z(n18011) );
  NAND2HSV0 U21068 ( .A1(\pe9/aot [12]), .A2(n23822), .ZN(n18013) );
  NAND2HSV0 U21069 ( .A1(\pe9/aot [15]), .A2(\pe9/bq[11] ), .ZN(n18012) );
  XOR2HSV0 U21070 ( .A1(n18013), .A2(n18012), .Z(n18017) );
  BUFHSV2 U21071 ( .I(\pe9/ti_1 ), .Z(n18498) );
  INHSV4 U21072 ( .I(n22116), .ZN(n28227) );
  CLKNAND2HSV0 U21073 ( .A1(n18498), .A2(n28227), .ZN(n18015) );
  NAND2HSV0 U21074 ( .A1(\pe9/aot [14]), .A2(\pe9/bq[12] ), .ZN(n18014) );
  XOR2HSV0 U21075 ( .A1(n18015), .A2(n18014), .Z(n18016) );
  XOR2HSV0 U21076 ( .A1(n18017), .A2(n18016), .Z(n18018) );
  INHSV2 U21077 ( .I(\pe9/got [11]), .ZN(n28085) );
  NOR2HSV2 U21078 ( .A1(n18481), .A2(n28085), .ZN(n18019) );
  XNOR2HSV4 U21079 ( .A1(n18020), .A2(n18019), .ZN(n18024) );
  NAND2HSV0 U21080 ( .A1(n28134), .A2(n28470), .ZN(n18023) );
  XNOR2HSV4 U21081 ( .A1(n18024), .A2(n18023), .ZN(n18031) );
  INHSV4 U21082 ( .I(n18076), .ZN(n25639) );
  INHSV1 U21083 ( .I(n18025), .ZN(n18026) );
  NAND2HSV2 U21084 ( .A1(n25639), .A2(n18026), .ZN(n18144) );
  CLKNAND2HSV1 U21085 ( .A1(n18107), .A2(n18029), .ZN(n18030) );
  INHSV2 U21086 ( .I(n18034), .ZN(n18032) );
  CLKNAND2HSV3 U21087 ( .A1(n18033), .A2(n18032), .ZN(n18037) );
  NAND2HSV4 U21088 ( .A1(n18037), .A2(n18036), .ZN(n18040) );
  INHSV3 U21089 ( .I(n18040), .ZN(n18038) );
  CLKNAND2HSV4 U21090 ( .A1(n18039), .A2(n18038), .ZN(n18192) );
  CLKNAND2HSV3 U21091 ( .A1(n18040), .A2(n18041), .ZN(n18191) );
  CLKNAND2HSV4 U21092 ( .A1(n18192), .A2(n18191), .ZN(n18223) );
  NAND2HSV2 U21093 ( .A1(n18180), .A2(n28081), .ZN(n23463) );
  NOR2HSV1 U21094 ( .A1(n23463), .A2(n18086), .ZN(n18045) );
  NAND2HSV2 U21095 ( .A1(n18042), .A2(n18045), .ZN(n18049) );
  INHSV2 U21096 ( .I(\pe9/ti_7t [4]), .ZN(n18051) );
  OAI21HSV4 U21097 ( .A1(n18051), .A2(n18611), .B(n19769), .ZN(n28949) );
  INHSV2 U21098 ( .I(n28949), .ZN(n18048) );
  NAND3HSV2 U21099 ( .A1(n18044), .A2(n18043), .A3(n18543), .ZN(n18087) );
  CLKNAND2HSV1 U21100 ( .A1(n18087), .A2(n18045), .ZN(n18046) );
  BUFHSV2 U21101 ( .I(n18050), .Z(n18611) );
  AOI21HSV2 U21102 ( .A1(n18051), .A2(n18545), .B(n18530), .ZN(n18052) );
  INHSV2 U21103 ( .I(\pe9/pvq [6]), .ZN(n18053) );
  NOR2HSV4 U21104 ( .A1(n18167), .A2(n18053), .ZN(n18055) );
  NAND2HSV0 U21105 ( .A1(\pe9/aot [15]), .A2(\pe9/bq[12] ), .ZN(n28039) );
  INHSV2 U21106 ( .I(n28039), .ZN(n18054) );
  XOR3HSV2 U21107 ( .A1(\pe9/phq [6]), .A2(n18055), .A3(n18054), .Z(n18059) );
  NAND2HSV0 U21108 ( .A1(n21761), .A2(\pe9/aot [12]), .ZN(n18057) );
  NAND2HSV0 U21109 ( .A1(\pe9/ti_1 ), .A2(\pe9/got [11]), .ZN(n18056) );
  XOR2HSV0 U21110 ( .A1(n18057), .A2(n18056), .Z(n18058) );
  XNOR2HSV4 U21111 ( .A1(n18059), .A2(n18058), .ZN(n18067) );
  NAND2HSV0 U21112 ( .A1(\pe9/aot [11]), .A2(\pe9/bq[16] ), .ZN(n18061) );
  NAND2HSV0 U21113 ( .A1(\pe9/aot [16]), .A2(\pe9/bq[11] ), .ZN(n18060) );
  XOR2HSV0 U21114 ( .A1(n18061), .A2(n18060), .Z(n18065) );
  NAND2HSV0 U21115 ( .A1(\pe9/aot [14]), .A2(\pe9/bq[13] ), .ZN(n18063) );
  NAND2HSV0 U21116 ( .A1(\pe9/aot [13]), .A2(\pe9/bq[14] ), .ZN(n18062) );
  XOR2HSV0 U21117 ( .A1(n18063), .A2(n18062), .Z(n18064) );
  XOR2HSV2 U21118 ( .A1(n18065), .A2(n18064), .Z(n18066) );
  XNOR2HSV4 U21119 ( .A1(n18067), .A2(n18066), .ZN(n18069) );
  NAND2HSV2 U21120 ( .A1(n18286), .A2(\pe9/got [12]), .ZN(n18068) );
  XNOR2HSV4 U21121 ( .A1(n18069), .A2(n18068), .ZN(n18071) );
  NAND2HSV2 U21122 ( .A1(n28470), .A2(\pe9/got [13]), .ZN(n18070) );
  XNOR2HSV4 U21123 ( .A1(n18071), .A2(n18070), .ZN(n18083) );
  NOR3HSV2 U21124 ( .A1(n18072), .A2(n18552), .A3(n18073), .ZN(n18074) );
  NAND2HSV2 U21125 ( .A1(n25639), .A2(n18074), .ZN(n18081) );
  CLKNAND2HSV0 U21126 ( .A1(n18147), .A2(n18078), .ZN(n18079) );
  NAND3HSV2 U21127 ( .A1(n18081), .A2(n18080), .A3(n18079), .ZN(n18082) );
  XOR2HSV4 U21128 ( .A1(n18083), .A2(n18082), .Z(n18084) );
  INHSV1 U21129 ( .I(n18087), .ZN(n18088) );
  NAND2HSV2 U21130 ( .A1(n18088), .A2(n22375), .ZN(n23464) );
  NOR2HSV2 U21131 ( .A1(n23463), .A2(n18623), .ZN(n18089) );
  CLKNAND2HSV3 U21132 ( .A1(n23464), .A2(n18089), .ZN(n18093) );
  NOR2HSV2 U21133 ( .A1(n18093), .A2(n23466), .ZN(n18091) );
  INHSV2 U21134 ( .I(n18090), .ZN(n23465) );
  INHSV2 U21135 ( .I(n18092), .ZN(n18103) );
  OAI21HSV4 U21136 ( .A1(n18097), .A2(n18096), .B(n18095), .ZN(n18222) );
  NAND2HSV2 U21137 ( .A1(n18310), .A2(n18558), .ZN(n18101) );
  CLKNAND2HSV1 U21138 ( .A1(n18225), .A2(n18398), .ZN(n18098) );
  OAI21HSV4 U21139 ( .A1(n18101), .A2(n18100), .B(n18099), .ZN(n18102) );
  NOR2HSV2 U21140 ( .A1(n18219), .A2(n18105), .ZN(n18106) );
  NOR2HSV4 U21141 ( .A1(n29001), .A2(n18106), .ZN(n18229) );
  INHSV2 U21142 ( .I(n18106), .ZN(n18376) );
  CLKNAND2HSV0 U21143 ( .A1(n18376), .A2(n18545), .ZN(n18227) );
  BUFHSV4 U21144 ( .I(n18107), .Z(n18400) );
  NAND2HSV2 U21145 ( .A1(n18400), .A2(\pe9/got [11]), .ZN(n18134) );
  NAND2HSV0 U21146 ( .A1(n18286), .A2(n14073), .ZN(n18132) );
  NAND2HSV0 U21147 ( .A1(n28227), .A2(n28470), .ZN(n18131) );
  CLKNAND2HSV0 U21148 ( .A1(\pe9/got [8]), .A2(n18498), .ZN(n18109) );
  NAND2HSV0 U21149 ( .A1(\pe9/aot [16]), .A2(\pe9/bq[8] ), .ZN(n18108) );
  XOR2HSV0 U21150 ( .A1(n18109), .A2(n18108), .Z(n18113) );
  NAND2HSV0 U21151 ( .A1(\pe9/aot [10]), .A2(\pe9/bq[14] ), .ZN(n18111) );
  NAND2HSV0 U21152 ( .A1(\pe9/aot [15]), .A2(\pe9/bq[9] ), .ZN(n18110) );
  XOR2HSV0 U21153 ( .A1(n18111), .A2(n18110), .Z(n18112) );
  XOR2HSV0 U21154 ( .A1(n18113), .A2(n18112), .Z(n18121) );
  CLKNAND2HSV1 U21155 ( .A1(n27078), .A2(\pe9/pvq [9]), .ZN(n18114) );
  XNOR2HSV1 U21156 ( .A1(n18114), .A2(\pe9/phq [9]), .ZN(n18119) );
  CLKNAND2HSV0 U21157 ( .A1(\pe9/aot [9]), .A2(\pe9/bq[13] ), .ZN(n18301) );
  CLKNHSV0 U21158 ( .I(\pe9/aot [9]), .ZN(n18407) );
  CLKNHSV1 U21159 ( .I(n21761), .ZN(n28026) );
  NAND2HSV0 U21160 ( .A1(\pe9/aot [11]), .A2(\pe9/bq[13] ), .ZN(n18115) );
  OAI21HSV2 U21161 ( .A1(n18407), .A2(n28026), .B(n18115), .ZN(n18116) );
  OAI21HSV0 U21162 ( .A1(n18301), .A2(n18117), .B(n18116), .ZN(n18118) );
  XOR2HSV0 U21163 ( .A1(n18119), .A2(n18118), .Z(n18120) );
  XNOR2HSV1 U21164 ( .A1(n18121), .A2(n18120), .ZN(n18129) );
  NAND2HSV0 U21165 ( .A1(\pe9/aot [12]), .A2(\pe9/bq[12] ), .ZN(n18123) );
  NAND2HSV0 U21166 ( .A1(\pe9/aot [14]), .A2(\pe9/bq[10] ), .ZN(n18122) );
  XOR2HSV0 U21167 ( .A1(n18123), .A2(n18122), .Z(n18127) );
  NAND2HSV0 U21168 ( .A1(\pe9/bq[11] ), .A2(\pe9/aot [13]), .ZN(n18125) );
  NAND2HSV0 U21169 ( .A1(\pe9/aot [8]), .A2(n28044), .ZN(n18124) );
  XOR2HSV0 U21170 ( .A1(n18125), .A2(n18124), .Z(n18126) );
  XOR2HSV0 U21171 ( .A1(n18127), .A2(n18126), .Z(n18128) );
  XNOR2HSV1 U21172 ( .A1(n18129), .A2(n18128), .ZN(n18130) );
  XOR3HSV1 U21173 ( .A1(n18132), .A2(n18131), .A3(n18130), .Z(n18133) );
  XNOR2HSV4 U21174 ( .A1(n18138), .A2(n18137), .ZN(n18140) );
  BUFHSV2 U21175 ( .I(\pe9/got [14]), .Z(n28928) );
  INHSV2 U21176 ( .I(n28928), .ZN(n18617) );
  INHSV2 U21177 ( .I(n18617), .ZN(n18464) );
  BUFHSV2 U21178 ( .I(\pe9/got [13]), .Z(n28137) );
  CLKNHSV0 U21179 ( .I(n18141), .ZN(n18481) );
  NOR2HSV2 U21180 ( .A1(n18481), .A2(n22116), .ZN(n18146) );
  NAND2HSV0 U21181 ( .A1(n18146), .A2(n18142), .ZN(n18154) );
  CLKNAND2HSV1 U21182 ( .A1(n18144), .A2(n18143), .ZN(n18153) );
  NOR2HSV0 U21183 ( .A1(n18146), .A2(n28016), .ZN(n18151) );
  CLKNHSV0 U21184 ( .I(n18146), .ZN(n18145) );
  NOR2HSV0 U21185 ( .A1(n18145), .A2(n28016), .ZN(n18149) );
  AOI21HSV0 U21186 ( .A1(n28134), .A2(n18147), .B(n18146), .ZN(n18148) );
  NOR2HSV1 U21187 ( .A1(n18149), .A2(n18148), .ZN(n18150) );
  NAND2HSV1 U21188 ( .A1(\pe9/aot [11]), .A2(n23822), .ZN(n18156) );
  NAND2HSV0 U21189 ( .A1(\pe9/aot [14]), .A2(\pe9/bq[11] ), .ZN(n18155) );
  XOR2HSV0 U21190 ( .A1(n18156), .A2(n18155), .Z(n18160) );
  NAND2HSV0 U21191 ( .A1(\pe9/aot [15]), .A2(\pe9/bq[10] ), .ZN(n18158) );
  NAND2HSV0 U21192 ( .A1(n21761), .A2(\pe9/aot [10]), .ZN(n18157) );
  XOR2HSV0 U21193 ( .A1(n18158), .A2(n18157), .Z(n18159) );
  XOR2HSV0 U21194 ( .A1(n18160), .A2(n18159), .Z(n18175) );
  BUFHSV2 U21195 ( .I(\pe9/ti_1 ), .Z(n28019) );
  NAND2HSV0 U21196 ( .A1(n14073), .A2(n28019), .ZN(n18162) );
  NAND2HSV0 U21197 ( .A1(\pe9/aot [16]), .A2(\pe9/bq[9] ), .ZN(n18161) );
  XOR2HSV0 U21198 ( .A1(n18162), .A2(n18161), .Z(n18166) );
  NAND2HSV0 U21199 ( .A1(\pe9/bq[16] ), .A2(\pe9/aot [9]), .ZN(n18164) );
  NAND2HSV0 U21200 ( .A1(\pe9/aot [12]), .A2(\pe9/bq[13] ), .ZN(n18163) );
  XOR2HSV0 U21201 ( .A1(n18164), .A2(n18163), .Z(n18165) );
  XOR2HSV0 U21202 ( .A1(n18166), .A2(n18165), .Z(n18172) );
  INHSV2 U21203 ( .I(n18167), .ZN(n23530) );
  NAND2HSV2 U21204 ( .A1(n23530), .A2(\pe9/pvq [8]), .ZN(n18168) );
  XNOR2HSV1 U21205 ( .A1(n18168), .A2(\pe9/phq [8]), .ZN(n18170) );
  CLKNHSV0 U21206 ( .I(\pe9/aot [13]), .ZN(n18169) );
  INHSV2 U21207 ( .I(\pe9/bq[12] ), .ZN(n27101) );
  NOR2HSV2 U21208 ( .A1(n18169), .A2(n27101), .ZN(n18568) );
  XNOR2HSV1 U21209 ( .A1(n18170), .A2(n18568), .ZN(n18171) );
  XNOR2HSV2 U21210 ( .A1(n18172), .A2(n18171), .ZN(n18174) );
  NAND2HSV0 U21211 ( .A1(n28110), .A2(\pe9/got [11]), .ZN(n18173) );
  XOR3HSV2 U21212 ( .A1(n18175), .A2(n18174), .A3(n18173), .Z(n18176) );
  XNOR2HSV4 U21213 ( .A1(n18177), .A2(n18176), .ZN(n18178) );
  XNOR2HSV4 U21214 ( .A1(n18179), .A2(n18178), .ZN(n18187) );
  CLKNAND2HSV1 U21215 ( .A1(n18180), .A2(n18464), .ZN(n18181) );
  NOR2HSV3 U21216 ( .A1(n18182), .A2(n18181), .ZN(n18183) );
  XNOR2HSV4 U21217 ( .A1(n18187), .A2(n18186), .ZN(n18199) );
  NAND2HSV2 U21218 ( .A1(n18199), .A2(n18530), .ZN(n18189) );
  CLKAND2HSV2 U21219 ( .A1(n18225), .A2(n25633), .Z(n18212) );
  AND2HSV2 U21220 ( .A1(n18212), .A2(n18543), .Z(n18188) );
  NAND3HSV3 U21221 ( .A1(n18206), .A2(n18189), .A3(n18188), .ZN(n18190) );
  BUFHSV8 U21222 ( .I(n18199), .Z(n25660) );
  CLKNAND2HSV2 U21223 ( .A1(n18192), .A2(n18191), .ZN(n18193) );
  CLKXOR2HSV4 U21224 ( .A1(n18193), .A2(n18222), .Z(n18211) );
  OAI21HSV2 U21225 ( .A1(n18199), .A2(n18214), .B(n18219), .ZN(n18198) );
  INHSV2 U21226 ( .I(n18198), .ZN(n18213) );
  CLKNHSV0 U21227 ( .I(n18199), .ZN(n18201) );
  NAND2HSV2 U21228 ( .A1(n18201), .A2(n18200), .ZN(n18215) );
  CLKAND2HSV4 U21229 ( .A1(n18213), .A2(n18215), .Z(n18203) );
  NAND3HSV2 U21230 ( .A1(n18210), .A2(n18216), .A3(n18203), .ZN(n18202) );
  NAND2HSV2 U21231 ( .A1(n18276), .A2(n25633), .ZN(n18205) );
  NOR2HSV2 U21232 ( .A1(n18208), .A2(n18207), .ZN(n18209) );
  CLKAND2HSV2 U21233 ( .A1(n18209), .A2(n18214), .Z(n18221) );
  CLKAND2HSV1 U21234 ( .A1(n18215), .A2(n18214), .Z(n18217) );
  NAND2HSV0 U21235 ( .A1(n18274), .A2(\pe9/got [15]), .ZN(n18220) );
  CLKAND2HSV2 U21236 ( .A1(n18225), .A2(n28928), .Z(n18226) );
  CLKNAND2HSV0 U21237 ( .A1(n18227), .A2(n28134), .ZN(n18228) );
  NOR2HSV2 U21238 ( .A1(n18229), .A2(n18228), .ZN(n18230) );
  CLKNAND2HSV1 U21239 ( .A1(n28227), .A2(n18400), .ZN(n18258) );
  NAND2HSV0 U21240 ( .A1(n18286), .A2(\pe9/got [8]), .ZN(n18256) );
  CLKNAND2HSV0 U21241 ( .A1(\pe9/got [7]), .A2(n28019), .ZN(n18233) );
  XOR2HSV0 U21242 ( .A1(n18233), .A2(n18232), .Z(n18237) );
  NAND2HSV0 U21243 ( .A1(\pe9/aot [8]), .A2(\pe9/bq[15] ), .ZN(n18235) );
  NAND2HSV0 U21244 ( .A1(\pe9/aot [9]), .A2(n23822), .ZN(n18234) );
  XOR2HSV0 U21245 ( .A1(n18235), .A2(n18234), .Z(n18236) );
  XOR2HSV0 U21246 ( .A1(n18237), .A2(n18236), .Z(n18245) );
  NAND2HSV0 U21247 ( .A1(\pe9/aot [12]), .A2(\pe9/bq[11] ), .ZN(n18239) );
  NAND2HSV0 U21248 ( .A1(\pe9/aot [10]), .A2(\pe9/bq[13] ), .ZN(n18238) );
  XOR2HSV0 U21249 ( .A1(n18239), .A2(n18238), .Z(n18243) );
  NAND2HSV0 U21250 ( .A1(\pe9/bq[10] ), .A2(\pe9/aot [13]), .ZN(n18241) );
  NAND2HSV0 U21251 ( .A1(\pe9/aot [11]), .A2(\pe9/bq[12] ), .ZN(n18240) );
  XOR2HSV0 U21252 ( .A1(n18241), .A2(n18240), .Z(n18242) );
  XOR2HSV0 U21253 ( .A1(n18243), .A2(n18242), .Z(n18244) );
  XOR2HSV0 U21254 ( .A1(n18245), .A2(n18244), .Z(n18255) );
  NAND2HSV0 U21255 ( .A1(\pe9/aot [14]), .A2(\pe9/bq[9] ), .ZN(n18251) );
  NAND2HSV2 U21256 ( .A1(n27093), .A2(\pe9/pvq [10]), .ZN(n18246) );
  XNOR2HSV1 U21257 ( .A1(n18246), .A2(\pe9/phq [10]), .ZN(n18250) );
  NAND2HSV0 U21258 ( .A1(\pe9/bq[16] ), .A2(\pe9/aot [7]), .ZN(n18248) );
  NAND2HSV0 U21259 ( .A1(\pe9/aot [15]), .A2(\pe9/bq[8] ), .ZN(n18247) );
  XOR2HSV0 U21260 ( .A1(n18248), .A2(n18247), .Z(n18249) );
  XOR3HSV2 U21261 ( .A1(n18251), .A2(n18250), .A3(n18249), .Z(n18254) );
  NAND2HSV0 U21262 ( .A1(\pe9/got [9]), .A2(n18252), .ZN(n18253) );
  XOR4HSV1 U21263 ( .A1(n18256), .A2(n18255), .A3(n18254), .A4(n18253), .Z(
        n18257) );
  XOR2HSV0 U21264 ( .A1(n18258), .A2(n18257), .Z(n18259) );
  XNOR2HSV1 U21265 ( .A1(n18260), .A2(n18259), .ZN(n18261) );
  INHSV2 U21266 ( .I(n18262), .ZN(n18263) );
  CLKNAND2HSV3 U21267 ( .A1(n18264), .A2(n18263), .ZN(n18265) );
  CLKNAND2HSV2 U21268 ( .A1(n18270), .A2(n18269), .ZN(n18271) );
  NAND2HSV2 U21269 ( .A1(n18613), .A2(\pe9/ti_7t [10]), .ZN(n18273) );
  AND2HSV2 U21270 ( .A1(n18276), .A2(\pe9/got [15]), .Z(n18277) );
  OAI21HSV1 U21271 ( .A1(n18280), .A2(n18278), .B(n18277), .ZN(n18279) );
  AOI31HSV2 U21272 ( .A1(n18439), .A2(n18336), .A3(n23244), .B(n18279), .ZN(
        n18284) );
  NAND2HSV0 U21273 ( .A1(n18558), .A2(n18280), .ZN(n18281) );
  NOR2HSV1 U21274 ( .A1(n18281), .A2(n18439), .ZN(n18282) );
  INHSV1 U21275 ( .I(n18282), .ZN(n18283) );
  NOR2HSV2 U21276 ( .A1(n18439), .A2(n18617), .ZN(n18321) );
  INHSV2 U21277 ( .I(n18383), .ZN(n18285) );
  NAND2HSV0 U21278 ( .A1(n28227), .A2(n28949), .ZN(n18307) );
  BUFHSV2 U21279 ( .I(n18400), .Z(n28804) );
  BUFHSV6 U21280 ( .I(n18286), .Z(n28688) );
  NAND2HSV0 U21281 ( .A1(\pe9/bq[9] ), .A2(\pe9/aot [13]), .ZN(n18288) );
  INHSV2 U21282 ( .I(\pe9/got [6]), .ZN(n28188) );
  NAND2HSV0 U21283 ( .A1(n18498), .A2(\pe9/got [6]), .ZN(n18287) );
  XOR2HSV0 U21284 ( .A1(n18288), .A2(n18287), .Z(n18292) );
  NAND2HSV0 U21285 ( .A1(\pe9/aot [14]), .A2(\pe9/bq[8] ), .ZN(n18290) );
  NAND2HSV0 U21286 ( .A1(\pe9/aot [12]), .A2(\pe9/bq[10] ), .ZN(n18289) );
  XOR2HSV0 U21287 ( .A1(n18290), .A2(n18289), .Z(n18291) );
  XOR2HSV0 U21288 ( .A1(n18292), .A2(n18291), .Z(n18300) );
  NAND2HSV0 U21289 ( .A1(\pe9/aot [6]), .A2(n28044), .ZN(n18294) );
  NAND2HSV0 U21290 ( .A1(\pe9/aot [15]), .A2(\pe9/bq[7] ), .ZN(n18293) );
  XOR2HSV0 U21291 ( .A1(n18294), .A2(n18293), .Z(n18298) );
  NAND2HSV0 U21292 ( .A1(\pe9/aot [11]), .A2(\pe9/bq[11] ), .ZN(n18296) );
  NAND2HSV0 U21293 ( .A1(n21761), .A2(\pe9/aot [7]), .ZN(n18295) );
  XOR2HSV0 U21294 ( .A1(n18296), .A2(n18295), .Z(n18297) );
  XOR2HSV0 U21295 ( .A1(n18298), .A2(n18297), .Z(n18299) );
  CLKNAND2HSV0 U21296 ( .A1(\pe9/aot [9]), .A2(\pe9/bq[6] ), .ZN(n22377) );
  INHSV2 U21297 ( .I(\pe9/bq[6] ), .ZN(n28199) );
  NAND2HSV0 U21298 ( .A1(\pe9/aot [8]), .A2(\pe9/bq[14] ), .ZN(n18421) );
  NAND2HSV0 U21299 ( .A1(\pe9/aot [10]), .A2(\pe9/bq[12] ), .ZN(n18303) );
  XOR2HSV0 U21300 ( .A1(n18421), .A2(n18303), .Z(n18304) );
  CLKNAND2HSV2 U21301 ( .A1(n29001), .A2(n18611), .ZN(n18377) );
  NAND2HSV2 U21302 ( .A1(n18377), .A2(n18376), .ZN(n28638) );
  INHSV2 U21303 ( .I(\pe9/got [11]), .ZN(n18308) );
  NAND2HSV2 U21304 ( .A1(n28638), .A2(n28423), .ZN(n18309) );
  BUFHSV8 U21305 ( .I(n18310), .Z(n28689) );
  NAND2HSV2 U21306 ( .A1(n18650), .A2(\pe9/ti_7t [7]), .ZN(n18339) );
  CLKNHSV0 U21307 ( .I(n18339), .ZN(n18312) );
  AOI21HSV2 U21308 ( .A1(n18194), .A2(n18339), .B(n18469), .ZN(n18311) );
  OA21HSV4 U21309 ( .A1(n29000), .A2(n18312), .B(n18311), .Z(n18314) );
  CLKNAND2HSV1 U21310 ( .A1(n18313), .A2(n18314), .ZN(n18318) );
  CLKNHSV1 U21311 ( .I(n18313), .ZN(n18316) );
  INHSV2 U21312 ( .I(n18314), .ZN(n18315) );
  CLKNAND2HSV1 U21313 ( .A1(n18316), .A2(n18315), .ZN(n18317) );
  NAND2HSV2 U21314 ( .A1(n18318), .A2(n18317), .ZN(n18319) );
  INHSV2 U21315 ( .I(n18322), .ZN(n18324) );
  INHSV4 U21316 ( .I(n18528), .ZN(n23449) );
  NAND2HSV0 U21317 ( .A1(n18330), .A2(n18326), .ZN(n18327) );
  NOR2HSV2 U21318 ( .A1(n23449), .A2(n18327), .ZN(n18329) );
  CLKAND2HSV1 U21319 ( .A1(n18462), .A2(\pe9/ti_7t [11]), .Z(n18328) );
  AOI21HSV2 U21320 ( .A1(n28795), .A2(n18329), .B(n18328), .ZN(n18333) );
  CLKAND2HSV2 U21321 ( .A1(n23449), .A2(n18330), .Z(n18331) );
  CLKNAND2HSV3 U21322 ( .A1(n18331), .A2(n23447), .ZN(n18332) );
  NAND2HSV4 U21323 ( .A1(n18333), .A2(n18332), .ZN(n19766) );
  INHSV6 U21324 ( .I(n19766), .ZN(n28146) );
  NOR2HSV4 U21325 ( .A1(n28146), .A2(n18469), .ZN(n18395) );
  INHSV2 U21326 ( .I(n18395), .ZN(n18393) );
  NAND2HSV2 U21327 ( .A1(\pe9/ti_7t [9]), .A2(n18194), .ZN(n18470) );
  NAND2HSV2 U21328 ( .A1(n19767), .A2(n28423), .ZN(n18387) );
  BUFHSV3 U21329 ( .I(n28952), .Z(n28264) );
  NAND2HSV0 U21330 ( .A1(n28264), .A2(n14073), .ZN(n18382) );
  NAND2HSV0 U21331 ( .A1(\pe9/aot [11]), .A2(\pe9/bq[7] ), .ZN(n22332) );
  NAND2HSV0 U21332 ( .A1(\pe9/aot [9]), .A2(\pe9/bq[9] ), .ZN(n28270) );
  XOR2HSV0 U21333 ( .A1(n22332), .A2(n28270), .Z(n18352) );
  NAND2HSV0 U21334 ( .A1(n27093), .A2(\pe9/pvq [15]), .ZN(n18341) );
  XOR2HSV0 U21335 ( .A1(n18341), .A2(\pe9/phq [15]), .Z(n18344) );
  CLKNAND2HSV0 U21336 ( .A1(\pe9/bq[2] ), .A2(\pe9/aot [4]), .ZN(n28308) );
  INHSV2 U21337 ( .I(\pe9/bq[2] ), .ZN(n28397) );
  CLKNHSV0 U21338 ( .I(\pe9/aot [4]), .ZN(n28194) );
  INHSV2 U21339 ( .I(\pe9/bq[14] ), .ZN(n22378) );
  OAI22HSV0 U21340 ( .A1(n23546), .A2(n28397), .B1(n28194), .B2(n22378), .ZN(
        n18342) );
  OAI21HSV1 U21341 ( .A1(n28308), .A2(n17939), .B(n18342), .ZN(n18343) );
  XNOR2HSV1 U21342 ( .A1(n18344), .A2(n18343), .ZN(n18351) );
  CLKNHSV0 U21343 ( .I(\pe9/aot [7]), .ZN(n18566) );
  CLKNHSV0 U21344 ( .I(\pe9/bq[11] ), .ZN(n23531) );
  NOR2HSV0 U21345 ( .A1(n18566), .A2(n23531), .ZN(n18346) );
  NAND2HSV0 U21346 ( .A1(\pe9/aot [6]), .A2(\pe9/bq[12] ), .ZN(n18345) );
  XOR2HSV0 U21347 ( .A1(n18346), .A2(n18345), .Z(n18349) );
  CLKNAND2HSV0 U21348 ( .A1(\pe9/bq[5] ), .A2(\pe9/aot [13]), .ZN(n22382) );
  NAND2HSV0 U21349 ( .A1(\pe9/aot [10]), .A2(\pe9/bq[8] ), .ZN(n18347) );
  XOR2HSV0 U21350 ( .A1(n22382), .A2(n18347), .Z(n18348) );
  XOR2HSV0 U21351 ( .A1(n18349), .A2(n18348), .Z(n18350) );
  XOR3HSV2 U21352 ( .A1(n18352), .A2(n18351), .A3(n18350), .Z(n18371) );
  NAND2HSV0 U21353 ( .A1(n28389), .A2(n11863), .ZN(n18370) );
  NAND2HSV0 U21354 ( .A1(n21761), .A2(\pe9/aot [3]), .ZN(n18354) );
  NAND2HSV0 U21355 ( .A1(n18498), .A2(n28654), .ZN(n18353) );
  XOR2HSV0 U21356 ( .A1(n18354), .A2(n18353), .Z(n18358) );
  NAND2HSV0 U21357 ( .A1(\pe9/aot [5]), .A2(\pe9/bq[13] ), .ZN(n18356) );
  NAND2HSV0 U21358 ( .A1(\pe9/aot [8]), .A2(\pe9/bq[10] ), .ZN(n18355) );
  XOR2HSV0 U21359 ( .A1(n18356), .A2(n18355), .Z(n18357) );
  XOR2HSV0 U21360 ( .A1(n18358), .A2(n18357), .Z(n18366) );
  NAND2HSV0 U21361 ( .A1(\pe9/aot [2]), .A2(n28044), .ZN(n18360) );
  NAND2HSV0 U21362 ( .A1(\pe9/aot [14]), .A2(\pe9/bq[4] ), .ZN(n18359) );
  XOR2HSV0 U21363 ( .A1(n18360), .A2(n18359), .Z(n18364) );
  NAND2HSV0 U21364 ( .A1(\pe9/aot [15]), .A2(\pe9/bq[3] ), .ZN(n18362) );
  NAND2HSV0 U21365 ( .A1(\pe9/aot [12]), .A2(\pe9/bq[6] ), .ZN(n18361) );
  XOR2HSV0 U21366 ( .A1(n18362), .A2(n18361), .Z(n18363) );
  XOR2HSV0 U21367 ( .A1(n18364), .A2(n18363), .Z(n18365) );
  XOR2HSV0 U21368 ( .A1(n18366), .A2(n18365), .Z(n18368) );
  BUFHSV2 U21369 ( .I(\pe9/got [3]), .Z(n28405) );
  NAND2HSV0 U21370 ( .A1(n28688), .A2(n28405), .ZN(n18367) );
  XNOR2HSV1 U21371 ( .A1(n18368), .A2(n18367), .ZN(n18369) );
  XOR3HSV2 U21372 ( .A1(n18371), .A2(n18370), .A3(n18369), .Z(n18373) );
  BUFHSV4 U21373 ( .I(\pe9/got [5]), .Z(n28643) );
  NAND2HSV0 U21374 ( .A1(n28643), .A2(n28804), .ZN(n18372) );
  XOR2HSV0 U21375 ( .A1(n18373), .A2(n18372), .Z(n18375) );
  NAND2HSV0 U21376 ( .A1(n28949), .A2(\pe9/got [6]), .ZN(n18374) );
  XOR2HSV0 U21377 ( .A1(n18375), .A2(n18374), .Z(n18380) );
  NAND2HSV0 U21378 ( .A1(n28689), .A2(\pe9/got [8]), .ZN(n18379) );
  CLKNAND2HSV2 U21379 ( .A1(n18377), .A2(n18376), .ZN(n28166) );
  NAND2HSV0 U21380 ( .A1(n28166), .A2(\pe9/got [7]), .ZN(n18378) );
  XOR3HSV1 U21381 ( .A1(n18380), .A2(n18379), .A3(n18378), .Z(n18381) );
  XNOR2HSV1 U21382 ( .A1(n18382), .A2(n18381), .ZN(n18385) );
  BUFHSV8 U21383 ( .I(n18439), .Z(n18604) );
  OR2HSV1 U21384 ( .A1(n18604), .A2(n22116), .Z(n18384) );
  XNOR2HSV4 U21385 ( .A1(n18385), .A2(n18384), .ZN(n18386) );
  CLKXOR2HSV4 U21386 ( .A1(n18387), .A2(n18386), .Z(n18389) );
  NOR2HSV2 U21387 ( .A1(n18389), .A2(n28016), .ZN(n18388) );
  INHSV4 U21388 ( .I(n18564), .ZN(n22373) );
  CLKNAND2HSV1 U21389 ( .A1(n18388), .A2(n28231), .ZN(n18391) );
  NAND2HSV2 U21390 ( .A1(n18391), .A2(n18390), .ZN(n18394) );
  INHSV2 U21391 ( .I(n18394), .ZN(n18392) );
  NAND2HSV2 U21392 ( .A1(n18395), .A2(n18394), .ZN(n18396) );
  CLKNAND2HSV1 U21393 ( .A1(n18399), .A2(\pe9/got [9]), .ZN(n18433) );
  NAND2HSV0 U21394 ( .A1(n18400), .A2(\pe9/got [8]), .ZN(n18431) );
  CLKNAND2HSV1 U21395 ( .A1(n28688), .A2(\pe9/got [6]), .ZN(n18429) );
  NAND2HSV0 U21396 ( .A1(\pe9/got [7]), .A2(n28470), .ZN(n18428) );
  NAND2HSV0 U21397 ( .A1(\pe9/aot [11]), .A2(\pe9/bq[10] ), .ZN(n18402) );
  NAND2HSV0 U21398 ( .A1(\pe9/aot [10]), .A2(\pe9/bq[11] ), .ZN(n18401) );
  XOR2HSV0 U21399 ( .A1(n18402), .A2(n18401), .Z(n18406) );
  NAND2HSV0 U21400 ( .A1(\pe9/aot [12]), .A2(\pe9/bq[9] ), .ZN(n18404) );
  NAND2HSV0 U21401 ( .A1(\pe9/aot [14]), .A2(\pe9/bq[7] ), .ZN(n18403) );
  XOR2HSV0 U21402 ( .A1(n18404), .A2(n18403), .Z(n18405) );
  XOR2HSV0 U21403 ( .A1(n18406), .A2(n18405), .Z(n18413) );
  CLKNHSV0 U21404 ( .I(\pe9/aot [6]), .ZN(n22330) );
  NAND2HSV0 U21405 ( .A1(\pe9/aot [6]), .A2(\pe9/bq[15] ), .ZN(n18409) );
  NAND2HSV0 U21406 ( .A1(\pe9/bq[8] ), .A2(\pe9/aot [13]), .ZN(n18408) );
  XOR2HSV0 U21407 ( .A1(n18409), .A2(n18408), .Z(n18410) );
  XOR2HSV0 U21408 ( .A1(n18411), .A2(n18410), .Z(n18412) );
  XOR2HSV0 U21409 ( .A1(n18413), .A2(n18412), .Z(n18426) );
  NAND2HSV0 U21410 ( .A1(n28019), .A2(n28643), .ZN(n18415) );
  XOR2HSV0 U21411 ( .A1(n18415), .A2(n18414), .Z(n18418) );
  XNOR2HSV1 U21412 ( .A1(n18418), .A2(n18417), .ZN(n18424) );
  NAND2HSV0 U21413 ( .A1(\pe9/aot [7]), .A2(\pe9/bq[13] ), .ZN(n18500) );
  NAND2HSV0 U21414 ( .A1(\pe9/aot [8]), .A2(\pe9/bq[13] ), .ZN(n18419) );
  OAI21HSV1 U21415 ( .A1(n18566), .A2(n22378), .B(n18419), .ZN(n18420) );
  OAI21HSV2 U21416 ( .A1(n18500), .A2(n18421), .B(n18420), .ZN(n18422) );
  NAND2HSV0 U21417 ( .A1(\pe9/aot [15]), .A2(\pe9/bq[6] ), .ZN(n18493) );
  XNOR2HSV1 U21418 ( .A1(n18422), .A2(n18493), .ZN(n18423) );
  XNOR2HSV1 U21419 ( .A1(n18424), .A2(n18423), .ZN(n18425) );
  XNOR2HSV1 U21420 ( .A1(n18426), .A2(n18425), .ZN(n18427) );
  XOR3HSV1 U21421 ( .A1(n18429), .A2(n18428), .A3(n18427), .Z(n18430) );
  XNOR2HSV1 U21422 ( .A1(n18431), .A2(n18430), .ZN(n18432) );
  XOR2HSV0 U21423 ( .A1(n18433), .A2(n18432), .Z(n18435) );
  NAND2HSV0 U21424 ( .A1(n28166), .A2(n28227), .ZN(n18434) );
  INHSV2 U21425 ( .I(n18470), .ZN(n18445) );
  INHSV2 U21426 ( .I(n18445), .ZN(n18466) );
  NAND3HSV2 U21427 ( .A1(n18467), .A2(n18447), .A3(n18466), .ZN(n18452) );
  INHSV2 U21428 ( .I(n18468), .ZN(n18646) );
  AOI21HSV2 U21429 ( .A1(n18470), .A2(n18646), .B(n18552), .ZN(n18446) );
  INHSV2 U21430 ( .I(n18446), .ZN(n18448) );
  NOR2HSV2 U21431 ( .A1(n18447), .A2(n18448), .ZN(n18444) );
  CLKAND2HSV1 U21432 ( .A1(n18446), .A2(n18445), .Z(n18449) );
  INHSV4 U21433 ( .I(n18528), .ZN(n18525) );
  NOR2HSV2 U21434 ( .A1(n18050), .A2(\pe9/ti_7t [11]), .ZN(n18553) );
  INHSV1 U21435 ( .I(n25633), .ZN(n23448) );
  OR2HSV1 U21436 ( .A1(n18553), .A2(n23448), .Z(n18457) );
  INHSV4 U21437 ( .I(n18535), .ZN(n18461) );
  INHSV2 U21438 ( .I(n18534), .ZN(n18460) );
  NAND2HSV2 U21439 ( .A1(n18462), .A2(\pe9/ti_7t [12]), .ZN(n18536) );
  INHSV2 U21440 ( .I(n18536), .ZN(n19808) );
  INHSV2 U21441 ( .I(n18648), .ZN(n23719) );
  CLKNAND2HSV3 U21442 ( .A1(n18467), .A2(n18466), .ZN(n18472) );
  CLKNHSV0 U21443 ( .I(n18468), .ZN(n18545) );
  AOI21HSV2 U21444 ( .A1(n18470), .A2(n18545), .B(n18469), .ZN(n18471) );
  CLKNAND2HSV1 U21445 ( .A1(n28952), .A2(n28423), .ZN(n18519) );
  NAND2HSV0 U21446 ( .A1(n28166), .A2(n14073), .ZN(n18515) );
  NAND2HSV0 U21447 ( .A1(\pe9/aot [4]), .A2(n28044), .ZN(n18474) );
  NAND2HSV0 U21448 ( .A1(\pe9/aot [16]), .A2(\pe9/bq[4] ), .ZN(n18473) );
  XOR2HSV0 U21449 ( .A1(n18474), .A2(n18473), .Z(n18477) );
  CLKNAND2HSV0 U21450 ( .A1(n27093), .A2(\pe9/pvq [13]), .ZN(n18475) );
  XNOR2HSV1 U21451 ( .A1(n18475), .A2(\pe9/phq [13]), .ZN(n18476) );
  XNOR2HSV1 U21452 ( .A1(n18477), .A2(n18476), .ZN(n18478) );
  AND2HSV2 U21453 ( .A1(n18478), .A2(\pe9/got [8]), .Z(n18480) );
  AOI21HSV0 U21454 ( .A1(\pe9/got [8]), .A2(n28949), .B(n18478), .ZN(n18479)
         );
  AOI21HSV2 U21455 ( .A1(n18480), .A2(n28059), .B(n18479), .ZN(n18513) );
  CLKNAND2HSV0 U21456 ( .A1(n28804), .A2(\pe9/got [7]), .ZN(n18511) );
  INHSV2 U21457 ( .I(\pe9/got [5]), .ZN(n28262) );
  NOR2HSV0 U21458 ( .A1(n18481), .A2(n28262), .ZN(n18509) );
  NAND2HSV0 U21459 ( .A1(\pe9/got [6]), .A2(n11863), .ZN(n18508) );
  NAND2HSV0 U21460 ( .A1(\pe9/aot [8]), .A2(\pe9/bq[12] ), .ZN(n18483) );
  NAND2HSV0 U21461 ( .A1(\pe9/aot [12]), .A2(\pe9/bq[8] ), .ZN(n18482) );
  XOR2HSV0 U21462 ( .A1(n18483), .A2(n18482), .Z(n18487) );
  NAND2HSV0 U21463 ( .A1(\pe9/aot [9]), .A2(\pe9/bq[11] ), .ZN(n18485) );
  NAND2HSV0 U21464 ( .A1(\pe9/bq[7] ), .A2(\pe9/aot [13]), .ZN(n18484) );
  XOR2HSV0 U21465 ( .A1(n18485), .A2(n18484), .Z(n18486) );
  XOR2HSV0 U21466 ( .A1(n18487), .A2(n18486), .Z(n18497) );
  NAND2HSV0 U21467 ( .A1(n21761), .A2(\pe9/aot [5]), .ZN(n18489) );
  NAND2HSV0 U21468 ( .A1(\pe9/aot [10]), .A2(\pe9/bq[10] ), .ZN(n18488) );
  XOR2HSV0 U21469 ( .A1(n18489), .A2(n18488), .Z(n18495) );
  CLKNAND2HSV0 U21470 ( .A1(\pe9/aot [14]), .A2(\pe9/bq[5] ), .ZN(n28089) );
  CLKNHSV0 U21471 ( .I(\pe9/aot [14]), .ZN(n18491) );
  NAND2HSV0 U21472 ( .A1(\pe9/aot [15]), .A2(\pe9/bq[5] ), .ZN(n18490) );
  OAI21HSV0 U21473 ( .A1(n18491), .A2(n28199), .B(n18490), .ZN(n18492) );
  OAI21HSV0 U21474 ( .A1(n18493), .A2(n28089), .B(n18492), .ZN(n18494) );
  XNOR2HSV1 U21475 ( .A1(n18495), .A2(n18494), .ZN(n18496) );
  XNOR2HSV1 U21476 ( .A1(n18497), .A2(n18496), .ZN(n18506) );
  NAND2HSV0 U21477 ( .A1(\pe9/got [4]), .A2(n18498), .ZN(n18499) );
  XOR2HSV0 U21478 ( .A1(n18500), .A2(n18499), .Z(n18504) );
  NAND2HSV0 U21479 ( .A1(\pe9/aot [11]), .A2(\pe9/bq[9] ), .ZN(n18502) );
  NAND2HSV0 U21480 ( .A1(\pe9/aot [6]), .A2(n23822), .ZN(n18501) );
  XOR2HSV0 U21481 ( .A1(n18502), .A2(n18501), .Z(n18503) );
  XOR2HSV0 U21482 ( .A1(n18504), .A2(n18503), .Z(n18505) );
  XNOR2HSV1 U21483 ( .A1(n18506), .A2(n18505), .ZN(n18507) );
  XOR3HSV1 U21484 ( .A1(n18509), .A2(n18508), .A3(n18507), .Z(n18510) );
  XNOR2HSV1 U21485 ( .A1(n18511), .A2(n18510), .ZN(n18512) );
  XOR2HSV0 U21486 ( .A1(n18513), .A2(n18512), .Z(n18514) );
  XNOR2HSV1 U21487 ( .A1(n18515), .A2(n18514), .ZN(n18517) );
  CLKNAND2HSV1 U21488 ( .A1(n28689), .A2(n28227), .ZN(n18516) );
  XNOR2HSV1 U21489 ( .A1(n18517), .A2(n18516), .ZN(n18518) );
  XNOR2HSV1 U21490 ( .A1(n18519), .A2(n18518), .ZN(n18521) );
  XNOR2HSV4 U21491 ( .A1(n18614), .A2(n18615), .ZN(n18533) );
  CLKNAND2HSV4 U21492 ( .A1(n18527), .A2(n18526), .ZN(n18620) );
  NAND2HSV2 U21493 ( .A1(n18529), .A2(n18528), .ZN(n18555) );
  OR2HSV1 U21494 ( .A1(n18553), .A2(n18530), .Z(n18618) );
  INHSV2 U21495 ( .I(n18618), .ZN(n18531) );
  CLKNAND2HSV2 U21496 ( .A1(n18555), .A2(n18531), .ZN(n18616) );
  NOR2HSV4 U21497 ( .A1(n18620), .A2(n18616), .ZN(n18532) );
  XNOR2HSV4 U21498 ( .A1(n18533), .A2(n18532), .ZN(n25683) );
  NAND2HSV2 U21499 ( .A1(\pe9/ti_7t [13]), .A2(n18641), .ZN(n18538) );
  XNOR2HSV4 U21500 ( .A1(n18535), .A2(n18534), .ZN(n28705) );
  NAND2HSV0 U21501 ( .A1(n18536), .A2(n18628), .ZN(n18537) );
  CLKNAND2HSV1 U21502 ( .A1(n18537), .A2(n28669), .ZN(n25682) );
  NOR2HSV0 U21503 ( .A1(n18539), .A2(n18330), .ZN(n18540) );
  INHSV2 U21504 ( .I(n18541), .ZN(n18542) );
  NOR2HSV2 U21505 ( .A1(n25682), .A2(n18462), .ZN(n18544) );
  CLKNAND2HSV1 U21506 ( .A1(n23719), .A2(n18546), .ZN(n18547) );
  INHSV2 U21507 ( .I(n18547), .ZN(n18638) );
  NAND2HSV2 U21508 ( .A1(n18648), .A2(n18549), .ZN(n18548) );
  CLKNAND2HSV2 U21509 ( .A1(n18548), .A2(n23244), .ZN(n18550) );
  NOR2HSV2 U21510 ( .A1(n18648), .A2(n18549), .ZN(n28343) );
  NAND2HSV4 U21511 ( .A1(n28133), .A2(n14039), .ZN(n18635) );
  NOR2HSV1 U21512 ( .A1(n23449), .A2(n18551), .ZN(n18557) );
  NOR2HSV0 U21513 ( .A1(n18553), .A2(n18552), .ZN(n18554) );
  CLKNAND2HSV0 U21514 ( .A1(n18555), .A2(n18554), .ZN(n18556) );
  AOI21HSV2 U21515 ( .A1(n18557), .A2(n18560), .B(n18556), .ZN(n18563) );
  CLKNAND2HSV1 U21516 ( .A1(n23449), .A2(n18558), .ZN(n18559) );
  OR2HSV1 U21517 ( .A1(n18560), .A2(n18559), .Z(n18561) );
  INHSV2 U21518 ( .I(n18561), .ZN(n18562) );
  INOR2HSV4 U21519 ( .A1(n18563), .B1(n18562), .ZN(n18610) );
  CLKNAND2HSV2 U21520 ( .A1(n19767), .A2(\pe9/got [12]), .ZN(n18608) );
  CLKNAND2HSV0 U21521 ( .A1(n28264), .A2(n28227), .ZN(n18603) );
  NAND2HSV0 U21522 ( .A1(n28804), .A2(\pe9/got [6]), .ZN(n18596) );
  NAND2HSV0 U21523 ( .A1(\pe9/aot [12]), .A2(\pe9/bq[7] ), .ZN(n18565) );
  XOR2HSV0 U21524 ( .A1(n28089), .A2(n18565), .Z(n18576) );
  NOR2HSV0 U21525 ( .A1(n18566), .A2(n28199), .ZN(n22343) );
  AOI22HSV0 U21526 ( .A1(\pe9/bq[6] ), .A2(\pe9/aot [13]), .B1(\pe9/bq[12] ), 
        .B2(\pe9/aot [7]), .ZN(n18567) );
  AOI21HSV0 U21527 ( .A1(n22343), .A2(n18568), .B(n18567), .ZN(n18569) );
  NAND2HSV0 U21528 ( .A1(\pe9/bq[11] ), .A2(\pe9/aot [8]), .ZN(n22333) );
  XOR2HSV0 U21529 ( .A1(n18569), .A2(n22333), .Z(n18575) );
  NAND2HSV0 U21530 ( .A1(\pe9/aot [3]), .A2(\pe9/bq[16] ), .ZN(n18571) );
  NAND2HSV0 U21531 ( .A1(\pe9/aot [4]), .A2(\pe9/bq[15] ), .ZN(n18570) );
  XOR2HSV0 U21532 ( .A1(n18571), .A2(n18570), .Z(n18573) );
  XOR2HSV0 U21533 ( .A1(n18573), .A2(n18572), .Z(n18574) );
  XOR3HSV2 U21534 ( .A1(n18576), .A2(n18575), .A3(n18574), .Z(n18594) );
  NAND2HSV0 U21535 ( .A1(n28110), .A2(n28643), .ZN(n18593) );
  NAND2HSV0 U21536 ( .A1(\pe9/aot [11]), .A2(\pe9/bq[8] ), .ZN(n18578) );
  NAND2HSV0 U21537 ( .A1(\pe9/aot [10]), .A2(\pe9/bq[9] ), .ZN(n18577) );
  XOR2HSV0 U21538 ( .A1(n18578), .A2(n18577), .Z(n18582) );
  NAND2HSV0 U21539 ( .A1(\pe9/aot [6]), .A2(\pe9/bq[13] ), .ZN(n18580) );
  NAND2HSV0 U21540 ( .A1(\pe9/aot [5]), .A2(n23822), .ZN(n18579) );
  XOR2HSV0 U21541 ( .A1(n18580), .A2(n18579), .Z(n18581) );
  XOR2HSV0 U21542 ( .A1(n18582), .A2(n18581), .Z(n18589) );
  NAND2HSV0 U21543 ( .A1(\pe9/aot [9]), .A2(\pe9/bq[10] ), .ZN(n18584) );
  XOR2HSV0 U21544 ( .A1(n18584), .A2(n18583), .Z(n18587) );
  NAND2HSV0 U21545 ( .A1(n27093), .A2(\pe9/pvq [14]), .ZN(n18585) );
  XOR2HSV0 U21546 ( .A1(n18585), .A2(\pe9/phq [14]), .Z(n18586) );
  XOR2HSV0 U21547 ( .A1(n18587), .A2(n18586), .Z(n18588) );
  XOR2HSV0 U21548 ( .A1(n18589), .A2(n18588), .Z(n18591) );
  BUFHSV2 U21549 ( .I(\pe9/got [4]), .Z(n28389) );
  NAND2HSV0 U21550 ( .A1(n28688), .A2(n28389), .ZN(n18590) );
  XNOR2HSV1 U21551 ( .A1(n18591), .A2(n18590), .ZN(n18592) );
  XOR3HSV2 U21552 ( .A1(n18594), .A2(n18593), .A3(n18592), .Z(n18595) );
  XOR2HSV0 U21553 ( .A1(n18596), .A2(n18595), .Z(n18598) );
  CLKNAND2HSV1 U21554 ( .A1(n28059), .A2(\pe9/got [7]), .ZN(n18597) );
  XOR2HSV0 U21555 ( .A1(n18598), .A2(n18597), .Z(n18601) );
  NAND2HSV0 U21556 ( .A1(n12295), .A2(n14073), .ZN(n18600) );
  NAND2HSV0 U21557 ( .A1(n28166), .A2(\pe9/got [8]), .ZN(n18599) );
  XOR3HSV2 U21558 ( .A1(n18601), .A2(n18600), .A3(n18599), .Z(n18602) );
  XNOR2HSV1 U21559 ( .A1(n18603), .A2(n18602), .ZN(n18606) );
  XNOR2HSV4 U21560 ( .A1(n18606), .A2(n18605), .ZN(n18607) );
  XNOR2HSV4 U21561 ( .A1(n18608), .A2(n18607), .ZN(n18609) );
  XNOR2HSV4 U21562 ( .A1(n18635), .A2(n18634), .ZN(n19814) );
  NOR2HSV2 U21563 ( .A1(n25683), .A2(n18646), .ZN(n18612) );
  NAND2HSV4 U21564 ( .A1(n28705), .A2(n18611), .ZN(n19809) );
  CLKNAND2HSV2 U21565 ( .A1(n18612), .A2(n18625), .ZN(n18633) );
  NAND2HSV2 U21566 ( .A1(n18613), .A2(\pe9/ti_7t [14]), .ZN(n23245) );
  BUFHSV2 U21567 ( .I(n23245), .Z(n19817) );
  NAND2HSV2 U21568 ( .A1(n18633), .A2(n19817), .ZN(n18626) );
  INHSV2 U21569 ( .I(n18614), .ZN(n18622) );
  NOR2HSV0 U21570 ( .A1(n18618), .A2(n18617), .ZN(n18619) );
  CLKNAND2HSV0 U21571 ( .A1(n18619), .A2(n28795), .ZN(n18621) );
  NOR2HSV4 U21572 ( .A1(n18625), .A2(n18624), .ZN(n18631) );
  NAND2HSV4 U21573 ( .A1(n18627), .A2(n19814), .ZN(n18644) );
  CLKNAND2HSV1 U21574 ( .A1(n23245), .A2(n18628), .ZN(n28340) );
  INOR2HSV1 U21575 ( .A1(n28340), .B1(n18629), .ZN(n18642) );
  CLKNAND2HSV4 U21576 ( .A1(n18644), .A2(n18642), .ZN(n18637) );
  CLKNHSV0 U21577 ( .I(\pe9/ti_7t [13]), .ZN(n18630) );
  NOR2HSV4 U21578 ( .A1(n18631), .A2(n13984), .ZN(n18632) );
  XNOR2HSV4 U21579 ( .A1(n18635), .A2(n18634), .ZN(n19816) );
  NOR2HSV8 U21580 ( .A1(n18636), .A2(n19816), .ZN(n18639) );
  NOR2HSV8 U21581 ( .A1(n18637), .A2(n18639), .ZN(n23720) );
  MUX2NHSV4 U21582 ( .I0(n18638), .I1(n28346), .S(n23720), .ZN(n25692) );
  INHSV2 U21583 ( .I(n18639), .ZN(n18640) );
  CLKNHSV2 U21584 ( .I(n18640), .ZN(n18654) );
  NAND2HSV2 U21585 ( .A1(\pe9/ti_7t [15]), .A2(n18641), .ZN(n18649) );
  AND2HSV2 U21586 ( .A1(n18642), .A2(n18649), .Z(n18643) );
  NOR2HSV4 U21587 ( .A1(n28344), .A2(n18646), .ZN(n18652) );
  CLKNAND2HSV2 U21588 ( .A1(n18648), .A2(n18647), .ZN(n28345) );
  OAI21HSV4 U21589 ( .A1(n28345), .A2(n18650), .B(n18649), .ZN(n18651) );
  OAI22HSV4 U21590 ( .A1(n18654), .A2(n18653), .B1(n18651), .B2(n18652), .ZN(
        n25691) );
  CLKNAND2HSV2 U21591 ( .A1(n25692), .A2(n25691), .ZN(n28943) );
  INHSV2 U21592 ( .I(n11929), .ZN(n19357) );
  INHSV2 U21593 ( .I(n28146), .ZN(n28419) );
  NAND2HSV2 U21594 ( .A1(n18655), .A2(n13998), .ZN(n18656) );
  CLKNAND2HSV0 U21595 ( .A1(n18716), .A2(n19940), .ZN(n18658) );
  BUFHSV2 U21596 ( .I(n16385), .Z(n27225) );
  CLKNHSV0 U21597 ( .I(\pe8/got [8]), .ZN(n25527) );
  NOR2HSV2 U21598 ( .A1(n27225), .A2(n25527), .ZN(n18683) );
  NAND2HSV0 U21599 ( .A1(\pe8/bq[8] ), .A2(\pe8/aot [15]), .ZN(n18660) );
  NAND2HSV0 U21600 ( .A1(\pe8/bq[9] ), .A2(\pe8/aot [14]), .ZN(n18659) );
  XOR2HSV0 U21601 ( .A1(n18660), .A2(n18659), .Z(n18664) );
  NAND2HSV0 U21602 ( .A1(\pe8/aot [8]), .A2(n25532), .ZN(n18662) );
  NAND2HSV0 U21603 ( .A1(\pe8/aot [10]), .A2(\pe8/bq[13] ), .ZN(n18661) );
  XOR2HSV0 U21604 ( .A1(n18662), .A2(n18661), .Z(n18663) );
  XOR2HSV0 U21605 ( .A1(n18664), .A2(n18663), .Z(n18672) );
  NOR2HSV1 U21606 ( .A1(n23869), .A2(n25531), .ZN(n18666) );
  NAND2HSV0 U21607 ( .A1(\pe8/aot [11]), .A2(\pe8/bq[12] ), .ZN(n18665) );
  NAND2HSV0 U21608 ( .A1(\pe8/aot [9]), .A2(n23627), .ZN(n18668) );
  NAND2HSV0 U21609 ( .A1(n28627), .A2(\pe8/bq[7] ), .ZN(n18667) );
  XOR2HSV0 U21610 ( .A1(n18668), .A2(n18667), .Z(n18669) );
  XOR2HSV0 U21611 ( .A1(n18672), .A2(n18671), .Z(n18682) );
  NAND2HSV0 U21612 ( .A1(\pe8/aot [12]), .A2(\pe8/bq[11] ), .ZN(n18679) );
  CLKNAND2HSV1 U21613 ( .A1(n23519), .A2(\pe8/pvq [10]), .ZN(n18674) );
  XNOR2HSV1 U21614 ( .A1(n18674), .A2(\pe8/phq [10]), .ZN(n18678) );
  NAND2HSV0 U21615 ( .A1(\pe8/bq[10] ), .A2(\pe8/aot [13]), .ZN(n18676) );
  NAND2HSV0 U21616 ( .A1(\pe8/aot [7]), .A2(n25539), .ZN(n18675) );
  XOR2HSV0 U21617 ( .A1(n18676), .A2(n18675), .Z(n18677) );
  XOR3HSV2 U21618 ( .A1(n18679), .A2(n18678), .A3(n18677), .Z(n18681) );
  CLKNAND2HSV1 U21619 ( .A1(n20009), .A2(\pe8/got [9]), .ZN(n18680) );
  XOR4HSV1 U21620 ( .A1(n18683), .A2(n18682), .A3(n18681), .A4(n18680), .Z(
        n18685) );
  NAND2HSV0 U21621 ( .A1(n18746), .A2(\pe8/got [10]), .ZN(n18684) );
  XOR2HSV0 U21622 ( .A1(n18685), .A2(n18684), .Z(n18687) );
  INAND2HSV2 U21623 ( .A1(n18823), .B1(n23653), .ZN(n18686) );
  XOR2HSV0 U21624 ( .A1(n18687), .A2(n18686), .Z(n18688) );
  NAND2HSV2 U21625 ( .A1(n18828), .A2(n22136), .ZN(n18692) );
  CLKXOR2HSV2 U21626 ( .A1(n18693), .A2(n18692), .Z(n18695) );
  NAND2HSV2 U21627 ( .A1(n18694), .A2(n18695), .ZN(n18699) );
  INHSV2 U21628 ( .I(n18694), .ZN(n18697) );
  INHSV2 U21629 ( .I(n18695), .ZN(n18696) );
  CLKNAND2HSV2 U21630 ( .A1(n18697), .A2(n18696), .ZN(n18698) );
  CLKNAND2HSV3 U21631 ( .A1(n18698), .A2(n18699), .ZN(n18702) );
  INHSV3 U21632 ( .I(n18702), .ZN(n18700) );
  CLKNAND2HSV2 U21633 ( .A1(n18703), .A2(n18702), .ZN(n18704) );
  INHSV2 U21634 ( .I(n18714), .ZN(n18707) );
  NAND3HSV3 U21635 ( .A1(n28815), .A2(n18709), .A3(n22125), .ZN(n18711) );
  OA21HSV2 U21636 ( .A1(n18787), .A2(\pe8/ti_7t [9]), .B(n19835), .Z(n18710)
         );
  XNOR2HSV4 U21637 ( .A1(n18774), .A2(n18713), .ZN(n19949) );
  CLKAND2HSV2 U21638 ( .A1(\pe8/ti_7t [8]), .A2(n18767), .Z(n18715) );
  CLKNAND2HSV0 U21639 ( .A1(n18716), .A2(n22136), .ZN(n18717) );
  CLKNAND2HSV1 U21640 ( .A1(n12404), .A2(n23653), .ZN(n18752) );
  NOR2HSV2 U21641 ( .A1(n27225), .A2(n23869), .ZN(n18745) );
  CLKNAND2HSV0 U21642 ( .A1(n23605), .A2(n20009), .ZN(n18744) );
  NAND2HSV0 U21643 ( .A1(\pe8/aot [13]), .A2(\pe8/bq[9] ), .ZN(n18719) );
  NAND2HSV0 U21644 ( .A1(\pe8/aot [12]), .A2(\pe8/bq[10] ), .ZN(n18718) );
  XOR2HSV0 U21645 ( .A1(n18719), .A2(n18718), .Z(n18724) );
  NAND2HSV0 U21646 ( .A1(\pe8/aot [6]), .A2(n25539), .ZN(n18722) );
  NAND2HSV0 U21647 ( .A1(\pe8/aot [7]), .A2(n18720), .ZN(n18721) );
  XOR2HSV0 U21648 ( .A1(n18722), .A2(n18721), .Z(n18723) );
  XOR2HSV0 U21649 ( .A1(n18724), .A2(n18723), .Z(n18732) );
  NAND2HSV0 U21650 ( .A1(\pe8/aot [14]), .A2(\pe8/bq[8] ), .ZN(n18726) );
  NAND2HSV0 U21651 ( .A1(\pe8/aot [11]), .A2(\pe8/bq[11] ), .ZN(n18725) );
  XOR2HSV0 U21652 ( .A1(n18726), .A2(n18725), .Z(n18730) );
  NAND2HSV0 U21653 ( .A1(\pe8/aot [15]), .A2(\pe8/bq[7] ), .ZN(n18728) );
  NAND2HSV0 U21654 ( .A1(\pe8/aot [10]), .A2(\pe8/bq[12] ), .ZN(n18727) );
  XOR2HSV0 U21655 ( .A1(n18728), .A2(n18727), .Z(n18729) );
  XOR2HSV0 U21656 ( .A1(n18730), .A2(n18729), .Z(n18731) );
  XOR2HSV0 U21657 ( .A1(n18732), .A2(n18731), .Z(n18742) );
  NAND2HSV0 U21658 ( .A1(\pe8/got [6]), .A2(n25624), .ZN(n18734) );
  NAND2HSV0 U21659 ( .A1(n28627), .A2(\pe8/bq[6] ), .ZN(n18733) );
  XOR2HSV0 U21660 ( .A1(n18734), .A2(n18733), .Z(n18737) );
  CLKNAND2HSV1 U21661 ( .A1(n23528), .A2(\pe8/pvq [11]), .ZN(n18735) );
  XNOR2HSV1 U21662 ( .A1(n18735), .A2(\pe8/phq [11]), .ZN(n18736) );
  XNOR2HSV1 U21663 ( .A1(n18737), .A2(n18736), .ZN(n18740) );
  NAND2HSV0 U21664 ( .A1(\pe8/aot [8]), .A2(\pe8/bq[14] ), .ZN(n22150) );
  NAND2HSV0 U21665 ( .A1(\pe8/aot [9]), .A2(\pe8/bq[13] ), .ZN(n18738) );
  XOR2HSV0 U21666 ( .A1(n22150), .A2(n18738), .Z(n18739) );
  XNOR2HSV1 U21667 ( .A1(n18740), .A2(n18739), .ZN(n18741) );
  XNOR2HSV1 U21668 ( .A1(n18742), .A2(n18741), .ZN(n18743) );
  XOR3HSV2 U21669 ( .A1(n18745), .A2(n18744), .A3(n18743), .Z(n18748) );
  NAND2HSV0 U21670 ( .A1(n18746), .A2(n23721), .ZN(n18747) );
  XNOR2HSV1 U21671 ( .A1(n18748), .A2(n18747), .ZN(n18750) );
  INAND2HSV2 U21672 ( .A1(n18823), .B1(\pe8/got [10]), .ZN(n18749) );
  XOR2HSV0 U21673 ( .A1(n18750), .A2(n18749), .Z(n18751) );
  XNOR2HSV1 U21674 ( .A1(n18752), .A2(n18751), .ZN(n18754) );
  XNOR2HSV4 U21675 ( .A1(n18756), .A2(n18755), .ZN(n18761) );
  CLKNHSV2 U21676 ( .I(n18761), .ZN(n18757) );
  INHSV2 U21677 ( .I(n18757), .ZN(n18758) );
  CLKNAND2HSV2 U21678 ( .A1(n18759), .A2(n18758), .ZN(n18764) );
  NOR2HSV2 U21679 ( .A1(n18761), .A2(n18760), .ZN(n18762) );
  NAND2HSV4 U21680 ( .A1(n18764), .A2(n18763), .ZN(n19943) );
  CLKBUFHSV4 U21681 ( .I(n19943), .Z(n18772) );
  INHSV2 U21682 ( .I(n18772), .ZN(n18765) );
  INAND2HSV2 U21683 ( .A1(n19943), .B1(n19835), .ZN(n19948) );
  BUFHSV2 U21684 ( .I(n28667), .Z(n19904) );
  CLKNAND2HSV2 U21685 ( .A1(n18772), .A2(n19904), .ZN(n19944) );
  NAND2HSV2 U21686 ( .A1(n18788), .A2(\pe8/ti_7t [9]), .ZN(n18785) );
  AOI21HSV2 U21687 ( .A1(n18785), .A2(n18767), .B(n18766), .ZN(n18776) );
  CLKNAND2HSV2 U21688 ( .A1(n19944), .A2(n18768), .ZN(n18769) );
  AOI21HSV4 U21689 ( .A1(n18771), .A2(n18770), .B(n18769), .ZN(n18782) );
  NOR2HSV2 U21690 ( .A1(n18774), .A2(n28667), .ZN(n19956) );
  INHSV3 U21691 ( .I(n19943), .ZN(n21320) );
  NOR2HSV0 U21692 ( .A1(n18788), .A2(n28667), .ZN(n18775) );
  NAND2HSV2 U21693 ( .A1(n19952), .A2(n18775), .ZN(n18777) );
  AOI21HSV2 U21694 ( .A1(n21320), .A2(n18777), .B(n21315), .ZN(n18778) );
  NAND2HSV2 U21695 ( .A1(n19969), .A2(\pe8/ti_7t [11]), .ZN(n19960) );
  CLKNAND2HSV4 U21696 ( .A1(n18780), .A2(n19960), .ZN(n18781) );
  NOR2HSV8 U21697 ( .A1(n18782), .A2(n18781), .ZN(n19900) );
  NAND2HSV2 U21698 ( .A1(n19992), .A2(n18784), .ZN(n18837) );
  CLKNAND2HSV2 U21699 ( .A1(n21322), .A2(n28599), .ZN(n18836) );
  INHSV2 U21700 ( .I(n22141), .ZN(n19994) );
  INHSV1 U21701 ( .I(\pe8/got [12]), .ZN(n18789) );
  NOR2HSV4 U21702 ( .A1(n19994), .A2(n18789), .ZN(n18832) );
  INHSV2 U21703 ( .I(n22310), .ZN(n28462) );
  NAND2HSV0 U21704 ( .A1(n28462), .A2(\pe8/got [10]), .ZN(n18827) );
  NAND2HSV0 U21705 ( .A1(n28796), .A2(\pe8/got [6]), .ZN(n18819) );
  NAND2HSV0 U21706 ( .A1(n20009), .A2(n14068), .ZN(n18818) );
  NAND2HSV0 U21707 ( .A1(\pe8/aot [11]), .A2(\pe8/bq[10] ), .ZN(n18791) );
  NAND2HSV0 U21708 ( .A1(\pe8/aot [10]), .A2(\pe8/bq[11] ), .ZN(n18790) );
  XOR2HSV0 U21709 ( .A1(n18791), .A2(n18790), .Z(n18795) );
  NAND2HSV0 U21710 ( .A1(\pe8/bq[6] ), .A2(\pe8/aot [15]), .ZN(n18793) );
  NAND2HSV0 U21711 ( .A1(\pe8/aot [6]), .A2(n25532), .ZN(n18792) );
  XOR2HSV0 U21712 ( .A1(n18793), .A2(n18792), .Z(n18794) );
  XOR2HSV0 U21713 ( .A1(n18795), .A2(n18794), .Z(n18801) );
  NAND2HSV0 U21714 ( .A1(\pe8/aot [12]), .A2(\pe8/bq[9] ), .ZN(n22284) );
  INHSV2 U21715 ( .I(\pe8/bq[5] ), .ZN(n23847) );
  INHSV2 U21716 ( .I(n23847), .ZN(n23529) );
  CLKNAND2HSV0 U21717 ( .A1(n28627), .A2(n23529), .ZN(n19847) );
  XOR2HSV0 U21718 ( .A1(n22284), .A2(n19847), .Z(n18799) );
  CLKNAND2HSV0 U21719 ( .A1(\pe8/got [5]), .A2(n25624), .ZN(n18797) );
  NAND2HSV0 U21720 ( .A1(\pe8/aot [7]), .A2(n23627), .ZN(n18796) );
  XOR2HSV0 U21721 ( .A1(n18797), .A2(n18796), .Z(n18798) );
  XOR2HSV0 U21722 ( .A1(n18799), .A2(n18798), .Z(n18800) );
  XOR2HSV0 U21723 ( .A1(n18801), .A2(n18800), .Z(n18816) );
  NAND2HSV0 U21724 ( .A1(\pe8/aot [5]), .A2(n25539), .ZN(n18803) );
  NAND2HSV0 U21725 ( .A1(\pe8/bq[8] ), .A2(\pe8/aot [13]), .ZN(n18802) );
  XOR2HSV0 U21726 ( .A1(n18803), .A2(n18802), .Z(n18806) );
  CLKNAND2HSV0 U21727 ( .A1(n23519), .A2(\pe8/pvq [12]), .ZN(n18804) );
  XNOR2HSV1 U21728 ( .A1(n18804), .A2(\pe8/phq [12]), .ZN(n18805) );
  XNOR2HSV1 U21729 ( .A1(n18806), .A2(n18805), .ZN(n18814) );
  CLKNHSV0 U21730 ( .I(\pe8/aot [14]), .ZN(n19845) );
  CLKNHSV0 U21731 ( .I(\pe8/bq[7] ), .ZN(n18808) );
  NAND2HSV0 U21732 ( .A1(\pe8/aot [9]), .A2(\pe8/bq[12] ), .ZN(n18807) );
  OAI21HSV2 U21733 ( .A1(n19845), .A2(n18808), .B(n18807), .ZN(n18809) );
  OAI21HSV0 U21734 ( .A1(n23727), .A2(n18810), .B(n18809), .ZN(n18812) );
  CLKNHSV0 U21735 ( .I(\pe8/bq[13] ), .ZN(n18811) );
  INHSV2 U21736 ( .I(n18811), .ZN(n25565) );
  NAND2HSV0 U21737 ( .A1(\pe8/aot [8]), .A2(n25565), .ZN(n23609) );
  XNOR2HSV1 U21738 ( .A1(n18812), .A2(n23609), .ZN(n18813) );
  XNOR2HSV1 U21739 ( .A1(n18814), .A2(n18813), .ZN(n18815) );
  XNOR2HSV1 U21740 ( .A1(n18816), .A2(n18815), .ZN(n18817) );
  XOR3HSV2 U21741 ( .A1(n18819), .A2(n18818), .A3(n18817), .Z(n18822) );
  INHSV2 U21742 ( .I(n18820), .ZN(n25578) );
  NAND2HSV0 U21743 ( .A1(n25578), .A2(n23605), .ZN(n18821) );
  XOR2HSV0 U21744 ( .A1(n18822), .A2(n18821), .Z(n18825) );
  BUFHSV4 U21745 ( .I(n18823), .Z(n23642) );
  INAND2HSV2 U21746 ( .A1(n23642), .B1(\pe8/got [9]), .ZN(n18824) );
  XOR2HSV0 U21747 ( .A1(n18825), .A2(n18824), .Z(n18826) );
  XNOR2HSV1 U21748 ( .A1(n18827), .A2(n18826), .ZN(n18830) );
  BUFHSV2 U21749 ( .I(\pe8/got [11]), .Z(n28618) );
  CLKNAND2HSV0 U21750 ( .A1(n18828), .A2(n28618), .ZN(n18829) );
  XNOR2HSV1 U21751 ( .A1(n18830), .A2(n18829), .ZN(n18831) );
  CLKXOR2HSV2 U21752 ( .A1(n18832), .A2(n18831), .Z(n18834) );
  XNOR2HSV4 U21753 ( .A1(n18834), .A2(n18833), .ZN(n18835) );
  XNOR2HSV4 U21754 ( .A1(n18836), .A2(n18835), .ZN(n18838) );
  CLKNAND2HSV3 U21755 ( .A1(n18837), .A2(n18838), .ZN(n18843) );
  INHSV4 U21756 ( .I(n18838), .ZN(n18841) );
  INHSV2 U21757 ( .I(n19901), .ZN(n18839) );
  NAND2HSV2 U21758 ( .A1(n19990), .A2(n19991), .ZN(pov8[12]) );
  NAND2HSV0 U21759 ( .A1(n28676), .A2(n28686), .ZN(n18845) );
  CLKNHSV0 U21760 ( .I(n18846), .ZN(n18848) );
  NAND3HSV0 U21761 ( .A1(n18849), .A2(n25420), .A3(n12297), .ZN(n18850) );
  NOR2HSV1 U21762 ( .A1(n18852), .A2(\pe6/ti_7t [11]), .ZN(n19129) );
  INHSV2 U21763 ( .I(n18853), .ZN(n18916) );
  CLKNAND2HSV0 U21764 ( .A1(\pe6/ti_7t [7]), .A2(n19068), .ZN(n18928) );
  CLKNHSV0 U21765 ( .I(n18928), .ZN(n18859) );
  AOI21HSV1 U21766 ( .A1(n18928), .A2(n19151), .B(n14217), .ZN(n18858) );
  CLKNHSV0 U21767 ( .I(\pe6/got [10]), .ZN(n18860) );
  NOR2HSV2 U21768 ( .A1(n12185), .A2(n18860), .ZN(n18894) );
  CLKNAND2HSV0 U21769 ( .A1(n18930), .A2(\pe6/got [7]), .ZN(n18862) );
  INHSV2 U21770 ( .I(n25785), .ZN(n25982) );
  NAND2HSV0 U21771 ( .A1(\pe6/ti_7[1] ), .A2(n25982), .ZN(n18861) );
  XNOR2HSV1 U21772 ( .A1(n18862), .A2(n18861), .ZN(n18888) );
  NAND2HSV0 U21773 ( .A1(\pe6/aot [5]), .A2(\pe6/bq[16] ), .ZN(n18864) );
  NAND2HSV0 U21774 ( .A1(\pe6/bq[9] ), .A2(\pe6/aot [12]), .ZN(n18863) );
  XOR2HSV0 U21775 ( .A1(n18864), .A2(n18863), .Z(n18868) );
  NAND2HSV0 U21776 ( .A1(\pe6/aot [10]), .A2(\pe6/bq[11] ), .ZN(n18865) );
  XOR2HSV0 U21777 ( .A1(n18866), .A2(n18865), .Z(n18867) );
  XOR2HSV0 U21778 ( .A1(n18868), .A2(n18867), .Z(n18870) );
  XOR2HSV0 U21779 ( .A1(n18870), .A2(n18869), .Z(n18886) );
  INHSV2 U21780 ( .I(n18871), .ZN(n21333) );
  INHSV2 U21781 ( .I(n21333), .ZN(n22109) );
  CLKNAND2HSV0 U21782 ( .A1(n22109), .A2(\pe6/pvq [12]), .ZN(n18872) );
  XNOR2HSV1 U21783 ( .A1(n18872), .A2(\pe6/phq [12]), .ZN(n18877) );
  NAND2HSV0 U21784 ( .A1(\pe6/aot [8]), .A2(\pe6/bq[8] ), .ZN(n23015) );
  CLKNHSV0 U21785 ( .I(\pe6/aot [8]), .ZN(n25963) );
  CLKNHSV0 U21786 ( .I(\pe6/bq[13] ), .ZN(n22107) );
  NAND2HSV0 U21787 ( .A1(\pe6/bq[8] ), .A2(\pe6/aot [13]), .ZN(n18873) );
  OAI21HSV0 U21788 ( .A1(n25963), .A2(n22107), .B(n18873), .ZN(n18874) );
  OAI21HSV0 U21789 ( .A1(n18875), .A2(n23015), .B(n18874), .ZN(n18876) );
  XOR2HSV0 U21790 ( .A1(n18877), .A2(n18876), .Z(n18884) );
  CLKNAND2HSV0 U21791 ( .A1(\pe6/aot [9]), .A2(\pe6/bq[10] ), .ZN(n19078) );
  CLKNHSV0 U21792 ( .I(\pe6/aot [9]), .ZN(n25790) );
  NAND2HSV0 U21793 ( .A1(\pe6/aot [11]), .A2(\pe6/bq[10] ), .ZN(n18878) );
  OAI21HSV0 U21794 ( .A1(n25790), .A2(n18879), .B(n18878), .ZN(n18880) );
  OAI21HSV1 U21795 ( .A1(n19078), .A2(n18881), .B(n18880), .ZN(n18882) );
  NAND2HSV2 U21796 ( .A1(n28681), .A2(\pe6/bq[5] ), .ZN(n25423) );
  XNOR2HSV1 U21797 ( .A1(n18882), .A2(n25423), .ZN(n18883) );
  XNOR2HSV1 U21798 ( .A1(n18884), .A2(n18883), .ZN(n18885) );
  XNOR2HSV1 U21799 ( .A1(n18886), .A2(n18885), .ZN(n18887) );
  XNOR2HSV1 U21800 ( .A1(n18888), .A2(n18887), .ZN(n18890) );
  XNOR2HSV1 U21801 ( .A1(n18890), .A2(n18889), .ZN(n18892) );
  CLKNAND2HSV0 U21802 ( .A1(n19109), .A2(\pe6/got [9]), .ZN(n18891) );
  XNOR2HSV1 U21803 ( .A1(n18892), .A2(n18891), .ZN(n18893) );
  XNOR2HSV1 U21804 ( .A1(n18894), .A2(n18893), .ZN(n18896) );
  CLKNAND2HSV1 U21805 ( .A1(n26033), .A2(n28586), .ZN(n18895) );
  XNOR2HSV1 U21806 ( .A1(n18896), .A2(n18895), .ZN(n18897) );
  XOR2HSV0 U21807 ( .A1(n18898), .A2(n18897), .Z(n18899) );
  NAND2HSV0 U21808 ( .A1(n28686), .A2(n28938), .ZN(n18901) );
  NAND2HSV0 U21809 ( .A1(n14285), .A2(n28938), .ZN(n18903) );
  INHSV1 U21810 ( .I(n18903), .ZN(n18904) );
  NAND2HSV2 U21811 ( .A1(n18904), .A2(n18908), .ZN(n18912) );
  CLKNHSV0 U21812 ( .I(n18997), .ZN(n18905) );
  CLKAND2HSV1 U21813 ( .A1(n18905), .A2(n25420), .Z(n18906) );
  OAI21HSV2 U21814 ( .A1(n18908), .A2(n18907), .B(n18906), .ZN(n18909) );
  INHSV2 U21815 ( .I(n18909), .ZN(n18911) );
  XNOR2HSV4 U21816 ( .A1(n18914), .A2(n18913), .ZN(n18919) );
  CLKNHSV1 U21817 ( .I(n18915), .ZN(n19068) );
  INHSV2 U21818 ( .I(n18916), .ZN(n18917) );
  INHSV2 U21819 ( .I(\pe6/ti_7t [12]), .ZN(n18993) );
  NAND2HSV2 U21820 ( .A1(n18921), .A2(n19138), .ZN(n18922) );
  CLKNAND2HSV1 U21821 ( .A1(n19068), .A2(\pe6/ti_7t [11]), .ZN(n19159) );
  CLKNHSV0 U21822 ( .I(n19159), .ZN(n18924) );
  AOI21HSV2 U21823 ( .A1(n19159), .A2(n19073), .B(n18855), .ZN(n18923) );
  NAND2HSV2 U21824 ( .A1(n19073), .A2(\pe6/ti_7t [10]), .ZN(n19072) );
  INHSV2 U21825 ( .I(n19072), .ZN(n18925) );
  INHSV2 U21826 ( .I(n18925), .ZN(n21742) );
  AOI21HSV2 U21827 ( .A1(n19073), .A2(n21742), .B(n14217), .ZN(n18926) );
  CLKNAND2HSV1 U21828 ( .A1(n19075), .A2(n18926), .ZN(n18983) );
  NAND2HSV4 U21829 ( .A1(n18929), .A2(n18928), .ZN(\pe6/ti_7[7] ) );
  NAND2HSV0 U21830 ( .A1(\pe6/ti_7[7] ), .A2(\pe6/got [9]), .ZN(n18977) );
  NAND2HSV0 U21831 ( .A1(n26033), .A2(\pe6/got [8]), .ZN(n18975) );
  INAND2HSV2 U21832 ( .A1(n14029), .B1(\pe6/got [7]), .ZN(n18973) );
  NAND2HSV0 U21833 ( .A1(n19076), .A2(\pe6/got [5]), .ZN(n18971) );
  BUFHSV3 U21834 ( .I(n18930), .Z(n25846) );
  NAND2HSV0 U21835 ( .A1(n25846), .A2(\pe6/got [4]), .ZN(n18948) );
  NAND2HSV0 U21836 ( .A1(\pe6/aot [11]), .A2(\pe6/bq[7] ), .ZN(n25709) );
  NAND2HSV0 U21837 ( .A1(\pe6/bq[4] ), .A2(\pe6/aot [14]), .ZN(n25427) );
  XOR2HSV0 U21838 ( .A1(n25709), .A2(n25427), .Z(n18946) );
  INHSV2 U21839 ( .I(n21333), .ZN(n23486) );
  CLKNAND2HSV0 U21840 ( .A1(n23486), .A2(\pe6/pvq [15]), .ZN(n18931) );
  XNOR2HSV1 U21841 ( .A1(n18931), .A2(\pe6/phq [15]), .ZN(n18937) );
  CLKNHSV0 U21842 ( .I(\pe6/aot [13]), .ZN(n18933) );
  CLKNHSV0 U21843 ( .I(\pe6/bq[5] ), .ZN(n18932) );
  NOR2HSV2 U21844 ( .A1(n18933), .A2(n18932), .ZN(n25716) );
  CLKNHSV0 U21845 ( .I(\pe6/bq[2] ), .ZN(n25990) );
  NOR2HSV0 U21846 ( .A1(n18934), .A2(n25990), .ZN(n18935) );
  CLKNAND2HSV0 U21847 ( .A1(\pe6/bq[2] ), .A2(\pe6/aot [13]), .ZN(n25841) );
  OAI22HSV1 U21848 ( .A1(n25716), .A2(n18935), .B1(n25423), .B2(n25841), .ZN(
        n18936) );
  XNOR2HSV1 U21849 ( .A1(n18937), .A2(n18936), .ZN(n18945) );
  NAND2HSV0 U21850 ( .A1(\pe6/aot [12]), .A2(\pe6/bq[6] ), .ZN(n18939) );
  NAND2HSV0 U21851 ( .A1(\pe6/aot [5]), .A2(\pe6/bq[13] ), .ZN(n18938) );
  XOR2HSV0 U21852 ( .A1(n18939), .A2(n18938), .Z(n18943) );
  NAND2HSV0 U21853 ( .A1(\pe6/aot [9]), .A2(\pe6/bq[9] ), .ZN(n18941) );
  NAND2HSV0 U21854 ( .A1(\pe6/aot [8]), .A2(\pe6/bq[10] ), .ZN(n18940) );
  XOR2HSV0 U21855 ( .A1(n18941), .A2(n18940), .Z(n18942) );
  XOR2HSV0 U21856 ( .A1(n18943), .A2(n18942), .Z(n18944) );
  XOR3HSV2 U21857 ( .A1(n18946), .A2(n18945), .A3(n18944), .Z(n18947) );
  XNOR2HSV1 U21858 ( .A1(n18948), .A2(n18947), .ZN(n18967) );
  NAND2HSV0 U21859 ( .A1(\pe6/aot [3]), .A2(\pe6/bq[15] ), .ZN(n18950) );
  NAND2HSV0 U21860 ( .A1(\pe6/aot [2]), .A2(n14028), .ZN(n18949) );
  XOR2HSV0 U21861 ( .A1(n18950), .A2(n18949), .Z(n18954) );
  NAND2HSV0 U21862 ( .A1(\pe6/aot [7]), .A2(\pe6/bq[11] ), .ZN(n18952) );
  NAND2HSV0 U21863 ( .A1(\pe6/aot [4]), .A2(\pe6/bq[14] ), .ZN(n18951) );
  XOR2HSV0 U21864 ( .A1(n18952), .A2(n18951), .Z(n18953) );
  XOR2HSV0 U21865 ( .A1(n18954), .A2(n18953), .Z(n18963) );
  NAND2HSV0 U21866 ( .A1(\pe6/got [2]), .A2(n19021), .ZN(n18957) );
  NAND2HSV0 U21867 ( .A1(\pe6/bq[8] ), .A2(\pe6/aot [10]), .ZN(n18956) );
  XOR2HSV0 U21868 ( .A1(n18957), .A2(n18956), .Z(n18961) );
  NAND2HSV0 U21869 ( .A1(\pe6/aot [6]), .A2(n25701), .ZN(n18959) );
  INHSV2 U21870 ( .I(\pe6/bq[3] ), .ZN(n25789) );
  NAND2HSV0 U21871 ( .A1(n28680), .A2(\pe6/bq[3] ), .ZN(n18958) );
  XOR2HSV0 U21872 ( .A1(n18959), .A2(n18958), .Z(n18960) );
  XOR2HSV0 U21873 ( .A1(n18961), .A2(n18960), .Z(n18962) );
  XOR2HSV0 U21874 ( .A1(n18963), .A2(n18962), .Z(n18965) );
  NOR2HSV0 U21875 ( .A1(n24963), .A2(n25932), .ZN(n18964) );
  XNOR2HSV1 U21876 ( .A1(n18965), .A2(n18964), .ZN(n18966) );
  XNOR2HSV1 U21877 ( .A1(n18967), .A2(n18966), .ZN(n18970) );
  CLKNHSV1 U21878 ( .I(n18968), .ZN(n28792) );
  NAND2HSV0 U21879 ( .A1(n28792), .A2(n25982), .ZN(n18969) );
  XOR3HSV2 U21880 ( .A1(n18971), .A2(n18970), .A3(n18969), .Z(n18972) );
  XOR2HSV0 U21881 ( .A1(n18973), .A2(n18972), .Z(n18974) );
  XNOR2HSV1 U21882 ( .A1(n18975), .A2(n18974), .ZN(n18976) );
  XNOR2HSV1 U21883 ( .A1(n18977), .A2(n18976), .ZN(n18979) );
  BUFHSV4 U21884 ( .I(n28940), .Z(n25764) );
  CLKNAND2HSV1 U21885 ( .A1(n25764), .A2(\pe6/got [10]), .ZN(n18978) );
  XOR2HSV0 U21886 ( .A1(n18979), .A2(n18978), .Z(n18981) );
  CLKBUFHSV4 U21887 ( .I(n19121), .Z(n25767) );
  NAND2HSV2 U21888 ( .A1(n25767), .A2(n14061), .ZN(n18980) );
  XNOR2HSV1 U21889 ( .A1(n18981), .A2(n18980), .ZN(n18982) );
  XNOR2HSV4 U21890 ( .A1(n18983), .A2(n18982), .ZN(n18984) );
  XNOR2HSV4 U21891 ( .A1(n18985), .A2(n18984), .ZN(n18988) );
  INHSV4 U21892 ( .I(n18988), .ZN(n18986) );
  CLKNAND2HSV2 U21893 ( .A1(n18987), .A2(n18986), .ZN(n18991) );
  NAND2HSV2 U21894 ( .A1(n18989), .A2(n18988), .ZN(n18990) );
  CLKNAND2HSV3 U21895 ( .A1(n18991), .A2(n18990), .ZN(n19062) );
  NAND3HSV2 U21896 ( .A1(n19132), .A2(n19131), .A3(n14369), .ZN(n18995) );
  INHSV2 U21897 ( .I(n25647), .ZN(n24962) );
  AOI21HSV2 U21898 ( .A1(n18993), .A2(n18992), .B(n24962), .ZN(n18994) );
  CLKNAND2HSV3 U21899 ( .A1(n18995), .A2(n18994), .ZN(n19058) );
  NOR2HSV2 U21900 ( .A1(n18997), .A2(n18996), .ZN(n18998) );
  NAND2HSV2 U21901 ( .A1(\pe6/ti_7[7] ), .A2(n14061), .ZN(n19036) );
  NAND2HSV0 U21902 ( .A1(\pe6/got [10]), .A2(n28526), .ZN(n19034) );
  INAND2HSV2 U21903 ( .A1(n22995), .B1(\pe6/got [9]), .ZN(n19032) );
  NAND2HSV0 U21904 ( .A1(n19076), .A2(\pe6/got [7]), .ZN(n19030) );
  NAND2HSV0 U21905 ( .A1(n25846), .A2(n25982), .ZN(n19000) );
  NOR2HSV0 U21906 ( .A1(n25455), .A2(n26014), .ZN(n18999) );
  XNOR2HSV1 U21907 ( .A1(n19000), .A2(n18999), .ZN(n19027) );
  NAND2HSV0 U21908 ( .A1(n28681), .A2(\pe6/bq[4] ), .ZN(n19002) );
  NAND2HSV0 U21909 ( .A1(\pe6/aot [12]), .A2(\pe6/bq[8] ), .ZN(n19001) );
  XOR2HSV0 U21910 ( .A1(n19002), .A2(n19001), .Z(n19006) );
  NAND2HSV0 U21911 ( .A1(\pe6/bq[10] ), .A2(\pe6/aot [10]), .ZN(n19004) );
  NAND2HSV0 U21912 ( .A1(\pe6/aot [7]), .A2(\pe6/bq[13] ), .ZN(n19003) );
  XOR2HSV0 U21913 ( .A1(n19004), .A2(n19003), .Z(n19005) );
  XOR2HSV0 U21914 ( .A1(n19006), .A2(n19005), .Z(n19014) );
  NAND2HSV0 U21915 ( .A1(\pe6/aot [13]), .A2(\pe6/bq[7] ), .ZN(n19008) );
  NAND2HSV0 U21916 ( .A1(\pe6/aot [9]), .A2(\pe6/bq[11] ), .ZN(n19007) );
  XOR2HSV0 U21917 ( .A1(n19008), .A2(n19007), .Z(n19012) );
  NAND2HSV0 U21918 ( .A1(\pe6/bq[16] ), .A2(\pe6/aot [4]), .ZN(n19010) );
  NAND2HSV0 U21919 ( .A1(\pe6/aot [11]), .A2(\pe6/bq[9] ), .ZN(n19009) );
  XOR2HSV0 U21920 ( .A1(n19010), .A2(n19009), .Z(n19011) );
  XOR2HSV0 U21921 ( .A1(n19012), .A2(n19011), .Z(n19013) );
  XOR2HSV0 U21922 ( .A1(n19014), .A2(n19013), .Z(n19025) );
  NAND2HSV0 U21923 ( .A1(\pe6/aot [8]), .A2(n25701), .ZN(n19016) );
  NAND2HSV0 U21924 ( .A1(\pe6/aot [5]), .A2(\pe6/bq[15] ), .ZN(n19015) );
  XOR2HSV0 U21925 ( .A1(n19016), .A2(n19015), .Z(n19020) );
  NAND2HSV0 U21926 ( .A1(\pe6/aot [6]), .A2(\pe6/bq[14] ), .ZN(n19018) );
  NAND2HSV0 U21927 ( .A1(\pe6/aot [14]), .A2(\pe6/bq[6] ), .ZN(n19017) );
  XOR2HSV0 U21928 ( .A1(n19018), .A2(n19017), .Z(n19019) );
  XOR2HSV0 U21929 ( .A1(n19020), .A2(n19019), .Z(n19023) );
  XOR2HSV0 U21930 ( .A1(n19023), .A2(n19022), .Z(n19024) );
  XOR2HSV0 U21931 ( .A1(n19025), .A2(n19024), .Z(n19026) );
  XNOR2HSV1 U21932 ( .A1(n19027), .A2(n19026), .ZN(n19029) );
  NAND2HSV0 U21933 ( .A1(n19109), .A2(\pe6/got [8]), .ZN(n19028) );
  XOR3HSV2 U21934 ( .A1(n19030), .A2(n19029), .A3(n19028), .Z(n19031) );
  XOR2HSV0 U21935 ( .A1(n19032), .A2(n19031), .Z(n19033) );
  XNOR2HSV1 U21936 ( .A1(n19034), .A2(n19033), .ZN(n19035) );
  XNOR2HSV4 U21937 ( .A1(n19036), .A2(n19035), .ZN(n19038) );
  NAND2HSV0 U21938 ( .A1(n28940), .A2(n28593), .ZN(n19037) );
  CLKXOR2HSV2 U21939 ( .A1(n19038), .A2(n19037), .Z(n19040) );
  XNOR2HSV4 U21940 ( .A1(n19042), .A2(n19041), .ZN(n19053) );
  CLKAND2HSV2 U21941 ( .A1(n19044), .A2(n19127), .Z(n19052) );
  INHSV2 U21942 ( .I(n19046), .ZN(n19130) );
  NAND3HSV2 U21943 ( .A1(n19047), .A2(n19046), .A3(n19127), .ZN(n19050) );
  NOR2HSV0 U21944 ( .A1(n19129), .A2(n19048), .ZN(n19049) );
  AOI21HSV4 U21945 ( .A1(n19052), .A2(n19130), .B(n19051), .ZN(n19054) );
  NAND2HSV2 U21946 ( .A1(\pe6/ti_7t [13]), .A2(n19055), .ZN(n25696) );
  BUFHSV2 U21947 ( .I(n25696), .Z(n19059) );
  AOI21HSV4 U21948 ( .A1(n19057), .A2(n19059), .B(n13983), .ZN(n19061) );
  INHSV2 U21949 ( .I(n19058), .ZN(n19156) );
  INHSV2 U21950 ( .I(n19070), .ZN(n19155) );
  CLKNAND2HSV3 U21951 ( .A1(n19061), .A2(n19060), .ZN(n19063) );
  INHSV3 U21952 ( .I(n19063), .ZN(n19064) );
  NOR2HSV2 U21953 ( .A1(n19070), .A2(n19138), .ZN(n19067) );
  CLKNAND2HSV2 U21954 ( .A1(n19070), .A2(n19069), .ZN(n19071) );
  NOR2HSV4 U21955 ( .A1(n22993), .A2(n19071), .ZN(n25519) );
  AOI21HSV2 U21956 ( .A1(n19073), .A2(n19072), .B(n18855), .ZN(n19074) );
  NAND2HSV0 U21957 ( .A1(\pe6/ti_7[7] ), .A2(\pe6/got [10]), .ZN(n19118) );
  NAND2HSV0 U21958 ( .A1(\pe6/got [9]), .A2(n26033), .ZN(n19116) );
  INAND2HSV2 U21959 ( .A1(n14029), .B1(\pe6/got [8]), .ZN(n19114) );
  NAND2HSV0 U21960 ( .A1(n19076), .A2(n25982), .ZN(n19112) );
  CLKNAND2HSV1 U21961 ( .A1(n25846), .A2(\pe6/got [5]), .ZN(n19090) );
  NAND2HSV0 U21962 ( .A1(n28680), .A2(\pe6/bq[4] ), .ZN(n19077) );
  XOR2HSV0 U21963 ( .A1(n19078), .A2(n19077), .Z(n19088) );
  NAND2HSV0 U21964 ( .A1(\pe6/aot [8]), .A2(\pe6/bq[11] ), .ZN(n26044) );
  XNOR2HSV1 U21965 ( .A1(n19079), .A2(n26044), .ZN(n19087) );
  NAND2HSV0 U21966 ( .A1(n28681), .A2(\pe6/bq[3] ), .ZN(n19081) );
  NAND2HSV0 U21967 ( .A1(\pe6/bq[15] ), .A2(\pe6/aot [4]), .ZN(n19080) );
  XOR2HSV0 U21968 ( .A1(n19081), .A2(n19080), .Z(n19085) );
  NAND2HSV0 U21969 ( .A1(\pe6/aot [3]), .A2(n14028), .ZN(n19083) );
  NAND2HSV0 U21970 ( .A1(\pe6/aot [6]), .A2(\pe6/bq[13] ), .ZN(n19082) );
  XOR2HSV0 U21971 ( .A1(n19083), .A2(n19082), .Z(n19084) );
  XOR2HSV0 U21972 ( .A1(n19085), .A2(n19084), .Z(n19086) );
  XOR3HSV2 U21973 ( .A1(n19088), .A2(n19087), .A3(n19086), .Z(n19089) );
  XNOR2HSV1 U21974 ( .A1(n19090), .A2(n19089), .ZN(n19108) );
  NAND2HSV0 U21975 ( .A1(\pe6/bq[7] ), .A2(\pe6/aot [12]), .ZN(n19092) );
  NAND2HSV0 U21976 ( .A1(n19021), .A2(n14008), .ZN(n19091) );
  XOR2HSV0 U21977 ( .A1(n19092), .A2(n19091), .Z(n19096) );
  NAND2HSV0 U21978 ( .A1(\pe6/aot [7]), .A2(\pe6/bq[12] ), .ZN(n19094) );
  NAND2HSV0 U21979 ( .A1(\pe6/aot [14]), .A2(\pe6/bq[5] ), .ZN(n19093) );
  XOR2HSV0 U21980 ( .A1(n19094), .A2(n19093), .Z(n19095) );
  XOR2HSV0 U21981 ( .A1(n19096), .A2(n19095), .Z(n19104) );
  NAND2HSV0 U21982 ( .A1(\pe6/bq[9] ), .A2(\pe6/aot [10]), .ZN(n19098) );
  NAND2HSV0 U21983 ( .A1(\pe6/bq[6] ), .A2(\pe6/aot [13]), .ZN(n19097) );
  XOR2HSV0 U21984 ( .A1(n19098), .A2(n19097), .Z(n19102) );
  NAND2HSV0 U21985 ( .A1(\pe6/aot [11]), .A2(\pe6/bq[8] ), .ZN(n19100) );
  NAND2HSV0 U21986 ( .A1(\pe6/aot [5]), .A2(\pe6/bq[14] ), .ZN(n19099) );
  XOR2HSV0 U21987 ( .A1(n19100), .A2(n19099), .Z(n19101) );
  XOR2HSV0 U21988 ( .A1(n19102), .A2(n19101), .Z(n19103) );
  XOR2HSV0 U21989 ( .A1(n19104), .A2(n19103), .Z(n19106) );
  NAND2HSV0 U21990 ( .A1(\pe6/ti_7[1] ), .A2(\pe6/got [4]), .ZN(n19105) );
  XNOR2HSV1 U21991 ( .A1(n19106), .A2(n19105), .ZN(n19107) );
  XNOR2HSV1 U21992 ( .A1(n19108), .A2(n19107), .ZN(n19111) );
  NAND2HSV0 U21993 ( .A1(n19109), .A2(\pe6/got [7]), .ZN(n19110) );
  XOR3HSV2 U21994 ( .A1(n19112), .A2(n19111), .A3(n19110), .Z(n19113) );
  XOR2HSV0 U21995 ( .A1(n19114), .A2(n19113), .Z(n19115) );
  XNOR2HSV1 U21996 ( .A1(n19116), .A2(n19115), .ZN(n19117) );
  XNOR2HSV1 U21997 ( .A1(n19118), .A2(n19117), .ZN(n19120) );
  INHSV2 U21998 ( .I(n28940), .ZN(n25057) );
  CLKNAND2HSV1 U21999 ( .A1(n23041), .A2(n28586), .ZN(n19119) );
  NAND2HSV0 U22000 ( .A1(n19121), .A2(n28593), .ZN(n19122) );
  CLKNAND2HSV1 U22001 ( .A1(n19130), .A2(n19127), .ZN(n19126) );
  XNOR2HSV4 U22002 ( .A1(n19144), .A2(n19134), .ZN(n19139) );
  NOR2HSV2 U22003 ( .A1(n25519), .A2(n19138), .ZN(n19150) );
  NAND2HSV2 U22004 ( .A1(n19142), .A2(\pe6/ti_7t [15]), .ZN(n19143) );
  INHSV4 U22005 ( .I(n28925), .ZN(n23997) );
  NAND2HSV2 U22006 ( .A1(n25784), .A2(\pe6/got [6]), .ZN(n19175) );
  CLKNHSV0 U22007 ( .I(\pe6/ti_7t [13]), .ZN(n19145) );
  AOI21HSV2 U22008 ( .A1(n19145), .A2(n19147), .B(n24962), .ZN(n19146) );
  NOR2HSV4 U22009 ( .A1(n25518), .A2(n25519), .ZN(n25520) );
  NOR2HSV4 U22010 ( .A1(n25520), .A2(n19147), .ZN(n19148) );
  CLKNAND2HSV3 U22011 ( .A1(n19148), .A2(n25521), .ZN(n19154) );
  INHSV2 U22012 ( .I(n25518), .ZN(n19149) );
  CLKNAND2HSV1 U22013 ( .A1(n19151), .A2(\pe6/ti_7t [14]), .ZN(n19152) );
  NAND3HSV4 U22014 ( .A1(n19154), .A2(n19153), .A3(n19152), .ZN(n25945) );
  INHSV2 U22015 ( .I(n26014), .ZN(n26065) );
  NAND2HSV0 U22016 ( .A1(n25950), .A2(n26065), .ZN(n19174) );
  NAND2HSV4 U22017 ( .A1(n25697), .A2(n25696), .ZN(n28699) );
  INHSV2 U22018 ( .I(\pe6/got [1]), .ZN(n21766) );
  INHSV2 U22019 ( .I(n21766), .ZN(n26083) );
  NAND2HSV0 U22020 ( .A1(\pe6/aot [3]), .A2(\pe6/bq[4] ), .ZN(n19162) );
  NAND2HSV0 U22021 ( .A1(\pe6/aot [1]), .A2(\pe6/bq[6] ), .ZN(n19161) );
  XOR2HSV0 U22022 ( .A1(n19162), .A2(n19161), .Z(n19166) );
  NAND2HSV0 U22023 ( .A1(\pe6/bq[3] ), .A2(\pe6/aot [6]), .ZN(n25956) );
  CLKNAND2HSV0 U22024 ( .A1(\pe6/aot [4]), .A2(\pe6/bq[1] ), .ZN(n23704) );
  CLKNHSV0 U22025 ( .I(\pe6/aot [4]), .ZN(n19163) );
  NAND2HSV0 U22026 ( .A1(\pe6/aot [6]), .A2(\pe6/bq[1] ), .ZN(n25923) );
  OAI21HSV0 U22027 ( .A1(n19163), .A2(n25789), .B(n25923), .ZN(n19164) );
  OAI21HSV1 U22028 ( .A1(n25956), .A2(n23704), .B(n19164), .ZN(n19165) );
  XNOR2HSV1 U22029 ( .A1(n19166), .A2(n19165), .ZN(n19168) );
  CLKNAND2HSV0 U22030 ( .A1(\pe6/bq[5] ), .A2(\pe6/aot [2]), .ZN(n26043) );
  NAND2HSV0 U22031 ( .A1(\pe6/aot [5]), .A2(\pe6/bq[2] ), .ZN(n19167) );
  XOR2HSV0 U22032 ( .A1(n19170), .A2(n19169), .Z(n19171) );
  INHSV2 U22033 ( .I(\pe7/phq [1]), .ZN(n19176) );
  NAND2HSV2 U22034 ( .A1(n19177), .A2(n12289), .ZN(n19180) );
  CLKBUFHSV4 U22035 ( .I(ctro7), .Z(n19267) );
  CLKNAND2HSV2 U22036 ( .A1(n19206), .A2(n19674), .ZN(n19182) );
  INAND2HSV2 U22037 ( .A1(n19674), .B1(\pe7/ti_7t [1]), .ZN(n19181) );
  NAND2HSV4 U22038 ( .A1(n19182), .A2(n19181), .ZN(n19226) );
  INHSV2 U22039 ( .I(n19512), .ZN(n19475) );
  INHSV4 U22040 ( .I(n19183), .ZN(n25641) );
  INHSV2 U22041 ( .I(\pe7/ctrq ), .ZN(n21763) );
  INHSV3 U22042 ( .I(n21763), .ZN(n23522) );
  INHSV2 U22043 ( .I(\pe7/bq[14] ), .ZN(n25278) );
  NOR2HSV2 U22044 ( .A1(n14077), .A2(n25278), .ZN(n19187) );
  NAND2HSV0 U22045 ( .A1(\pe7/bq[15] ), .A2(\pe7/aot [15]), .ZN(n19186) );
  XOR2HSV2 U22046 ( .A1(n19187), .A2(n19186), .Z(n19213) );
  XNOR2HSV4 U22047 ( .A1(n19214), .A2(n19213), .ZN(n19235) );
  CLKNHSV0 U22048 ( .I(n19235), .ZN(n19188) );
  CLKNAND2HSV2 U22049 ( .A1(n25641), .A2(n19188), .ZN(n19239) );
  INHSV4 U22050 ( .I(n19226), .ZN(n25309) );
  BUFHSV2 U22051 ( .I(ctro7), .Z(n19262) );
  OR2HSV1 U22052 ( .A1(n19262), .A2(n19512), .Z(n19189) );
  INHSV4 U22053 ( .I(n19279), .ZN(n19526) );
  NAND2HSV2 U22054 ( .A1(n19526), .A2(n23138), .ZN(n19191) );
  INHSV2 U22055 ( .I(n19191), .ZN(n19195) );
  CLKNAND2HSV1 U22056 ( .A1(n19192), .A2(\pe7/phq [2]), .ZN(n19196) );
  CLKNAND2HSV1 U22057 ( .A1(n19194), .A2(n19196), .ZN(n19193) );
  INAND2HSV2 U22058 ( .A1(n19195), .B1(n19193), .ZN(n19202) );
  NAND3HSV2 U22059 ( .A1(n19196), .A2(n19195), .A3(n19194), .ZN(n19201) );
  NAND2HSV2 U22060 ( .A1(n19202), .A2(n19201), .ZN(n19200) );
  NAND2HSV2 U22061 ( .A1(n12688), .A2(\pe7/pvq [2]), .ZN(n19197) );
  CLKNAND2HSV2 U22062 ( .A1(n19204), .A2(n19203), .ZN(n19207) );
  INHSV2 U22063 ( .I(n19207), .ZN(n25629) );
  INHSV4 U22064 ( .I(\pe7/got [16]), .ZN(n19264) );
  AOI21HSV2 U22065 ( .A1(n28610), .A2(n19206), .B(n19466), .ZN(n19205) );
  NAND2HSV4 U22066 ( .A1(n25629), .A2(n19205), .ZN(n19256) );
  BUFHSV2 U22067 ( .I(ctro7), .Z(n19613) );
  INHSV4 U22068 ( .I(n19206), .ZN(n19253) );
  NOR2HSV4 U22069 ( .A1(n25499), .A2(n19264), .ZN(n19366) );
  INHSV2 U22070 ( .I(n19366), .ZN(n19456) );
  NOR2HSV4 U22071 ( .A1(n19253), .A2(n19456), .ZN(n19208) );
  AOI22HSV4 U22072 ( .A1(n19613), .A2(\pe7/ti_7t [2]), .B1(n19208), .B2(n19207), .ZN(n19255) );
  CLKNAND2HSV4 U22073 ( .A1(n19256), .A2(n19255), .ZN(n19263) );
  NAND2HSV4 U22074 ( .A1(n28610), .A2(n19263), .ZN(n25642) );
  INHSV2 U22075 ( .I(n19512), .ZN(n23120) );
  NOR2HSV2 U22076 ( .A1(n25642), .A2(n25339), .ZN(n19210) );
  INHSV2 U22077 ( .I(n19279), .ZN(n19365) );
  CLKAND2HSV2 U22078 ( .A1(n19282), .A2(n19365), .Z(n19209) );
  AOI21HSV2 U22079 ( .A1(n19211), .A2(n19210), .B(n19209), .ZN(n19220) );
  AND2HSV2 U22080 ( .A1(n25642), .A2(n19365), .Z(n19218) );
  XNOR2HSV4 U22081 ( .A1(n19214), .A2(n19213), .ZN(n25640) );
  INHSV2 U22082 ( .I(n19253), .ZN(n28797) );
  INHSV2 U22083 ( .I(n19262), .ZN(n19215) );
  OA21HSV4 U22084 ( .A1(n25640), .A2(n28797), .B(n19215), .Z(n19232) );
  NOR2HSV2 U22085 ( .A1(n25640), .A2(n19475), .ZN(n19216) );
  AOI21HSV4 U22086 ( .A1(n25641), .A2(n25640), .B(n19216), .ZN(n19233) );
  NAND2HSV2 U22087 ( .A1(n19232), .A2(n19233), .ZN(n19269) );
  INHSV1 U22088 ( .I(n19269), .ZN(n19217) );
  NAND2HSV2 U22089 ( .A1(n19218), .A2(n19217), .ZN(n19219) );
  NAND2HSV4 U22090 ( .A1(n19220), .A2(n19219), .ZN(n19318) );
  BUFHSV6 U22091 ( .I(n19263), .Z(n19348) );
  CLKNAND2HSV2 U22092 ( .A1(n19348), .A2(n11929), .ZN(n19230) );
  NAND2HSV0 U22093 ( .A1(\pe7/bq[12] ), .A2(\pe7/aot [16]), .ZN(n19222) );
  NAND2HSV0 U22094 ( .A1(\pe7/bq[14] ), .A2(\pe7/aot [14]), .ZN(n19221) );
  XOR2HSV0 U22095 ( .A1(n19222), .A2(n19221), .Z(n19223) );
  CLKNHSV3 U22096 ( .I(\pe7/ctrq ), .ZN(n27085) );
  INHSV4 U22097 ( .I(n27085), .ZN(n27104) );
  NAND2HSV0 U22098 ( .A1(\pe7/aot [13]), .A2(\pe7/bq[15] ), .ZN(n19224) );
  CLKNHSV2 U22099 ( .I(n19224), .ZN(n19225) );
  INHSV4 U22100 ( .I(n19226), .ZN(n19429) );
  NOR2HSV4 U22101 ( .A1(n19429), .A2(n19242), .ZN(n19227) );
  XNOR2HSV4 U22102 ( .A1(n19228), .A2(n19227), .ZN(n19229) );
  XNOR2HSV4 U22103 ( .A1(n19230), .A2(n19229), .ZN(n19317) );
  XNOR2HSV4 U22104 ( .A1(n19318), .A2(n19317), .ZN(n19376) );
  INHSV2 U22105 ( .I(n19765), .ZN(n23180) );
  INHSV2 U22106 ( .I(n19231), .ZN(n19274) );
  NAND3HSV3 U22107 ( .A1(n25642), .A2(n19233), .A3(n19232), .ZN(n19281) );
  AOI21HSV2 U22108 ( .A1(n19235), .A2(n19512), .B(n19262), .ZN(n19234) );
  NAND2HSV0 U22109 ( .A1(n25309), .A2(n19235), .ZN(n19236) );
  CLKNAND2HSV1 U22110 ( .A1(n19236), .A2(n28610), .ZN(n19237) );
  INHSV2 U22111 ( .I(n19237), .ZN(n19238) );
  NAND3HSV4 U22112 ( .A1(n19240), .A2(n19239), .A3(n19238), .ZN(n19284) );
  CLKNAND2HSV3 U22113 ( .A1(n12688), .A2(\pe7/pvq [4]), .ZN(n19241) );
  NAND2HSV0 U22114 ( .A1(\pe7/bq[13] ), .A2(\pe7/aot [16]), .ZN(n19494) );
  NAND2HSV0 U22115 ( .A1(\pe7/aot [15]), .A2(\pe7/bq[14] ), .ZN(n19245) );
  XNOR2HSV4 U22116 ( .A1(n19245), .A2(n19244), .ZN(n19251) );
  XNOR2HSV4 U22117 ( .A1(n19249), .A2(n19248), .ZN(n19250) );
  XNOR2HSV4 U22118 ( .A1(n19251), .A2(n19250), .ZN(n19254) );
  INHSV2 U22119 ( .I(ctro7), .ZN(n25494) );
  OAI21HSV1 U22120 ( .A1(n25494), .A2(\pe7/ti_7t [1]), .B(n11929), .ZN(n19252)
         );
  AOI21HSV2 U22121 ( .A1(n19256), .A2(n19255), .B(n19279), .ZN(n19258) );
  INHSV2 U22122 ( .I(n19258), .ZN(n19259) );
  NAND2HSV2 U22123 ( .A1(n19262), .A2(\pe7/ti_7t [4]), .ZN(n19358) );
  NAND2HSV4 U22124 ( .A1(n19370), .A2(n19358), .ZN(n19275) );
  CLKBUFHSV4 U22125 ( .I(ctro7), .Z(n23188) );
  NOR2HSV2 U22126 ( .A1(n28610), .A2(n23188), .ZN(n19372) );
  NAND2HSV2 U22127 ( .A1(n19270), .A2(n19269), .ZN(n19271) );
  CLKNAND2HSV2 U22128 ( .A1(n19272), .A2(n19271), .ZN(n19273) );
  INHSV4 U22129 ( .I(n23844), .ZN(n19359) );
  NAND2HSV4 U22130 ( .A1(n19273), .A2(n19359), .ZN(n19371) );
  NOR2HSV4 U22131 ( .A1(n19275), .A2(n19362), .ZN(n19308) );
  INHSV4 U22132 ( .I(n19308), .ZN(n21326) );
  NOR2HSV4 U22133 ( .A1(n19362), .A2(n19275), .ZN(n19316) );
  INHSV2 U22134 ( .I(n23188), .ZN(n28789) );
  CLKAND2HSV2 U22135 ( .A1(n19316), .A2(n28789), .Z(n19277) );
  CLKNHSV2 U22136 ( .I(n19376), .ZN(n19276) );
  NAND3HSV4 U22137 ( .A1(n19278), .A2(n19322), .A3(n19319), .ZN(n24960) );
  INHSV2 U22138 ( .I(n19279), .ZN(n28816) );
  INHSV2 U22139 ( .I(n28816), .ZN(n19684) );
  NOR2HSV4 U22140 ( .A1(n19308), .A2(n19684), .ZN(n19280) );
  INHSV4 U22141 ( .I(n19280), .ZN(n19315) );
  INHSV2 U22142 ( .I(n19281), .ZN(n19283) );
  NOR2HSV4 U22143 ( .A1(n19283), .A2(n19282), .ZN(n19328) );
  BUFHSV4 U22144 ( .I(n19284), .Z(n19327) );
  INHSV2 U22145 ( .I(n11929), .ZN(n25338) );
  AOI21HSV2 U22146 ( .A1(n19328), .A2(n19327), .B(n25338), .ZN(n19307) );
  NAND2HSV0 U22147 ( .A1(\pe7/aot [15]), .A2(\pe7/bq[12] ), .ZN(n19286) );
  NAND2HSV0 U22148 ( .A1(\pe7/aot [11]), .A2(\pe7/bq[16] ), .ZN(n19285) );
  XOR2HSV0 U22149 ( .A1(n19286), .A2(n19285), .Z(n19297) );
  INHSV2 U22150 ( .I(n19243), .ZN(n25299) );
  NAND2HSV0 U22151 ( .A1(\pe7/got [11]), .A2(n25299), .ZN(n19287) );
  XNOR2HSV4 U22152 ( .A1(n19288), .A2(n19287), .ZN(n19296) );
  NAND2HSV0 U22153 ( .A1(\pe7/aot [12]), .A2(\pe7/bq[15] ), .ZN(n19290) );
  NAND2HSV0 U22154 ( .A1(\pe7/bq[11] ), .A2(\pe7/aot [16]), .ZN(n19289) );
  XOR2HSV0 U22155 ( .A1(n19290), .A2(n19289), .Z(n19294) );
  NAND2HSV0 U22156 ( .A1(\pe7/aot [14]), .A2(\pe7/bq[13] ), .ZN(n19292) );
  NAND2HSV0 U22157 ( .A1(\pe7/bq[14] ), .A2(\pe7/aot [13]), .ZN(n19291) );
  XOR2HSV0 U22158 ( .A1(n19292), .A2(n19291), .Z(n19293) );
  XOR2HSV0 U22159 ( .A1(n19294), .A2(n19293), .Z(n19295) );
  XOR3HSV2 U22160 ( .A1(n19297), .A2(n19296), .A3(n19295), .Z(n19299) );
  NOR2HSV2 U22161 ( .A1(n19429), .A2(n24321), .ZN(n19298) );
  XNOR2HSV4 U22162 ( .A1(n19299), .A2(n19298), .ZN(n19301) );
  NAND2HSV2 U22163 ( .A1(n19348), .A2(\pe7/got [13]), .ZN(n19300) );
  XNOR2HSV4 U22164 ( .A1(n19301), .A2(n19300), .ZN(n19302) );
  INHSV2 U22165 ( .I(n19302), .ZN(n19306) );
  NOR2HSV4 U22166 ( .A1(n19302), .A2(n25338), .ZN(n19304) );
  CLKNAND2HSV1 U22167 ( .A1(n19327), .A2(n19328), .ZN(n19303) );
  CLKNAND2HSV2 U22168 ( .A1(n19304), .A2(n19303), .ZN(n19305) );
  OAI21HSV4 U22169 ( .A1(n19307), .A2(n19306), .B(n19305), .ZN(n19312) );
  NAND2HSV0 U22170 ( .A1(n19312), .A2(n19308), .ZN(n19309) );
  CLKNAND2HSV1 U22171 ( .A1(n19309), .A2(n19674), .ZN(n19310) );
  NOR2HSV2 U22172 ( .A1(n19684), .A2(n19316), .ZN(n19314) );
  INHSV4 U22173 ( .I(n19312), .ZN(n19313) );
  MUX2NHSV4 U22174 ( .I0(n19315), .I1(n19314), .S(n19313), .ZN(n24961) );
  INHSV2 U22175 ( .I(n19316), .ZN(n19739) );
  XNOR2HSV4 U22176 ( .A1(n19318), .A2(n19317), .ZN(n22091) );
  INHSV2 U22177 ( .I(n19466), .ZN(n19699) );
  NAND2HSV2 U22178 ( .A1(n19319), .A2(n19699), .ZN(n19320) );
  NAND2HSV2 U22179 ( .A1(n19765), .A2(\pe7/ti_7t [6]), .ZN(n19323) );
  OAI21HSV4 U22180 ( .A1(n24961), .A2(n19324), .B(n19323), .ZN(n19325) );
  AOI21HSV4 U22181 ( .A1(n24960), .A2(n19326), .B(n19325), .ZN(n19478) );
  INHSV4 U22182 ( .I(n19478), .ZN(n19422) );
  CLKNAND2HSV4 U22183 ( .A1(n19422), .A2(n28610), .ZN(n27215) );
  INHSV4 U22184 ( .I(n27215), .ZN(n19474) );
  NAND2HSV4 U22185 ( .A1(n19328), .A2(n19327), .ZN(n19405) );
  INHSV2 U22186 ( .I(n19242), .ZN(n24181) );
  NAND2HSV2 U22187 ( .A1(n19405), .A2(n24181), .ZN(n19351) );
  NAND2HSV2 U22188 ( .A1(\pe7/got [10]), .A2(n25299), .ZN(n19330) );
  NAND2HSV0 U22189 ( .A1(\pe7/aot [12]), .A2(\pe7/bq[14] ), .ZN(n19329) );
  XOR2HSV0 U22190 ( .A1(n19330), .A2(n19329), .Z(n19333) );
  NAND2HSV2 U22191 ( .A1(n27104), .A2(\pe7/pvq [7]), .ZN(n19331) );
  XNOR2HSV1 U22192 ( .A1(n19331), .A2(\pe7/phq [7]), .ZN(n19332) );
  XNOR2HSV4 U22193 ( .A1(n19333), .A2(n19332), .ZN(n19337) );
  NAND2HSV0 U22194 ( .A1(\pe7/aot [13]), .A2(\pe7/bq[13] ), .ZN(n19335) );
  NAND2HSV0 U22195 ( .A1(\pe7/aot [10]), .A2(n25273), .ZN(n19334) );
  XOR2HSV0 U22196 ( .A1(n19335), .A2(n19334), .Z(n19336) );
  XNOR2HSV4 U22197 ( .A1(n19337), .A2(n19336), .ZN(n19345) );
  NAND2HSV0 U22198 ( .A1(\pe7/aot [14]), .A2(\pe7/bq[12] ), .ZN(n19339) );
  NAND2HSV0 U22199 ( .A1(\pe7/aot [11]), .A2(\pe7/bq[15] ), .ZN(n19338) );
  XOR2HSV0 U22200 ( .A1(n19339), .A2(n19338), .Z(n19343) );
  NAND2HSV0 U22201 ( .A1(\pe7/aot [15]), .A2(\pe7/bq[11] ), .ZN(n19341) );
  NAND2HSV0 U22202 ( .A1(\pe7/bq[10] ), .A2(\pe7/aot [16]), .ZN(n19340) );
  XOR2HSV0 U22203 ( .A1(n19341), .A2(n19340), .Z(n19342) );
  XOR2HSV0 U22204 ( .A1(n19343), .A2(n19342), .Z(n19344) );
  XNOR2HSV4 U22205 ( .A1(n19345), .A2(n19344), .ZN(n19347) );
  INHSV2 U22206 ( .I(n19429), .ZN(\pe7/ti_7[1] ) );
  NAND2HSV2 U22207 ( .A1(\pe7/ti_7[1] ), .A2(\pe7/got [11]), .ZN(n19346) );
  XNOR2HSV4 U22208 ( .A1(n19347), .A2(n19346), .ZN(n19350) );
  BUFHSV8 U22209 ( .I(n19348), .Z(n28808) );
  NAND2HSV2 U22210 ( .A1(n28808), .A2(\pe7/got [12]), .ZN(n19349) );
  XNOR2HSV4 U22211 ( .A1(n19350), .A2(n19349), .ZN(n19352) );
  NAND2HSV2 U22212 ( .A1(n19351), .A2(n19352), .ZN(n19356) );
  INHSV2 U22213 ( .I(n19351), .ZN(n19354) );
  INHSV4 U22214 ( .I(n19352), .ZN(n19353) );
  OAI22HSV2 U22215 ( .A1(n19360), .A2(n19359), .B1(n25338), .B2(n19358), .ZN(
        n19361) );
  AOI21HSV2 U22216 ( .A1(n24271), .A2(n19362), .B(n19361), .ZN(n19363) );
  XNOR2HSV4 U22217 ( .A1(n19364), .A2(n19363), .ZN(n19379) );
  IAO21HSV4 U22218 ( .A1(n19379), .A2(n19365), .B(n19695), .ZN(n19378) );
  INHSV2 U22219 ( .I(n19379), .ZN(n27214) );
  NAND2HSV0 U22220 ( .A1(n19371), .A2(n19370), .ZN(n19367) );
  CLKNAND2HSV2 U22221 ( .A1(n19367), .A2(n19366), .ZN(n19368) );
  INHSV4 U22222 ( .I(n19369), .ZN(n19667) );
  CLKNHSV0 U22223 ( .I(n19370), .ZN(n19374) );
  NAND2HSV2 U22224 ( .A1(n19371), .A2(n19699), .ZN(n19373) );
  INHSV2 U22225 ( .I(n19372), .ZN(n19420) );
  OAI21HSV2 U22226 ( .A1(n19374), .A2(n19373), .B(n19420), .ZN(n19375) );
  CLKNAND2HSV3 U22227 ( .A1(n19376), .A2(n19375), .ZN(n19666) );
  NAND2HSV4 U22228 ( .A1(n19667), .A2(n19666), .ZN(n19507) );
  INHSV4 U22229 ( .I(n19507), .ZN(n19380) );
  CLKNAND2HSV3 U22230 ( .A1(n19378), .A2(n19377), .ZN(n19417) );
  NAND2HSV3 U22231 ( .A1(n19667), .A2(n19666), .ZN(n28657) );
  INHSV2 U22232 ( .I(n19379), .ZN(n19381) );
  NOR2HSV4 U22233 ( .A1(n27213), .A2(n19381), .ZN(n19416) );
  NOR2HSV4 U22234 ( .A1(n19417), .A2(n19416), .ZN(n19472) );
  INHSV4 U22235 ( .I(n19380), .ZN(n19529) );
  NOR2HSV4 U22236 ( .A1(n19383), .A2(n19382), .ZN(n19415) );
  CLKNAND2HSV2 U22237 ( .A1(n27215), .A2(n19415), .ZN(n19457) );
  NAND2HSV2 U22238 ( .A1(n19613), .A2(\pe7/ti_7t [7]), .ZN(n19470) );
  NAND3HSV3 U22239 ( .A1(n19458), .A2(n19457), .A3(n19470), .ZN(n19527) );
  NAND2HSV2 U22240 ( .A1(n19527), .A2(n24271), .ZN(n19460) );
  INHSV2 U22241 ( .I(n19242), .ZN(n25334) );
  NAND2HSV0 U22242 ( .A1(n25292), .A2(\pe7/got [9]), .ZN(n19408) );
  NAND2HSV0 U22243 ( .A1(\pe7/bq[9] ), .A2(\pe7/aot [14]), .ZN(n19584) );
  NAND2HSV0 U22244 ( .A1(\pe7/bq[8] ), .A2(\pe7/aot [16]), .ZN(n19491) );
  NAND2HSV0 U22245 ( .A1(\pe7/bq[7] ), .A2(\pe7/aot [15]), .ZN(n19588) );
  NOR2HSV0 U22246 ( .A1(n19491), .A2(n19588), .ZN(n19385) );
  AOI22HSV0 U22247 ( .A1(\pe7/aot [15]), .A2(\pe7/bq[8] ), .B1(n14078), .B2(
        \pe7/bq[7] ), .ZN(n19384) );
  NOR2HSV2 U22248 ( .A1(n19385), .A2(n19384), .ZN(n19389) );
  NAND2HSV0 U22249 ( .A1(n25273), .A2(\pe7/aot [7]), .ZN(n19387) );
  NAND2HSV0 U22250 ( .A1(\pe7/aot [10]), .A2(\pe7/bq[13] ), .ZN(n19386) );
  XOR2HSV0 U22251 ( .A1(n19387), .A2(n19386), .Z(n19388) );
  XOR3HSV2 U22252 ( .A1(n19584), .A2(n19389), .A3(n19388), .Z(n19404) );
  NOR2HSV2 U22253 ( .A1(n25309), .A2(n19479), .ZN(n19403) );
  NAND2HSV0 U22254 ( .A1(\pe7/aot [11]), .A2(\pe7/bq[12] ), .ZN(n19391) );
  NAND2HSV0 U22255 ( .A1(\pe7/aot [9]), .A2(\pe7/bq[14] ), .ZN(n19390) );
  XOR2HSV0 U22256 ( .A1(n19391), .A2(n19390), .Z(n19395) );
  NAND2HSV0 U22257 ( .A1(\pe7/got [7]), .A2(n25299), .ZN(n19393) );
  NAND2HSV0 U22258 ( .A1(n14050), .A2(\pe7/bq[10] ), .ZN(n19392) );
  XOR2HSV0 U22259 ( .A1(n19393), .A2(n19392), .Z(n19394) );
  XOR2HSV0 U22260 ( .A1(n19395), .A2(n19394), .Z(n19401) );
  NAND2HSV0 U22261 ( .A1(\pe7/aot [8]), .A2(\pe7/bq[15] ), .ZN(n19397) );
  NAND2HSV0 U22262 ( .A1(\pe7/aot [12]), .A2(\pe7/bq[11] ), .ZN(n19396) );
  XOR2HSV0 U22263 ( .A1(n19397), .A2(n19396), .Z(n19399) );
  CLKNHSV1 U22264 ( .I(n27085), .ZN(n27082) );
  XOR2HSV0 U22265 ( .A1(n19399), .A2(n19398), .Z(n19400) );
  XOR2HSV0 U22266 ( .A1(n19401), .A2(n19400), .Z(n19402) );
  XOR3HSV2 U22267 ( .A1(n19404), .A2(n19403), .A3(n19402), .Z(n19407) );
  NAND2HSV2 U22268 ( .A1(n28621), .A2(n24214), .ZN(n19406) );
  XOR3HSV2 U22269 ( .A1(n19408), .A2(n19407), .A3(n19406), .Z(n19410) );
  NAND2HSV0 U22270 ( .A1(n21326), .A2(\pe7/got [11]), .ZN(n19409) );
  CLKXOR2HSV2 U22271 ( .A1(n19410), .A2(n19409), .Z(n19412) );
  NAND2HSV0 U22272 ( .A1(n28657), .A2(\pe7/got [12]), .ZN(n19411) );
  INHSV4 U22273 ( .I(n19517), .ZN(n25664) );
  INHSV3 U22274 ( .I(n19415), .ZN(n19469) );
  NOR2HSV2 U22275 ( .A1(n19417), .A2(n19416), .ZN(n19418) );
  INHSV2 U22276 ( .I(n19478), .ZN(n28466) );
  OAI21HSV4 U22277 ( .A1(n19469), .A2(n19579), .B(n19419), .ZN(n19421) );
  NAND2HSV4 U22278 ( .A1(n19421), .A2(n19420), .ZN(n19462) );
  NAND2HSV2 U22279 ( .A1(n19422), .A2(n19526), .ZN(n19452) );
  INHSV2 U22280 ( .I(n19452), .ZN(n19449) );
  NAND2HSV0 U22281 ( .A1(n21326), .A2(n25334), .ZN(n19446) );
  NAND2HSV0 U22282 ( .A1(\pe7/aot [15]), .A2(\pe7/bq[10] ), .ZN(n19424) );
  NAND2HSV0 U22283 ( .A1(\pe7/aot [12]), .A2(\pe7/bq[13] ), .ZN(n19423) );
  XOR2HSV0 U22284 ( .A1(n19424), .A2(n19423), .Z(n19428) );
  NAND2HSV0 U22285 ( .A1(\pe7/bq[9] ), .A2(\pe7/aot [16]), .ZN(n19426) );
  NAND2HSV0 U22286 ( .A1(\pe7/aot [9]), .A2(n25273), .ZN(n19425) );
  XOR2HSV0 U22287 ( .A1(n19426), .A2(n19425), .Z(n19427) );
  XOR2HSV0 U22288 ( .A1(n19428), .A2(n19427), .Z(n19438) );
  INHSV2 U22289 ( .I(\pe7/got [10]), .ZN(n24084) );
  NOR2HSV2 U22290 ( .A1(n19429), .A2(n24084), .ZN(n19437) );
  CLKNHSV1 U22291 ( .I(\pe7/aot [11]), .ZN(n19492) );
  NAND2HSV0 U22292 ( .A1(\pe7/aot [13]), .A2(\pe7/bq[12] ), .ZN(n19431) );
  NAND2HSV0 U22293 ( .A1(\pe7/got [9]), .A2(n25299), .ZN(n19430) );
  XOR2HSV0 U22294 ( .A1(n19431), .A2(n19430), .Z(n19432) );
  XOR2HSV0 U22295 ( .A1(n19433), .A2(n19432), .Z(n19435) );
  INHSV2 U22296 ( .I(n12688), .ZN(n19552) );
  INHSV2 U22297 ( .I(n19552), .ZN(n27096) );
  XNOR2HSV1 U22298 ( .A1(n19435), .A2(n19434), .ZN(n19436) );
  XOR3HSV2 U22299 ( .A1(n19438), .A2(n19437), .A3(n19436), .Z(n19440) );
  NAND2HSV2 U22300 ( .A1(n28808), .A2(\pe7/got [11]), .ZN(n19439) );
  XNOR2HSV1 U22301 ( .A1(n19440), .A2(n19439), .ZN(n19441) );
  NAND3HSV2 U22302 ( .A1(n19441), .A2(n12288), .A3(\pe7/got [12]), .ZN(n19444)
         );
  INHSV2 U22303 ( .I(n12288), .ZN(n23477) );
  INHSV1 U22304 ( .I(n19441), .ZN(n19442) );
  OAI21HSV2 U22305 ( .A1(n23477), .A2(n24321), .B(n19442), .ZN(n19443) );
  CLKNAND2HSV1 U22306 ( .A1(n19444), .A2(n19443), .ZN(n19445) );
  CLKXOR2HSV4 U22307 ( .A1(n19446), .A2(n19445), .Z(n19448) );
  NAND2HSV2 U22308 ( .A1(n19507), .A2(n24271), .ZN(n19447) );
  XNOR2HSV4 U22309 ( .A1(n19448), .A2(n19447), .ZN(n19450) );
  CLKNAND2HSV2 U22310 ( .A1(n19449), .A2(n19450), .ZN(n19454) );
  INHSV2 U22311 ( .I(n19450), .ZN(n19451) );
  CLKNAND2HSV4 U22312 ( .A1(n19454), .A2(n19453), .ZN(n22089) );
  INHSV4 U22313 ( .I(n22089), .ZN(n19455) );
  AOI21HSV4 U22314 ( .A1(n19458), .A2(n19457), .B(n19456), .ZN(n19459) );
  CLKNAND2HSV1 U22315 ( .A1(n19765), .A2(\pe7/ti_7t [8]), .ZN(n27133) );
  CLKNAND2HSV4 U22316 ( .A1(n19670), .A2(n28816), .ZN(n19518) );
  NAND2HSV0 U22317 ( .A1(n19565), .A2(n22089), .ZN(n19465) );
  CLKNHSV0 U22318 ( .I(n19462), .ZN(n19463) );
  AOI21HSV1 U22319 ( .A1(n19565), .A2(n19463), .B(n19512), .ZN(n19464) );
  OAI21HSV2 U22320 ( .A1(n19467), .A2(n19515), .B(n19623), .ZN(n19468) );
  AOI21HSV2 U22321 ( .A1(n25664), .A2(n19518), .B(n19468), .ZN(n19614) );
  NAND3HSV2 U22322 ( .A1(n19469), .A2(n27215), .A3(n19470), .ZN(n19477) );
  CLKNHSV0 U22323 ( .I(n19470), .ZN(n19471) );
  NOR2HSV2 U22324 ( .A1(n19472), .A2(n19471), .ZN(n19473) );
  NAND2HSV2 U22325 ( .A1(n19474), .A2(n19473), .ZN(n19476) );
  NAND3HSV4 U22326 ( .A1(n19477), .A2(n19476), .A3(n19475), .ZN(n19567) );
  INHSV2 U22327 ( .I(n19478), .ZN(n25270) );
  NAND2HSV2 U22328 ( .A1(n28808), .A2(\pe7/got [10]), .ZN(n19504) );
  CLKNHSV1 U22329 ( .I(\pe7/aot [10]), .ZN(n24105) );
  NAND2HSV0 U22330 ( .A1(\pe7/got [8]), .A2(n25622), .ZN(n19481) );
  NAND2HSV0 U22331 ( .A1(\pe7/aot [15]), .A2(\pe7/bq[9] ), .ZN(n19480) );
  XOR2HSV0 U22332 ( .A1(n19481), .A2(n19480), .Z(n19482) );
  XOR2HSV0 U22333 ( .A1(n19483), .A2(n19482), .Z(n19501) );
  INHSV2 U22334 ( .I(\pe7/got [9]), .ZN(n24213) );
  NOR2HSV2 U22335 ( .A1(n25309), .A2(n24213), .ZN(n19500) );
  BUFHSV2 U22336 ( .I(\pe7/bq[15] ), .Z(n27083) );
  NAND2HSV0 U22337 ( .A1(\pe7/aot [9]), .A2(n27083), .ZN(n19485) );
  NAND2HSV0 U22338 ( .A1(\pe7/aot [14]), .A2(\pe7/bq[10] ), .ZN(n19484) );
  XOR2HSV0 U22339 ( .A1(n19485), .A2(n19484), .Z(n19489) );
  NAND2HSV0 U22340 ( .A1(\pe7/aot [13]), .A2(\pe7/bq[11] ), .ZN(n19487) );
  NAND2HSV0 U22341 ( .A1(\pe7/aot [12]), .A2(\pe7/bq[12] ), .ZN(n19486) );
  XOR2HSV0 U22342 ( .A1(n19487), .A2(n19486), .Z(n19488) );
  XOR2HSV0 U22343 ( .A1(n19489), .A2(n19488), .Z(n19498) );
  INHSV2 U22344 ( .I(n19552), .ZN(n27087) );
  NAND2HSV2 U22345 ( .A1(n27087), .A2(\pe7/pvq [9]), .ZN(n19490) );
  XOR2HSV0 U22346 ( .A1(n19490), .A2(\pe7/phq [9]), .Z(n19496) );
  CLKNAND2HSV0 U22347 ( .A1(\pe7/aot [11]), .A2(\pe7/bq[8] ), .ZN(n19713) );
  OAI21HSV0 U22348 ( .A1(n19713), .A2(n19494), .B(n19493), .ZN(n19495) );
  XOR2HSV0 U22349 ( .A1(n19496), .A2(n19495), .Z(n19497) );
  XNOR2HSV1 U22350 ( .A1(n19498), .A2(n19497), .ZN(n19499) );
  XOR3HSV2 U22351 ( .A1(n19501), .A2(n19500), .A3(n19499), .Z(n19503) );
  NAND2HSV2 U22352 ( .A1(n12288), .A2(\pe7/got [11]), .ZN(n19502) );
  XOR3HSV2 U22353 ( .A1(n19504), .A2(n19503), .A3(n19502), .Z(n19506) );
  NAND2HSV0 U22354 ( .A1(n21326), .A2(\pe7/got [12]), .ZN(n19505) );
  XOR2HSV2 U22355 ( .A1(n19506), .A2(n19505), .Z(n19508) );
  XOR2HSV4 U22356 ( .A1(n19567), .A2(n19566), .Z(n19510) );
  NAND2HSV2 U22357 ( .A1(n19565), .A2(n19569), .ZN(n19509) );
  XNOR2HSV4 U22358 ( .A1(n19510), .A2(n19509), .ZN(n19511) );
  NAND2HSV2 U22359 ( .A1(n25499), .A2(\pe7/ti_7t [10]), .ZN(n19678) );
  INHSV2 U22360 ( .I(n19512), .ZN(n19702) );
  INHSV2 U22361 ( .I(n19515), .ZN(n19516) );
  INHSV4 U22362 ( .I(n19519), .ZN(n19520) );
  INHSV4 U22363 ( .I(n19522), .ZN(n19525) );
  NAND2HSV2 U22364 ( .A1(n19215), .A2(n19523), .ZN(n19524) );
  NOR2HSV8 U22365 ( .A1(n19525), .A2(n19524), .ZN(n19615) );
  INHSV2 U22366 ( .I(n19527), .ZN(n19528) );
  INHSV4 U22367 ( .I(n19528), .ZN(n19711) );
  INHSV2 U22368 ( .I(\pe7/got [10]), .ZN(n19710) );
  CLKBUFHSV4 U22369 ( .I(n28621), .Z(n24250) );
  NAND2HSV0 U22370 ( .A1(n24250), .A2(\pe7/got [8]), .ZN(n19530) );
  XNOR2HSV4 U22371 ( .A1(n19531), .A2(n19530), .ZN(n19564) );
  NAND2HSV0 U22372 ( .A1(n21326), .A2(\pe7/got [9]), .ZN(n19562) );
  NAND2HSV0 U22373 ( .A1(n11858), .A2(\pe7/got [6]), .ZN(n19560) );
  BUFHSV2 U22374 ( .I(\pe7/got [7]), .Z(n25271) );
  NAND2HSV0 U22375 ( .A1(n28808), .A2(n25271), .ZN(n19559) );
  NAND2HSV0 U22376 ( .A1(\pe7/aot [9]), .A2(\pe7/bq[12] ), .ZN(n19534) );
  NAND2HSV0 U22377 ( .A1(\pe7/aot [6]), .A2(\pe7/bq[15] ), .ZN(n19533) );
  XOR2HSV0 U22378 ( .A1(n19534), .A2(n19533), .Z(n19538) );
  NAND2HSV0 U22379 ( .A1(\pe7/aot [5]), .A2(n25273), .ZN(n19536) );
  NAND2HSV0 U22380 ( .A1(\pe7/aot [12]), .A2(\pe7/bq[9] ), .ZN(n19535) );
  XOR2HSV0 U22381 ( .A1(n19536), .A2(n19535), .Z(n19537) );
  XOR2HSV0 U22382 ( .A1(n19538), .A2(n19537), .Z(n19545) );
  NAND2HSV0 U22383 ( .A1(\pe7/got [5]), .A2(n25299), .ZN(n19540) );
  NAND2HSV0 U22384 ( .A1(\pe7/aot [15]), .A2(\pe7/bq[6] ), .ZN(n19539) );
  XOR2HSV0 U22385 ( .A1(n19540), .A2(n19539), .Z(n19543) );
  NAND2HSV0 U22386 ( .A1(n14050), .A2(\pe7/bq[8] ), .ZN(n19585) );
  NAND2HSV0 U22387 ( .A1(\pe7/aot [10]), .A2(\pe7/bq[11] ), .ZN(n19541) );
  XOR2HSV0 U22388 ( .A1(n19585), .A2(n19541), .Z(n19542) );
  XOR2HSV0 U22389 ( .A1(n19543), .A2(n19542), .Z(n19544) );
  XOR2HSV0 U22390 ( .A1(n19545), .A2(n19544), .Z(n19557) );
  NAND2HSV0 U22391 ( .A1(\pe7/bq[7] ), .A2(\pe7/aot [14]), .ZN(n19547) );
  NAND2HSV0 U22392 ( .A1(\pe7/aot [8]), .A2(\pe7/bq[13] ), .ZN(n19546) );
  XOR2HSV0 U22393 ( .A1(n19547), .A2(n19546), .Z(n19551) );
  NAND2HSV0 U22394 ( .A1(\pe7/aot [7]), .A2(\pe7/bq[14] ), .ZN(n19549) );
  NAND2HSV0 U22395 ( .A1(\pe7/aot [11]), .A2(\pe7/bq[10] ), .ZN(n19548) );
  XOR2HSV0 U22396 ( .A1(n19549), .A2(n19548), .Z(n19550) );
  XOR2HSV0 U22397 ( .A1(n19551), .A2(n19550), .Z(n19555) );
  INHSV2 U22398 ( .I(n19552), .ZN(n27099) );
  CLKNHSV0 U22399 ( .I(\pe7/bq[5] ), .ZN(n27097) );
  NOR2HSV1 U22400 ( .A1(n11855), .A2(n27097), .ZN(n19651) );
  XNOR2HSV1 U22401 ( .A1(n19553), .A2(n19651), .ZN(n19554) );
  XNOR2HSV1 U22402 ( .A1(n19555), .A2(n19554), .ZN(n19556) );
  XNOR2HSV1 U22403 ( .A1(n19557), .A2(n19556), .ZN(n19558) );
  XOR3HSV1 U22404 ( .A1(n19560), .A2(n19559), .A3(n19558), .Z(n19561) );
  XNOR2HSV1 U22405 ( .A1(n19562), .A2(n19561), .ZN(n19563) );
  INHSV2 U22406 ( .I(n19570), .ZN(n27132) );
  NAND2HSV2 U22407 ( .A1(n27132), .A2(n23180), .ZN(n19568) );
  XNOR2HSV4 U22408 ( .A1(n19567), .A2(n19566), .ZN(n27135) );
  NOR2HSV4 U22409 ( .A1(n19568), .A2(n27135), .ZN(n19575) );
  OAI21HSV4 U22410 ( .A1(n19571), .A2(n19570), .B(n27135), .ZN(n19573) );
  CLKNAND2HSV1 U22411 ( .A1(n19613), .A2(\pe7/ti_7t [9]), .ZN(n19572) );
  NAND2HSV2 U22412 ( .A1(n19711), .A2(n24181), .ZN(n19609) );
  CLKNAND2HSV1 U22413 ( .A1(n27082), .A2(\pe7/pvq [11]), .ZN(n19580) );
  XNOR2HSV1 U22414 ( .A1(n19580), .A2(\pe7/phq [11]), .ZN(n19587) );
  CLKNHSV0 U22415 ( .I(\pe7/aot [14]), .ZN(n19582) );
  CLKNHSV0 U22416 ( .I(\pe7/bq[8] ), .ZN(n23497) );
  NAND2HSV0 U22417 ( .A1(n14050), .A2(\pe7/bq[9] ), .ZN(n19581) );
  OAI21HSV1 U22418 ( .A1(n19582), .A2(n23497), .B(n19581), .ZN(n19583) );
  OAI21HSV1 U22419 ( .A1(n19585), .A2(n19584), .B(n19583), .ZN(n19586) );
  XNOR2HSV1 U22420 ( .A1(n19587), .A2(n19586), .ZN(n19590) );
  NAND2HSV0 U22421 ( .A1(\pe7/aot [11]), .A2(\pe7/bq[11] ), .ZN(n24241) );
  XOR2HSV0 U22422 ( .A1(n19588), .A2(n24241), .Z(n19589) );
  NAND2HSV0 U22423 ( .A1(\pe7/got [6]), .A2(n23138), .ZN(n19592) );
  NAND2HSV0 U22424 ( .A1(\pe7/aot [9]), .A2(\pe7/bq[13] ), .ZN(n19591) );
  XOR2HSV0 U22425 ( .A1(n19592), .A2(n19591), .Z(n19596) );
  NAND2HSV0 U22426 ( .A1(\pe7/aot [10]), .A2(\pe7/bq[12] ), .ZN(n19594) );
  NAND2HSV0 U22427 ( .A1(\pe7/aot [8]), .A2(\pe7/bq[14] ), .ZN(n19593) );
  XOR2HSV0 U22428 ( .A1(n19594), .A2(n19593), .Z(n19595) );
  XOR2HSV0 U22429 ( .A1(n19596), .A2(n19595), .Z(n19604) );
  NAND2HSV0 U22430 ( .A1(\pe7/bq[6] ), .A2(\pe7/aot [16]), .ZN(n19598) );
  NAND2HSV0 U22431 ( .A1(\pe7/aot [6]), .A2(n25273), .ZN(n19597) );
  XOR2HSV0 U22432 ( .A1(n19598), .A2(n19597), .Z(n19602) );
  NAND2HSV0 U22433 ( .A1(\pe7/aot [7]), .A2(n27083), .ZN(n19600) );
  NAND2HSV0 U22434 ( .A1(\pe7/aot [12]), .A2(\pe7/bq[10] ), .ZN(n19599) );
  XOR2HSV0 U22435 ( .A1(n19600), .A2(n19599), .Z(n19601) );
  XOR2HSV0 U22436 ( .A1(n19602), .A2(n19601), .Z(n19603) );
  NAND2HSV2 U22437 ( .A1(n28657), .A2(n14022), .ZN(n19605) );
  XOR2HSV0 U22438 ( .A1(n19606), .A2(n19605), .Z(n19607) );
  CLKNHSV2 U22439 ( .I(n19671), .ZN(n23901) );
  CLKNAND2HSV3 U22440 ( .A1(n19614), .A2(n25665), .ZN(n19679) );
  NAND2HSV2 U22441 ( .A1(n25673), .A2(n23901), .ZN(n19703) );
  INHSV2 U22442 ( .I(\pe7/ti_7t [11]), .ZN(n19689) );
  AOI21HSV1 U22443 ( .A1(n19689), .A2(n19695), .B(n27134), .ZN(n25344) );
  CLKNHSV0 U22444 ( .I(n25344), .ZN(n19621) );
  NOR2HSV1 U22445 ( .A1(n19621), .A2(n23188), .ZN(n19622) );
  CLKNAND2HSV4 U22446 ( .A1(n19693), .A2(n19692), .ZN(n23111) );
  NOR2HSV2 U22447 ( .A1(n25347), .A2(n19695), .ZN(n19628) );
  INHSV2 U22448 ( .I(n19696), .ZN(n19694) );
  CLKNHSV1 U22449 ( .I(n19694), .ZN(n19627) );
  INHSV2 U22450 ( .I(n25346), .ZN(n19626) );
  AND2HSV2 U22451 ( .A1(n19694), .A2(n25344), .Z(n19624) );
  CLKNAND2HSV2 U22452 ( .A1(n25345), .A2(n19624), .ZN(n19625) );
  OAI22HSV4 U22453 ( .A1(n19628), .A2(n19627), .B1(n19626), .B2(n19625), .ZN(
        n19759) );
  NAND2HSV4 U22454 ( .A1(n23111), .A2(n19759), .ZN(n23210) );
  CLKNHSV0 U22455 ( .I(n23210), .ZN(n25495) );
  BUFHSV2 U22456 ( .I(\pe7/got [5]), .Z(n25375) );
  NAND2HSV0 U22457 ( .A1(n11858), .A2(n25375), .ZN(n19661) );
  NAND2HSV0 U22458 ( .A1(n25292), .A2(\pe7/got [6]), .ZN(n19660) );
  INHSV2 U22459 ( .I(\pe7/got [4]), .ZN(n23839) );
  NAND2HSV0 U22460 ( .A1(\pe7/got [4]), .A2(n23138), .ZN(n19630) );
  NAND2HSV0 U22461 ( .A1(\pe7/aot [7]), .A2(\pe7/bq[13] ), .ZN(n19629) );
  XOR2HSV0 U22462 ( .A1(n19630), .A2(n19629), .Z(n19634) );
  NAND2HSV0 U22463 ( .A1(n14050), .A2(\pe7/bq[7] ), .ZN(n19632) );
  NAND2HSV0 U22464 ( .A1(\pe7/aot [6]), .A2(\pe7/bq[14] ), .ZN(n19631) );
  XOR2HSV0 U22465 ( .A1(n19632), .A2(n19631), .Z(n19633) );
  XOR2HSV0 U22466 ( .A1(n19634), .A2(n19633), .Z(n19641) );
  NAND2HSV0 U22467 ( .A1(\pe7/aot [9]), .A2(\pe7/bq[11] ), .ZN(n19636) );
  NAND2HSV0 U22468 ( .A1(\pe7/aot [12]), .A2(\pe7/bq[8] ), .ZN(n19635) );
  XOR2HSV0 U22469 ( .A1(n19636), .A2(n19635), .Z(n19639) );
  NAND2HSV0 U22470 ( .A1(\pe7/bq[6] ), .A2(\pe7/aot [14]), .ZN(n25280) );
  NAND2HSV0 U22471 ( .A1(\pe7/aot [11]), .A2(\pe7/bq[9] ), .ZN(n19637) );
  XOR2HSV0 U22472 ( .A1(n25280), .A2(n19637), .Z(n19638) );
  XOR2HSV0 U22473 ( .A1(n19639), .A2(n19638), .Z(n19640) );
  XOR2HSV0 U22474 ( .A1(n19641), .A2(n19640), .Z(n19658) );
  NAND2HSV0 U22475 ( .A1(\pe7/aot [5]), .A2(n27083), .ZN(n19643) );
  NAND2HSV0 U22476 ( .A1(\pe7/aot [8]), .A2(\pe7/bq[12] ), .ZN(n19642) );
  XOR2HSV0 U22477 ( .A1(n19643), .A2(n19642), .Z(n19647) );
  NAND2HSV0 U22478 ( .A1(\pe7/aot [10]), .A2(\pe7/bq[10] ), .ZN(n19645) );
  NAND2HSV0 U22479 ( .A1(\pe7/aot [4]), .A2(n25273), .ZN(n19644) );
  XNOR2HSV1 U22480 ( .A1(n19645), .A2(n19644), .ZN(n19646) );
  XNOR2HSV1 U22481 ( .A1(n19647), .A2(n19646), .ZN(n19656) );
  NAND2HSV0 U22482 ( .A1(n27087), .A2(\pe7/pvq [13]), .ZN(n19648) );
  XOR2HSV0 U22483 ( .A1(n19648), .A2(\pe7/phq [13]), .Z(n19654) );
  CLKNAND2HSV0 U22484 ( .A1(n14078), .A2(\pe7/bq[4] ), .ZN(n23125) );
  NAND2HSV0 U22485 ( .A1(\pe7/aot [15]), .A2(\pe7/bq[5] ), .ZN(n19652) );
  CLKNHSV0 U22486 ( .I(\pe7/aot [15]), .ZN(n19650) );
  NOR2HSV2 U22487 ( .A1(n19650), .A2(n19649), .ZN(n19714) );
  AOI22HSV1 U22488 ( .A1(n23125), .A2(n19652), .B1(n19651), .B2(n19714), .ZN(
        n19653) );
  XOR2HSV0 U22489 ( .A1(n19654), .A2(n19653), .Z(n19655) );
  XNOR2HSV1 U22490 ( .A1(n19656), .A2(n19655), .ZN(n19657) );
  XNOR2HSV1 U22491 ( .A1(n19658), .A2(n19657), .ZN(n19659) );
  XOR3HSV2 U22492 ( .A1(n19661), .A2(n19660), .A3(n19659), .Z(n19663) );
  NAND2HSV0 U22493 ( .A1(n24250), .A2(n25271), .ZN(n19662) );
  XNOR2HSV1 U22494 ( .A1(n19663), .A2(n19662), .ZN(n19665) );
  NAND2HSV0 U22495 ( .A1(n11936), .A2(\pe7/got [8]), .ZN(n19664) );
  XOR2HSV0 U22496 ( .A1(n19665), .A2(n19664), .Z(n19669) );
  NAND2HSV4 U22497 ( .A1(n19667), .A2(n19666), .ZN(n25318) );
  NAND2HSV0 U22498 ( .A1(n25318), .A2(\pe7/got [9]), .ZN(n19668) );
  INHSV4 U22499 ( .I(n19670), .ZN(n19709) );
  INHSV4 U22500 ( .I(n19709), .ZN(n28587) );
  CLKBUFHSV4 U22501 ( .I(n19671), .Z(n28430) );
  NAND2HSV2 U22502 ( .A1(n28430), .A2(n24181), .ZN(n19672) );
  NOR2HSV2 U22503 ( .A1(n19677), .A2(n19706), .ZN(n19681) );
  CLKNHSV0 U22504 ( .I(n19688), .ZN(n19680) );
  INHSV2 U22505 ( .I(n19703), .ZN(n19685) );
  NOR2HSV2 U22506 ( .A1(n19685), .A2(n19684), .ZN(n19686) );
  NAND2HSV2 U22507 ( .A1(n19704), .A2(n19686), .ZN(n19687) );
  CLKNHSV2 U22508 ( .I(n19687), .ZN(n19691) );
  NOR2HSV2 U22509 ( .A1(n19215), .A2(n19689), .ZN(n19707) );
  INOR2HSV1 U22510 ( .A1(n25344), .B1(n19696), .ZN(n19697) );
  AND2HSV2 U22511 ( .A1(n25496), .A2(n19699), .Z(n19700) );
  CLKNAND2HSV2 U22512 ( .A1(n25498), .A2(n19700), .ZN(n19701) );
  AOI21HSV2 U22513 ( .A1(n25495), .A2(n23116), .B(n19701), .ZN(n19757) );
  NAND2HSV4 U22514 ( .A1(n28926), .A2(n19702), .ZN(n19764) );
  INHSV4 U22515 ( .I(n19708), .ZN(n25377) );
  INHSV4 U22516 ( .I(n19709), .ZN(n25325) );
  NAND2HSV2 U22517 ( .A1(n25325), .A2(n14022), .ZN(n19749) );
  NAND2HSV0 U22518 ( .A1(n19711), .A2(\pe7/got [10]), .ZN(n19747) );
  NAND2HSV0 U22519 ( .A1(\pe7/got [9]), .A2(n28466), .ZN(n19745) );
  NAND2HSV0 U22520 ( .A1(\pe7/aot [10]), .A2(\pe7/bq[9] ), .ZN(n19712) );
  XOR2HSV0 U22521 ( .A1(n19713), .A2(n19712), .Z(n19723) );
  NAND2HSV0 U22522 ( .A1(\pe7/aot [5]), .A2(\pe7/bq[14] ), .ZN(n19716) );
  NAND2HSV0 U22523 ( .A1(\pe7/aot [4]), .A2(\pe7/bq[15] ), .ZN(n19715) );
  XOR2HSV0 U22524 ( .A1(n19716), .A2(n19715), .Z(n19720) );
  NAND2HSV0 U22525 ( .A1(n14050), .A2(\pe7/bq[6] ), .ZN(n19718) );
  NAND2HSV0 U22526 ( .A1(\pe7/aot [9]), .A2(\pe7/bq[10] ), .ZN(n19717) );
  XOR2HSV0 U22527 ( .A1(n19718), .A2(n19717), .Z(n19719) );
  XOR2HSV0 U22528 ( .A1(n19720), .A2(n19719), .Z(n19721) );
  NAND2HSV0 U22529 ( .A1(\pe7/bq[5] ), .A2(\pe7/aot [14]), .ZN(n19725) );
  NAND2HSV0 U22530 ( .A1(\pe7/aot [7]), .A2(\pe7/bq[12] ), .ZN(n19724) );
  XOR2HSV0 U22531 ( .A1(n19725), .A2(n19724), .Z(n19729) );
  NAND2HSV0 U22532 ( .A1(n14078), .A2(\pe7/bq[3] ), .ZN(n19727) );
  NAND2HSV0 U22533 ( .A1(\pe7/aot [8]), .A2(\pe7/bq[11] ), .ZN(n19726) );
  XOR2HSV0 U22534 ( .A1(n19727), .A2(n19726), .Z(n19728) );
  XOR2HSV0 U22535 ( .A1(n19729), .A2(n19728), .Z(n19737) );
  NAND2HSV0 U22536 ( .A1(\pe7/aot [3]), .A2(n25273), .ZN(n19731) );
  NAND2HSV0 U22537 ( .A1(\pe7/aot [12]), .A2(\pe7/bq[7] ), .ZN(n19730) );
  XOR2HSV0 U22538 ( .A1(n19731), .A2(n19730), .Z(n19735) );
  NAND2HSV0 U22539 ( .A1(\pe7/got [3]), .A2(n25299), .ZN(n19733) );
  NAND2HSV0 U22540 ( .A1(\pe7/aot [6]), .A2(\pe7/bq[13] ), .ZN(n19732) );
  XOR2HSV0 U22541 ( .A1(n19733), .A2(n19732), .Z(n19734) );
  XOR2HSV0 U22542 ( .A1(n19735), .A2(n19734), .Z(n19736) );
  NAND2HSV0 U22543 ( .A1(\pe7/ti_7[1] ), .A2(n25272), .ZN(n19738) );
  NAND2HSV0 U22544 ( .A1(n19739), .A2(n25271), .ZN(n19740) );
  XNOR2HSV1 U22545 ( .A1(n19741), .A2(n19740), .ZN(n19743) );
  NAND2HSV0 U22546 ( .A1(n25318), .A2(\pe7/got [8]), .ZN(n19742) );
  XOR2HSV0 U22547 ( .A1(n19743), .A2(n19742), .Z(n19744) );
  XOR2HSV0 U22548 ( .A1(n19745), .A2(n19744), .Z(n19746) );
  XNOR2HSV1 U22549 ( .A1(n19749), .A2(n19748), .ZN(n19751) );
  XNOR2HSV2 U22550 ( .A1(n19751), .A2(n19750), .ZN(n19752) );
  XNOR2HSV4 U22551 ( .A1(n19753), .A2(n19752), .ZN(n19754) );
  XOR2HSV2 U22552 ( .A1(n19764), .A2(n19763), .Z(n19756) );
  NAND2HSV4 U22553 ( .A1(n19757), .A2(n19756), .ZN(n24075) );
  NAND2HSV2 U22554 ( .A1(n23210), .A2(n25496), .ZN(n19758) );
  OAI21HSV2 U22555 ( .A1(n19758), .A2(n23115), .B(n28789), .ZN(n19762) );
  NAND3HSV2 U22556 ( .A1(n23111), .A2(n19759), .A3(n25496), .ZN(n19760) );
  NOR2HSV2 U22557 ( .A1(n23116), .A2(n19760), .ZN(n19761) );
  NOR2HSV4 U22558 ( .A1(n19762), .A2(n19761), .ZN(n23108) );
  XNOR2HSV4 U22559 ( .A1(n19764), .A2(n19763), .ZN(n25500) );
  NAND2HSV4 U22560 ( .A1(n23108), .A2(n25500), .ZN(n24074) );
  CLKNAND2HSV1 U22561 ( .A1(n19765), .A2(\pe7/ti_7t [14]), .ZN(n24073) );
  INHSV2 U22562 ( .I(n19766), .ZN(n28368) );
  NOR2HSV2 U22563 ( .A1(n28368), .A2(n28067), .ZN(n19807) );
  CLKNAND2HSV0 U22564 ( .A1(n28317), .A2(\pe9/got [8]), .ZN(n19805) );
  INHSV2 U22565 ( .I(n19767), .ZN(n22374) );
  NAND2HSV0 U22566 ( .A1(n28437), .A2(\pe9/got [7]), .ZN(n19803) );
  NAND2HSV0 U22567 ( .A1(n28264), .A2(n28643), .ZN(n19799) );
  NAND2HSV0 U22568 ( .A1(n22375), .A2(\pe9/got [2]), .ZN(n19793) );
  NAND2HSV0 U22569 ( .A1(\pe9/got [1]), .A2(n28804), .ZN(n19791) );
  NAND2HSV0 U22570 ( .A1(\pe9/aot [11]), .A2(\pe9/bq[3] ), .ZN(n19771) );
  NAND2HSV0 U22571 ( .A1(\pe9/aot [6]), .A2(\pe9/bq[8] ), .ZN(n19770) );
  XOR2HSV0 U22572 ( .A1(n19771), .A2(n19770), .Z(n19775) );
  NAND2HSV0 U22573 ( .A1(\pe9/aot [3]), .A2(\pe9/bq[11] ), .ZN(n19773) );
  NAND2HSV0 U22574 ( .A1(\pe9/aot [8]), .A2(\pe9/bq[6] ), .ZN(n19772) );
  XOR2HSV0 U22575 ( .A1(n19773), .A2(n19772), .Z(n19774) );
  XOR2HSV0 U22576 ( .A1(n19775), .A2(n19774), .Z(n19782) );
  NAND2HSV0 U22577 ( .A1(\pe9/aot [10]), .A2(\pe9/bq[4] ), .ZN(n19777) );
  NAND2HSV0 U22578 ( .A1(\pe9/aot [7]), .A2(\pe9/bq[7] ), .ZN(n19776) );
  XOR2HSV0 U22579 ( .A1(n19777), .A2(n19776), .Z(n19780) );
  NAND2HSV0 U22580 ( .A1(\pe9/aot [9]), .A2(\pe9/bq[1] ), .ZN(n28265) );
  AO22HSV2 U22581 ( .A1(\pe9/bq[1] ), .A2(\pe9/aot [13]), .B1(\pe9/aot [9]), 
        .B2(\pe9/bq[5] ), .Z(n19778) );
  OAI21HSV0 U22582 ( .A1(n22382), .A2(n28265), .B(n19778), .ZN(n19779) );
  XNOR2HSV1 U22583 ( .A1(n19780), .A2(n19779), .ZN(n19781) );
  XNOR2HSV1 U22584 ( .A1(n19782), .A2(n19781), .ZN(n19789) );
  NAND2HSV0 U22585 ( .A1(\pe9/aot [1]), .A2(\pe9/bq[13] ), .ZN(n22379) );
  CLKNHSV0 U22586 ( .I(\pe9/aot [5]), .ZN(n28200) );
  NOR2HSV0 U22587 ( .A1(n28200), .A2(n27101), .ZN(n28041) );
  INHSV2 U22588 ( .I(\pe9/aot [2]), .ZN(n28398) );
  INHSV2 U22589 ( .I(\pe9/bq[9] ), .ZN(n28266) );
  NOR2HSV0 U22590 ( .A1(n28398), .A2(n28266), .ZN(n28191) );
  AOI22HSV0 U22591 ( .A1(\pe9/aot [5]), .A2(\pe9/bq[9] ), .B1(\pe9/bq[12] ), 
        .B2(\pe9/aot [2]), .ZN(n19783) );
  AOI21HSV2 U22592 ( .A1(n28041), .A2(n28191), .B(n19783), .ZN(n19787) );
  NAND2HSV0 U22593 ( .A1(\pe9/aot [12]), .A2(\pe9/bq[2] ), .ZN(n19785) );
  NAND2HSV0 U22594 ( .A1(\pe9/aot [4]), .A2(\pe9/bq[10] ), .ZN(n19784) );
  XOR2HSV0 U22595 ( .A1(n19785), .A2(n19784), .Z(n19786) );
  XOR3HSV2 U22596 ( .A1(n22379), .A2(n19787), .A3(n19786), .Z(n19788) );
  XNOR2HSV1 U22597 ( .A1(n19789), .A2(n19788), .ZN(n19790) );
  XNOR2HSV1 U22598 ( .A1(n19791), .A2(n19790), .ZN(n19792) );
  XNOR2HSV1 U22599 ( .A1(n19793), .A2(n19792), .ZN(n19797) );
  CLKNAND2HSV0 U22600 ( .A1(n28189), .A2(n28389), .ZN(n19796) );
  NAND2HSV0 U22601 ( .A1(n28638), .A2(\pe9/got [3]), .ZN(n19795) );
  XOR3HSV2 U22602 ( .A1(n19797), .A2(n19796), .A3(n19795), .Z(n19798) );
  XNOR2HSV1 U22603 ( .A1(n19799), .A2(n19798), .ZN(n19801) );
  CLKNHSV2 U22604 ( .I(n28790), .ZN(n28214) );
  OR2HSV1 U22605 ( .A1(n28214), .A2(n28188), .Z(n19800) );
  XNOR2HSV1 U22606 ( .A1(n19801), .A2(n19800), .ZN(n19802) );
  XNOR2HSV1 U22607 ( .A1(n19803), .A2(n19802), .ZN(n19804) );
  XNOR2HSV1 U22608 ( .A1(n19805), .A2(n19804), .ZN(n19806) );
  XOR2HSV2 U22609 ( .A1(n19807), .A2(n19806), .Z(n19811) );
  NAND2HSV4 U22610 ( .A1(n19809), .A2(n18463), .ZN(n28580) );
  NAND2HSV0 U22611 ( .A1(n28580), .A2(n28227), .ZN(n19810) );
  XOR2HSV0 U22612 ( .A1(n19811), .A2(n19810), .Z(n19813) );
  CLKNAND2HSV0 U22613 ( .A1(n28394), .A2(n28423), .ZN(n19812) );
  INAND2HSV4 U22614 ( .A1(n19814), .B1(n12268), .ZN(n23243) );
  INHSV4 U22615 ( .I(n28140), .ZN(n28080) );
  INHSV4 U22616 ( .I(n28080), .ZN(n28404) );
  INHSV2 U22617 ( .I(n28340), .ZN(n28184) );
  INHSV2 U22618 ( .I(n28184), .ZN(n28412) );
  NAND3HSV2 U22619 ( .A1(n28404), .A2(n28134), .A3(n28412), .ZN(n19819) );
  NOR2HSV0 U22620 ( .A1(n20058), .A2(n18773), .ZN(n19945) );
  NOR2HSV0 U22621 ( .A1(n28667), .A2(n25602), .ZN(n19821) );
  AOI22HSV0 U22622 ( .A1(n19940), .A2(n19822), .B1(n19945), .B2(n19821), .ZN(
        n19823) );
  OR2HSV1 U22623 ( .A1(n19900), .A2(n19823), .Z(n19829) );
  NOR2HSV2 U22624 ( .A1(n22129), .A2(\pe8/ti_7t [12]), .ZN(n19988) );
  NAND3HSV0 U22625 ( .A1(n22138), .A2(n13998), .A3(\pe8/ti_7t [12]), .ZN(
        n19824) );
  CLKNHSV2 U22626 ( .I(n19824), .ZN(n19825) );
  CLKNHSV2 U22627 ( .I(n19826), .ZN(n19827) );
  NOR2HSV0 U22628 ( .A1(n19940), .A2(n19835), .ZN(n19836) );
  CLKNHSV0 U22629 ( .I(n19836), .ZN(n19837) );
  INHSV2 U22630 ( .I(n19945), .ZN(n19953) );
  CLKNHSV1 U22631 ( .I(n19953), .ZN(n19838) );
  CLKNAND2HSV1 U22632 ( .A1(n21322), .A2(\pe8/got [12]), .ZN(n19893) );
  INHSV4 U22633 ( .I(n22081), .ZN(n22140) );
  NAND2HSV2 U22634 ( .A1(n22140), .A2(\pe8/got [11]), .ZN(n19891) );
  INHSV2 U22635 ( .I(n22141), .ZN(n25528) );
  NOR2HSV2 U22636 ( .A1(n25528), .A2(n19841), .ZN(n19889) );
  CLKNAND2HSV0 U22637 ( .A1(n28462), .A2(n23605), .ZN(n19882) );
  NAND2HSV0 U22638 ( .A1(n20009), .A2(\pe8/got [5]), .ZN(n19859) );
  NAND2HSV0 U22639 ( .A1(\pe8/aot [5]), .A2(\pe8/bq[14] ), .ZN(n19843) );
  NAND2HSV0 U22640 ( .A1(\pe8/bq[6] ), .A2(\pe8/aot [13]), .ZN(n19842) );
  XOR2HSV0 U22641 ( .A1(n19843), .A2(n19842), .Z(n19857) );
  NAND2HSV0 U22642 ( .A1(\pe8/aot [14]), .A2(\pe8/bq[3] ), .ZN(n25554) );
  NAND2HSV0 U22643 ( .A1(n28627), .A2(\pe8/bq[3] ), .ZN(n19844) );
  OAI21HSV0 U22644 ( .A1(n19845), .A2(n23847), .B(n19844), .ZN(n19846) );
  OAI21HSV2 U22645 ( .A1(n25554), .A2(n19847), .B(n19846), .ZN(n19848) );
  NAND2HSV0 U22646 ( .A1(\pe8/aot [12]), .A2(\pe8/bq[7] ), .ZN(n25560) );
  XNOR2HSV1 U22647 ( .A1(n19848), .A2(n25560), .ZN(n19856) );
  NAND2HSV0 U22648 ( .A1(\pe8/bq[4] ), .A2(\pe8/aot [15]), .ZN(n19850) );
  NAND2HSV0 U22649 ( .A1(\pe8/aot [6]), .A2(n25565), .ZN(n19849) );
  XOR2HSV0 U22650 ( .A1(n19850), .A2(n19849), .Z(n19854) );
  NAND2HSV0 U22651 ( .A1(\pe8/aot [7]), .A2(\pe8/bq[12] ), .ZN(n19852) );
  NAND2HSV0 U22652 ( .A1(\pe8/got [3]), .A2(n25624), .ZN(n19851) );
  XOR2HSV0 U22653 ( .A1(n19852), .A2(n19851), .Z(n19853) );
  XOR2HSV0 U22654 ( .A1(n19854), .A2(n19853), .Z(n19855) );
  XOR3HSV2 U22655 ( .A1(n19857), .A2(n19856), .A3(n19855), .Z(n19858) );
  XNOR2HSV1 U22656 ( .A1(n19859), .A2(n19858), .ZN(n19876) );
  NAND2HSV0 U22657 ( .A1(\pe8/aot [4]), .A2(n25532), .ZN(n19861) );
  NAND2HSV0 U22658 ( .A1(\pe8/aot [8]), .A2(\pe8/bq[11] ), .ZN(n19860) );
  XOR2HSV0 U22659 ( .A1(n19861), .A2(n19860), .Z(n19865) );
  NAND2HSV0 U22660 ( .A1(\pe8/aot [9]), .A2(\pe8/bq[10] ), .ZN(n19863) );
  NAND2HSV0 U22661 ( .A1(\pe8/aot [3]), .A2(n25539), .ZN(n19862) );
  XOR2HSV0 U22662 ( .A1(n19863), .A2(n19862), .Z(n19864) );
  XOR2HSV0 U22663 ( .A1(n19865), .A2(n19864), .Z(n19872) );
  NAND2HSV0 U22664 ( .A1(\pe8/aot [11]), .A2(\pe8/bq[8] ), .ZN(n19867) );
  NAND2HSV0 U22665 ( .A1(\pe8/aot [10]), .A2(\pe8/bq[9] ), .ZN(n19866) );
  XOR2HSV0 U22666 ( .A1(n19867), .A2(n19866), .Z(n19870) );
  NAND2HSV0 U22667 ( .A1(n14036), .A2(\pe8/pvq [14]), .ZN(n19868) );
  XOR2HSV0 U22668 ( .A1(n19868), .A2(\pe8/phq [14]), .Z(n19869) );
  XOR2HSV0 U22669 ( .A1(n19870), .A2(n19869), .Z(n19871) );
  XOR2HSV0 U22670 ( .A1(n19872), .A2(n19871), .Z(n19874) );
  NOR2HSV0 U22671 ( .A1(n27225), .A2(n22230), .ZN(n19873) );
  XNOR2HSV1 U22672 ( .A1(n19874), .A2(n19873), .ZN(n19875) );
  XNOR2HSV1 U22673 ( .A1(n19876), .A2(n19875), .ZN(n19878) );
  NAND2HSV0 U22674 ( .A1(n25578), .A2(\pe8/got [6]), .ZN(n19877) );
  XOR2HSV0 U22675 ( .A1(n19878), .A2(n19877), .Z(n19880) );
  INAND2HSV2 U22676 ( .A1(n23642), .B1(n14060), .ZN(n19879) );
  XOR2HSV0 U22677 ( .A1(n19880), .A2(n19879), .Z(n19881) );
  XNOR2HSV1 U22678 ( .A1(n19882), .A2(n19881), .ZN(n19887) );
  XNOR2HSV1 U22679 ( .A1(n19887), .A2(n19886), .ZN(n19888) );
  XOR2HSV0 U22680 ( .A1(n19889), .A2(n19888), .Z(n19890) );
  XOR2HSV0 U22681 ( .A1(n19891), .A2(n19890), .Z(n19892) );
  XOR2HSV2 U22682 ( .A1(n19893), .A2(n19892), .Z(n19895) );
  NAND2HSV0 U22683 ( .A1(n22136), .A2(n19992), .ZN(n19894) );
  INHSV2 U22684 ( .I(n19979), .ZN(n19976) );
  INHSV2 U22685 ( .I(n19976), .ZN(n19896) );
  OAI21HSV2 U22686 ( .A1(n19975), .A2(n19980), .B(n19896), .ZN(n19899) );
  NOR2HSV4 U22687 ( .A1(n19975), .A2(n19896), .ZN(n19897) );
  CLKNAND2HSV3 U22688 ( .A1(n19899), .A2(n19898), .ZN(n23423) );
  NAND2HSV2 U22689 ( .A1(n22128), .A2(n23423), .ZN(n19974) );
  XNOR2HSV4 U22690 ( .A1(n19901), .A2(n19900), .ZN(n19903) );
  CLKNAND2HSV4 U22691 ( .A1(n19903), .A2(n19902), .ZN(n22119) );
  NOR2HSV2 U22692 ( .A1(n19988), .A2(n19904), .ZN(n19967) );
  NAND2HSV4 U22693 ( .A1(n22119), .A2(n19967), .ZN(n23444) );
  NAND2HSV2 U22694 ( .A1(n22140), .A2(\pe8/got [12]), .ZN(n19937) );
  NOR2HSV2 U22695 ( .A1(n19994), .A2(n19905), .ZN(n19935) );
  NAND2HSV0 U22696 ( .A1(n12007), .A2(n23721), .ZN(n19930) );
  NAND2HSV0 U22697 ( .A1(n28796), .A2(\pe8/got [5]), .ZN(n19924) );
  CLKNAND2HSV0 U22698 ( .A1(n28788), .A2(\pe8/got [6]), .ZN(n19923) );
  NAND2HSV0 U22699 ( .A1(\pe8/aot [9]), .A2(\pe8/bq[11] ), .ZN(n19907) );
  NAND2HSV0 U22700 ( .A1(\pe8/aot [14]), .A2(\pe8/bq[6] ), .ZN(n19906) );
  NAND2HSV0 U22701 ( .A1(\pe8/aot [13]), .A2(\pe8/bq[7] ), .ZN(n19909) );
  NAND2HSV0 U22702 ( .A1(\pe8/aot [4]), .A2(n25539), .ZN(n19908) );
  NAND2HSV0 U22703 ( .A1(\pe8/aot [5]), .A2(n25532), .ZN(n19911) );
  NAND2HSV0 U22704 ( .A1(\pe8/aot [12]), .A2(\pe8/bq[8] ), .ZN(n19910) );
  XOR2HSV0 U22705 ( .A1(n19911), .A2(n19910), .Z(n19913) );
  NAND2HSV0 U22706 ( .A1(\pe8/bq[10] ), .A2(\pe8/aot [10]), .ZN(n22252) );
  INHSV2 U22707 ( .I(n22230), .ZN(n25203) );
  NAND2HSV0 U22708 ( .A1(\pe8/aot [11]), .A2(\pe8/bq[9] ), .ZN(n19915) );
  NAND2HSV0 U22709 ( .A1(n28627), .A2(\pe8/bq[4] ), .ZN(n19914) );
  NAND2HSV0 U22710 ( .A1(\pe8/aot [8]), .A2(\pe8/bq[12] ), .ZN(n19917) );
  NAND2HSV0 U22711 ( .A1(\pe8/aot [7]), .A2(\pe8/bq[13] ), .ZN(n19916) );
  CLKNAND2HSV0 U22712 ( .A1(n23519), .A2(\pe8/pvq [13]), .ZN(n19918) );
  CLKNAND2HSV0 U22713 ( .A1(\pe8/aot [6]), .A2(n23529), .ZN(n23731) );
  NAND2HSV0 U22714 ( .A1(\pe8/aot [6]), .A2(\pe8/bq[14] ), .ZN(n19919) );
  OAI21HSV0 U22715 ( .A1(n19995), .A2(n23847), .B(n19919), .ZN(n19920) );
  XOR3HSV2 U22716 ( .A1(n19924), .A2(n19923), .A3(n19922), .Z(n19926) );
  NAND2HSV0 U22717 ( .A1(n25578), .A2(n14060), .ZN(n19925) );
  XOR2HSV0 U22718 ( .A1(n19926), .A2(n19925), .Z(n19928) );
  INAND2HSV2 U22719 ( .A1(n23642), .B1(n23605), .ZN(n19927) );
  XOR2HSV0 U22720 ( .A1(n19928), .A2(n19927), .Z(n19929) );
  XNOR2HSV1 U22721 ( .A1(n19930), .A2(n19929), .ZN(n19933) );
  NAND2HSV0 U22722 ( .A1(\pe8/got [10]), .A2(n19931), .ZN(n19932) );
  XNOR2HSV1 U22723 ( .A1(n19933), .A2(n19932), .ZN(n19934) );
  XNOR2HSV1 U22724 ( .A1(n19935), .A2(n19934), .ZN(n19936) );
  XNOR2HSV4 U22725 ( .A1(n19942), .A2(n19941), .ZN(n19966) );
  INHSV2 U22726 ( .I(n19944), .ZN(n19947) );
  CLKNAND2HSV1 U22727 ( .A1(n21315), .A2(n19945), .ZN(n19946) );
  CLKNHSV0 U22728 ( .I(n19948), .ZN(n19950) );
  NAND2HSV0 U22729 ( .A1(n19950), .A2(n19949), .ZN(n19951) );
  CLKNAND2HSV1 U22730 ( .A1(n18774), .A2(n21320), .ZN(n19955) );
  NOR2HSV1 U22731 ( .A1(n21315), .A2(n19953), .ZN(n19954) );
  CLKAND2HSV2 U22732 ( .A1(n19955), .A2(n19954), .Z(n19959) );
  INAND2HSV2 U22733 ( .A1(n28667), .B1(n18765), .ZN(n19957) );
  OAI21HSV2 U22734 ( .A1(n21320), .A2(n19956), .B(n19957), .ZN(n19958) );
  NAND2HSV2 U22735 ( .A1(n19959), .A2(n19958), .ZN(n19962) );
  OR2HSV1 U22736 ( .A1(n19960), .A2(n20058), .Z(n19961) );
  NAND3HSV4 U22737 ( .A1(n19963), .A2(n19962), .A3(n19961), .ZN(n19965) );
  XNOR2HSV4 U22738 ( .A1(n19966), .A2(n19965), .ZN(n22126) );
  NOR2HSV4 U22739 ( .A1(n22126), .A2(n18657), .ZN(n19964) );
  NOR2HSV4 U22740 ( .A1(n23443), .A2(n22118), .ZN(n19968) );
  AOI22HSV4 U22741 ( .A1(n19969), .A2(\pe8/ti_7t [13]), .B1(n19968), .B2(
        n22119), .ZN(n19970) );
  INHSV4 U22742 ( .I(n20052), .ZN(n22199) );
  INHSV4 U22743 ( .I(n22199), .ZN(n23846) );
  AOI21HSV2 U22744 ( .A1(n28685), .A2(n18773), .B(n19972), .ZN(n19973) );
  OAI21HSV4 U22745 ( .A1(n19974), .A2(n23846), .B(n19973), .ZN(n20054) );
  NOR2HSV1 U22746 ( .A1(n19980), .A2(n19979), .ZN(n19982) );
  CLKNAND2HSV1 U22747 ( .A1(n19982), .A2(n19981), .ZN(n19983) );
  INHSV2 U22748 ( .I(n19986), .ZN(n22137) );
  OR2HSV1 U22749 ( .A1(n19988), .A2(n19987), .Z(n19989) );
  NAND2HSV0 U22750 ( .A1(\pe8/got [12]), .A2(n19992), .ZN(n20046) );
  CLKNAND2HSV1 U22751 ( .A1(n21322), .A2(n28618), .ZN(n20043) );
  NAND2HSV2 U22752 ( .A1(n22140), .A2(\pe8/got [10]), .ZN(n20041) );
  NOR2HSV2 U22753 ( .A1(n19994), .A2(n19993), .ZN(n20039) );
  NAND2HSV0 U22754 ( .A1(n14060), .A2(n12007), .ZN(n20035) );
  INHSV2 U22755 ( .I(n19995), .ZN(n28641) );
  NAND2HSV0 U22756 ( .A1(n28641), .A2(\pe8/bq[3] ), .ZN(n25557) );
  XOR2HSV0 U22757 ( .A1(n23615), .A2(n25557), .Z(n20008) );
  NAND2HSV0 U22758 ( .A1(\pe8/aot [14]), .A2(\pe8/bq[4] ), .ZN(n19997) );
  INHSV2 U22759 ( .I(\pe8/bq[2] ), .ZN(n25555) );
  INHSV2 U22760 ( .I(n25555), .ZN(n21762) );
  NAND2HSV0 U22761 ( .A1(n28627), .A2(n21762), .ZN(n19996) );
  XOR2HSV0 U22762 ( .A1(n19997), .A2(n19996), .Z(n19999) );
  XNOR2HSV1 U22763 ( .A1(n19999), .A2(n19998), .ZN(n20007) );
  NAND2HSV0 U22764 ( .A1(\pe8/aot [9]), .A2(\pe8/bq[9] ), .ZN(n20001) );
  NAND2HSV0 U22765 ( .A1(\pe8/aot [4]), .A2(\pe8/bq[14] ), .ZN(n20000) );
  XOR2HSV0 U22766 ( .A1(n20001), .A2(n20000), .Z(n20005) );
  NAND2HSV0 U22767 ( .A1(\pe8/got [2]), .A2(n25624), .ZN(n20003) );
  NAND2HSV0 U22768 ( .A1(\pe8/aot [3]), .A2(n25532), .ZN(n20002) );
  XOR2HSV0 U22769 ( .A1(n20003), .A2(n20002), .Z(n20004) );
  XOR2HSV0 U22770 ( .A1(n20005), .A2(n20004), .Z(n20006) );
  XOR3HSV2 U22771 ( .A1(n20008), .A2(n20007), .A3(n20006), .Z(n20011) );
  NAND2HSV0 U22772 ( .A1(n25203), .A2(n20009), .ZN(n20010) );
  XOR2HSV0 U22773 ( .A1(n20011), .A2(n20010), .Z(n20029) );
  NAND2HSV0 U22774 ( .A1(\pe8/aot [5]), .A2(n25565), .ZN(n20013) );
  NAND2HSV0 U22775 ( .A1(\pe8/aot [12]), .A2(\pe8/bq[6] ), .ZN(n20012) );
  XOR2HSV0 U22776 ( .A1(n20013), .A2(n20012), .Z(n20017) );
  NAND2HSV0 U22777 ( .A1(\pe8/aot [7]), .A2(\pe8/bq[11] ), .ZN(n20015) );
  NAND2HSV0 U22778 ( .A1(\pe8/aot [2]), .A2(n25539), .ZN(n20014) );
  XOR2HSV0 U22779 ( .A1(n20015), .A2(n20014), .Z(n20016) );
  XOR2HSV0 U22780 ( .A1(n20017), .A2(n20016), .Z(n20025) );
  NAND2HSV0 U22781 ( .A1(\pe8/aot [13]), .A2(\pe8/bq[5] ), .ZN(n20019) );
  NAND2HSV0 U22782 ( .A1(\pe8/aot [8]), .A2(\pe8/bq[10] ), .ZN(n20018) );
  XOR2HSV0 U22783 ( .A1(n20019), .A2(n20018), .Z(n20023) );
  NAND2HSV0 U22784 ( .A1(\pe8/aot [6]), .A2(\pe8/bq[12] ), .ZN(n20021) );
  NAND2HSV0 U22785 ( .A1(\pe8/aot [10]), .A2(\pe8/bq[8] ), .ZN(n20020) );
  XOR2HSV0 U22786 ( .A1(n20021), .A2(n20020), .Z(n20022) );
  XOR2HSV0 U22787 ( .A1(n20023), .A2(n20022), .Z(n20024) );
  XOR2HSV0 U22788 ( .A1(n20025), .A2(n20024), .Z(n20027) );
  NAND2HSV0 U22789 ( .A1(n28796), .A2(\pe8/got [3]), .ZN(n20026) );
  XNOR2HSV1 U22790 ( .A1(n20027), .A2(n20026), .ZN(n20028) );
  XNOR2HSV1 U22791 ( .A1(n20029), .A2(n20028), .ZN(n20031) );
  NAND2HSV0 U22792 ( .A1(n25578), .A2(\pe8/got [5]), .ZN(n20030) );
  XNOR2HSV1 U22793 ( .A1(n20031), .A2(n20030), .ZN(n20033) );
  INAND2HSV0 U22794 ( .A1(n23642), .B1(\pe8/got [6]), .ZN(n20032) );
  XNOR2HSV1 U22795 ( .A1(n20033), .A2(n20032), .ZN(n20034) );
  XNOR2HSV1 U22796 ( .A1(n20035), .A2(n20034), .ZN(n20037) );
  XNOR2HSV1 U22797 ( .A1(n20037), .A2(n20036), .ZN(n20038) );
  XOR2HSV0 U22798 ( .A1(n20039), .A2(n20038), .Z(n20040) );
  XNOR2HSV1 U22799 ( .A1(n20041), .A2(n20040), .ZN(n20042) );
  XOR2HSV2 U22800 ( .A1(n20043), .A2(n20042), .Z(n20045) );
  XNOR3HSV2 U22801 ( .A1(n20046), .A2(n20045), .A3(n20044), .ZN(n20047) );
  XNOR2HSV4 U22802 ( .A1(n20048), .A2(n20047), .ZN(n23866) );
  NOR2HSV2 U22803 ( .A1(n23866), .A2(n20049), .ZN(n20050) );
  INHSV2 U22804 ( .I(n22137), .ZN(n22138) );
  INHSV3 U22805 ( .I(n23866), .ZN(n20055) );
  INHSV3 U22806 ( .I(n20052), .ZN(n21004) );
  INHSV2 U22807 ( .I(\pe8/ti_7t [15]), .ZN(n23870) );
  NOR2HSV1 U22808 ( .A1(n18783), .A2(n23870), .ZN(n25524) );
  INHSV2 U22809 ( .I(n25524), .ZN(n20053) );
  AOI21HSV2 U22810 ( .A1(n12218), .A2(n20055), .B(n20054), .ZN(n20062) );
  CLKNAND2HSV0 U22811 ( .A1(n21004), .A2(n23866), .ZN(n20056) );
  CLKAND2HSV2 U22812 ( .A1(n20057), .A2(n20056), .Z(n20061) );
  IOA21HSV2 U22813 ( .A1(n23866), .A2(n20058), .B(n22128), .ZN(n20059) );
  INHSV2 U22814 ( .I(n20059), .ZN(n20060) );
  NAND3HSV4 U22815 ( .A1(n20062), .A2(n20061), .A3(n20060), .ZN(n25522) );
  INHSV4 U22816 ( .I(n25522), .ZN(n20063) );
  NOR2HSV4 U22817 ( .A1(n20064), .A2(n20063), .ZN(n22198) );
  INHSV4 U22818 ( .I(n22198), .ZN(n28420) );
  INHSV4 U22819 ( .I(n23717), .ZN(n28475) );
  NOR2HSV1 U22820 ( .A1(n20066), .A2(n20065), .ZN(n20067) );
  INHSV2 U22821 ( .I(n20069), .ZN(n20071) );
  NAND2HSV2 U22822 ( .A1(n20073), .A2(n20072), .ZN(n22509) );
  CLKNAND2HSV1 U22823 ( .A1(n22509), .A2(n16759), .ZN(n20122) );
  NAND2HSV0 U22824 ( .A1(n28644), .A2(n26094), .ZN(n20120) );
  INHSV1 U22825 ( .I(n20074), .ZN(n26159) );
  INHSV2 U22826 ( .I(\pe10/got [9]), .ZN(n25214) );
  NOR2HSV2 U22827 ( .A1(n26159), .A2(n25214), .ZN(n20118) );
  NAND2HSV0 U22828 ( .A1(n28794), .A2(\pe10/got [7]), .ZN(n20114) );
  NAND2HSV0 U22829 ( .A1(n22458), .A2(\pe10/got [3]), .ZN(n20076) );
  NAND2HSV0 U22830 ( .A1(\pe10/aot [4]), .A2(n16897), .ZN(n20075) );
  XOR2HSV0 U22831 ( .A1(n20076), .A2(n20075), .Z(n20092) );
  CLKNAND2HSV0 U22832 ( .A1(\pe10/bq[8] ), .A2(\pe10/aot [9]), .ZN(n26161) );
  CLKNHSV0 U22833 ( .I(\pe10/aot [9]), .ZN(n20078) );
  OAI21HSV0 U22834 ( .A1(n22722), .A2(n20078), .B(n20077), .ZN(n20079) );
  OAI21HSV0 U22835 ( .A1(n20080), .A2(n26161), .B(n20079), .ZN(n20082) );
  CLKNHSV0 U22836 ( .I(\pe10/aot [10]), .ZN(n22719) );
  NOR2HSV0 U22837 ( .A1(n22719), .A2(n20081), .ZN(n25223) );
  XNOR2HSV1 U22838 ( .A1(n20082), .A2(n25223), .ZN(n20091) );
  NAND2HSV0 U22839 ( .A1(n20083), .A2(\pe10/bq[3] ), .ZN(n20085) );
  NAND2HSV0 U22840 ( .A1(\pe10/aot [7]), .A2(\pe10/bq[12] ), .ZN(n20084) );
  XOR2HSV0 U22841 ( .A1(n20085), .A2(n20084), .Z(n20089) );
  NAND2HSV0 U22842 ( .A1(\pe10/bq[5] ), .A2(\pe10/aot [14]), .ZN(n20087) );
  NAND2HSV0 U22843 ( .A1(\pe10/aot [6]), .A2(\pe10/bq[13] ), .ZN(n20086) );
  XOR2HSV0 U22844 ( .A1(n20087), .A2(n20086), .Z(n20088) );
  XOR2HSV0 U22845 ( .A1(n20089), .A2(n20088), .Z(n20090) );
  XOR3HSV2 U22846 ( .A1(n20092), .A2(n20091), .A3(n20090), .Z(n20110) );
  CLKNAND2HSV0 U22847 ( .A1(n16850), .A2(\pe10/got [5]), .ZN(n20109) );
  NAND2HSV0 U22848 ( .A1(\pe10/aot [8]), .A2(\pe10/bq[11] ), .ZN(n20094) );
  NAND2HSV0 U22849 ( .A1(\pe10/aot [3]), .A2(n17084), .ZN(n20093) );
  XOR2HSV0 U22850 ( .A1(n20094), .A2(n20093), .Z(n20098) );
  NAND2HSV0 U22851 ( .A1(\pe10/aot [5]), .A2(\pe10/bq[14] ), .ZN(n20096) );
  NAND2HSV0 U22852 ( .A1(\pe10/aot [13]), .A2(\pe10/bq[6] ), .ZN(n20095) );
  XOR2HSV0 U22853 ( .A1(n20096), .A2(n20095), .Z(n20097) );
  XOR2HSV0 U22854 ( .A1(n20098), .A2(n20097), .Z(n20105) );
  NAND2HSV0 U22855 ( .A1(n16973), .A2(\pe10/bq[4] ), .ZN(n20100) );
  NAND2HSV0 U22856 ( .A1(\pe10/aot [12]), .A2(\pe10/bq[7] ), .ZN(n20099) );
  XOR2HSV0 U22857 ( .A1(n20100), .A2(n20099), .Z(n20103) );
  NAND2HSV0 U22858 ( .A1(n23544), .A2(\pe10/pvq [14]), .ZN(n20101) );
  XOR2HSV0 U22859 ( .A1(n20101), .A2(\pe10/phq [14]), .Z(n20102) );
  XOR2HSV0 U22860 ( .A1(n20103), .A2(n20102), .Z(n20104) );
  XOR2HSV0 U22861 ( .A1(n20105), .A2(n20104), .Z(n20107) );
  NAND2HSV0 U22862 ( .A1(n26189), .A2(\pe10/got [4]), .ZN(n20106) );
  XNOR2HSV1 U22863 ( .A1(n20107), .A2(n20106), .ZN(n20108) );
  XOR3HSV2 U22864 ( .A1(n20110), .A2(n20109), .A3(n20108), .Z(n20112) );
  NAND2HSV0 U22865 ( .A1(n23474), .A2(\pe10/got [6]), .ZN(n20111) );
  XNOR2HSV1 U22866 ( .A1(n20112), .A2(n20111), .ZN(n20113) );
  XNOR2HSV1 U22867 ( .A1(n20114), .A2(n20113), .ZN(n20116) );
  NAND2HSV0 U22868 ( .A1(n26131), .A2(n28642), .ZN(n20115) );
  XNOR2HSV1 U22869 ( .A1(n20116), .A2(n20115), .ZN(n20117) );
  XOR2HSV0 U22870 ( .A1(n20118), .A2(n20117), .Z(n20119) );
  XNOR2HSV1 U22871 ( .A1(n20120), .A2(n20119), .ZN(n20121) );
  NAND2HSV0 U22872 ( .A1(n21741), .A2(n26212), .ZN(n20123) );
  XNOR2HSV1 U22873 ( .A1(n20124), .A2(n20123), .ZN(n20127) );
  NAND2HSV2 U22874 ( .A1(n20125), .A2(n28479), .ZN(n20126) );
  AND2HSV2 U22875 ( .A1(n20133), .A2(n20128), .Z(n20129) );
  CLKNAND2HSV2 U22876 ( .A1(n20130), .A2(n20129), .ZN(n20141) );
  INHSV2 U22877 ( .I(n22432), .ZN(n20131) );
  INAND2HSV2 U22878 ( .A1(n20133), .B1(n20142), .ZN(n22430) );
  INHSV2 U22879 ( .I(n20134), .ZN(n20135) );
  CLKNAND2HSV3 U22880 ( .A1(n20137), .A2(n20136), .ZN(n20138) );
  CLKNAND2HSV2 U22881 ( .A1(n20138), .A2(n20139), .ZN(n20140) );
  NAND2HSV2 U22882 ( .A1(n25685), .A2(n20142), .ZN(n20143) );
  OAI21HSV2 U22883 ( .A1(n25685), .A2(n20145), .B(n28988), .ZN(n20146) );
  CLKNAND2HSV2 U22884 ( .A1(n20147), .A2(n20146), .ZN(n22440) );
  NOR2HSV1 U22885 ( .A1(n28810), .A2(n20148), .ZN(n25258) );
  AOI22HSV2 U22886 ( .A1(n20149), .A2(\pe10/ti_7t [14]), .B1(n25685), .B2(
        n25258), .ZN(n25689) );
  INHSV4 U22887 ( .I(ctro11), .ZN(n20207) );
  BUFHSV2 U22888 ( .I(n20207), .Z(n20636) );
  CLKBUFHSV4 U22889 ( .I(n20207), .Z(n20559) );
  CLKNAND2HSV1 U22890 ( .A1(n20302), .A2(\pe11/ti_7t [15]), .ZN(n24884) );
  NAND2HSV2 U22891 ( .A1(n20302), .A2(\pe11/ti_7t [7]), .ZN(n20403) );
  INHSV2 U22892 ( .I(n20403), .ZN(n20458) );
  CLKBUFHSV4 U22893 ( .I(\pe11/got [16]), .Z(n20182) );
  INHSV2 U22894 ( .I(n20182), .ZN(n20370) );
  INHSV3 U22895 ( .I(n20370), .ZN(n25488) );
  CLKBUFHSV4 U22896 ( .I(\pe11/got [14]), .Z(n20613) );
  INHSV2 U22897 ( .I(\pe11/phq [3]), .ZN(n20150) );
  CLKNAND2HSV1 U22898 ( .A1(n20152), .A2(n20153), .ZN(n20156) );
  INHSV2 U22899 ( .I(n20152), .ZN(n20155) );
  INHSV2 U22900 ( .I(\pe11/aot [16]), .ZN(n20336) );
  CLKAND2HSV2 U22901 ( .A1(n20157), .A2(\pe11/bq[14] ), .Z(n20159) );
  INHSV2 U22902 ( .I(n20164), .ZN(n20470) );
  NAND2HSV2 U22903 ( .A1(n20470), .A2(\pe11/pvq [3]), .ZN(n20158) );
  XNOR2HSV4 U22904 ( .A1(n20159), .A2(n20158), .ZN(n20160) );
  INHSV2 U22905 ( .I(n11851), .ZN(n20255) );
  BUFHSV8 U22906 ( .I(n20207), .Z(n25512) );
  INHSV2 U22907 ( .I(n25512), .ZN(n20620) );
  CLKXOR2HSV4 U22908 ( .A1(n20161), .A2(n20160), .Z(n25505) );
  NAND2HSV2 U22909 ( .A1(n25505), .A2(n20187), .ZN(n20162) );
  INHSV2 U22910 ( .I(n20219), .ZN(n20184) );
  INHSV6 U22911 ( .I(n20164), .ZN(n20408) );
  NOR2HSV4 U22912 ( .A1(n20165), .A2(n20166), .ZN(n20168) );
  CLKNAND2HSV3 U22913 ( .A1(n20408), .A2(\pe11/pvq [2]), .ZN(n20167) );
  AOI22HSV4 U22914 ( .A1(n20408), .A2(n20168), .B1(n20167), .B2(n20165), .ZN(
        n20170) );
  NAND2HSV0 U22915 ( .A1(\pe11/bq[15] ), .A2(\pe11/aot [16]), .ZN(n20169) );
  XNOR2HSV4 U22916 ( .A1(n20170), .A2(n20169), .ZN(n20175) );
  CLKNAND2HSV1 U22917 ( .A1(n20329), .A2(n20171), .ZN(n20173) );
  NAND2HSV0 U22918 ( .A1(\pe11/aot [15]), .A2(\pe11/bq[16] ), .ZN(n20172) );
  XNOR2HSV4 U22919 ( .A1(n20175), .A2(n20174), .ZN(n25490) );
  INHSV2 U22920 ( .I(n20565), .ZN(n20689) );
  NOR2HSV4 U22921 ( .A1(n20176), .A2(n20215), .ZN(n20177) );
  CLKNHSV0 U22922 ( .I(ctro11), .ZN(n20543) );
  BUFHSV2 U22923 ( .I(n20179), .Z(n20450) );
  INHSV2 U22924 ( .I(n20450), .ZN(n20561) );
  NAND2HSV2 U22925 ( .A1(n20543), .A2(n20561), .ZN(n20367) );
  NOR2HSV4 U22926 ( .A1(n25502), .A2(n20367), .ZN(n20285) );
  CLKAND2HSV2 U22927 ( .A1(n20302), .A2(\pe11/ti_7t [2]), .Z(n20284) );
  AOI21HSV2 U22928 ( .A1(n25490), .A2(n20285), .B(n20284), .ZN(n20180) );
  INHSV2 U22929 ( .I(n25502), .ZN(n20185) );
  INHSV2 U22930 ( .I(n20182), .ZN(n20619) );
  NAND3HSV3 U22931 ( .A1(n20184), .A2(n20186), .A3(n20183), .ZN(n20253) );
  CLKNAND2HSV0 U22932 ( .A1(n20253), .A2(n20636), .ZN(n20194) );
  NOR2HSV3 U22933 ( .A1(n20188), .A2(n20185), .ZN(n20221) );
  NOR2HSV2 U22934 ( .A1(n20188), .A2(\pe11/got [15]), .ZN(n20189) );
  INHSV2 U22935 ( .I(n20189), .ZN(n20190) );
  INHSV2 U22936 ( .I(n20222), .ZN(n20192) );
  NAND2HSV4 U22937 ( .A1(n20193), .A2(n20192), .ZN(n20254) );
  INHSV3 U22938 ( .I(n20254), .ZN(n20214) );
  NOR2HSV2 U22939 ( .A1(n20194), .A2(n20214), .ZN(n20317) );
  INHSV2 U22940 ( .I(n20195), .ZN(n20218) );
  CLKNAND2HSV1 U22941 ( .A1(\pe11/aot [15]), .A2(\pe11/bq[14] ), .ZN(n20197)
         );
  NAND2HSV2 U22942 ( .A1(\pe11/bq[15] ), .A2(\pe11/aot [14]), .ZN(n20196) );
  XOR2HSV0 U22943 ( .A1(n20197), .A2(n20196), .Z(n20200) );
  NAND2HSV0 U22944 ( .A1(\pe11/aot [13]), .A2(\pe11/bq[16] ), .ZN(n20199) );
  CLKNAND2HSV0 U22945 ( .A1(\pe11/bq[13] ), .A2(\pe11/aot [16]), .ZN(n20198)
         );
  CLKNAND2HSV1 U22946 ( .A1(n20470), .A2(\pe11/pvq [4]), .ZN(n20202) );
  CLKXOR2HSV2 U22947 ( .A1(n20203), .A2(n20202), .Z(n20204) );
  XNOR2HSV4 U22948 ( .A1(n20205), .A2(n20204), .ZN(n20209) );
  BUFHSV2 U22949 ( .I(n20207), .Z(n25515) );
  BUFHSV2 U22950 ( .I(\pe11/got [14]), .Z(n20354) );
  OAI21HSV1 U22951 ( .A1(n25515), .A2(\pe11/ti_7t [1]), .B(n20354), .ZN(n20206) );
  AOI21HSV4 U22952 ( .A1(n12291), .A2(n20285), .B(n20284), .ZN(n20279) );
  NAND2HSV2 U22953 ( .A1(n20228), .A2(\pe11/got [15]), .ZN(n20210) );
  XNOR2HSV4 U22954 ( .A1(n20211), .A2(n20210), .ZN(n20314) );
  BUFHSV2 U22955 ( .I(n20314), .Z(n20318) );
  INHSV2 U22956 ( .I(n20559), .ZN(n20308) );
  NOR2HSV2 U22957 ( .A1(n20308), .A2(n20255), .ZN(n20456) );
  INHSV2 U22958 ( .I(n20456), .ZN(n20556) );
  NOR2HSV2 U22959 ( .A1(n20314), .A2(n20556), .ZN(n20212) );
  INHSV2 U22960 ( .I(n20212), .ZN(n20216) );
  CLKNHSV1 U22961 ( .I(n20253), .ZN(n20213) );
  NOR2HSV2 U22962 ( .A1(n20214), .A2(n20213), .ZN(n20315) );
  NAND2HSV2 U22963 ( .A1(n20215), .A2(\pe11/ti_7t [4]), .ZN(n20313) );
  OAI22HSV2 U22964 ( .A1(n20216), .A2(n20315), .B1(n20255), .B2(n20313), .ZN(
        n20217) );
  AOI21HSV4 U22965 ( .A1(n20218), .A2(n20318), .B(n20217), .ZN(n20307) );
  CLKNHSV0 U22966 ( .I(n20344), .ZN(n20220) );
  NAND2HSV2 U22967 ( .A1(n20620), .A2(\pe11/ti_7t [3]), .ZN(n20348) );
  INHSV2 U22968 ( .I(n20450), .ZN(n20775) );
  NAND2HSV4 U22969 ( .A1(n20228), .A2(n20775), .ZN(n20345) );
  CLKBUFHSV4 U22970 ( .I(n20345), .Z(n25508) );
  INHSV2 U22971 ( .I(n20354), .ZN(n20402) );
  AOI31HSV2 U22972 ( .A1(n20220), .A2(n20348), .A3(n25508), .B(n20402), .ZN(
        n20226) );
  INHSV2 U22973 ( .I(n20348), .ZN(n20256) );
  NOR2HSV2 U22974 ( .A1(n25508), .A2(n20256), .ZN(n20224) );
  NOR2HSV3 U22975 ( .A1(n20222), .A2(n20221), .ZN(n20347) );
  INHSV1 U22976 ( .I(n20347), .ZN(n20223) );
  CLKNAND2HSV1 U22977 ( .A1(n20224), .A2(n20223), .ZN(n20225) );
  CLKNAND2HSV1 U22978 ( .A1(n20226), .A2(n20225), .ZN(n20246) );
  BUFHSV2 U22979 ( .I(\pe11/got [13]), .Z(n20292) );
  BUFHSV8 U22980 ( .I(n20228), .Z(n20505) );
  CLKNHSV2 U22981 ( .I(n20707), .ZN(n20229) );
  NAND2HSV0 U22982 ( .A1(\pe11/bq[11] ), .A2(\pe11/aot [16]), .ZN(n20231) );
  CLKNAND2HSV0 U22983 ( .A1(\pe11/bq[13] ), .A2(\pe11/aot [14]), .ZN(n20230)
         );
  XOR2HSV0 U22984 ( .A1(n20231), .A2(n20230), .Z(n20235) );
  CLKNHSV1 U22985 ( .I(\pe11/aot [15]), .ZN(n20385) );
  NOR2HSV2 U22986 ( .A1(n20267), .A2(n20385), .ZN(n20233) );
  NAND2HSV0 U22987 ( .A1(\pe11/bq[14] ), .A2(\pe11/aot [13]), .ZN(n20232) );
  XOR2HSV0 U22988 ( .A1(n20233), .A2(n20232), .Z(n20234) );
  XOR2HSV0 U22989 ( .A1(n20235), .A2(n20234), .Z(n20242) );
  CLKNAND2HSV0 U22990 ( .A1(n20470), .A2(\pe11/pvq [6]), .ZN(n20236) );
  NAND2HSV0 U22991 ( .A1(\pe11/bq[16] ), .A2(\pe11/aot [11]), .ZN(n20238) );
  NAND2HSV0 U22992 ( .A1(\pe11/bq[15] ), .A2(\pe11/aot [12]), .ZN(n20237) );
  XOR2HSV0 U22993 ( .A1(n20238), .A2(n20237), .Z(n20239) );
  CLKNAND2HSV2 U22994 ( .A1(n28629), .A2(\pe11/got [12]), .ZN(n20240) );
  XOR3HSV2 U22995 ( .A1(n20242), .A2(n20241), .A3(n20240), .Z(n20243) );
  MUX2NHSV2 U22996 ( .I0(n20245), .I1(n20244), .S(n20243), .ZN(n20247) );
  NAND2HSV2 U22997 ( .A1(n20246), .A2(n20247), .ZN(n20251) );
  INHSV2 U22998 ( .I(n20246), .ZN(n20249) );
  CLKNHSV2 U22999 ( .I(n20247), .ZN(n20248) );
  CLKNAND2HSV2 U23000 ( .A1(n20249), .A2(n20248), .ZN(n20250) );
  NAND2HSV4 U23001 ( .A1(n20251), .A2(n20250), .ZN(n20306) );
  XNOR2HSV4 U23002 ( .A1(n20307), .A2(n20306), .ZN(n20459) );
  CLKNAND2HSV3 U23003 ( .A1(n20459), .A2(n24889), .ZN(n20252) );
  INHSV4 U23004 ( .I(n20252), .ZN(n20371) );
  NOR2HSV2 U23005 ( .A1(n20345), .A2(n20255), .ZN(n20258) );
  CLKAND2HSV1 U23006 ( .A1(n20256), .A2(n25504), .Z(n20257) );
  AOI21HSV2 U23007 ( .A1(n20347), .A2(n20258), .B(n20257), .ZN(n20262) );
  NAND2HSV0 U23008 ( .A1(n20345), .A2(n25504), .ZN(n20259) );
  CLKNHSV1 U23009 ( .I(n20259), .ZN(n20260) );
  CLKNAND2HSV1 U23010 ( .A1(n20260), .A2(n20344), .ZN(n20261) );
  INHSV2 U23011 ( .I(\pe11/aot [12]), .ZN(n20263) );
  NOR2HSV2 U23012 ( .A1(n20326), .A2(n20263), .ZN(n20266) );
  XNOR2HSV4 U23013 ( .A1(n20266), .A2(n20265), .ZN(n20271) );
  CLKNAND2HSV1 U23014 ( .A1(\pe11/bq[12] ), .A2(\pe11/aot [16]), .ZN(n20269)
         );
  XNOR2HSV4 U23015 ( .A1(n20271), .A2(n20270), .ZN(n20281) );
  CLKNAND2HSV1 U23016 ( .A1(n20329), .A2(\pe11/got [12]), .ZN(n20274) );
  XNOR2HSV4 U23017 ( .A1(n20274), .A2(n20273), .ZN(n20277) );
  NAND2HSV2 U23018 ( .A1(\pe11/aot [13]), .A2(\pe11/bq[15] ), .ZN(n20275) );
  XNOR2HSV1 U23019 ( .A1(n20275), .A2(\pe11/phq [5]), .ZN(n20276) );
  XNOR2HSV4 U23020 ( .A1(n20277), .A2(n20276), .ZN(n20280) );
  XOR2HSV0 U23021 ( .A1(n20281), .A2(n20280), .Z(n20278) );
  NAND2HSV2 U23022 ( .A1(n12293), .A2(n20278), .ZN(n20283) );
  CLKNHSV2 U23023 ( .I(n20279), .ZN(n20282) );
  XNOR2HSV4 U23024 ( .A1(n20281), .A2(n20280), .ZN(n20286) );
  OAI22HSV2 U23025 ( .A1(n20283), .A2(n20282), .B1(n20354), .B2(n20286), .ZN(
        n20291) );
  AOI21HSV0 U23026 ( .A1(n12291), .A2(n20285), .B(n20284), .ZN(n20289) );
  CLKNAND2HSV0 U23027 ( .A1(n20286), .A2(n20354), .ZN(n20287) );
  AOI21HSV2 U23028 ( .A1(n20289), .A2(n12292), .B(n20287), .ZN(n20290) );
  NOR2HSV4 U23029 ( .A1(n20291), .A2(n20290), .ZN(n20294) );
  NAND2HSV2 U23030 ( .A1(n20292), .A2(n25489), .ZN(n20293) );
  XNOR2HSV4 U23031 ( .A1(n20294), .A2(n20293), .ZN(n20296) );
  INHSV3 U23032 ( .I(n20295), .ZN(n20298) );
  INHSV2 U23033 ( .I(n20296), .ZN(n20297) );
  NAND2HSV4 U23034 ( .A1(n20298), .A2(n20297), .ZN(n20299) );
  CLKNAND2HSV8 U23035 ( .A1(n20300), .A2(n20299), .ZN(n23468) );
  AOI22HSV4 U23036 ( .A1(\pe11/ti_7t [5]), .A2(n20302), .B1(n20301), .B2(
        n23468), .ZN(n20369) );
  INHSV2 U23037 ( .I(n25513), .ZN(n20303) );
  NAND2HSV2 U23038 ( .A1(n20565), .A2(n20303), .ZN(n20305) );
  NOR2HSV4 U23039 ( .A1(n23468), .A2(n25032), .ZN(n20304) );
  CLKNAND2HSV4 U23040 ( .A1(n20305), .A2(n20304), .ZN(n20368) );
  INHSV2 U23041 ( .I(n28668), .ZN(n24831) );
  CLKNAND2HSV3 U23042 ( .A1(n20371), .A2(n24831), .ZN(n20312) );
  XNOR2HSV4 U23043 ( .A1(n20307), .A2(n20306), .ZN(n20309) );
  NOR2HSV4 U23044 ( .A1(n20309), .A2(n20308), .ZN(n20374) );
  NAND2HSV2 U23045 ( .A1(n20374), .A2(n28668), .ZN(n20311) );
  NOR2HSV2 U23046 ( .A1(n20636), .A2(\pe11/ti_7t [6]), .ZN(n20464) );
  NOR2HSV2 U23047 ( .A1(n20464), .A2(n20619), .ZN(n20310) );
  OAI21HSV2 U23048 ( .A1(n20315), .A2(n20314), .B(n20313), .ZN(n20316) );
  AOI21HSV4 U23049 ( .A1(n20318), .A2(n20317), .B(n20316), .ZN(n21941) );
  NOR2HSV1 U23050 ( .A1(n21941), .A2(n20402), .ZN(n20353) );
  NAND2HSV0 U23051 ( .A1(n20320), .A2(n20319), .ZN(n20321) );
  NAND2HSV0 U23052 ( .A1(n20321), .A2(\pe11/got [11]), .ZN(n20322) );
  XNOR2HSV4 U23053 ( .A1(n20323), .A2(n20322), .ZN(n20343) );
  NAND2HSV0 U23054 ( .A1(\pe11/aot [12]), .A2(\pe11/bq[14] ), .ZN(n20325) );
  NAND2HSV0 U23055 ( .A1(n20470), .A2(\pe11/pvq [7]), .ZN(n20324) );
  XOR2HSV0 U23056 ( .A1(n20325), .A2(n20324), .Z(n20341) );
  NAND2HSV0 U23057 ( .A1(\pe11/bq[13] ), .A2(\pe11/aot [13]), .ZN(n20328) );
  INHSV2 U23058 ( .I(n20326), .ZN(n27058) );
  NAND2HSV0 U23059 ( .A1(n27058), .A2(\pe11/aot [10]), .ZN(n20327) );
  XOR2HSV0 U23060 ( .A1(n20328), .A2(n20327), .Z(n20332) );
  NAND2HSV0 U23061 ( .A1(n20329), .A2(\pe11/got [10]), .ZN(n20330) );
  XNOR2HSV1 U23062 ( .A1(n20330), .A2(\pe11/phq [7]), .ZN(n20331) );
  XNOR2HSV1 U23063 ( .A1(n20332), .A2(n20331), .ZN(n20340) );
  CLKNHSV0 U23064 ( .I(\pe11/aot [14]), .ZN(n20333) );
  INHSV2 U23065 ( .I(n20333), .ZN(n24771) );
  NAND2HSV0 U23066 ( .A1(\pe11/bq[12] ), .A2(n24771), .ZN(n20335) );
  BUFHSV4 U23067 ( .I(\pe11/bq[15] ), .Z(n24997) );
  NAND2HSV0 U23068 ( .A1(n24997), .A2(\pe11/aot [11]), .ZN(n20334) );
  XOR2HSV0 U23069 ( .A1(n20335), .A2(n20334), .Z(n20338) );
  CLKNHSV0 U23070 ( .I(\pe11/bq[11] ), .ZN(n24314) );
  XOR2HSV0 U23071 ( .A1(n20338), .A2(n20337), .Z(n20339) );
  XOR3HSV2 U23072 ( .A1(n20341), .A2(n20340), .A3(n20339), .Z(n20342) );
  XNOR2HSV4 U23073 ( .A1(n20343), .A2(n20342), .ZN(n20352) );
  INHSV2 U23074 ( .I(n20345), .ZN(n20346) );
  NAND2HSV2 U23075 ( .A1(n20347), .A2(n20346), .ZN(n20349) );
  NAND3HSV3 U23076 ( .A1(n20350), .A2(n20349), .A3(n20348), .ZN(n28807) );
  XNOR2HSV4 U23077 ( .A1(n20352), .A2(n20351), .ZN(n20357) );
  NAND2HSV2 U23078 ( .A1(n20353), .A2(n20357), .ZN(n20360) );
  CLKNHSV0 U23079 ( .I(n25028), .ZN(n20356) );
  INHSV3 U23080 ( .I(n20357), .ZN(n20358) );
  XNOR2HSV4 U23081 ( .A1(n20362), .A2(n20361), .ZN(n20400) );
  INHSV2 U23082 ( .I(n20400), .ZN(n20363) );
  CLKNAND2HSV2 U23083 ( .A1(n20364), .A2(n20363), .ZN(n20366) );
  NAND2HSV2 U23084 ( .A1(n20401), .A2(n20400), .ZN(n20365) );
  CLKNAND2HSV3 U23085 ( .A1(n20366), .A2(n20365), .ZN(n20446) );
  INHSV2 U23086 ( .I(n20367), .ZN(n20844) );
  AOI22HSV4 U23087 ( .A1(n20458), .A2(n25488), .B1(n20446), .B2(n20844), .ZN(
        n20394) );
  NAND2HSV4 U23088 ( .A1(n20369), .A2(n20368), .ZN(n28668) );
  NAND2HSV4 U23089 ( .A1(n28668), .A2(n20182), .ZN(n20462) );
  CLKNAND2HSV1 U23090 ( .A1(n20462), .A2(n20371), .ZN(n20438) );
  NOR2HSV1 U23091 ( .A1(n20464), .A2(n20372), .ZN(n20373) );
  INHSV4 U23092 ( .I(n20462), .ZN(n20461) );
  NAND2HSV2 U23093 ( .A1(n20461), .A2(n20374), .ZN(n20440) );
  NAND2HSV2 U23094 ( .A1(n20505), .A2(\pe11/got [11]), .ZN(n20376) );
  NAND2HSV0 U23095 ( .A1(n25489), .A2(\pe11/got [10]), .ZN(n20375) );
  NAND2HSV0 U23096 ( .A1(\pe11/bq[14] ), .A2(\pe11/aot [11]), .ZN(n20378) );
  NAND2HSV0 U23097 ( .A1(\pe11/aot [9]), .A2(n27058), .ZN(n20377) );
  XOR2HSV0 U23098 ( .A1(n20378), .A2(n20377), .Z(n20382) );
  NAND2HSV0 U23099 ( .A1(\pe11/bq[12] ), .A2(\pe11/aot [13]), .ZN(n20380) );
  CLKNAND2HSV0 U23100 ( .A1(n20157), .A2(\pe11/bq[9] ), .ZN(n20379) );
  XOR2HSV0 U23101 ( .A1(n20380), .A2(n20379), .Z(n20381) );
  XOR2HSV0 U23102 ( .A1(n20382), .A2(n20381), .Z(n20388) );
  CLKNHSV1 U23103 ( .I(n20587), .ZN(n22112) );
  INHSV2 U23104 ( .I(n22112), .ZN(n24975) );
  XNOR2HSV1 U23105 ( .A1(n20383), .A2(\pe11/phq [8]), .ZN(n20386) );
  NOR2HSV2 U23106 ( .A1(n20384), .A2(n20385), .ZN(n20662) );
  XNOR2HSV1 U23107 ( .A1(n20386), .A2(n20662), .ZN(n20387) );
  INHSV4 U23108 ( .I(n21941), .ZN(n20467) );
  INHSV2 U23109 ( .I(n20707), .ZN(n25027) );
  NAND2HSV2 U23110 ( .A1(n20601), .A2(n20613), .ZN(n20391) );
  NAND2HSV2 U23111 ( .A1(n20394), .A2(n20452), .ZN(n20397) );
  INHSV2 U23112 ( .I(n20394), .ZN(n20395) );
  INHSV4 U23113 ( .I(n20452), .ZN(n20448) );
  NAND2HSV2 U23114 ( .A1(\pe11/ti_7t [8]), .A2(n20637), .ZN(n20552) );
  OR2HSV1 U23115 ( .A1(n20552), .A2(n20372), .Z(n20398) );
  XNOR2HSV4 U23116 ( .A1(n20401), .A2(n20400), .ZN(n20457) );
  AOI21HSV2 U23117 ( .A1(n23470), .A2(n20403), .B(n20402), .ZN(n20404) );
  IOA21HSV4 U23118 ( .A1(n23460), .A2(n20403), .B(n20404), .ZN(n20444) );
  NAND2HSV0 U23119 ( .A1(n28629), .A2(\pe11/got [8]), .ZN(n20405) );
  XNOR2HSV1 U23120 ( .A1(n20406), .A2(n20405), .ZN(n20430) );
  NAND2HSV0 U23121 ( .A1(n24975), .A2(\pe11/got [7]), .ZN(n20407) );
  XNOR2HSV1 U23122 ( .A1(n20407), .A2(\pe11/phq [10]), .ZN(n20410) );
  BUFHSV2 U23123 ( .I(n20470), .Z(n24980) );
  NAND2HSV2 U23124 ( .A1(n24980), .A2(\pe11/pvq [10]), .ZN(n20409) );
  XNOR2HSV1 U23125 ( .A1(n20410), .A2(n20409), .ZN(n20428) );
  NAND2HSV0 U23126 ( .A1(\pe11/bq[10] ), .A2(n12011), .ZN(n20412) );
  NAND2HSV0 U23127 ( .A1(\pe11/bq[9] ), .A2(n24771), .ZN(n20411) );
  XOR2HSV0 U23128 ( .A1(n20412), .A2(n20411), .Z(n20416) );
  NAND2HSV0 U23129 ( .A1(n24997), .A2(\pe11/aot [8]), .ZN(n20414) );
  NAND2HSV0 U23130 ( .A1(\pe11/bq[12] ), .A2(\pe11/aot [11]), .ZN(n20413) );
  XOR2HSV0 U23131 ( .A1(n20414), .A2(n20413), .Z(n20415) );
  XOR2HSV0 U23132 ( .A1(n20416), .A2(n20415), .Z(n20427) );
  NAND2HSV0 U23133 ( .A1(\pe11/bq[13] ), .A2(\pe11/aot [10]), .ZN(n20418) );
  NAND2HSV0 U23134 ( .A1(n27058), .A2(\pe11/aot [7]), .ZN(n20417) );
  XOR2HSV0 U23135 ( .A1(n20418), .A2(n20417), .Z(n20426) );
  NAND2HSV0 U23136 ( .A1(\pe11/bq[14] ), .A2(\pe11/aot [9]), .ZN(n20420) );
  NAND2HSV0 U23137 ( .A1(\pe11/bq[11] ), .A2(\pe11/aot [12]), .ZN(n20419) );
  XOR2HSV0 U23138 ( .A1(n20420), .A2(n20419), .Z(n20424) );
  BUFHSV2 U23139 ( .I(\pe11/aot [15]), .Z(n24994) );
  NAND2HSV0 U23140 ( .A1(\pe11/bq[8] ), .A2(n24994), .ZN(n20422) );
  NAND2HSV0 U23141 ( .A1(\pe11/bq[7] ), .A2(n20157), .ZN(n20421) );
  XOR2HSV0 U23142 ( .A1(n20422), .A2(n20421), .Z(n20423) );
  XOR2HSV0 U23143 ( .A1(n20424), .A2(n20423), .Z(n20425) );
  XOR4HSV1 U23144 ( .A1(n20428), .A2(n20427), .A3(n20426), .A4(n20425), .Z(
        n20429) );
  XNOR2HSV1 U23145 ( .A1(n20430), .A2(n20429), .ZN(n20433) );
  INHSV2 U23146 ( .I(n28807), .ZN(n20536) );
  CLKNHSV0 U23147 ( .I(n20536), .ZN(n20431) );
  NAND2HSV0 U23148 ( .A1(n20431), .A2(\pe11/got [10]), .ZN(n20432) );
  XNOR2HSV1 U23149 ( .A1(n20433), .A2(n20432), .ZN(n20435) );
  NAND2HSV0 U23150 ( .A1(n14043), .A2(n14049), .ZN(n20436) );
  XNOR2HSV4 U23151 ( .A1(n20437), .A2(n20436), .ZN(n20442) );
  NOR2HSV0 U23152 ( .A1(n20464), .A2(n20229), .ZN(n20439) );
  NAND3HSV2 U23153 ( .A1(n20438), .A2(n20440), .A3(n20439), .ZN(n20441) );
  XNOR2HSV4 U23154 ( .A1(n20442), .A2(n20441), .ZN(n20443) );
  XNOR2HSV4 U23155 ( .A1(n20444), .A2(n20443), .ZN(n20560) );
  INHSV2 U23156 ( .I(n20559), .ZN(n25032) );
  INHSV2 U23157 ( .I(n25032), .ZN(n20463) );
  CLKNAND2HSV3 U23158 ( .A1(n20446), .A2(n20463), .ZN(n20547) );
  CLKNAND2HSV1 U23159 ( .A1(n20547), .A2(n20463), .ZN(n20447) );
  INHSV2 U23160 ( .I(n20447), .ZN(n20449) );
  CLKNAND2HSV1 U23161 ( .A1(n20449), .A2(n20448), .ZN(n20455) );
  INHSV2 U23162 ( .I(n20636), .ZN(n23470) );
  OAI21HSV2 U23163 ( .A1(\pe11/ti_7t [8]), .A2(n20698), .B(n20565), .ZN(n20451) );
  AOI21HSV2 U23164 ( .A1(n20453), .A2(n20452), .B(n20451), .ZN(n20454) );
  AOI22HSV2 U23165 ( .A1(n25504), .A2(n20458), .B1(n20457), .B2(n20456), .ZN(
        n20498) );
  CLKBUFHSV4 U23166 ( .I(n20459), .Z(n20460) );
  MUX2NHSV4 U23167 ( .I0(n20462), .I1(n20461), .S(n20460), .ZN(n25516) );
  CLKNHSV0 U23168 ( .I(n21785), .ZN(n20466) );
  OR2HSV1 U23169 ( .A1(n20464), .A2(n25028), .Z(n20465) );
  AOI21HSV4 U23170 ( .A1(n25516), .A2(n20466), .B(n20465), .ZN(n20496) );
  NAND2HSV2 U23171 ( .A1(n20467), .A2(n14049), .ZN(n20492) );
  NAND2HSV0 U23172 ( .A1(n20505), .A2(\pe11/got [10]), .ZN(n20469) );
  CLKNAND2HSV0 U23173 ( .A1(n28629), .A2(\pe11/got [9]), .ZN(n20468) );
  CLKNAND2HSV0 U23174 ( .A1(\pe11/aot [14]), .A2(\pe11/bq[10] ), .ZN(n24770)
         );
  NAND2HSV0 U23175 ( .A1(n20470), .A2(\pe11/pvq [9]), .ZN(n20471) );
  XOR2HSV0 U23176 ( .A1(n24770), .A2(n20471), .Z(n20481) );
  NAND2HSV0 U23177 ( .A1(\pe11/bq[9] ), .A2(n24994), .ZN(n20473) );
  NAND2HSV0 U23178 ( .A1(\pe11/bq[14] ), .A2(\pe11/aot [10]), .ZN(n20472) );
  XOR2HSV0 U23179 ( .A1(n20473), .A2(n20472), .Z(n20480) );
  INHSV2 U23180 ( .I(\pe11/aot [8]), .ZN(n20811) );
  NOR2HSV1 U23181 ( .A1(n20326), .A2(n20811), .ZN(n20475) );
  NAND2HSV0 U23182 ( .A1(n24997), .A2(\pe11/aot [9]), .ZN(n20474) );
  XOR2HSV0 U23183 ( .A1(n20475), .A2(n20474), .Z(n20478) );
  NAND2HSV0 U23184 ( .A1(n20587), .A2(\pe11/got [8]), .ZN(n20476) );
  XOR2HSV0 U23185 ( .A1(n20476), .A2(\pe11/phq [9]), .Z(n20477) );
  XOR2HSV0 U23186 ( .A1(n20478), .A2(n20477), .Z(n20479) );
  XOR3HSV2 U23187 ( .A1(n20481), .A2(n20480), .A3(n20479), .Z(n20487) );
  NAND2HSV0 U23188 ( .A1(\pe11/bq[13] ), .A2(\pe11/aot [11]), .ZN(n20483) );
  NAND2HSV0 U23189 ( .A1(\pe11/bq[11] ), .A2(n12011), .ZN(n20482) );
  XOR2HSV0 U23190 ( .A1(n20483), .A2(n20482), .Z(n20485) );
  NAND2HSV0 U23191 ( .A1(\pe11/bq[8] ), .A2(n20157), .ZN(n20731) );
  NAND2HSV0 U23192 ( .A1(\pe11/bq[12] ), .A2(\pe11/aot [12]), .ZN(n20711) );
  XNOR2HSV1 U23193 ( .A1(n20731), .A2(n20711), .ZN(n20484) );
  XNOR2HSV1 U23194 ( .A1(n20485), .A2(n20484), .ZN(n20486) );
  XNOR2HSV1 U23195 ( .A1(n20487), .A2(n20486), .ZN(n20488) );
  NAND2HSV0 U23196 ( .A1(n28807), .A2(\pe11/got [11]), .ZN(n20489) );
  XNOR2HSV4 U23197 ( .A1(n20490), .A2(n20489), .ZN(n20491) );
  XNOR2HSV4 U23198 ( .A1(n20492), .A2(n20491), .ZN(n20494) );
  NAND2HSV0 U23199 ( .A1(n28668), .A2(n20707), .ZN(n20493) );
  XOR2HSV2 U23200 ( .A1(n20494), .A2(n20493), .Z(n20495) );
  XNOR2HSV4 U23201 ( .A1(n20496), .A2(n20495), .ZN(n20497) );
  XNOR2HSV4 U23202 ( .A1(n20498), .A2(n20497), .ZN(n20500) );
  NAND2HSV2 U23203 ( .A1(n20499), .A2(n20500), .ZN(n20504) );
  INHSV3 U23204 ( .I(n20500), .ZN(n20501) );
  CLKNAND2HSV4 U23205 ( .A1(n20504), .A2(n20503), .ZN(n20611) );
  NAND2HSV2 U23206 ( .A1(n23470), .A2(\pe11/ti_7t [9]), .ZN(n20690) );
  XNOR2HSV4 U23207 ( .A1(n20693), .A2(n20691), .ZN(n20630) );
  NAND2HSV2 U23208 ( .A1(n20562), .A2(n25488), .ZN(n20629) );
  AOI21HSV4 U23209 ( .A1(n20630), .A2(n25512), .B(n20629), .ZN(n20628) );
  INHSV2 U23210 ( .I(n20505), .ZN(n20568) );
  NAND2HSV0 U23211 ( .A1(n20506), .A2(\pe11/got [8]), .ZN(n20508) );
  NAND2HSV0 U23212 ( .A1(n25489), .A2(\pe11/got [7]), .ZN(n20507) );
  XOR2HSV0 U23213 ( .A1(n20508), .A2(n20507), .Z(n20535) );
  NAND2HSV0 U23214 ( .A1(n24994), .A2(\pe11/bq[7] ), .ZN(n20510) );
  NAND2HSV0 U23215 ( .A1(\pe11/aot [10]), .A2(\pe11/bq[12] ), .ZN(n20509) );
  XOR2HSV0 U23216 ( .A1(n20510), .A2(n20509), .Z(n20514) );
  NAND2HSV0 U23217 ( .A1(n27058), .A2(\pe11/aot [6]), .ZN(n20512) );
  NAND2HSV0 U23218 ( .A1(\pe11/bq[13] ), .A2(\pe11/aot [9]), .ZN(n20511) );
  XOR2HSV0 U23219 ( .A1(n20512), .A2(n20511), .Z(n20513) );
  XOR2HSV0 U23220 ( .A1(n20514), .A2(n20513), .Z(n20522) );
  NAND2HSV0 U23221 ( .A1(\pe11/bq[8] ), .A2(n24771), .ZN(n20516) );
  NAND2HSV0 U23222 ( .A1(\pe11/bq[14] ), .A2(\pe11/aot [8]), .ZN(n20515) );
  XOR2HSV0 U23223 ( .A1(n20516), .A2(n20515), .Z(n20520) );
  NAND2HSV0 U23224 ( .A1(\pe11/bq[11] ), .A2(\pe11/aot [11]), .ZN(n20518) );
  NAND2HSV0 U23225 ( .A1(\pe11/bq[10] ), .A2(\pe11/aot [12]), .ZN(n20517) );
  XOR2HSV0 U23226 ( .A1(n20518), .A2(n20517), .Z(n20519) );
  XOR2HSV0 U23227 ( .A1(n20520), .A2(n20519), .Z(n20521) );
  XOR2HSV0 U23228 ( .A1(n20522), .A2(n20521), .Z(n20533) );
  NAND2HSV0 U23229 ( .A1(n24997), .A2(\pe11/aot [7]), .ZN(n20524) );
  NAND2HSV0 U23230 ( .A1(n20157), .A2(\pe11/bq[6] ), .ZN(n20523) );
  XOR2HSV0 U23231 ( .A1(n20524), .A2(n20523), .Z(n20527) );
  NAND2HSV0 U23232 ( .A1(n20587), .A2(\pe11/got [6]), .ZN(n20525) );
  XNOR2HSV1 U23233 ( .A1(n20525), .A2(\pe11/phq [11]), .ZN(n20526) );
  XNOR2HSV1 U23234 ( .A1(n20527), .A2(n20526), .ZN(n20531) );
  CLKNAND2HSV1 U23235 ( .A1(n20650), .A2(\pe11/pvq [11]), .ZN(n20529) );
  NAND2HSV0 U23236 ( .A1(\pe11/bq[9] ), .A2(n12011), .ZN(n20528) );
  XOR2HSV0 U23237 ( .A1(n20529), .A2(n20528), .Z(n20530) );
  XNOR2HSV1 U23238 ( .A1(n20531), .A2(n20530), .ZN(n20532) );
  XNOR2HSV1 U23239 ( .A1(n20533), .A2(n20532), .ZN(n20534) );
  XOR2HSV0 U23240 ( .A1(n20535), .A2(n20534), .Z(n20538) );
  INHSV2 U23241 ( .I(n20536), .ZN(n25008) );
  NAND2HSV0 U23242 ( .A1(n25008), .A2(\pe11/got [9]), .ZN(n20537) );
  XNOR2HSV1 U23243 ( .A1(n20538), .A2(n20537), .ZN(n20540) );
  CLKNAND2HSV1 U23244 ( .A1(n20467), .A2(\pe11/got [10]), .ZN(n20539) );
  XNOR2HSV1 U23245 ( .A1(n20540), .A2(n20539), .ZN(n20542) );
  NAND2HSV0 U23246 ( .A1(n11852), .A2(\pe11/got [11]), .ZN(n20541) );
  XOR2HSV0 U23247 ( .A1(n20542), .A2(n20541), .Z(n20550) );
  CLKNAND2HSV1 U23248 ( .A1(n25516), .A2(n20543), .ZN(n20546) );
  CLKNHSV0 U23249 ( .I(\pe11/ti_7t [6]), .ZN(n20544) );
  CLKNAND2HSV1 U23250 ( .A1(n21785), .A2(n20544), .ZN(n20545) );
  NAND2HSV2 U23251 ( .A1(n20546), .A2(n20545), .ZN(n20708) );
  INHSV2 U23252 ( .I(n20708), .ZN(n20784) );
  NAND2HSV2 U23253 ( .A1(n20784), .A2(n14049), .ZN(n20549) );
  NAND2HSV2 U23254 ( .A1(n20547), .A2(n20403), .ZN(n28791) );
  NAND2HSV2 U23255 ( .A1(n28791), .A2(n20227), .ZN(n20548) );
  XOR3HSV2 U23256 ( .A1(n20550), .A2(n20549), .A3(n20548), .Z(n20555) );
  INHSV2 U23257 ( .I(n20552), .ZN(n20608) );
  AOI21HSV2 U23258 ( .A1(n20552), .A2(n20637), .B(n25028), .ZN(n20553) );
  OAI21HSV2 U23259 ( .A1(n23458), .A2(n20608), .B(n20553), .ZN(n20554) );
  XNOR2HSV4 U23260 ( .A1(n20555), .A2(n20554), .ZN(n20558) );
  XNOR2HSV4 U23261 ( .A1(n20628), .A2(n20631), .ZN(n20639) );
  CLKNAND2HSV3 U23262 ( .A1(n23458), .A2(n20559), .ZN(n20682) );
  XNOR2HSV4 U23263 ( .A1(n20560), .A2(n20682), .ZN(n20622) );
  NOR2HSV2 U23264 ( .A1(n20561), .A2(ctro11), .ZN(n20621) );
  NAND2HSV2 U23265 ( .A1(n20622), .A2(n20621), .ZN(n20564) );
  INHSV2 U23266 ( .I(n20624), .ZN(n20563) );
  NOR2HSV3 U23267 ( .A1(n20639), .A2(n20566), .ZN(n20618) );
  INHSV2 U23268 ( .I(n28791), .ZN(n21910) );
  INHSV2 U23269 ( .I(n21910), .ZN(n20783) );
  NAND2HSV0 U23270 ( .A1(n20783), .A2(n14049), .ZN(n20607) );
  NAND2HSV0 U23271 ( .A1(n20784), .A2(\pe11/got [11]), .ZN(n20605) );
  NAND2HSV0 U23272 ( .A1(n20506), .A2(\pe11/got [7]), .ZN(n20570) );
  NAND2HSV0 U23273 ( .A1(n28629), .A2(\pe11/got [6]), .ZN(n20569) );
  XOR2HSV0 U23274 ( .A1(n20570), .A2(n20569), .Z(n20596) );
  NAND2HSV0 U23275 ( .A1(n27058), .A2(\pe11/aot [5]), .ZN(n20572) );
  NAND2HSV0 U23276 ( .A1(\pe11/bq[5] ), .A2(n20157), .ZN(n20571) );
  XOR2HSV0 U23277 ( .A1(n20572), .A2(n20571), .Z(n20576) );
  NAND2HSV0 U23278 ( .A1(n24997), .A2(\pe11/aot [6]), .ZN(n20574) );
  NAND2HSV0 U23279 ( .A1(\pe11/bq[11] ), .A2(\pe11/aot [10]), .ZN(n20573) );
  XOR2HSV0 U23280 ( .A1(n20574), .A2(n20573), .Z(n20575) );
  XOR2HSV0 U23281 ( .A1(n20576), .A2(n20575), .Z(n20584) );
  NAND2HSV0 U23282 ( .A1(\pe11/bq[7] ), .A2(n24771), .ZN(n20578) );
  NAND2HSV0 U23283 ( .A1(\pe11/bq[8] ), .A2(n12011), .ZN(n20577) );
  XOR2HSV0 U23284 ( .A1(n20578), .A2(n20577), .Z(n20582) );
  NAND2HSV0 U23285 ( .A1(n20650), .A2(\pe11/pvq [12]), .ZN(n20580) );
  NAND2HSV0 U23286 ( .A1(\pe11/bq[10] ), .A2(\pe11/aot [11]), .ZN(n20579) );
  XOR2HSV0 U23287 ( .A1(n20580), .A2(n20579), .Z(n20581) );
  XOR2HSV0 U23288 ( .A1(n20582), .A2(n20581), .Z(n20583) );
  XOR2HSV0 U23289 ( .A1(n20584), .A2(n20583), .Z(n20594) );
  NAND2HSV0 U23290 ( .A1(\pe11/bq[13] ), .A2(\pe11/aot [8]), .ZN(n20586) );
  NAND2HSV0 U23291 ( .A1(\pe11/bq[6] ), .A2(n24994), .ZN(n20585) );
  XOR2HSV0 U23292 ( .A1(n20586), .A2(n20585), .Z(n20590) );
  NAND2HSV0 U23293 ( .A1(n20587), .A2(\pe11/got [5]), .ZN(n20588) );
  XNOR2HSV1 U23294 ( .A1(n20588), .A2(\pe11/phq [12]), .ZN(n20589) );
  XNOR2HSV1 U23295 ( .A1(n20590), .A2(n20589), .ZN(n20592) );
  NAND2HSV0 U23296 ( .A1(\pe11/bq[9] ), .A2(\pe11/aot [9]), .ZN(n20786) );
  NAND2HSV0 U23297 ( .A1(\pe11/bq[14] ), .A2(\pe11/aot [7]), .ZN(n24765) );
  XNOR2HSV1 U23298 ( .A1(n20592), .A2(n20591), .ZN(n20593) );
  XNOR2HSV1 U23299 ( .A1(n20594), .A2(n20593), .ZN(n20595) );
  XOR2HSV0 U23300 ( .A1(n20596), .A2(n20595), .Z(n20598) );
  NAND2HSV0 U23301 ( .A1(n25008), .A2(\pe11/got [8]), .ZN(n20597) );
  XNOR2HSV1 U23302 ( .A1(n20598), .A2(n20597), .ZN(n20600) );
  CLKNAND2HSV0 U23303 ( .A1(n20467), .A2(\pe11/got [9]), .ZN(n20599) );
  XNOR2HSV1 U23304 ( .A1(n20600), .A2(n20599), .ZN(n20603) );
  NAND2HSV0 U23305 ( .A1(n14043), .A2(\pe11/got [10]), .ZN(n20602) );
  XOR2HSV0 U23306 ( .A1(n20603), .A2(n20602), .Z(n20604) );
  XOR2HSV0 U23307 ( .A1(n20605), .A2(n20604), .Z(n20606) );
  XOR2HSV0 U23308 ( .A1(n20607), .A2(n20606), .Z(n20610) );
  INHSV2 U23309 ( .I(n20608), .ZN(n20681) );
  NAND2HSV2 U23310 ( .A1(n20682), .A2(n20681), .ZN(n28935) );
  CLKNAND2HSV1 U23311 ( .A1(n28935), .A2(n20707), .ZN(n20609) );
  XNOR2HSV1 U23312 ( .A1(n20610), .A2(n20609), .ZN(n20615) );
  CLKBUFHSV4 U23313 ( .I(n20611), .Z(n20685) );
  INHSV2 U23314 ( .I(n20687), .ZN(n20612) );
  OAI21HSV4 U23315 ( .A1(n20685), .A2(n20308), .B(n20612), .ZN(n21787) );
  BUFHSV2 U23316 ( .I(n20613), .Z(n25030) );
  NAND2HSV2 U23317 ( .A1(n21787), .A2(n25030), .ZN(n20614) );
  XNOR2HSV4 U23318 ( .A1(n20615), .A2(n20614), .ZN(n23452) );
  CLKNAND2HSV1 U23319 ( .A1(n20616), .A2(n23452), .ZN(n20617) );
  NOR2HSV4 U23320 ( .A1(n20618), .A2(n20617), .ZN(n20760) );
  NOR2HSV0 U23321 ( .A1(n20620), .A2(n20619), .ZN(n20778) );
  CLKNAND2HSV1 U23322 ( .A1(n20622), .A2(n20621), .ZN(n20626) );
  NAND2HSV0 U23323 ( .A1(n20624), .A2(n20623), .ZN(n20625) );
  CLKNAND2HSV1 U23324 ( .A1(n20626), .A2(n20625), .ZN(n20627) );
  NAND2HSV2 U23325 ( .A1(n20637), .A2(\pe11/ti_7t [12]), .ZN(n20633) );
  AO21HSV1 U23326 ( .A1(n20630), .A2(n25512), .B(n20629), .Z(n20632) );
  CLKAND2HSV1 U23327 ( .A1(n23451), .A2(n20565), .Z(n20634) );
  CLKAND2HSV2 U23328 ( .A1(n20634), .A2(n20633), .Z(n20635) );
  INHSV2 U23329 ( .I(n23450), .ZN(n20782) );
  AOI21HSV2 U23330 ( .A1(n20782), .A2(n20637), .B(n20372), .ZN(n20638) );
  OAI21HSV4 U23331 ( .A1(n20639), .A2(n23450), .B(n20638), .ZN(n20700) );
  NAND2HSV0 U23332 ( .A1(n20783), .A2(\pe11/got [11]), .ZN(n20680) );
  NAND2HSV0 U23333 ( .A1(n20784), .A2(\pe11/got [10]), .ZN(n20678) );
  NAND2HSV0 U23334 ( .A1(n20506), .A2(\pe11/got [6]), .ZN(n20641) );
  NAND2HSV0 U23335 ( .A1(n28629), .A2(\pe11/got [5]), .ZN(n20640) );
  XOR2HSV0 U23336 ( .A1(n20641), .A2(n20640), .Z(n20670) );
  NAND2HSV0 U23337 ( .A1(\pe11/bq[7] ), .A2(n12011), .ZN(n20643) );
  NAND2HSV0 U23338 ( .A1(n27058), .A2(\pe11/aot [4]), .ZN(n20642) );
  XOR2HSV0 U23339 ( .A1(n20643), .A2(n20642), .Z(n20647) );
  NAND2HSV0 U23340 ( .A1(\pe11/bq[11] ), .A2(\pe11/aot [9]), .ZN(n20645) );
  NAND2HSV0 U23341 ( .A1(\pe11/bq[13] ), .A2(\pe11/aot [7]), .ZN(n20644) );
  XOR2HSV0 U23342 ( .A1(n20645), .A2(n20644), .Z(n20646) );
  XOR2HSV0 U23343 ( .A1(n20647), .A2(n20646), .Z(n20656) );
  NAND2HSV0 U23344 ( .A1(\pe11/bq[6] ), .A2(n24771), .ZN(n20649) );
  NAND2HSV0 U23345 ( .A1(n20157), .A2(\pe11/bq[4] ), .ZN(n20648) );
  XOR2HSV0 U23346 ( .A1(n20649), .A2(n20648), .Z(n20654) );
  NAND2HSV0 U23347 ( .A1(n20650), .A2(\pe11/pvq [13]), .ZN(n20652) );
  NAND2HSV0 U23348 ( .A1(\pe11/bq[8] ), .A2(\pe11/aot [12]), .ZN(n20651) );
  XOR2HSV0 U23349 ( .A1(n20652), .A2(n20651), .Z(n20653) );
  XOR2HSV0 U23350 ( .A1(n20654), .A2(n20653), .Z(n20655) );
  XOR2HSV0 U23351 ( .A1(n20656), .A2(n20655), .Z(n20668) );
  XNOR2HSV1 U23352 ( .A1(n20658), .A2(n20657), .ZN(n20666) );
  NAND2HSV0 U23353 ( .A1(n24975), .A2(\pe11/got [4]), .ZN(n20659) );
  XOR2HSV0 U23354 ( .A1(n20659), .A2(\pe11/phq [13]), .Z(n20664) );
  INHSV2 U23355 ( .I(\pe11/bq[5] ), .ZN(n20714) );
  CLKNHSV0 U23356 ( .I(\pe11/aot [10]), .ZN(n20660) );
  NOR2HSV0 U23357 ( .A1(n20714), .A2(n20660), .ZN(n21932) );
  AOI22HSV0 U23358 ( .A1(n24994), .A2(\pe11/bq[5] ), .B1(\pe11/bq[10] ), .B2(
        \pe11/aot [10]), .ZN(n20661) );
  AOI21HSV0 U23359 ( .A1(n20662), .A2(n21932), .B(n20661), .ZN(n20663) );
  XOR2HSV0 U23360 ( .A1(n20664), .A2(n20663), .Z(n20665) );
  XNOR2HSV1 U23361 ( .A1(n20666), .A2(n20665), .ZN(n20667) );
  XNOR2HSV1 U23362 ( .A1(n20668), .A2(n20667), .ZN(n20669) );
  XOR2HSV0 U23363 ( .A1(n20670), .A2(n20669), .Z(n20672) );
  NAND2HSV0 U23364 ( .A1(n25008), .A2(\pe11/got [7]), .ZN(n20671) );
  XNOR2HSV1 U23365 ( .A1(n20672), .A2(n20671), .ZN(n20674) );
  NAND2HSV0 U23366 ( .A1(n24966), .A2(\pe11/got [8]), .ZN(n20673) );
  XNOR2HSV1 U23367 ( .A1(n20674), .A2(n20673), .ZN(n20676) );
  NAND2HSV0 U23368 ( .A1(n11852), .A2(\pe11/got [9]), .ZN(n20675) );
  XOR2HSV0 U23369 ( .A1(n20676), .A2(n20675), .Z(n20677) );
  XOR2HSV0 U23370 ( .A1(n20678), .A2(n20677), .Z(n20679) );
  XNOR2HSV1 U23371 ( .A1(n20680), .A2(n20679), .ZN(n20684) );
  CLKNAND2HSV3 U23372 ( .A1(n20682), .A2(n20681), .ZN(n25138) );
  NAND2HSV0 U23373 ( .A1(n25138), .A2(n14049), .ZN(n20683) );
  INHSV2 U23374 ( .I(n20685), .ZN(n23457) );
  AOI21HSV0 U23375 ( .A1(n20690), .A2(n23470), .B(n20229), .ZN(n20686) );
  OAI21HSV2 U23376 ( .A1(n23457), .A2(n20687), .B(n20686), .ZN(n20688) );
  AOI21HSV0 U23377 ( .A1(n20690), .A2(n25032), .B(n20689), .ZN(n20692) );
  NAND2HSV2 U23378 ( .A1(\pe11/ti_7t [10]), .A2(n20770), .ZN(n20694) );
  INHSV2 U23379 ( .I(n20694), .ZN(n20706) );
  AOI21HSV2 U23380 ( .A1(n20694), .A2(n25032), .B(n25028), .ZN(n20695) );
  OAI21HSV4 U23381 ( .A1(n25352), .A2(n20706), .B(n20695), .ZN(n20696) );
  XNOR2HSV4 U23382 ( .A1(n20697), .A2(n20696), .ZN(n20699) );
  XNOR2HSV4 U23383 ( .A1(n20700), .A2(n20699), .ZN(n21734) );
  NOR2HSV4 U23384 ( .A1(n21734), .A2(n20770), .ZN(n20702) );
  INAND2HSV4 U23385 ( .A1(n20760), .B1(n20761), .ZN(n25026) );
  INHSV2 U23386 ( .I(\pe11/ti_7t [13]), .ZN(n21784) );
  NAND2HSV2 U23387 ( .A1(n21784), .A2(n20637), .ZN(n25029) );
  CLKNAND2HSV1 U23388 ( .A1(n25029), .A2(n25488), .ZN(n20701) );
  CLKNHSV0 U23389 ( .I(n20782), .ZN(n20705) );
  CLKNHSV0 U23390 ( .I(\pe11/got [14]), .ZN(n25028) );
  AOI21HSV2 U23391 ( .A1(n20782), .A2(n21785), .B(n25028), .ZN(n20704) );
  OAI21HSV2 U23392 ( .A1(n20705), .A2(n23454), .B(n20704), .ZN(n20759) );
  NAND2HSV0 U23393 ( .A1(n28935), .A2(\pe11/got [11]), .ZN(n20753) );
  NAND2HSV0 U23394 ( .A1(n20783), .A2(\pe11/got [10]), .ZN(n20751) );
  INHSV2 U23395 ( .I(n20708), .ZN(n28471) );
  NAND2HSV0 U23396 ( .A1(n20506), .A2(\pe11/got [5]), .ZN(n20723) );
  NAND2HSV0 U23397 ( .A1(\pe11/bq[14] ), .A2(\pe11/aot [5]), .ZN(n20710) );
  NAND2HSV0 U23398 ( .A1(\pe11/bq[13] ), .A2(\pe11/aot [6]), .ZN(n20709) );
  XOR2HSV0 U23399 ( .A1(n20710), .A2(n20709), .Z(n20721) );
  NAND2HSV0 U23400 ( .A1(\pe11/aot [7]), .A2(\pe11/bq[7] ), .ZN(n24715) );
  NAND2HSV0 U23401 ( .A1(\pe11/bq[11] ), .A2(\pe11/aot [8]), .ZN(n20713) );
  NAND2HSV0 U23402 ( .A1(n24994), .A2(\pe11/bq[4] ), .ZN(n20712) );
  XOR2HSV0 U23403 ( .A1(n20713), .A2(n20712), .Z(n20718) );
  INHSV2 U23404 ( .I(n20714), .ZN(n22106) );
  NAND2HSV0 U23405 ( .A1(n22106), .A2(n24771), .ZN(n20716) );
  NAND2HSV0 U23406 ( .A1(\pe11/bq[6] ), .A2(n12011), .ZN(n20715) );
  XOR2HSV0 U23407 ( .A1(n20716), .A2(n20715), .Z(n20717) );
  XOR2HSV0 U23408 ( .A1(n20718), .A2(n20717), .Z(n20719) );
  XOR3HSV2 U23409 ( .A1(n20721), .A2(n20720), .A3(n20719), .Z(n20722) );
  XNOR2HSV1 U23410 ( .A1(n20723), .A2(n20722), .ZN(n20741) );
  NAND2HSV0 U23411 ( .A1(\pe11/aot [3]), .A2(\pe11/bq[16] ), .ZN(n20725) );
  NAND2HSV0 U23412 ( .A1(\pe11/bq[9] ), .A2(\pe11/aot [10]), .ZN(n20724) );
  XOR2HSV0 U23413 ( .A1(n20725), .A2(n20724), .Z(n20729) );
  NAND2HSV0 U23414 ( .A1(n24997), .A2(\pe11/aot [4]), .ZN(n20727) );
  NAND2HSV0 U23415 ( .A1(\pe11/bq[10] ), .A2(\pe11/aot [9]), .ZN(n20726) );
  XOR2HSV0 U23416 ( .A1(n20727), .A2(n20726), .Z(n20728) );
  XOR2HSV0 U23417 ( .A1(n20729), .A2(n20728), .Z(n20737) );
  NAND2HSV0 U23418 ( .A1(n24975), .A2(\pe11/got [3]), .ZN(n20730) );
  XNOR2HSV1 U23419 ( .A1(n20730), .A2(\pe11/phq [14]), .ZN(n20735) );
  NAND2HSV0 U23420 ( .A1(\pe11/bq[3] ), .A2(\pe11/aot [11]), .ZN(n24720) );
  NOR2HSV0 U23421 ( .A1(n20731), .A2(n24720), .ZN(n20733) );
  AOI22HSV0 U23422 ( .A1(\pe11/bq[8] ), .A2(\pe11/aot [11]), .B1(n20157), .B2(
        \pe11/bq[3] ), .ZN(n20732) );
  NOR2HSV2 U23423 ( .A1(n20733), .A2(n20732), .ZN(n20734) );
  XNOR2HSV1 U23424 ( .A1(n20735), .A2(n20734), .ZN(n20736) );
  XNOR2HSV1 U23425 ( .A1(n20737), .A2(n20736), .ZN(n20739) );
  NAND2HSV0 U23426 ( .A1(n25489), .A2(\pe11/got [4]), .ZN(n20738) );
  XOR2HSV0 U23427 ( .A1(n20739), .A2(n20738), .Z(n20740) );
  XNOR2HSV1 U23428 ( .A1(n20741), .A2(n20740), .ZN(n20743) );
  NAND2HSV0 U23429 ( .A1(n25008), .A2(\pe11/got [6]), .ZN(n20742) );
  XNOR2HSV1 U23430 ( .A1(n20743), .A2(n20742), .ZN(n20745) );
  NAND2HSV0 U23431 ( .A1(n20467), .A2(\pe11/got [7]), .ZN(n20744) );
  XOR2HSV0 U23432 ( .A1(n20745), .A2(n20744), .Z(n20747) );
  NAND2HSV0 U23433 ( .A1(n14043), .A2(\pe11/got [8]), .ZN(n20746) );
  XOR2HSV0 U23434 ( .A1(n20747), .A2(n20746), .Z(n20748) );
  XOR2HSV0 U23435 ( .A1(n20751), .A2(n20750), .Z(n20752) );
  CLKNAND2HSV0 U23436 ( .A1(n21787), .A2(\pe11/got [12]), .ZN(n20754) );
  XOR2HSV0 U23437 ( .A1(n20755), .A2(n20754), .Z(n20756) );
  CLKXOR2HSV2 U23438 ( .A1(n20757), .A2(n20756), .Z(n20758) );
  XNOR2HSV4 U23439 ( .A1(n20759), .A2(n20758), .ZN(n20762) );
  INHSV4 U23440 ( .I(n20760), .ZN(n20774) );
  INHSV3 U23441 ( .I(n20766), .ZN(n20763) );
  CLKNHSV0 U23442 ( .I(n20182), .ZN(n20767) );
  NOR2HSV2 U23443 ( .A1(n20768), .A2(n20767), .ZN(n20769) );
  NAND2HSV4 U23444 ( .A1(n20779), .A2(n20775), .ZN(n25034) );
  INHSV2 U23445 ( .I(n25034), .ZN(n25040) );
  INHSV2 U23446 ( .I(n20776), .ZN(n25045) );
  CLKNAND2HSV0 U23447 ( .A1(n25029), .A2(n25504), .ZN(n20777) );
  OAI21HSV2 U23448 ( .A1(n25040), .A2(n20781), .B(n20780), .ZN(n20846) );
  CLKNAND2HSV1 U23449 ( .A1(n21321), .A2(n14049), .ZN(n20836) );
  NAND2HSV0 U23450 ( .A1(n28935), .A2(\pe11/got [10]), .ZN(n20832) );
  NAND2HSV0 U23451 ( .A1(n20783), .A2(\pe11/got [9]), .ZN(n20830) );
  NAND2HSV0 U23452 ( .A1(n20784), .A2(\pe11/got [8]), .ZN(n20828) );
  NAND2HSV0 U23453 ( .A1(n25008), .A2(\pe11/got [5]), .ZN(n20824) );
  NAND2HSV0 U23454 ( .A1(n24980), .A2(\pe11/pvq [15]), .ZN(n20785) );
  XOR2HSV0 U23455 ( .A1(n20786), .A2(n20785), .Z(n20800) );
  NAND2HSV0 U23456 ( .A1(\pe11/bq[6] ), .A2(\pe11/aot [12]), .ZN(n20788) );
  NAND2HSV0 U23457 ( .A1(\pe11/bq[8] ), .A2(\pe11/aot [10]), .ZN(n20787) );
  XOR2HSV0 U23458 ( .A1(n20788), .A2(n20787), .Z(n20791) );
  NAND2HSV0 U23459 ( .A1(\pe11/bq[12] ), .A2(\pe11/aot [6]), .ZN(n20789) );
  XNOR2HSV1 U23460 ( .A1(n20789), .A2(\pe11/phq [15]), .ZN(n20790) );
  XNOR2HSV1 U23461 ( .A1(n20791), .A2(n20790), .ZN(n20799) );
  NAND2HSV0 U23462 ( .A1(\pe11/aot [2]), .A2(\pe11/bq[16] ), .ZN(n20793) );
  NAND2HSV0 U23463 ( .A1(\pe11/bq[14] ), .A2(\pe11/aot [4]), .ZN(n20792) );
  XOR2HSV0 U23464 ( .A1(n20793), .A2(n20792), .Z(n20797) );
  NAND2HSV0 U23465 ( .A1(\pe11/got [2]), .A2(n24975), .ZN(n20795) );
  NAND2HSV0 U23466 ( .A1(n24997), .A2(\pe11/aot [3]), .ZN(n20794) );
  XOR2HSV0 U23467 ( .A1(n20795), .A2(n20794), .Z(n20796) );
  XOR2HSV0 U23468 ( .A1(n20797), .A2(n20796), .Z(n20798) );
  XOR3HSV2 U23469 ( .A1(n20800), .A2(n20799), .A3(n20798), .Z(n20802) );
  NAND2HSV0 U23470 ( .A1(n20506), .A2(\pe11/got [4]), .ZN(n20801) );
  XNOR2HSV1 U23471 ( .A1(n20802), .A2(n20801), .ZN(n20821) );
  NAND2HSV0 U23472 ( .A1(\pe11/bq[7] ), .A2(\pe11/aot [11]), .ZN(n20804) );
  NAND2HSV0 U23473 ( .A1(\pe11/bq[13] ), .A2(\pe11/aot [5]), .ZN(n20803) );
  XOR2HSV0 U23474 ( .A1(n20804), .A2(n20803), .Z(n20808) );
  NAND2HSV0 U23475 ( .A1(\pe11/bq[11] ), .A2(\pe11/aot [7]), .ZN(n20806) );
  NAND2HSV0 U23476 ( .A1(\pe11/bq[3] ), .A2(n24994), .ZN(n20805) );
  XOR2HSV0 U23477 ( .A1(n20806), .A2(n20805), .Z(n20807) );
  XOR2HSV0 U23478 ( .A1(n20808), .A2(n20807), .Z(n20817) );
  NAND2HSV0 U23479 ( .A1(\pe11/bq[4] ), .A2(n24771), .ZN(n20810) );
  NAND2HSV0 U23480 ( .A1(\pe11/bq[5] ), .A2(n12011), .ZN(n20809) );
  XOR2HSV0 U23481 ( .A1(n20810), .A2(n20809), .Z(n20815) );
  NOR2HSV0 U23482 ( .A1(n20384), .A2(n20811), .ZN(n20813) );
  NAND2HSV0 U23483 ( .A1(\pe11/bq[2] ), .A2(n20157), .ZN(n20812) );
  XOR2HSV0 U23484 ( .A1(n20813), .A2(n20812), .Z(n20814) );
  XOR2HSV0 U23485 ( .A1(n20815), .A2(n20814), .Z(n20816) );
  XOR2HSV0 U23486 ( .A1(n20817), .A2(n20816), .Z(n20819) );
  NAND2HSV0 U23487 ( .A1(n25489), .A2(\pe11/got [3]), .ZN(n20818) );
  XNOR2HSV1 U23488 ( .A1(n20819), .A2(n20818), .ZN(n20820) );
  XNOR2HSV1 U23489 ( .A1(n20821), .A2(n20820), .ZN(n20823) );
  NAND2HSV0 U23490 ( .A1(n11804), .A2(\pe11/got [6]), .ZN(n20822) );
  XOR3HSV2 U23491 ( .A1(n20824), .A2(n20823), .A3(n20822), .Z(n20826) );
  NAND2HSV0 U23492 ( .A1(n11852), .A2(\pe11/got [7]), .ZN(n20825) );
  XOR2HSV0 U23493 ( .A1(n20826), .A2(n20825), .Z(n20827) );
  XOR2HSV0 U23494 ( .A1(n20828), .A2(n20827), .Z(n20829) );
  XOR2HSV0 U23495 ( .A1(n20830), .A2(n20829), .Z(n20831) );
  XNOR2HSV1 U23496 ( .A1(n20832), .A2(n20831), .ZN(n20834) );
  NAND2HSV0 U23497 ( .A1(n21787), .A2(\pe11/got [11]), .ZN(n20833) );
  XOR2HSV0 U23498 ( .A1(n20834), .A2(n20833), .Z(n20835) );
  XNOR2HSV1 U23499 ( .A1(n20836), .A2(n20835), .ZN(n20837) );
  CLKNHSV0 U23500 ( .I(n20837), .ZN(n20838) );
  NOR2HSV2 U23501 ( .A1(n20838), .A2(n20229), .ZN(n20839) );
  CLKBUFHSV4 U23502 ( .I(n28918), .Z(n24965) );
  CLKNAND2HSV1 U23503 ( .A1(n20839), .A2(n24965), .ZN(n20840) );
  NAND2HSV2 U23504 ( .A1(n13976), .A2(n20840), .ZN(n20842) );
  NAND2HSV2 U23505 ( .A1(n25026), .A2(n25030), .ZN(n20841) );
  CLKNAND2HSV3 U23506 ( .A1(n24883), .A2(n24884), .ZN(n20843) );
  NAND2HSV2 U23507 ( .A1(n24881), .A2(n20844), .ZN(n24887) );
  INHSV2 U23508 ( .I(n24887), .ZN(n20847) );
  XNOR2HSV4 U23509 ( .A1(n20845), .A2(n20846), .ZN(n25415) );
  INHSV2 U23510 ( .I(n20985), .ZN(n20850) );
  CLKNHSV0 U23511 ( .I(n20855), .ZN(n20852) );
  INAND2HSV2 U23512 ( .A1(n20983), .B1(n20985), .ZN(n20857) );
  NAND3HSV2 U23513 ( .A1(n20919), .A2(n20852), .A3(n20857), .ZN(n20853) );
  CLKNAND2HSV2 U23514 ( .A1(n20854), .A2(n20853), .ZN(n20864) );
  NOR2HSV0 U23515 ( .A1(n20855), .A2(n21345), .ZN(n20856) );
  CLKNAND2HSV1 U23516 ( .A1(n20857), .A2(n20856), .ZN(n20859) );
  INHSV2 U23517 ( .I(n20919), .ZN(n20858) );
  NOR2HSV2 U23518 ( .A1(n20859), .A2(n20858), .ZN(n20861) );
  NAND2HSV2 U23519 ( .A1(n20861), .A2(n20860), .ZN(n20863) );
  NAND3HSV4 U23520 ( .A1(n20864), .A2(n20863), .A3(n20862), .ZN(n23266) );
  XNOR2HSV4 U23521 ( .A1(n20865), .A2(n23266), .ZN(n20867) );
  CLKNAND2HSV1 U23522 ( .A1(n28989), .A2(n14526), .ZN(n20872) );
  NAND2HSV0 U23523 ( .A1(n20870), .A2(\pe5/ti_7t [8]), .ZN(n20871) );
  CLKNAND2HSV2 U23524 ( .A1(n20872), .A2(n20871), .ZN(n28800) );
  CLKAND2HSV2 U23525 ( .A1(n28800), .A2(\pe5/got [12]), .Z(n20915) );
  NAND2HSV2 U23526 ( .A1(n21523), .A2(n20977), .ZN(n20913) );
  NOR2HSV2 U23527 ( .A1(n20931), .A2(n24685), .ZN(n20909) );
  NAND2HSV0 U23528 ( .A1(n28614), .A2(n28645), .ZN(n20907) );
  NAND2HSV0 U23529 ( .A1(n28647), .A2(n28594), .ZN(n20874) );
  XNOR2HSV1 U23530 ( .A1(n20874), .A2(n20873), .ZN(n20904) );
  NAND2HSV0 U23531 ( .A1(\pe5/aot [8]), .A2(n23909), .ZN(n20876) );
  NAND2HSV0 U23532 ( .A1(n25626), .A2(\pe5/got [4]), .ZN(n20875) );
  XOR2HSV0 U23533 ( .A1(n20876), .A2(n20875), .Z(n20880) );
  NAND2HSV0 U23534 ( .A1(\pe5/aot [10]), .A2(\pe5/bq[10] ), .ZN(n20878) );
  NAND2HSV0 U23535 ( .A1(\pe5/aot [11]), .A2(\pe5/bq[9] ), .ZN(n20877) );
  XOR2HSV0 U23536 ( .A1(n20878), .A2(n20877), .Z(n20879) );
  XOR2HSV0 U23537 ( .A1(n20880), .A2(n20879), .Z(n20886) );
  XOR2HSV0 U23538 ( .A1(n21470), .A2(n20881), .Z(n20884) );
  NAND2HSV0 U23539 ( .A1(\pe5/bq[8] ), .A2(\pe5/aot [12]), .ZN(n20933) );
  INHSV2 U23540 ( .I(\pe5/bq[4] ), .ZN(n21532) );
  NAND2HSV0 U23541 ( .A1(n21488), .A2(\pe5/bq[4] ), .ZN(n20882) );
  XOR2HSV0 U23542 ( .A1(n20933), .A2(n20882), .Z(n20883) );
  XOR2HSV0 U23543 ( .A1(n20884), .A2(n20883), .Z(n20885) );
  XOR2HSV0 U23544 ( .A1(n20886), .A2(n20885), .Z(n20902) );
  NAND2HSV0 U23545 ( .A1(\pe5/aot [14]), .A2(\pe5/bq[6] ), .ZN(n20888) );
  NAND2HSV0 U23546 ( .A1(\pe5/aot [4]), .A2(n25349), .ZN(n20887) );
  XOR2HSV0 U23547 ( .A1(n20888), .A2(n20887), .Z(n20893) );
  NAND2HSV0 U23548 ( .A1(n21374), .A2(\pe5/aot [5]), .ZN(n20891) );
  INHSV2 U23549 ( .I(n20889), .ZN(n23507) );
  NAND2HSV0 U23550 ( .A1(\pe5/aot [6]), .A2(n23507), .ZN(n20890) );
  XOR2HSV0 U23551 ( .A1(n20891), .A2(n20890), .Z(n20892) );
  XOR2HSV0 U23552 ( .A1(n20893), .A2(n20892), .Z(n20900) );
  NAND2HSV0 U23553 ( .A1(\pe5/aot [13]), .A2(\pe5/bq[7] ), .ZN(n20895) );
  NAND2HSV0 U23554 ( .A1(\pe5/aot [7]), .A2(\pe5/bq[13] ), .ZN(n20894) );
  XOR2HSV0 U23555 ( .A1(n20895), .A2(n20894), .Z(n20898) );
  NAND2HSV0 U23556 ( .A1(n28682), .A2(\pe5/pvq [13]), .ZN(n20896) );
  XOR2HSV0 U23557 ( .A1(n20896), .A2(\pe5/phq [13]), .Z(n20897) );
  XOR2HSV0 U23558 ( .A1(n20898), .A2(n20897), .Z(n20899) );
  XOR2HSV0 U23559 ( .A1(n20900), .A2(n20899), .Z(n20901) );
  XOR2HSV0 U23560 ( .A1(n20902), .A2(n20901), .Z(n20903) );
  XOR2HSV0 U23561 ( .A1(n20904), .A2(n20903), .Z(n20906) );
  NOR2HSV0 U23562 ( .A1(n14630), .A2(n24683), .ZN(n20905) );
  XOR3HSV2 U23563 ( .A1(n20907), .A2(n20906), .A3(n20905), .Z(n20908) );
  XNOR2HSV1 U23564 ( .A1(n20909), .A2(n20908), .ZN(n20911) );
  NAND2HSV0 U23565 ( .A1(n21504), .A2(n24637), .ZN(n20910) );
  XOR2HSV0 U23566 ( .A1(n20911), .A2(n20910), .Z(n20912) );
  XNOR2HSV1 U23567 ( .A1(n20913), .A2(n20912), .ZN(n20914) );
  XNOR2HSV4 U23568 ( .A1(n20915), .A2(n20914), .ZN(n20923) );
  NAND2HSV0 U23569 ( .A1(n20987), .A2(\pe5/got [14]), .ZN(n20916) );
  NOR2HSV1 U23570 ( .A1(n20917), .A2(n20916), .ZN(n20918) );
  CLKNAND2HSV1 U23571 ( .A1(n20919), .A2(n20918), .ZN(n20921) );
  NOR2HSV2 U23572 ( .A1(n20921), .A2(n20920), .ZN(n20922) );
  XOR3HSV2 U23573 ( .A1(n20924), .A2(n20923), .A3(n20922), .Z(n20925) );
  INHSV2 U23574 ( .I(n20927), .ZN(n20929) );
  INHSV1 U23575 ( .I(n21338), .ZN(n21348) );
  CLKNAND2HSV0 U23576 ( .A1(n21348), .A2(n14482), .ZN(n20930) );
  CLKNAND2HSV1 U23577 ( .A1(\pe5/ti_7t [12]), .A2(n20870), .ZN(n21413) );
  INHSV2 U23578 ( .I(n21413), .ZN(n21423) );
  NAND2HSV0 U23579 ( .A1(n21465), .A2(n24637), .ZN(n20976) );
  NOR2HSV1 U23580 ( .A1(n20931), .A2(n24683), .ZN(n20972) );
  NAND2HSV0 U23581 ( .A1(n28682), .A2(\pe5/pvq [14]), .ZN(n20932) );
  XNOR2HSV1 U23582 ( .A1(n20932), .A2(\pe5/phq [14]), .ZN(n20937) );
  NAND2HSV0 U23583 ( .A1(\pe5/aot [11]), .A2(\pe5/bq[7] ), .ZN(n21356) );
  NOR2HSV1 U23584 ( .A1(n20933), .A2(n21356), .ZN(n20935) );
  AOI22HSV0 U23585 ( .A1(\pe5/aot [12]), .A2(\pe5/bq[7] ), .B1(\pe5/aot [11]), 
        .B2(\pe5/bq[8] ), .ZN(n20934) );
  NOR2HSV2 U23586 ( .A1(n20935), .A2(n20934), .ZN(n20936) );
  XNOR2HSV1 U23587 ( .A1(n20937), .A2(n20936), .ZN(n20946) );
  INAND2HSV0 U23588 ( .A1(n14766), .B1(\pe5/aot [7]), .ZN(n20938) );
  XOR2HSV0 U23589 ( .A1(n20939), .A2(n20938), .Z(n20943) );
  NAND2HSV0 U23590 ( .A1(\pe5/aot [3]), .A2(n25349), .ZN(n20941) );
  NAND2HSV0 U23591 ( .A1(\pe5/bq[5] ), .A2(\pe5/aot [14]), .ZN(n20940) );
  XOR2HSV0 U23592 ( .A1(n20941), .A2(n20940), .Z(n20942) );
  XOR2HSV0 U23593 ( .A1(n20943), .A2(n20942), .Z(n20945) );
  NOR2HSV0 U23594 ( .A1(n27191), .A2(n24414), .ZN(n20944) );
  XOR3HSV2 U23595 ( .A1(n20946), .A2(n20945), .A3(n20944), .Z(n20968) );
  NAND2HSV0 U23596 ( .A1(n14072), .A2(n28594), .ZN(n20965) );
  NAND2HSV0 U23597 ( .A1(\pe5/aot [10]), .A2(\pe5/bq[9] ), .ZN(n20948) );
  NAND2HSV0 U23598 ( .A1(\pe5/aot [4]), .A2(n24647), .ZN(n20947) );
  XOR2HSV0 U23599 ( .A1(n20948), .A2(n20947), .Z(n20952) );
  NAND2HSV0 U23600 ( .A1(\pe5/aot [5]), .A2(\pe5/bq[14] ), .ZN(n20950) );
  NAND2HSV0 U23601 ( .A1(\pe5/aot [13]), .A2(\pe5/bq[6] ), .ZN(n20949) );
  XOR2HSV0 U23602 ( .A1(n20950), .A2(n20949), .Z(n20951) );
  XOR2HSV0 U23603 ( .A1(n20952), .A2(n20951), .Z(n20963) );
  NAND2HSV0 U23604 ( .A1(\pe5/aot [6]), .A2(\pe5/bq[3] ), .ZN(n23255) );
  AOI22HSV0 U23605 ( .A1(n21488), .A2(\pe5/bq[3] ), .B1(\pe5/bq[13] ), .B2(
        \pe5/aot [6]), .ZN(n20954) );
  NOR2HSV2 U23606 ( .A1(n20955), .A2(n20954), .ZN(n20957) );
  NAND2HSV0 U23607 ( .A1(n14031), .A2(\pe5/bq[4] ), .ZN(n20956) );
  XNOR2HSV1 U23608 ( .A1(n20957), .A2(n20956), .ZN(n20961) );
  NAND2HSV0 U23609 ( .A1(\pe5/aot [8]), .A2(\pe5/bq[11] ), .ZN(n20959) );
  NAND2HSV0 U23610 ( .A1(\pe5/aot [9]), .A2(\pe5/bq[10] ), .ZN(n20958) );
  XOR2HSV0 U23611 ( .A1(n20959), .A2(n20958), .Z(n20960) );
  XOR2HSV0 U23612 ( .A1(n20961), .A2(n20960), .Z(n20962) );
  XOR2HSV0 U23613 ( .A1(n20963), .A2(n20962), .Z(n20964) );
  XNOR2HSV1 U23614 ( .A1(n20965), .A2(n20964), .ZN(n20967) );
  NAND2HSV0 U23615 ( .A1(n28614), .A2(n28647), .ZN(n20966) );
  XOR3HSV2 U23616 ( .A1(n20968), .A2(n20967), .A3(n20966), .Z(n20970) );
  NAND2HSV0 U23617 ( .A1(n24674), .A2(n28645), .ZN(n20969) );
  XNOR2HSV1 U23618 ( .A1(n20970), .A2(n20969), .ZN(n20971) );
  XNOR2HSV1 U23619 ( .A1(n20972), .A2(n20971), .ZN(n20974) );
  NAND2HSV0 U23620 ( .A1(n21504), .A2(n14069), .ZN(n20973) );
  XOR2HSV0 U23621 ( .A1(n20974), .A2(n20973), .Z(n20975) );
  XNOR2HSV1 U23622 ( .A1(n20976), .A2(n20975), .ZN(n20982) );
  CLKAND2HSV2 U23623 ( .A1(n28800), .A2(n20977), .Z(n20981) );
  INHSV2 U23624 ( .I(n20978), .ZN(n21554) );
  INHSV2 U23625 ( .I(n21554), .ZN(n21614) );
  NOR2HSV2 U23626 ( .A1(n24686), .A2(n20979), .ZN(n20980) );
  XOR3HSV2 U23627 ( .A1(n20982), .A2(n20981), .A3(n20980), .Z(n20991) );
  CLKNHSV0 U23628 ( .I(n20987), .ZN(n20988) );
  NOR2HSV2 U23629 ( .A1(n20988), .A2(n14544), .ZN(n20989) );
  XNOR2HSV4 U23630 ( .A1(n20991), .A2(n20990), .ZN(n20992) );
  INHSV2 U23631 ( .I(n20992), .ZN(n20993) );
  NAND2HSV2 U23632 ( .A1(n21159), .A2(\pe2/ti_7t [8]), .ZN(n21290) );
  INHSV2 U23633 ( .I(n21290), .ZN(n21292) );
  NAND2HSV4 U23634 ( .A1(n21005), .A2(n27123), .ZN(n21109) );
  CLKNAND2HSV2 U23635 ( .A1(n21006), .A2(n22085), .ZN(n21020) );
  INHSV2 U23636 ( .I(n21008), .ZN(n21014) );
  NAND2HSV2 U23637 ( .A1(n17813), .A2(n21010), .ZN(n21108) );
  NOR2HSV1 U23638 ( .A1(n17773), .A2(n21235), .ZN(n21692) );
  BUFHSV2 U23639 ( .I(n21011), .Z(n23445) );
  CLKAND2HSV2 U23640 ( .A1(n27121), .A2(n23445), .Z(n21015) );
  INHSV2 U23641 ( .I(n21013), .ZN(n27122) );
  AOI21HSV4 U23642 ( .A1(n21015), .A2(n27122), .B(n21014), .ZN(n21016) );
  OAI21HSV4 U23643 ( .A1(n21018), .A2(n21017), .B(n21016), .ZN(n21107) );
  NAND3HSV2 U23644 ( .A1(n21108), .A2(n21107), .A3(n21702), .ZN(n21019) );
  INHSV2 U23645 ( .I(n21813), .ZN(n21643) );
  INHSV2 U23646 ( .I(n21643), .ZN(n21714) );
  NAND2HSV2 U23647 ( .A1(n27571), .A2(\pe2/ti_7t [6]), .ZN(n21106) );
  CLKNHSV1 U23648 ( .I(n21106), .ZN(n21024) );
  AOI21HSV2 U23649 ( .A1(n21106), .A2(n21159), .B(n21880), .ZN(n21023) );
  OAI21HSV4 U23650 ( .A1(n29041), .A2(n21024), .B(n21023), .ZN(n21059) );
  NOR2HSV1 U23651 ( .A1(n21278), .A2(n17781), .ZN(n21051) );
  INHSV4 U23652 ( .I(\pe2/got [10]), .ZN(n27394) );
  NOR2HSV4 U23653 ( .A1(n21260), .A2(n27394), .ZN(n21026) );
  BUFHSV2 U23654 ( .I(\pe2/got [9]), .Z(n28636) );
  CLKNAND2HSV0 U23655 ( .A1(n21065), .A2(n28636), .ZN(n21025) );
  XNOR2HSV4 U23656 ( .A1(n21026), .A2(n21025), .ZN(n21049) );
  NAND2HSV0 U23657 ( .A1(\pe2/aot [15]), .A2(\pe2/bq[9] ), .ZN(n21028) );
  NAND2HSV0 U23658 ( .A1(\pe2/aot [14]), .A2(\pe2/bq[10] ), .ZN(n21027) );
  XOR2HSV0 U23659 ( .A1(n21028), .A2(n21027), .Z(n21032) );
  NAND2HSV0 U23660 ( .A1(\pe2/aot [13]), .A2(\pe2/bq[11] ), .ZN(n21030) );
  INAND2HSV0 U23661 ( .A1(n27322), .B1(\pe2/aot [8]), .ZN(n21029) );
  XOR2HSV0 U23662 ( .A1(n21030), .A2(n21029), .Z(n21031) );
  XOR2HSV0 U23663 ( .A1(n21032), .A2(n21031), .Z(n21039) );
  NAND2HSV0 U23664 ( .A1(\pe2/aot [12]), .A2(\pe2/bq[12] ), .ZN(n21034) );
  NAND2HSV0 U23665 ( .A1(\pe2/aot [11]), .A2(\pe2/bq[13] ), .ZN(n21033) );
  XOR2HSV0 U23666 ( .A1(n21034), .A2(n21033), .Z(n21037) );
  CLKNAND2HSV1 U23667 ( .A1(n21253), .A2(\pe2/pvq [9]), .ZN(n21035) );
  XOR2HSV0 U23668 ( .A1(n21035), .A2(\pe2/phq [9]), .Z(n21036) );
  XOR2HSV0 U23669 ( .A1(n21037), .A2(n21036), .Z(n21038) );
  XOR2HSV0 U23670 ( .A1(n21039), .A2(n21038), .Z(n21047) );
  NAND2HSV0 U23671 ( .A1(\pe2/aot [10]), .A2(\pe2/bq[14] ), .ZN(n21041) );
  NAND2HSV0 U23672 ( .A1(\pe2/bq[8] ), .A2(n11953), .ZN(n21040) );
  XOR2HSV0 U23673 ( .A1(n21041), .A2(n21040), .Z(n21045) );
  NAND2HSV0 U23674 ( .A1(\pe2/aot [9]), .A2(\pe2/bq[15] ), .ZN(n21043) );
  CLKBUFHSV4 U23675 ( .I(n21269), .Z(n27321) );
  CLKNAND2HSV1 U23676 ( .A1(\pe2/got [8]), .A2(n27321), .ZN(n21042) );
  XOR2HSV0 U23677 ( .A1(n21043), .A2(n21042), .Z(n21044) );
  XOR2HSV0 U23678 ( .A1(n21045), .A2(n21044), .Z(n21046) );
  XNOR2HSV1 U23679 ( .A1(n21047), .A2(n21046), .ZN(n21048) );
  CLKXOR2HSV2 U23680 ( .A1(n21049), .A2(n21048), .Z(n21050) );
  XNOR2HSV1 U23681 ( .A1(n21051), .A2(n21050), .ZN(n21053) );
  CLKNHSV0 U23682 ( .I(n21052), .ZN(n21055) );
  CLKNHSV0 U23683 ( .I(n21053), .ZN(n21054) );
  CLKNAND2HSV1 U23684 ( .A1(n21055), .A2(n21054), .ZN(n21056) );
  XNOR2HSV4 U23685 ( .A1(n21059), .A2(n21058), .ZN(n21061) );
  INHSV4 U23686 ( .I(n21061), .ZN(n21062) );
  INHSV4 U23687 ( .I(n21239), .ZN(n21232) );
  INHSV2 U23688 ( .I(n21232), .ZN(n21064) );
  INHSV2 U23689 ( .I(n21292), .ZN(n21148) );
  NAND2HSV2 U23690 ( .A1(n12624), .A2(n27544), .ZN(n21115) );
  NAND2HSV0 U23691 ( .A1(n21817), .A2(\pe2/got [8]), .ZN(n21101) );
  BUFHSV2 U23692 ( .I(n21278), .Z(n27452) );
  NOR2HSV1 U23693 ( .A1(n27452), .A2(n27572), .ZN(n21099) );
  BUFHSV2 U23694 ( .I(n21065), .Z(n28697) );
  NAND2HSV0 U23695 ( .A1(n28697), .A2(\pe2/got [5]), .ZN(n21097) );
  BUFHSV2 U23696 ( .I(n21066), .Z(n27423) );
  NOR2HSV2 U23697 ( .A1(n27423), .A2(n27498), .ZN(n21096) );
  NAND2HSV0 U23698 ( .A1(\pe2/aot [12]), .A2(\pe2/bq[8] ), .ZN(n21068) );
  NAND2HSV0 U23699 ( .A1(\pe2/aot [10]), .A2(\pe2/bq[10] ), .ZN(n21067) );
  XOR2HSV0 U23700 ( .A1(n21068), .A2(n21067), .Z(n21072) );
  NAND2HSV0 U23701 ( .A1(\pe2/bq[5] ), .A2(\pe2/aot [15]), .ZN(n21070) );
  NAND2HSV0 U23702 ( .A1(\pe2/bq[6] ), .A2(\pe2/aot [14]), .ZN(n21069) );
  XOR2HSV0 U23703 ( .A1(n21070), .A2(n21069), .Z(n21071) );
  XOR2HSV0 U23704 ( .A1(n21072), .A2(n21071), .Z(n21081) );
  NAND2HSV0 U23705 ( .A1(\pe2/aot [5]), .A2(\pe2/bq[15] ), .ZN(n21074) );
  NAND2HSV0 U23706 ( .A1(\pe2/aot [7]), .A2(\pe2/bq[13] ), .ZN(n21073) );
  XOR2HSV0 U23707 ( .A1(n21074), .A2(n21073), .Z(n21079) );
  NAND2HSV0 U23708 ( .A1(\pe2/aot [9]), .A2(\pe2/bq[11] ), .ZN(n21077) );
  CLKNHSV0 U23709 ( .I(\pe2/bq[14] ), .ZN(n21075) );
  NAND2HSV0 U23710 ( .A1(\pe2/aot [6]), .A2(n27312), .ZN(n21076) );
  XOR2HSV0 U23711 ( .A1(n21077), .A2(n21076), .Z(n21078) );
  XOR2HSV0 U23712 ( .A1(n21079), .A2(n21078), .Z(n21080) );
  XOR2HSV0 U23713 ( .A1(n21081), .A2(n21080), .Z(n21094) );
  NAND2HSV0 U23714 ( .A1(\pe2/aot [4]), .A2(n21842), .ZN(n21083) );
  NAND2HSV0 U23715 ( .A1(\pe2/aot [13]), .A2(\pe2/bq[7] ), .ZN(n21082) );
  XOR2HSV0 U23716 ( .A1(n21083), .A2(n21082), .Z(n21087) );
  NAND2HSV0 U23717 ( .A1(\pe2/aot [8]), .A2(\pe2/bq[12] ), .ZN(n21085) );
  NAND2HSV0 U23718 ( .A1(\pe2/got [4]), .A2(n27321), .ZN(n21084) );
  XOR2HSV0 U23719 ( .A1(n21085), .A2(n21084), .Z(n21086) );
  XNOR2HSV1 U23720 ( .A1(n21087), .A2(n21086), .ZN(n21092) );
  BUFHSV2 U23721 ( .I(n22114), .Z(n23539) );
  NAND2HSV0 U23722 ( .A1(n11953), .A2(\pe2/bq[4] ), .ZN(n21088) );
  NAND2HSV0 U23723 ( .A1(\pe2/aot [11]), .A2(\pe2/bq[9] ), .ZN(n27502) );
  CLKNHSV0 U23724 ( .I(\pe2/aot [11]), .ZN(n27462) );
  INHSV2 U23725 ( .I(\pe2/bq[4] ), .ZN(n27692) );
  NOR2HSV0 U23726 ( .A1(n27462), .A2(n27692), .ZN(n27417) );
  AOI22HSV0 U23727 ( .A1(n21088), .A2(n27502), .B1(n21130), .B2(n27417), .ZN(
        n21089) );
  XOR2HSV0 U23728 ( .A1(n21090), .A2(n21089), .Z(n21091) );
  XNOR2HSV1 U23729 ( .A1(n21092), .A2(n21091), .ZN(n21093) );
  XNOR2HSV1 U23730 ( .A1(n21094), .A2(n21093), .ZN(n21095) );
  XOR3HSV2 U23731 ( .A1(n21097), .A2(n21096), .A3(n21095), .Z(n21098) );
  XOR2HSV0 U23732 ( .A1(n21099), .A2(n21098), .Z(n21100) );
  XNOR2HSV1 U23733 ( .A1(n21101), .A2(n21100), .ZN(n21105) );
  CLKNHSV4 U23734 ( .I(n21102), .ZN(n27524) );
  INHSV2 U23735 ( .I(n21103), .ZN(n27647) );
  CLKNAND2HSV0 U23736 ( .A1(n27524), .A2(n27647), .ZN(n21104) );
  XNOR2HSV1 U23737 ( .A1(n21105), .A2(n21104), .ZN(n21113) );
  BUFHSV3 U23738 ( .I(n28942), .Z(n27271) );
  NOR2HSV2 U23739 ( .A1(n27527), .A2(n27394), .ZN(n21112) );
  CLKNAND2HSV3 U23740 ( .A1(n21110), .A2(n21109), .ZN(n21145) );
  INHSV3 U23741 ( .I(n21145), .ZN(n21324) );
  INHSV4 U23742 ( .I(n21324), .ZN(n27432) );
  NAND2HSV0 U23743 ( .A1(n27432), .A2(n27543), .ZN(n21111) );
  XOR3HSV2 U23744 ( .A1(n21113), .A2(n21112), .A3(n21111), .Z(n21114) );
  XNOR2HSV4 U23745 ( .A1(n21115), .A2(n21114), .ZN(n21306) );
  CLKNAND2HSV2 U23746 ( .A1(n21239), .A2(n23445), .ZN(n21242) );
  NOR2HSV2 U23747 ( .A1(n21713), .A2(\pe2/ti_7t [9]), .ZN(n21236) );
  NOR2HSV4 U23748 ( .A1(n21153), .A2(n21152), .ZN(n21222) );
  INHSV2 U23749 ( .I(n21241), .ZN(n21147) );
  NAND2HSV0 U23750 ( .A1(n27543), .A2(n21817), .ZN(n21143) );
  NOR2HSV1 U23751 ( .A1(n21118), .A2(n27394), .ZN(n21141) );
  NAND2HSV0 U23752 ( .A1(n28697), .A2(\pe2/got [8]), .ZN(n21139) );
  NAND2HSV0 U23753 ( .A1(\pe2/aot [13]), .A2(\pe2/bq[10] ), .ZN(n21120) );
  NAND2HSV0 U23754 ( .A1(\pe2/aot [11]), .A2(\pe2/bq[12] ), .ZN(n21119) );
  XOR2HSV0 U23755 ( .A1(n21120), .A2(n21119), .Z(n21122) );
  XOR2HSV0 U23756 ( .A1(n21122), .A2(n21121), .Z(n21127) );
  CLKNHSV2 U23757 ( .I(\pe2/aot [7]), .ZN(n27580) );
  BUFHSV4 U23758 ( .I(n22114), .Z(n23537) );
  NAND2HSV2 U23759 ( .A1(n22114), .A2(\pe2/pvq [10]), .ZN(n21123) );
  XOR2HSV0 U23760 ( .A1(n21123), .A2(\pe2/phq [10]), .Z(n21124) );
  CLKNHSV0 U23761 ( .I(\pe2/aot [14]), .ZN(n21128) );
  INHSV2 U23762 ( .I(\pe2/bq[7] ), .ZN(n27461) );
  NOR2HSV2 U23763 ( .A1(n21128), .A2(n27461), .ZN(n21268) );
  AOI22HSV0 U23764 ( .A1(n17785), .A2(\pe2/bq[7] ), .B1(\pe2/aot [14]), .B2(
        \pe2/bq[9] ), .ZN(n21129) );
  AOI21HSV2 U23765 ( .A1(n21130), .A2(n21268), .B(n21129), .ZN(n21134) );
  NAND2HSV0 U23766 ( .A1(\pe2/aot [12]), .A2(\pe2/bq[11] ), .ZN(n21132) );
  NAND2HSV0 U23767 ( .A1(n27312), .A2(\pe2/aot [9]), .ZN(n21131) );
  XOR2HSV0 U23768 ( .A1(n21132), .A2(n21131), .Z(n21133) );
  XOR3HSV2 U23769 ( .A1(n27299), .A2(n21134), .A3(n21133), .Z(n21135) );
  XNOR2HSV4 U23770 ( .A1(n21136), .A2(n21135), .ZN(n21138) );
  INHSV2 U23771 ( .I(\pe2/got [9]), .ZN(n27610) );
  NOR2HSV2 U23772 ( .A1(n21260), .A2(n27610), .ZN(n21137) );
  XOR3HSV2 U23773 ( .A1(n21139), .A2(n21138), .A3(n21137), .Z(n21140) );
  XNOR2HSV1 U23774 ( .A1(n21141), .A2(n21140), .ZN(n21142) );
  OAI21HSV2 U23775 ( .A1(n22086), .A2(n28421), .B(n21713), .ZN(n21146) );
  AOI21HSV4 U23776 ( .A1(n21154), .A2(n21147), .B(n21146), .ZN(n21221) );
  CLKNAND2HSV2 U23777 ( .A1(n21151), .A2(n21150), .ZN(n21223) );
  NAND2HSV2 U23778 ( .A1(n21701), .A2(\pe2/ti_7t [10]), .ZN(n21867) );
  BUFHSV2 U23779 ( .I(n21867), .Z(n21163) );
  NOR2HSV2 U23780 ( .A1(n12270), .A2(n21152), .ZN(n21218) );
  INHSV2 U23781 ( .I(n21241), .ZN(n21231) );
  NAND2HSV2 U23782 ( .A1(n21150), .A2(n21231), .ZN(n21165) );
  NAND3HSV2 U23783 ( .A1(n21154), .A2(n17774), .A3(n21241), .ZN(n21162) );
  INHSV2 U23784 ( .I(n21156), .ZN(n21158) );
  AOI21HSV2 U23785 ( .A1(n21160), .A2(n21225), .B(n21159), .ZN(n21161) );
  CLKNAND2HSV1 U23786 ( .A1(n27344), .A2(n21144), .ZN(n21308) );
  CLKNAND2HSV3 U23787 ( .A1(n21166), .A2(n21165), .ZN(n21217) );
  INHSV2 U23788 ( .I(n21221), .ZN(n21169) );
  OAI22HSV4 U23789 ( .A1(n21170), .A2(n21169), .B1(n21168), .B2(n21867), .ZN(
        n21171) );
  NAND2HSV0 U23790 ( .A1(n21241), .A2(\pe2/got [16]), .ZN(n21173) );
  INHSV2 U23791 ( .I(n21173), .ZN(n21179) );
  CLKAND2HSV2 U23792 ( .A1(n21232), .A2(n23445), .Z(n21178) );
  NOR2HSV1 U23793 ( .A1(n21236), .A2(n21225), .ZN(n21175) );
  CLKAND2HSV1 U23794 ( .A1(n21175), .A2(n28693), .Z(n21174) );
  CLKNAND2HSV1 U23795 ( .A1(n22084), .A2(n21174), .ZN(n21177) );
  CLKNAND2HSV1 U23796 ( .A1(n21242), .A2(n21175), .ZN(n21176) );
  NAND2HSV2 U23797 ( .A1(n21145), .A2(n28429), .ZN(n21214) );
  NAND2HSV0 U23798 ( .A1(\pe2/got [10]), .A2(n21817), .ZN(n21209) );
  NAND2HSV0 U23799 ( .A1(n28697), .A2(\pe2/got [7]), .ZN(n21205) );
  NAND2HSV0 U23800 ( .A1(\pe2/aot [10]), .A2(\pe2/bq[12] ), .ZN(n21181) );
  NAND2HSV0 U23801 ( .A1(\pe2/aot [9]), .A2(\pe2/bq[13] ), .ZN(n21180) );
  XOR2HSV0 U23802 ( .A1(n21181), .A2(n21180), .Z(n21183) );
  XOR2HSV0 U23803 ( .A1(n21183), .A2(n21182), .Z(n21191) );
  NAND2HSV0 U23804 ( .A1(\pe2/aot [15]), .A2(\pe2/bq[7] ), .ZN(n21185) );
  NAND2HSV0 U23805 ( .A1(\pe2/aot [14]), .A2(\pe2/bq[8] ), .ZN(n21184) );
  XOR2HSV0 U23806 ( .A1(n21185), .A2(n21184), .Z(n21189) );
  NAND2HSV0 U23807 ( .A1(\pe2/aot [11]), .A2(\pe2/bq[11] ), .ZN(n21187) );
  NAND2HSV0 U23808 ( .A1(n17785), .A2(\pe2/bq[6] ), .ZN(n21186) );
  XOR2HSV0 U23809 ( .A1(n21187), .A2(n21186), .Z(n21188) );
  XOR2HSV0 U23810 ( .A1(n21189), .A2(n21188), .Z(n21190) );
  XOR2HSV0 U23811 ( .A1(n21191), .A2(n21190), .Z(n21202) );
  NAND2HSV0 U23812 ( .A1(\pe2/aot [8]), .A2(n27312), .ZN(n21193) );
  NAND2HSV0 U23813 ( .A1(\pe2/aot [12]), .A2(\pe2/bq[10] ), .ZN(n21192) );
  XOR2HSV0 U23814 ( .A1(n21193), .A2(n21192), .Z(n21196) );
  CLKNAND2HSV1 U23815 ( .A1(n21253), .A2(\pe2/pvq [11]), .ZN(n21194) );
  XNOR2HSV1 U23816 ( .A1(n21194), .A2(\pe2/phq [11]), .ZN(n21195) );
  XNOR2HSV1 U23817 ( .A1(n21196), .A2(n21195), .ZN(n21200) );
  NAND2HSV0 U23818 ( .A1(\pe2/aot [13]), .A2(\pe2/bq[9] ), .ZN(n21198) );
  CLKNAND2HSV0 U23819 ( .A1(\pe2/got [6]), .A2(n27321), .ZN(n21197) );
  XOR2HSV0 U23820 ( .A1(n21198), .A2(n21197), .Z(n21199) );
  XNOR2HSV1 U23821 ( .A1(n21200), .A2(n21199), .ZN(n21201) );
  XNOR2HSV1 U23822 ( .A1(n21202), .A2(n21201), .ZN(n21204) );
  INHSV2 U23823 ( .I(\pe2/got [8]), .ZN(n27645) );
  NOR2HSV0 U23824 ( .A1(n27423), .A2(n27645), .ZN(n21203) );
  XOR3HSV2 U23825 ( .A1(n21205), .A2(n21204), .A3(n21203), .Z(n21207) );
  NOR2HSV0 U23826 ( .A1(n21278), .A2(n27610), .ZN(n21206) );
  XOR2HSV0 U23827 ( .A1(n21207), .A2(n21206), .Z(n21208) );
  XNOR2HSV1 U23828 ( .A1(n21209), .A2(n21208), .ZN(n21211) );
  NAND2HSV0 U23829 ( .A1(n27543), .A2(n27524), .ZN(n21210) );
  XNOR2HSV1 U23830 ( .A1(n21211), .A2(n21210), .ZN(n21212) );
  XNOR2HSV4 U23831 ( .A1(n21213), .A2(n21214), .ZN(n21215) );
  XNOR2HSV4 U23832 ( .A1(n21640), .A2(n21639), .ZN(n28950) );
  NAND2HSV4 U23833 ( .A1(n21879), .A2(n22085), .ZN(n21310) );
  XNOR2HSV4 U23834 ( .A1(n25361), .A2(n21310), .ZN(n21636) );
  INHSV2 U23835 ( .I(n21696), .ZN(n21301) );
  INHSV2 U23836 ( .I(n21217), .ZN(n21220) );
  CLKNAND2HSV1 U23837 ( .A1(n21220), .A2(n21219), .ZN(n21230) );
  NOR2HSV1 U23838 ( .A1(n21867), .A2(n21225), .ZN(n21226) );
  AOI21HSV4 U23839 ( .A1(n21228), .A2(n21227), .B(n21226), .ZN(n21229) );
  INHSV2 U23840 ( .I(n21231), .ZN(n21816) );
  CLKAND2HSV1 U23841 ( .A1(n21232), .A2(n21696), .Z(n21233) );
  NAND2HSV2 U23842 ( .A1(n21816), .A2(n21233), .ZN(n21245) );
  NOR2HSV0 U23843 ( .A1(n21235), .A2(n21234), .ZN(n21703) );
  CLKNHSV0 U23844 ( .I(n21236), .ZN(n21237) );
  NAND2HSV0 U23845 ( .A1(n21237), .A2(n17767), .ZN(n21238) );
  OAI21HSV0 U23846 ( .A1(n21242), .A2(n21241), .B(n21240), .ZN(n21243) );
  CLKNHSV0 U23847 ( .I(n21243), .ZN(n21244) );
  NAND2HSV0 U23848 ( .A1(\pe2/aot [13]), .A2(\pe2/bq[8] ), .ZN(n21248) );
  NAND2HSV0 U23849 ( .A1(\pe2/aot [8]), .A2(\pe2/bq[13] ), .ZN(n21247) );
  XOR2HSV0 U23850 ( .A1(n21248), .A2(n21247), .Z(n21252) );
  NAND2HSV0 U23851 ( .A1(\pe2/aot [7]), .A2(n27312), .ZN(n21250) );
  NAND2HSV0 U23852 ( .A1(\pe2/aot [15]), .A2(\pe2/bq[6] ), .ZN(n21249) );
  XOR2HSV0 U23853 ( .A1(n21250), .A2(n21249), .Z(n21251) );
  XOR2HSV0 U23854 ( .A1(n21252), .A2(n21251), .Z(n21257) );
  CLKNHSV0 U23855 ( .I(\pe2/bq[5] ), .ZN(n23538) );
  NOR2HSV0 U23856 ( .A1(n21254), .A2(n23538), .ZN(n27298) );
  XNOR2HSV1 U23857 ( .A1(n21255), .A2(n27298), .ZN(n21256) );
  XNOR2HSV1 U23858 ( .A1(n21257), .A2(n21256), .ZN(n21259) );
  NAND2HSV0 U23859 ( .A1(n28697), .A2(n14006), .ZN(n21258) );
  XOR2HSV0 U23860 ( .A1(n21259), .A2(n21258), .Z(n21281) );
  NOR2HSV1 U23861 ( .A1(n21260), .A2(n27572), .ZN(n21277) );
  NAND2HSV0 U23862 ( .A1(\pe2/aot [12]), .A2(\pe2/bq[9] ), .ZN(n21262) );
  NAND2HSV0 U23863 ( .A1(\pe2/aot [10]), .A2(\pe2/bq[11] ), .ZN(n21261) );
  XOR2HSV0 U23864 ( .A1(n21262), .A2(n21261), .Z(n21266) );
  NAND2HSV0 U23865 ( .A1(\pe2/aot [6]), .A2(\pe2/bq[15] ), .ZN(n21264) );
  NAND2HSV0 U23866 ( .A1(\pe2/aot [5]), .A2(n21842), .ZN(n21263) );
  XOR2HSV0 U23867 ( .A1(n21264), .A2(n21263), .Z(n21265) );
  XOR2HSV0 U23868 ( .A1(n21266), .A2(n21265), .Z(n21275) );
  NAND2HSV0 U23869 ( .A1(\pe2/aot [11]), .A2(\pe2/bq[10] ), .ZN(n21267) );
  XOR2HSV0 U23870 ( .A1(n21268), .A2(n21267), .Z(n21273) );
  NAND2HSV0 U23871 ( .A1(\pe2/got [5]), .A2(n21269), .ZN(n21271) );
  NAND2HSV0 U23872 ( .A1(\pe2/aot [9]), .A2(\pe2/bq[12] ), .ZN(n21270) );
  XOR2HSV0 U23873 ( .A1(n21271), .A2(n21270), .Z(n21272) );
  XOR2HSV0 U23874 ( .A1(n21273), .A2(n21272), .Z(n21274) );
  XOR2HSV0 U23875 ( .A1(n21275), .A2(n21274), .Z(n21276) );
  XOR2HSV0 U23876 ( .A1(n21277), .A2(n21276), .Z(n21280) );
  NOR2HSV0 U23877 ( .A1(n21278), .A2(n27645), .ZN(n21279) );
  XOR3HSV2 U23878 ( .A1(n21281), .A2(n21280), .A3(n21279), .Z(n21282) );
  XNOR2HSV1 U23879 ( .A1(n21283), .A2(n21282), .ZN(n21285) );
  NAND2HSV0 U23880 ( .A1(n27524), .A2(\pe2/got [10]), .ZN(n21284) );
  XNOR2HSV1 U23881 ( .A1(n21285), .A2(n21284), .ZN(n21286) );
  NAND2HSV2 U23882 ( .A1(n27432), .A2(n27544), .ZN(n21287) );
  AOI21HSV0 U23883 ( .A1(n21290), .A2(n21289), .B(n21305), .ZN(n21291) );
  OAI21HSV2 U23884 ( .A1(n14033), .A2(n21292), .B(n21291), .ZN(n21293) );
  INHSV2 U23885 ( .I(n21708), .ZN(n21296) );
  NAND2HSV2 U23886 ( .A1(n21297), .A2(n21296), .ZN(n21300) );
  CLKNAND2HSV2 U23887 ( .A1(n21298), .A2(n21708), .ZN(n21299) );
  INHSV2 U23888 ( .I(n21632), .ZN(n25366) );
  NOR2HSV2 U23889 ( .A1(n25357), .A2(n28950), .ZN(n23446) );
  CLKNHSV1 U23890 ( .I(n21301), .ZN(n21302) );
  NAND2HSV2 U23891 ( .A1(n23446), .A2(n21302), .ZN(n25364) );
  CLKNAND2HSV0 U23892 ( .A1(n25364), .A2(n21714), .ZN(n21303) );
  NOR2HSV2 U23893 ( .A1(n25366), .A2(n21303), .ZN(n21304) );
  XNOR2HSV1 U23894 ( .A1(n21309), .A2(n21308), .ZN(n21311) );
  AOI21HSV4 U23895 ( .A1(n21629), .A2(n21628), .B(n21630), .ZN(n27295) );
  CLKNAND2HSV2 U23896 ( .A1(n27294), .A2(n27295), .ZN(n28590) );
  NAND2HSV2 U23897 ( .A1(n21313), .A2(\pe3/ti_7t [12]), .ZN(n23384) );
  NAND2HSV4 U23898 ( .A1(n21314), .A2(n23384), .ZN(n26349) );
  INHSV2 U23899 ( .I(n26349), .ZN(n26730) );
  INHSV1 U23900 ( .I(n26730), .ZN(n28939) );
  INHSV2 U23901 ( .I(n23871), .ZN(n28665) );
  BUFHSV2 U23902 ( .I(n21315), .Z(n21319) );
  BUFHSV2 U23903 ( .I(n21316), .Z(n21318) );
  NAND2HSV4 U23904 ( .A1(n21318), .A2(n21317), .ZN(n28457) );
  INHSV2 U23905 ( .I(n21322), .ZN(n22139) );
  INHSV2 U23906 ( .I(n22139), .ZN(n28631) );
  INHSV1 U23907 ( .I(n21323), .ZN(n28589) );
  CLKNHSV0 U23908 ( .I(n21324), .ZN(n28617) );
  CLKNHSV1 U23909 ( .I(n21325), .ZN(n28478) );
  BUFHSV2 U23910 ( .I(\pe4/got [3]), .Z(n28626) );
  CLKNHSV1 U23911 ( .I(n21327), .ZN(n28635) );
  XOR2HSV0 U23912 ( .A1(n21329), .A2(n21328), .Z(n21331) );
  XNOR2HSV0 U23913 ( .A1(n21331), .A2(n21330), .ZN(n29010) );
  MUX2HSV1 U23914 ( .I0(bo4[16]), .I1(n22834), .S(n27076), .Z(n28854) );
  INHSV2 U23915 ( .I(n20164), .ZN(n28639) );
  MUX2HSV1 U23916 ( .I0(bo11[14]), .I1(\pe11/bq[14] ), .S(n23499), .Z(n28717)
         );
  INHSV1 U23917 ( .I(n21332), .ZN(n27076) );
  MUX2HSV1 U23918 ( .I0(bo4[12]), .I1(\pe4/bq[12] ), .S(n27076), .Z(n28760) );
  MUX2HSV1 U23919 ( .I0(bo6[12]), .I1(n25701), .S(n28867), .Z(n28871) );
  MUX2HSV2 U23920 ( .I0(bo9[6]), .I1(\pe9/bq[6] ), .S(n27093), .Z(n28898) );
  INHSV1 U23921 ( .I(n28682), .ZN(n21758) );
  MUX2HSV1 U23922 ( .I0(\pe5/bq[13] ), .I1(bo5[13]), .S(n21758), .Z(n28710) );
  MUX2HSV1 U23923 ( .I0(bo3[16]), .I1(n23336), .S(n23520), .Z(n28838) );
  MUX2HSV1 U23924 ( .I0(bo9[16]), .I1(n28044), .S(n27078), .Z(n28753) );
  MUX2HSV1 U23925 ( .I0(bo9[2]), .I1(\pe9/bq[2] ), .S(n21760), .Z(n28779) );
  XOR2HSV4 U23926 ( .A1(n21337), .A2(n21336), .Z(n21341) );
  INHSV2 U23927 ( .I(n21341), .ZN(n21340) );
  MUX2NHSV2 U23928 ( .I0(n21341), .I1(n21340), .S(n21718), .ZN(n21343) );
  CLKNHSV0 U23929 ( .I(\pe5/ti_7t [14]), .ZN(n21344) );
  AOI21HSV0 U23930 ( .A1(n21345), .A2(n21344), .B(n27190), .ZN(n21715) );
  AND2HSV2 U23931 ( .A1(n21346), .A2(n21715), .Z(n21461) );
  CLKNAND2HSV1 U23932 ( .A1(n21348), .A2(n14820), .ZN(n21417) );
  NAND2HSV2 U23933 ( .A1(n28803), .A2(\pe5/got [13]), .ZN(n21410) );
  NAND2HSV2 U23934 ( .A1(n21003), .A2(\pe5/ti_7t [10]), .ZN(n21424) );
  CLKNHSV0 U23935 ( .I(n21424), .ZN(n21351) );
  AOI21HSV2 U23936 ( .A1(n21424), .A2(n21003), .B(n21349), .ZN(n21350) );
  OAI21HSV2 U23937 ( .A1(pov5[10]), .A2(n21351), .B(n21350), .ZN(n21408) );
  CLKNAND2HSV0 U23938 ( .A1(n11931), .A2(n14071), .ZN(n21402) );
  INHSV2 U23939 ( .I(n21352), .ZN(n25350) );
  CLKNHSV0 U23940 ( .I(\pe5/got [7]), .ZN(n24420) );
  NOR2HSV1 U23941 ( .A1(n25350), .A2(n24420), .ZN(n21398) );
  NAND2HSV0 U23942 ( .A1(n13999), .A2(n28594), .ZN(n21373) );
  NAND2HSV0 U23943 ( .A1(\pe5/aot [12]), .A2(\pe5/bq[6] ), .ZN(n21354) );
  NAND2HSV0 U23944 ( .A1(\pe5/aot [7]), .A2(\pe5/bq[11] ), .ZN(n21353) );
  XOR2HSV0 U23945 ( .A1(n21354), .A2(n21353), .Z(n21371) );
  NAND2HSV0 U23946 ( .A1(n28682), .A2(\pe5/pvq [15]), .ZN(n21355) );
  XNOR2HSV1 U23947 ( .A1(n21355), .A2(\pe5/phq [15]), .ZN(n21362) );
  CLKNHSV0 U23948 ( .I(n21356), .ZN(n21360) );
  CLKNHSV0 U23949 ( .I(\pe5/aot [5]), .ZN(n24440) );
  NOR2HSV0 U23950 ( .A1(n24440), .A2(n21357), .ZN(n21359) );
  NAND2HSV0 U23951 ( .A1(\pe5/aot [5]), .A2(\pe5/bq[7] ), .ZN(n21436) );
  OAI22HSV0 U23952 ( .A1(n21360), .A2(n21359), .B1(n21358), .B2(n21436), .ZN(
        n21361) );
  XNOR2HSV1 U23953 ( .A1(n21362), .A2(n21361), .ZN(n21370) );
  NAND2HSV0 U23954 ( .A1(\pe5/aot [4]), .A2(\pe5/bq[14] ), .ZN(n21364) );
  NAND2HSV0 U23955 ( .A1(\pe5/aot [8]), .A2(\pe5/bq[10] ), .ZN(n21363) );
  XOR2HSV0 U23956 ( .A1(n21364), .A2(n21363), .Z(n21368) );
  NAND2HSV0 U23957 ( .A1(\pe5/bq[4] ), .A2(\pe5/aot [14]), .ZN(n21366) );
  NAND2HSV0 U23958 ( .A1(\pe5/aot [13]), .A2(\pe5/bq[5] ), .ZN(n21365) );
  XOR2HSV0 U23959 ( .A1(n21366), .A2(n21365), .Z(n21367) );
  XOR2HSV0 U23960 ( .A1(n21368), .A2(n21367), .Z(n21369) );
  XOR3HSV2 U23961 ( .A1(n21371), .A2(n21370), .A3(n21369), .Z(n21372) );
  XNOR2HSV1 U23962 ( .A1(n21373), .A2(n21372), .ZN(n21392) );
  NAND2HSV0 U23963 ( .A1(n21374), .A2(\pe5/aot [3]), .ZN(n21376) );
  NAND2HSV0 U23964 ( .A1(\pe5/aot [10]), .A2(\pe5/bq[8] ), .ZN(n21375) );
  XOR2HSV0 U23965 ( .A1(n21376), .A2(n21375), .Z(n21380) );
  NAND2HSV0 U23966 ( .A1(n14031), .A2(\pe5/bq[3] ), .ZN(n21378) );
  NAND2HSV0 U23967 ( .A1(\pe5/aot [9]), .A2(\pe5/bq[9] ), .ZN(n21377) );
  XOR2HSV0 U23968 ( .A1(n21378), .A2(n21377), .Z(n21379) );
  XOR2HSV0 U23969 ( .A1(n21380), .A2(n21379), .Z(n21388) );
  NAND2HSV0 U23970 ( .A1(n25626), .A2(\pe5/got [2]), .ZN(n21382) );
  CLKNHSV0 U23971 ( .I(\pe5/aot [2]), .ZN(n21573) );
  NAND2HSV0 U23972 ( .A1(\pe5/aot [2]), .A2(n25349), .ZN(n21381) );
  XOR2HSV0 U23973 ( .A1(n21382), .A2(n21381), .Z(n21386) );
  INHSV2 U23974 ( .I(\pe5/bq[2] ), .ZN(n24439) );
  INHSV2 U23975 ( .I(n24439), .ZN(n27053) );
  NAND2HSV0 U23976 ( .A1(n21488), .A2(n27053), .ZN(n21384) );
  NAND2HSV0 U23977 ( .A1(\pe5/aot [6]), .A2(n23909), .ZN(n21383) );
  XOR2HSV0 U23978 ( .A1(n21384), .A2(n21383), .Z(n21385) );
  XOR2HSV0 U23979 ( .A1(n21386), .A2(n21385), .Z(n21387) );
  XOR2HSV0 U23980 ( .A1(n21388), .A2(n21387), .Z(n21390) );
  XNOR2HSV1 U23981 ( .A1(n21390), .A2(n21389), .ZN(n21391) );
  XNOR2HSV1 U23982 ( .A1(n21392), .A2(n21391), .ZN(n21394) );
  NAND2HSV0 U23983 ( .A1(n28614), .A2(n14072), .ZN(n21393) );
  XNOR2HSV1 U23984 ( .A1(n21394), .A2(n21393), .ZN(n21396) );
  NAND2HSV0 U23985 ( .A1(n24674), .A2(n28647), .ZN(n21395) );
  XNOR2HSV1 U23986 ( .A1(n21396), .A2(n21395), .ZN(n21397) );
  XNOR2HSV1 U23987 ( .A1(n21398), .A2(n21397), .ZN(n21400) );
  NAND2HSV0 U23988 ( .A1(n21504), .A2(n24340), .ZN(n21399) );
  XOR2HSV0 U23989 ( .A1(n21400), .A2(n21399), .Z(n21401) );
  XNOR2HSV1 U23990 ( .A1(n21402), .A2(n21401), .ZN(n21406) );
  CLKNHSV1 U23991 ( .I(n28800), .ZN(n21613) );
  NOR2HSV2 U23992 ( .A1(n21613), .A2(n21510), .ZN(n21405) );
  NOR2HSV0 U23993 ( .A1(n21614), .A2(n14535), .ZN(n21403) );
  INHSV2 U23994 ( .I(n21403), .ZN(n21404) );
  XOR3HSV2 U23995 ( .A1(n21406), .A2(n21405), .A3(n21404), .Z(n21407) );
  XNOR2HSV1 U23996 ( .A1(n21408), .A2(n21407), .ZN(n21409) );
  XNOR2HSV4 U23997 ( .A1(n21410), .A2(n21409), .ZN(n21416) );
  AOI21HSV2 U23998 ( .A1(n21413), .A2(n21412), .B(n21411), .ZN(n21414) );
  XNOR2HSV4 U23999 ( .A1(n21416), .A2(n21415), .ZN(n21420) );
  INHSV2 U24000 ( .I(n23275), .ZN(n23277) );
  NAND2HSV4 U24001 ( .A1(n21464), .A2(n21463), .ZN(n27106) );
  INHSV2 U24002 ( .I(n21423), .ZN(n21521) );
  NAND2HSV0 U24003 ( .A1(n24341), .A2(n24340), .ZN(n21456) );
  NAND2HSV0 U24004 ( .A1(\pe5/ti_7[10] ), .A2(n28647), .ZN(n21451) );
  NAND2HSV0 U24005 ( .A1(n21523), .A2(\pe5/got [3]), .ZN(n21446) );
  NAND2HSV0 U24006 ( .A1(\pe5/aot [9]), .A2(\pe5/bq[3] ), .ZN(n21426) );
  NAND2HSV0 U24007 ( .A1(\pe5/aot [4]), .A2(\pe5/bq[8] ), .ZN(n21425) );
  XOR2HSV0 U24008 ( .A1(n21426), .A2(n21425), .Z(n21430) );
  NAND2HSV0 U24009 ( .A1(\pe5/aot [3]), .A2(\pe5/bq[9] ), .ZN(n21428) );
  NAND2HSV0 U24010 ( .A1(\pe5/aot [10]), .A2(\pe5/bq[2] ), .ZN(n21427) );
  XOR2HSV0 U24011 ( .A1(n21428), .A2(n21427), .Z(n21429) );
  XOR2HSV0 U24012 ( .A1(n21430), .A2(n21429), .Z(n21435) );
  NAND2HSV0 U24013 ( .A1(\pe5/aot [2]), .A2(\pe5/bq[10] ), .ZN(n21432) );
  NAND2HSV0 U24014 ( .A1(\pe5/aot [1]), .A2(\pe5/bq[11] ), .ZN(n21431) );
  XOR2HSV0 U24015 ( .A1(n21432), .A2(n21431), .Z(n21433) );
  NAND2HSV0 U24016 ( .A1(\pe5/bq[1] ), .A2(\pe5/aot [11]), .ZN(n23916) );
  XNOR2HSV1 U24017 ( .A1(n21433), .A2(n23916), .ZN(n21434) );
  XNOR2HSV1 U24018 ( .A1(n21435), .A2(n21434), .ZN(n21441) );
  NAND2HSV0 U24019 ( .A1(\pe5/aot [6]), .A2(\pe5/bq[6] ), .ZN(n21560) );
  XOR2HSV0 U24020 ( .A1(n21436), .A2(n21560), .Z(n21439) );
  CLKNHSV0 U24021 ( .I(\pe5/aot [8]), .ZN(n21437) );
  NOR2HSV0 U24022 ( .A1(n21437), .A2(n21532), .ZN(n21469) );
  NAND2HSV0 U24023 ( .A1(\pe5/bq[5] ), .A2(\pe5/aot [7]), .ZN(n21558) );
  XOR2HSV0 U24024 ( .A1(n21469), .A2(n21558), .Z(n21438) );
  XOR2HSV0 U24025 ( .A1(n21439), .A2(n21438), .Z(n21440) );
  XNOR2HSV1 U24026 ( .A1(n21441), .A2(n21440), .ZN(n21444) );
  CLKNHSV0 U24027 ( .I(\pe5/got [1]), .ZN(n24638) );
  NOR2HSV0 U24028 ( .A1(n25350), .A2(n24638), .ZN(n21443) );
  NAND2HSV0 U24029 ( .A1(n21504), .A2(\pe5/got [2]), .ZN(n21442) );
  XOR3HSV1 U24030 ( .A1(n21444), .A2(n21443), .A3(n21442), .Z(n21445) );
  XNOR2HSV1 U24031 ( .A1(n21446), .A2(n21445), .ZN(n21449) );
  NOR2HSV0 U24032 ( .A1(n21613), .A2(n24414), .ZN(n21448) );
  CLKNHSV0 U24033 ( .I(\pe5/got [5]), .ZN(n24677) );
  OR2HSV1 U24034 ( .A1(n21614), .A2(n24677), .Z(n21447) );
  XOR3HSV1 U24035 ( .A1(n21449), .A2(n21448), .A3(n21447), .Z(n21450) );
  XNOR2HSV1 U24036 ( .A1(n21451), .A2(n21450), .ZN(n21454) );
  CLKNAND2HSV0 U24037 ( .A1(n21452), .A2(n28645), .ZN(n21453) );
  XNOR2HSV1 U24038 ( .A1(n21454), .A2(n21453), .ZN(n21455) );
  XOR2HSV0 U24039 ( .A1(n21456), .A2(n21455), .Z(n21457) );
  XOR2HSV0 U24040 ( .A1(n21458), .A2(n21457), .Z(n21459) );
  CLKNAND2HSV1 U24041 ( .A1(n27112), .A2(n14045), .ZN(n21520) );
  NAND2HSV0 U24042 ( .A1(n24341), .A2(\pe5/got [13]), .ZN(n21518) );
  NAND2HSV0 U24043 ( .A1(\pe5/ti_7[10] ), .A2(\pe5/got [11]), .ZN(n21515) );
  NAND2HSV0 U24044 ( .A1(n21465), .A2(n24340), .ZN(n21509) );
  NAND2HSV0 U24045 ( .A1(n28594), .A2(\pe5/got [3]), .ZN(n21485) );
  NAND2HSV0 U24046 ( .A1(\pe5/aot [1]), .A2(\pe5/bq[16] ), .ZN(n21467) );
  NAND2HSV0 U24047 ( .A1(\pe5/aot [6]), .A2(\pe5/bq[11] ), .ZN(n21466) );
  XOR2HSV0 U24048 ( .A1(n21467), .A2(n21466), .Z(n21483) );
  AOI22HSV0 U24049 ( .A1(\pe5/aot [13]), .A2(\pe5/bq[4] ), .B1(\pe5/bq[9] ), 
        .B2(\pe5/aot [8]), .ZN(n21468) );
  AOI21HSV0 U24050 ( .A1(n24388), .A2(n21469), .B(n21468), .ZN(n21474) );
  NAND2HSV0 U24051 ( .A1(\pe5/bq[2] ), .A2(\pe5/aot [12]), .ZN(n23919) );
  NOR2HSV0 U24052 ( .A1(n21470), .A2(n23919), .ZN(n21472) );
  AOI22HSV0 U24053 ( .A1(n14031), .A2(n27053), .B1(\pe5/aot [12]), .B2(
        \pe5/bq[5] ), .ZN(n21471) );
  NOR2HSV1 U24054 ( .A1(n21472), .A2(n21471), .ZN(n21473) );
  XOR2HSV0 U24055 ( .A1(n21474), .A2(n21473), .Z(n21482) );
  NAND2HSV0 U24056 ( .A1(n24647), .A2(\pe5/aot [2]), .ZN(n21476) );
  NAND2HSV0 U24057 ( .A1(\pe5/aot [7]), .A2(\pe5/bq[10] ), .ZN(n21475) );
  XOR2HSV0 U24058 ( .A1(n21476), .A2(n21475), .Z(n21480) );
  NAND2HSV0 U24059 ( .A1(\pe5/aot [5]), .A2(n23909), .ZN(n21478) );
  XOR2HSV0 U24060 ( .A1(n21478), .A2(n21477), .Z(n21479) );
  XOR2HSV0 U24061 ( .A1(n21480), .A2(n21479), .Z(n21481) );
  XOR3HSV2 U24062 ( .A1(n21483), .A2(n21482), .A3(n21481), .Z(n21484) );
  XNOR2HSV1 U24063 ( .A1(n21485), .A2(n21484), .ZN(n21499) );
  NAND2HSV0 U24064 ( .A1(n28682), .A2(\pe5/pq ), .ZN(n21487) );
  NAND2HSV0 U24065 ( .A1(\pe5/aot [4]), .A2(\pe5/bq[13] ), .ZN(n21486) );
  XOR2HSV0 U24066 ( .A1(n21487), .A2(n21486), .Z(n21492) );
  NAND2HSV0 U24067 ( .A1(\pe5/aot [3]), .A2(\pe5/bq[14] ), .ZN(n21490) );
  NAND2HSV0 U24068 ( .A1(n21488), .A2(\pe5/bq[1] ), .ZN(n21489) );
  XOR2HSV0 U24069 ( .A1(n21490), .A2(n21489), .Z(n21491) );
  XOR2HSV0 U24070 ( .A1(n21492), .A2(n21491), .Z(n21495) );
  XOR2HSV0 U24071 ( .A1(n21495), .A2(n21494), .Z(n21497) );
  NOR2HSV0 U24072 ( .A1(n27191), .A2(n23260), .ZN(n21496) );
  XNOR2HSV1 U24073 ( .A1(n21497), .A2(n21496), .ZN(n21498) );
  XNOR2HSV1 U24074 ( .A1(n21499), .A2(n21498), .ZN(n21501) );
  NAND2HSV0 U24075 ( .A1(n28614), .A2(n13993), .ZN(n21500) );
  XNOR2HSV1 U24076 ( .A1(n21501), .A2(n21500), .ZN(n21503) );
  NAND2HSV0 U24077 ( .A1(n24674), .A2(n14072), .ZN(n21502) );
  XNOR2HSV1 U24078 ( .A1(n21503), .A2(n21502), .ZN(n21507) );
  CLKNHSV0 U24079 ( .I(\pe5/got [6]), .ZN(n23940) );
  NOR2HSV0 U24080 ( .A1(n25350), .A2(n23940), .ZN(n21506) );
  NAND2HSV0 U24081 ( .A1(n21504), .A2(n28645), .ZN(n21505) );
  XOR3HSV1 U24082 ( .A1(n21507), .A2(n21506), .A3(n21505), .Z(n21508) );
  XNOR2HSV1 U24083 ( .A1(n21509), .A2(n21508), .ZN(n21513) );
  NOR2HSV0 U24084 ( .A1(n21613), .A2(n24685), .ZN(n21512) );
  OR2HSV1 U24085 ( .A1(n21614), .A2(n21510), .Z(n21511) );
  XOR3HSV1 U24086 ( .A1(n21513), .A2(n21512), .A3(n21511), .Z(n21514) );
  XNOR2HSV1 U24087 ( .A1(n21515), .A2(n21514), .ZN(n21517) );
  NAND2HSV0 U24088 ( .A1(n21452), .A2(n24636), .ZN(n21516) );
  NAND2HSV4 U24089 ( .A1(n21522), .A2(n21521), .ZN(n28473) );
  NAND2HSV0 U24090 ( .A1(n28473), .A2(n28647), .ZN(n21549) );
  NAND2HSV0 U24091 ( .A1(\pe5/ti_7[10] ), .A2(n13993), .ZN(n21545) );
  NAND2HSV0 U24092 ( .A1(n21523), .A2(n28640), .ZN(n21540) );
  NAND2HSV0 U24093 ( .A1(\pe5/aot [3]), .A2(\pe5/bq[7] ), .ZN(n21525) );
  NAND2HSV0 U24094 ( .A1(\pe5/aot [4]), .A2(\pe5/bq[6] ), .ZN(n21524) );
  XOR2HSV0 U24095 ( .A1(n21525), .A2(n21524), .Z(n21529) );
  NAND2HSV0 U24096 ( .A1(\pe5/aot [1]), .A2(\pe5/bq[9] ), .ZN(n21527) );
  NAND2HSV0 U24097 ( .A1(\pe5/aot [9]), .A2(\pe5/bq[1] ), .ZN(n21526) );
  XOR2HSV0 U24098 ( .A1(n21527), .A2(n21526), .Z(n21528) );
  XOR2HSV0 U24099 ( .A1(n21529), .A2(n21528), .Z(n21538) );
  NAND2HSV0 U24100 ( .A1(\pe5/aot [7]), .A2(\pe5/bq[3] ), .ZN(n23254) );
  NAND2HSV0 U24101 ( .A1(\pe5/aot [5]), .A2(\pe5/bq[8] ), .ZN(n21601) );
  CLKNAND2HSV0 U24102 ( .A1(\pe5/aot [2]), .A2(\pe5/bq[5] ), .ZN(n24443) );
  NOR2HSV0 U24103 ( .A1(n21601), .A2(n24443), .ZN(n21531) );
  AOI22HSV0 U24104 ( .A1(\pe5/aot [5]), .A2(\pe5/bq[5] ), .B1(\pe5/bq[8] ), 
        .B2(\pe5/aot [2]), .ZN(n21530) );
  NOR2HSV2 U24105 ( .A1(n21531), .A2(n21530), .ZN(n21536) );
  CLKNHSV0 U24106 ( .I(\pe5/aot [6]), .ZN(n23924) );
  NOR2HSV0 U24107 ( .A1(n23924), .A2(n21532), .ZN(n21534) );
  NAND2HSV0 U24108 ( .A1(\pe5/aot [8]), .A2(\pe5/bq[2] ), .ZN(n21533) );
  XOR2HSV0 U24109 ( .A1(n21534), .A2(n21533), .Z(n21535) );
  XOR3HSV2 U24110 ( .A1(n23254), .A2(n21536), .A3(n21535), .Z(n21537) );
  XOR2HSV0 U24111 ( .A1(n21538), .A2(n21537), .Z(n21539) );
  XNOR2HSV1 U24112 ( .A1(n21540), .A2(n21539), .ZN(n21543) );
  CLKNHSV2 U24113 ( .I(n28800), .ZN(n24684) );
  NOR2HSV1 U24114 ( .A1(n24684), .A2(n23260), .ZN(n21542) );
  OR2HSV1 U24115 ( .A1(n21614), .A2(n24364), .Z(n21541) );
  XOR3HSV2 U24116 ( .A1(n21543), .A2(n21542), .A3(n21541), .Z(n21544) );
  XNOR2HSV1 U24117 ( .A1(n21545), .A2(n21544), .ZN(n21547) );
  NAND2HSV0 U24118 ( .A1(n21452), .A2(\pe5/got [5]), .ZN(n21546) );
  XNOR2HSV1 U24119 ( .A1(n21547), .A2(n21546), .ZN(n21548) );
  XOR2HSV0 U24120 ( .A1(n21549), .A2(n21548), .Z(n21550) );
  NAND2HSV0 U24121 ( .A1(n12517), .A2(\pe5/got [5]), .ZN(n21567) );
  NAND2HSV0 U24122 ( .A1(n28473), .A2(n13993), .ZN(n21565) );
  NAND2HSV0 U24123 ( .A1(\pe5/aot [4]), .A2(\pe5/bq[4] ), .ZN(n21556) );
  NAND2HSV0 U24124 ( .A1(\pe5/aot [1]), .A2(\pe5/bq[7] ), .ZN(n21555) );
  CLKNAND2HSV1 U24125 ( .A1(\pe5/aot [3]), .A2(\pe5/bq[1] ), .ZN(n24329) );
  AO22HSV2 U24126 ( .A1(\pe5/aot [7]), .A2(\pe5/bq[1] ), .B1(\pe5/bq[5] ), 
        .B2(\pe5/aot [3]), .Z(n21557) );
  OAI21HSV0 U24127 ( .A1(n21558), .A2(n24329), .B(n21557), .ZN(n21559) );
  NOR2HSV0 U24128 ( .A1(n23924), .A2(n24439), .ZN(n24389) );
  CLKNHSV0 U24129 ( .I(\pe5/bq[6] ), .ZN(n24346) );
  CLKNAND2HSV1 U24130 ( .A1(\pe5/aot [2]), .A2(\pe5/bq[2] ), .ZN(n23233) );
  NAND2HSV0 U24131 ( .A1(\pe5/aot [5]), .A2(\pe5/bq[3] ), .ZN(n24328) );
  NAND2HSV0 U24132 ( .A1(n21452), .A2(\pe5/got [3]), .ZN(n21562) );
  XNOR2HSV1 U24133 ( .A1(n21563), .A2(n21562), .ZN(n21564) );
  XOR2HSV0 U24134 ( .A1(n21565), .A2(n21564), .Z(n21566) );
  XOR2HSV0 U24135 ( .A1(n21567), .A2(n21566), .Z(n21568) );
  NAND2HSV0 U24136 ( .A1(n12517), .A2(\pe5/got [2]), .ZN(n21581) );
  NAND2HSV0 U24137 ( .A1(n28473), .A2(n28640), .ZN(n21579) );
  CLKNAND2HSV0 U24138 ( .A1(\pe5/bq[1] ), .A2(\pe5/aot [4]), .ZN(n24390) );
  NAND2HSV0 U24139 ( .A1(\pe5/bq[4] ), .A2(\pe5/aot [1]), .ZN(n24323) );
  XOR2HSV0 U24140 ( .A1(n24390), .A2(n24323), .Z(n21577) );
  NOR2HSV1 U24141 ( .A1(n21573), .A2(n21572), .ZN(n21575) );
  NAND2HSV0 U24142 ( .A1(\pe5/aot [3]), .A2(\pe5/bq[2] ), .ZN(n21574) );
  XOR2HSV0 U24143 ( .A1(n21575), .A2(n21574), .Z(n21576) );
  XOR2HSV0 U24144 ( .A1(n21577), .A2(n21576), .Z(n21578) );
  XOR2HSV0 U24145 ( .A1(n21579), .A2(n21578), .Z(n21580) );
  NAND2HSV0 U24146 ( .A1(n24341), .A2(n14069), .ZN(n21623) );
  NAND2HSV0 U24147 ( .A1(\pe5/ti_7[10] ), .A2(n28645), .ZN(n21619) );
  NAND2HSV0 U24148 ( .A1(n11931), .A2(n13993), .ZN(n21612) );
  NAND2HSV0 U24149 ( .A1(n24674), .A2(n28640), .ZN(n21607) );
  NAND2HSV0 U24150 ( .A1(\pe5/aot [3]), .A2(\pe5/bq[10] ), .ZN(n21585) );
  NAND2HSV0 U24151 ( .A1(\pe5/aot [8]), .A2(\pe5/bq[5] ), .ZN(n21584) );
  XOR2HSV0 U24152 ( .A1(n21585), .A2(n21584), .Z(n21589) );
  NAND2HSV0 U24153 ( .A1(\pe5/aot [9]), .A2(\pe5/bq[4] ), .ZN(n21587) );
  INAND2HSV0 U24154 ( .A1(n14766), .B1(\pe5/aot [1]), .ZN(n21586) );
  XOR2HSV0 U24155 ( .A1(n21587), .A2(n21586), .Z(n21588) );
  XOR2HSV0 U24156 ( .A1(n21589), .A2(n21588), .Z(n21597) );
  NAND2HSV0 U24157 ( .A1(\pe5/aot [10]), .A2(\pe5/bq[3] ), .ZN(n21591) );
  NAND2HSV0 U24158 ( .A1(\pe5/aot [6]), .A2(\pe5/bq[7] ), .ZN(n21590) );
  XOR2HSV0 U24159 ( .A1(n21591), .A2(n21590), .Z(n21595) );
  NAND2HSV0 U24160 ( .A1(\pe5/aot [12]), .A2(\pe5/bq[1] ), .ZN(n21593) );
  NAND2HSV0 U24161 ( .A1(\pe5/aot [2]), .A2(\pe5/bq[11] ), .ZN(n21592) );
  XOR2HSV0 U24162 ( .A1(n21593), .A2(n21592), .Z(n21594) );
  XOR2HSV0 U24163 ( .A1(n21595), .A2(n21594), .Z(n21596) );
  XOR2HSV0 U24164 ( .A1(n21597), .A2(n21596), .Z(n21605) );
  NAND2HSV0 U24165 ( .A1(\pe5/aot [11]), .A2(\pe5/bq[2] ), .ZN(n21599) );
  NAND2HSV0 U24166 ( .A1(\pe5/aot [4]), .A2(\pe5/bq[9] ), .ZN(n21598) );
  XOR2HSV0 U24167 ( .A1(n21599), .A2(n21598), .Z(n21603) );
  NAND2HSV0 U24168 ( .A1(\pe5/aot [7]), .A2(\pe5/bq[6] ), .ZN(n21600) );
  XOR2HSV0 U24169 ( .A1(n21601), .A2(n21600), .Z(n21602) );
  XOR2HSV0 U24170 ( .A1(n21603), .A2(n21602), .Z(n21604) );
  XNOR2HSV1 U24171 ( .A1(n21605), .A2(n21604), .ZN(n21606) );
  XNOR2HSV1 U24172 ( .A1(n21607), .A2(n21606), .ZN(n21610) );
  NOR2HSV0 U24173 ( .A1(n25350), .A2(n23260), .ZN(n21609) );
  NAND2HSV0 U24174 ( .A1(n28478), .A2(\pe5/got [3]), .ZN(n21608) );
  XOR3HSV1 U24175 ( .A1(n21610), .A2(n21609), .A3(n21608), .Z(n21611) );
  XNOR2HSV1 U24176 ( .A1(n21612), .A2(n21611), .ZN(n21617) );
  NOR2HSV0 U24177 ( .A1(n21613), .A2(n24677), .ZN(n21616) );
  OR2HSV1 U24178 ( .A1(n21614), .A2(n23940), .Z(n21615) );
  XOR3HSV1 U24179 ( .A1(n21617), .A2(n21616), .A3(n21615), .Z(n21618) );
  XNOR2HSV1 U24180 ( .A1(n21619), .A2(n21618), .ZN(n21621) );
  NAND2HSV0 U24181 ( .A1(n21452), .A2(n24340), .ZN(n21620) );
  XNOR2HSV1 U24182 ( .A1(n21621), .A2(n21620), .ZN(n21622) );
  XOR2HSV0 U24183 ( .A1(n21623), .A2(n21622), .Z(n21624) );
  XOR2HSV0 U24184 ( .A1(n21625), .A2(n21624), .Z(n21626) );
  AND2HSV2 U24185 ( .A1(n21630), .A2(n28693), .Z(n21631) );
  CLKNHSV0 U24186 ( .I(n25364), .ZN(n21634) );
  NOR2HSV2 U24187 ( .A1(n21634), .A2(n21633), .ZN(n21635) );
  NAND2HSV2 U24188 ( .A1(n21636), .A2(n21635), .ZN(n21637) );
  XNOR2HSV4 U24189 ( .A1(n21640), .A2(n21639), .ZN(n21693) );
  CLKNAND2HSV1 U24190 ( .A1(n21701), .A2(\pe2/ti_7t [11]), .ZN(n22079) );
  CLKNAND2HSV1 U24191 ( .A1(n12624), .A2(n27543), .ZN(n21687) );
  NAND2HSV0 U24192 ( .A1(n14046), .A2(n21817), .ZN(n21680) );
  NOR2HSV1 U24193 ( .A1(n27452), .A2(n27498), .ZN(n21678) );
  INHSV2 U24194 ( .I(\pe2/got [5]), .ZN(n27663) );
  NOR2HSV0 U24195 ( .A1(n27423), .A2(n27663), .ZN(n21658) );
  INAND2HSV0 U24196 ( .A1(n27322), .B1(\pe2/aot [3]), .ZN(n21647) );
  NAND2HSV0 U24197 ( .A1(\pe2/aot [15]), .A2(\pe2/bq[4] ), .ZN(n21646) );
  XOR2HSV0 U24198 ( .A1(n21647), .A2(n21646), .Z(n21656) );
  NAND2HSV0 U24199 ( .A1(\pe2/aot [7]), .A2(\pe2/bq[12] ), .ZN(n21649) );
  NAND2HSV0 U24200 ( .A1(\pe2/aot [9]), .A2(\pe2/bq[10] ), .ZN(n21648) );
  XOR2HSV0 U24201 ( .A1(n21649), .A2(n21648), .Z(n21653) );
  NAND2HSV0 U24202 ( .A1(\pe2/aot [14]), .A2(\pe2/bq[5] ), .ZN(n21651) );
  NAND2HSV0 U24203 ( .A1(\pe2/aot [13]), .A2(\pe2/bq[6] ), .ZN(n21650) );
  XOR2HSV0 U24204 ( .A1(n21651), .A2(n21650), .Z(n21652) );
  XOR2HSV0 U24205 ( .A1(n21653), .A2(n21652), .Z(n21654) );
  XOR3HSV2 U24206 ( .A1(n21656), .A2(n21655), .A3(n21654), .Z(n21657) );
  XOR2HSV0 U24207 ( .A1(n21658), .A2(n21657), .Z(n21676) );
  NAND2HSV0 U24208 ( .A1(\pe2/got [3]), .A2(n27321), .ZN(n21660) );
  NAND2HSV0 U24209 ( .A1(\pe2/aot [4]), .A2(\pe2/bq[15] ), .ZN(n21659) );
  XOR2HSV0 U24210 ( .A1(n21660), .A2(n21659), .Z(n21664) );
  NAND2HSV0 U24211 ( .A1(\pe2/aot [6]), .A2(\pe2/bq[13] ), .ZN(n21662) );
  NAND2HSV0 U24212 ( .A1(\pe2/aot [5]), .A2(n27312), .ZN(n21661) );
  XOR2HSV0 U24213 ( .A1(n21662), .A2(n21661), .Z(n21663) );
  XOR2HSV0 U24214 ( .A1(n21664), .A2(n21663), .Z(n21672) );
  NAND2HSV0 U24215 ( .A1(\pe2/aot [11]), .A2(\pe2/bq[8] ), .ZN(n21666) );
  NAND2HSV0 U24216 ( .A1(\pe2/aot [10]), .A2(\pe2/bq[9] ), .ZN(n21665) );
  XOR2HSV0 U24217 ( .A1(n21666), .A2(n21665), .Z(n21670) );
  NAND2HSV0 U24218 ( .A1(n11953), .A2(\pe2/bq[3] ), .ZN(n21668) );
  NAND2HSV0 U24219 ( .A1(\pe2/aot [12]), .A2(\pe2/bq[7] ), .ZN(n21667) );
  XOR2HSV0 U24220 ( .A1(n21668), .A2(n21667), .Z(n21669) );
  XOR2HSV0 U24221 ( .A1(n21670), .A2(n21669), .Z(n21671) );
  XOR2HSV0 U24222 ( .A1(n21672), .A2(n21671), .Z(n21674) );
  BUFHSV2 U24223 ( .I(\pe2/got [4]), .Z(n28634) );
  NAND2HSV0 U24224 ( .A1(n28697), .A2(n28634), .ZN(n21673) );
  XNOR2HSV1 U24225 ( .A1(n21674), .A2(n21673), .ZN(n21675) );
  XOR2HSV0 U24226 ( .A1(n21676), .A2(n21675), .Z(n21677) );
  XOR2HSV0 U24227 ( .A1(n21678), .A2(n21677), .Z(n21679) );
  XNOR2HSV1 U24228 ( .A1(n21680), .A2(n21679), .ZN(n21682) );
  NAND2HSV0 U24229 ( .A1(n27485), .A2(\pe2/got [8]), .ZN(n21681) );
  XNOR2HSV1 U24230 ( .A1(n21682), .A2(n21681), .ZN(n21685) );
  NAND2HSV0 U24231 ( .A1(n27432), .A2(\pe2/got [10]), .ZN(n21683) );
  XOR3HSV2 U24232 ( .A1(n21685), .A2(n21684), .A3(n21683), .Z(n21686) );
  INHSV2 U24233 ( .I(n21692), .ZN(n21905) );
  NOR2HSV1 U24234 ( .A1(n25357), .A2(n21905), .ZN(n21695) );
  CLKNHSV0 U24235 ( .I(n21693), .ZN(n21694) );
  CLKNAND2HSV1 U24236 ( .A1(n21695), .A2(n21694), .ZN(n21711) );
  AND2HSV2 U24237 ( .A1(n21696), .A2(n28421), .Z(n21697) );
  CLKNAND2HSV1 U24238 ( .A1(n27344), .A2(n21702), .ZN(n21700) );
  CLKNHSV0 U24239 ( .I(n21703), .ZN(n21698) );
  NOR2HSV1 U24240 ( .A1(n21708), .A2(n21698), .ZN(n21699) );
  CLKNAND2HSV1 U24241 ( .A1(n21700), .A2(n21699), .ZN(n21710) );
  CLKNAND2HSV1 U24242 ( .A1(n21701), .A2(\pe2/ti_7t [12]), .ZN(n21704) );
  CLKNHSV0 U24243 ( .I(n21704), .ZN(n21707) );
  NAND2HSV0 U24244 ( .A1(n21703), .A2(n21702), .ZN(n21705) );
  OAI21HSV2 U24245 ( .A1(n21868), .A2(n21705), .B(n21704), .ZN(n21706) );
  OAI21HSV2 U24246 ( .A1(n21708), .A2(n21707), .B(n21706), .ZN(n21709) );
  CLKNAND2HSV2 U24247 ( .A1(n21710), .A2(n21709), .ZN(n25362) );
  XNOR2HSV4 U24248 ( .A1(n21712), .A2(n21814), .ZN(n28967) );
  CLKNAND2HSV2 U24249 ( .A1(n28967), .A2(n21713), .ZN(n27290) );
  NAND2HSV2 U24250 ( .A1(n28932), .A2(\pe2/ti_7t [14]), .ZN(n27289) );
  CLKNAND2HSV2 U24251 ( .A1(pov4[13]), .A2(n26923), .ZN(n22928) );
  CLKNAND2HSV1 U24252 ( .A1(n27976), .A2(\pe4/ti_7t [13]), .ZN(n22927) );
  CLKNAND2HSV3 U24253 ( .A1(n22928), .A2(n22927), .ZN(n28480) );
  CLKNHSV0 U24254 ( .I(\pe3/ti_7t [12]), .ZN(n21721) );
  AOI21HSV2 U24255 ( .A1(n21721), .A2(n21720), .B(n21719), .ZN(n23397) );
  NAND3HSV2 U24256 ( .A1(n23395), .A2(n23397), .A3(n21722), .ZN(n21723) );
  INOR2HSV2 U24257 ( .A1(n23400), .B1(n21723), .ZN(n21726) );
  OR2HSV1 U24258 ( .A1(n23372), .A2(n21724), .Z(n23403) );
  INHSV2 U24259 ( .I(n23403), .ZN(n21725) );
  AOI21HSV4 U24260 ( .A1(n21726), .A2(n21732), .B(n21725), .ZN(n23815) );
  INHSV2 U24261 ( .I(n23397), .ZN(n21728) );
  INHSV2 U24262 ( .I(n21728), .ZN(n27125) );
  NAND2HSV2 U24263 ( .A1(n21727), .A2(n27125), .ZN(n23390) );
  NOR2HSV0 U24264 ( .A1(n26291), .A2(n21728), .ZN(n21729) );
  CLKNAND2HSV1 U24265 ( .A1(n21730), .A2(n21729), .ZN(n23392) );
  NAND3HSV2 U24266 ( .A1(n23390), .A2(n15333), .A3(n23392), .ZN(n21731) );
  INHSV2 U24267 ( .I(n21731), .ZN(n21733) );
  INHSV3 U24268 ( .I(n21732), .ZN(n27127) );
  CLKNAND2HSV3 U24269 ( .A1(n21733), .A2(n27127), .ZN(n23814) );
  NAND2HSV4 U24270 ( .A1(n23815), .A2(n23814), .ZN(n28652) );
  NOR2HSV2 U24271 ( .A1(n23437), .A2(n25515), .ZN(n21735) );
  NOR2HSV1 U24272 ( .A1(n21736), .A2(n25688), .ZN(n21740) );
  CLKNHSV0 U24273 ( .I(n21737), .ZN(n25244) );
  IOA21HSV4 U24274 ( .A1(n21740), .A2(n25244), .B(n21739), .ZN(n28996) );
  INHSV2 U24275 ( .I(n21741), .ZN(n22490) );
  NAND2HSV4 U24276 ( .A1(n21743), .A2(n21742), .ZN(n28662) );
  CLKNHSV0 U24277 ( .I(n27277), .ZN(n28805) );
  NAND2HSV0 U24278 ( .A1(n12267), .A2(n15813), .ZN(n21746) );
  INAND2HSV0 U24279 ( .A1(n21746), .B1(n27877), .ZN(n21747) );
  CLKNAND2HSV1 U24280 ( .A1(n21748), .A2(n21747), .ZN(pov4[10]) );
  XNOR2HSV0 U24281 ( .A1(n21750), .A2(n21749), .ZN(n21751) );
  XNOR2HSV0 U24282 ( .A1(n21752), .A2(n21751), .ZN(n29047) );
  INHSV2 U24283 ( .I(n21753), .ZN(n28427) );
  CLKNAND2HSV0 U24284 ( .A1(n21755), .A2(n21754), .ZN(n28649) );
  CLKNHSV0 U24285 ( .I(\pe5/bq[11] ), .ZN(n21756) );
  INHSV1 U24286 ( .I(n21756), .ZN(n21757) );
  MUX2HSV2 U24287 ( .I0(n21757), .I1(bo5[11]), .S(n21758), .Z(n28711) );
  MUX2HSV2 U24288 ( .I0(\pe5/bq[1] ), .I1(bo5[1]), .S(n21758), .Z(n28866) );
  MUX2HSV1 U24289 ( .I0(bo4[13]), .I1(n26961), .S(n21759), .Z(n28856) );
  BUFHSV2 U24290 ( .I(n22114), .Z(n27311) );
  BUFHSV2 U24291 ( .I(n27311), .Z(n23503) );
  MUX2HSV1 U24292 ( .I0(bo2[16]), .I1(n21842), .S(n23503), .Z(n28822) );
  MUX2HSV1 U24293 ( .I0(bo11[15]), .I1(n24997), .S(n22111), .Z(n28725) );
  MUX2HSV1 U24294 ( .I0(bo9[15]), .I1(n21761), .S(n21760), .Z(n28730) );
  MUX2HSV2 U24295 ( .I0(bo8[2]), .I1(n21762), .S(n25625), .Z(n28896) );
  INHSV2 U24296 ( .I(n26940), .ZN(n28433) );
  CLKNHSV0 U24297 ( .I(n21763), .ZN(n28876) );
  MUX2HSV1 U24298 ( .I0(bo7[13]), .I1(\pe7/bq[13] ), .S(n28876), .Z(n28784) );
  MUX2HSV1 U24299 ( .I0(bo3[13]), .I1(\pe3/bq[13] ), .S(n23516), .Z(n28839) );
  CLKNHSV0 U24300 ( .I(\pe6/bq[1] ), .ZN(n25964) );
  MUX2HSV1 U24301 ( .I0(bo6[1]), .I1(\pe6/bq[1] ), .S(n12437), .Z(n28773) );
  INHSV2 U24302 ( .I(\pe4/got [1]), .ZN(n23986) );
  INHSV2 U24303 ( .I(\pe10/got [1]), .ZN(n26186) );
  CLKNHSV0 U24304 ( .I(n26186), .ZN(n28633) );
  NAND2HSV2 U24305 ( .A1(n25784), .A2(n26065), .ZN(n21783) );
  NAND2HSV0 U24306 ( .A1(n22078), .A2(\pe6/got [2]), .ZN(n21777) );
  NOR2HSV2 U24307 ( .A1(n25818), .A2(n21766), .ZN(n21775) );
  NAND2HSV0 U24308 ( .A1(\pe6/aot [4]), .A2(\pe6/bq[2] ), .ZN(n21773) );
  CLKNAND2HSV0 U24309 ( .A1(\pe6/bq[3] ), .A2(\pe6/aot [5]), .ZN(n25924) );
  NAND2HSV0 U24310 ( .A1(\pe6/aot [3]), .A2(\pe6/bq[1] ), .ZN(n24000) );
  NOR2HSV0 U24311 ( .A1(n25924), .A2(n24000), .ZN(n21768) );
  AOI22HSV0 U24312 ( .A1(\pe6/aot [5]), .A2(\pe6/bq[1] ), .B1(\pe6/bq[3] ), 
        .B2(\pe6/aot [3]), .ZN(n21767) );
  NOR2HSV2 U24313 ( .A1(n21768), .A2(n21767), .ZN(n21772) );
  NAND2HSV0 U24314 ( .A1(\pe6/aot [2]), .A2(\pe6/bq[4] ), .ZN(n21770) );
  NAND2HSV0 U24315 ( .A1(\pe6/aot [1]), .A2(\pe6/bq[5] ), .ZN(n21769) );
  XOR2HSV0 U24316 ( .A1(n21770), .A2(n21769), .Z(n21771) );
  XOR3HSV2 U24317 ( .A1(n21773), .A2(n21772), .A3(n21771), .Z(n21774) );
  XOR2HSV0 U24318 ( .A1(n21775), .A2(n21774), .Z(n21776) );
  XOR2HSV0 U24319 ( .A1(n21777), .A2(n21776), .Z(n21778) );
  XOR2HSV0 U24320 ( .A1(n21779), .A2(n21778), .Z(n21780) );
  NAND2HSV2 U24321 ( .A1(n25414), .A2(\pe11/got [6]), .ZN(n21810) );
  INHSV2 U24322 ( .I(n21785), .ZN(n23436) );
  CLKNAND2HSV1 U24323 ( .A1(n21785), .A2(n21784), .ZN(n21786) );
  NAND2HSV2 U24324 ( .A1(n24893), .A2(\pe11/got [5]), .ZN(n21808) );
  BUFHSV8 U24325 ( .I(n28918), .Z(n25137) );
  NAND2HSV0 U24326 ( .A1(n25137), .A2(\pe11/got [3]), .ZN(n21804) );
  NAND2HSV0 U24327 ( .A1(n14064), .A2(\pe11/got [2]), .ZN(n21802) );
  CLKNHSV0 U24328 ( .I(n21787), .ZN(n23300) );
  CLKNHSV1 U24329 ( .I(n23300), .ZN(n25169) );
  NAND2HSV0 U24330 ( .A1(n25169), .A2(\pe11/got [1]), .ZN(n21800) );
  NAND2HSV0 U24331 ( .A1(\pe11/bq[4] ), .A2(\pe11/aot [4]), .ZN(n21789) );
  NAND2HSV0 U24332 ( .A1(\pe11/bq[5] ), .A2(\pe11/aot [3]), .ZN(n21788) );
  XOR2HSV0 U24333 ( .A1(n21789), .A2(n21788), .Z(n21793) );
  NAND2HSV0 U24334 ( .A1(\pe11/bq[1] ), .A2(\pe11/aot [7]), .ZN(n21791) );
  NAND2HSV0 U24335 ( .A1(\pe11/bq[3] ), .A2(\pe11/aot [5]), .ZN(n21790) );
  XOR2HSV0 U24336 ( .A1(n21791), .A2(n21790), .Z(n21792) );
  XOR2HSV0 U24337 ( .A1(n21793), .A2(n21792), .Z(n21798) );
  NAND2HSV0 U24338 ( .A1(\pe11/bq[6] ), .A2(\pe11/aot [2]), .ZN(n21795) );
  NAND2HSV0 U24339 ( .A1(\pe11/bq[7] ), .A2(\pe11/aot [1]), .ZN(n21794) );
  XOR2HSV0 U24340 ( .A1(n21795), .A2(n21794), .Z(n21796) );
  NAND2HSV0 U24341 ( .A1(\pe11/bq[2] ), .A2(\pe11/aot [6]), .ZN(n24769) );
  XNOR2HSV1 U24342 ( .A1(n21796), .A2(n24769), .ZN(n21797) );
  XNOR2HSV1 U24343 ( .A1(n21798), .A2(n21797), .ZN(n21799) );
  XOR2HSV0 U24344 ( .A1(n21800), .A2(n21799), .Z(n21801) );
  XOR2HSV0 U24345 ( .A1(n21802), .A2(n21801), .Z(n21803) );
  XNOR2HSV1 U24346 ( .A1(n21804), .A2(n21803), .ZN(n21806) );
  XNOR2HSV4 U24347 ( .A1(n21810), .A2(n21809), .ZN(n21812) );
  CLKNAND2HSV1 U24348 ( .A1(n28927), .A2(\pe11/got [7]), .ZN(n21811) );
  XOR2HSV0 U24349 ( .A1(n21812), .A2(n21811), .Z(\pe11/poht [9]) );
  OAI21HSV1 U24350 ( .A1(n21813), .A2(\pe2/ti_7t [14]), .B(\pe2/got [16]), 
        .ZN(n23434) );
  NOR2HSV2 U24351 ( .A1(n27277), .A2(n17781), .ZN(n21865) );
  CLKNAND2HSV1 U24352 ( .A1(n21816), .A2(\pe2/got [10]), .ZN(n21863) );
  NAND2HSV0 U24353 ( .A1(n14003), .A2(n21817), .ZN(n21856) );
  INHSV2 U24354 ( .I(n27452), .ZN(n28954) );
  BUFHSV2 U24355 ( .I(\pe2/got [5]), .Z(n27719) );
  NAND2HSV0 U24356 ( .A1(n28954), .A2(n27719), .ZN(n21854) );
  INHSV2 U24357 ( .I(\pe2/got [4]), .ZN(n27718) );
  NOR2HSV0 U24358 ( .A1(n27423), .A2(n27718), .ZN(n21833) );
  NAND2HSV0 U24359 ( .A1(\pe2/bq[6] ), .A2(\pe2/aot [12]), .ZN(n27499) );
  NAND2HSV0 U24360 ( .A1(\pe2/aot [11]), .A2(\pe2/bq[7] ), .ZN(n27463) );
  XOR2HSV0 U24361 ( .A1(n27499), .A2(n27463), .Z(n21831) );
  NAND2HSV0 U24362 ( .A1(\pe2/bq[2] ), .A2(n11953), .ZN(n21819) );
  NAND2HSV0 U24363 ( .A1(\pe2/aot [13]), .A2(\pe2/bq[5] ), .ZN(n21818) );
  XOR2HSV0 U24364 ( .A1(n21819), .A2(n21818), .Z(n21822) );
  CLKNAND2HSV0 U24365 ( .A1(n27311), .A2(\pe2/pvq [15]), .ZN(n21820) );
  XNOR2HSV1 U24366 ( .A1(n21820), .A2(\pe2/phq [15]), .ZN(n21821) );
  XNOR2HSV1 U24367 ( .A1(n21822), .A2(n21821), .ZN(n21830) );
  NAND2HSV0 U24368 ( .A1(\pe2/bq[4] ), .A2(\pe2/aot [14]), .ZN(n21824) );
  NAND2HSV0 U24369 ( .A1(\pe2/aot [10]), .A2(\pe2/bq[8] ), .ZN(n21823) );
  XOR2HSV0 U24370 ( .A1(n21824), .A2(n21823), .Z(n21828) );
  NAND2HSV0 U24371 ( .A1(\pe2/aot [4]), .A2(\pe2/bq[14] ), .ZN(n21826) );
  NAND2HSV0 U24372 ( .A1(\pe2/aot [3]), .A2(\pe2/bq[15] ), .ZN(n21825) );
  XOR2HSV0 U24373 ( .A1(n21826), .A2(n21825), .Z(n21827) );
  XOR2HSV0 U24374 ( .A1(n21828), .A2(n21827), .Z(n21829) );
  XOR3HSV2 U24375 ( .A1(n21831), .A2(n21830), .A3(n21829), .Z(n21832) );
  XOR2HSV0 U24376 ( .A1(n21833), .A2(n21832), .Z(n21852) );
  NAND2HSV0 U24377 ( .A1(\pe2/aot [6]), .A2(\pe2/bq[12] ), .ZN(n21835) );
  NAND2HSV0 U24378 ( .A1(\pe2/aot [8]), .A2(\pe2/bq[10] ), .ZN(n21834) );
  XOR2HSV0 U24379 ( .A1(n21835), .A2(n21834), .Z(n21839) );
  NAND2HSV0 U24380 ( .A1(\pe2/aot [9]), .A2(\pe2/bq[9] ), .ZN(n21837) );
  NAND2HSV0 U24381 ( .A1(\pe2/aot [5]), .A2(\pe2/bq[13] ), .ZN(n21836) );
  XOR2HSV0 U24382 ( .A1(n21837), .A2(n21836), .Z(n21838) );
  XOR2HSV0 U24383 ( .A1(n21839), .A2(n21838), .Z(n21848) );
  NAND2HSV0 U24384 ( .A1(\pe2/aot [7]), .A2(\pe2/bq[11] ), .ZN(n21841) );
  NAND2HSV0 U24385 ( .A1(\pe2/aot [15]), .A2(\pe2/bq[3] ), .ZN(n21840) );
  XOR2HSV0 U24386 ( .A1(n21841), .A2(n21840), .Z(n21846) );
  NAND2HSV0 U24387 ( .A1(\pe2/got [2]), .A2(n27321), .ZN(n21844) );
  NAND2HSV0 U24388 ( .A1(\pe2/aot [2]), .A2(n21842), .ZN(n21843) );
  XOR2HSV0 U24389 ( .A1(n21844), .A2(n21843), .Z(n21845) );
  XOR2HSV0 U24390 ( .A1(n21846), .A2(n21845), .Z(n21847) );
  XOR2HSV0 U24391 ( .A1(n21848), .A2(n21847), .Z(n21850) );
  NAND2HSV0 U24392 ( .A1(n28697), .A2(n14052), .ZN(n21849) );
  XNOR2HSV1 U24393 ( .A1(n21850), .A2(n21849), .ZN(n21851) );
  XNOR2HSV1 U24394 ( .A1(n21852), .A2(n21851), .ZN(n21853) );
  XOR2HSV0 U24395 ( .A1(n21854), .A2(n21853), .Z(n21855) );
  XNOR2HSV1 U24396 ( .A1(n21856), .A2(n21855), .ZN(n21858) );
  NAND2HSV0 U24397 ( .A1(n14046), .A2(n27524), .ZN(n21857) );
  XNOR2HSV1 U24398 ( .A1(n21858), .A2(n21857), .ZN(n21861) );
  NOR2HSV2 U24399 ( .A1(n27527), .A2(n27645), .ZN(n21860) );
  NAND2HSV0 U24400 ( .A1(n28617), .A2(n27647), .ZN(n21859) );
  XOR3HSV2 U24401 ( .A1(n21861), .A2(n21860), .A3(n21859), .Z(n21862) );
  XNOR2HSV1 U24402 ( .A1(n21865), .A2(n21864), .ZN(n21872) );
  INHSV1 U24403 ( .I(n21866), .ZN(n21870) );
  CLKNAND2HSV2 U24404 ( .A1(n21868), .A2(n21867), .ZN(n21869) );
  INHSV3 U24405 ( .I(n23453), .ZN(n27439) );
  XNOR2HSV4 U24406 ( .A1(n21872), .A2(n21871), .ZN(n21874) );
  CLKNAND2HSV1 U24407 ( .A1(n21873), .A2(n21874), .ZN(n21878) );
  INHSV3 U24408 ( .I(n21874), .ZN(n21875) );
  CLKNAND2HSV4 U24409 ( .A1(n21878), .A2(n21877), .ZN(n21890) );
  NOR2HSV4 U24410 ( .A1(n11853), .A2(n21880), .ZN(n21882) );
  CLKNAND2HSV1 U24411 ( .A1(n25362), .A2(n17767), .ZN(n21883) );
  NAND3HSV4 U24412 ( .A1(n21885), .A2(n21884), .A3(n21883), .ZN(n21889) );
  XNOR2HSV4 U24413 ( .A1(n21890), .A2(n21889), .ZN(n23435) );
  CLKXOR2HSV2 U24414 ( .A1(n21886), .A2(n23435), .Z(n21888) );
  NOR2HSV2 U24415 ( .A1(n27731), .A2(n21235), .ZN(n21887) );
  CLKNAND2HSV4 U24416 ( .A1(n21888), .A2(n21887), .ZN(n23230) );
  NOR2HSV0 U24417 ( .A1(n22085), .A2(n21643), .ZN(n21898) );
  CLKNAND2HSV1 U24418 ( .A1(n21904), .A2(n21898), .ZN(n21896) );
  XNOR2HSV4 U24419 ( .A1(n21892), .A2(n21891), .ZN(n23433) );
  CLKNHSV0 U24420 ( .I(n23434), .ZN(n21899) );
  AND2HSV2 U24421 ( .A1(n21899), .A2(n21898), .Z(n21894) );
  NOR2HSV1 U24422 ( .A1(n21905), .A2(n21899), .ZN(n21893) );
  AOI21HSV2 U24423 ( .A1(n12285), .A2(n21894), .B(n21893), .ZN(n21895) );
  OAI22HSV2 U24424 ( .A1(n21896), .A2(n23433), .B1(n23435), .B2(n21895), .ZN(
        n21897) );
  OR2HSV1 U24425 ( .A1(n21905), .A2(n23434), .Z(n21906) );
  NOR2HSV4 U24426 ( .A1(n21908), .A2(n21907), .ZN(n23229) );
  CLKNAND2HSV1 U24427 ( .A1(n23230), .A2(n23229), .ZN(n28456) );
  NAND2HSV2 U24428 ( .A1(n24902), .A2(n20227), .ZN(n21963) );
  INHSV2 U24429 ( .I(n21909), .ZN(n24903) );
  CLKNAND2HSV1 U24430 ( .A1(n24893), .A2(\pe11/got [12]), .ZN(n21961) );
  NAND2HSV0 U24431 ( .A1(n25137), .A2(\pe11/got [10]), .ZN(n21957) );
  NAND2HSV0 U24432 ( .A1(n14063), .A2(\pe11/got [9]), .ZN(n21955) );
  NAND2HSV0 U24433 ( .A1(n25138), .A2(\pe11/got [7]), .ZN(n21951) );
  CLKNHSV1 U24434 ( .I(n21910), .ZN(n25139) );
  NAND2HSV0 U24435 ( .A1(n25139), .A2(\pe11/got [6]), .ZN(n21949) );
  NAND2HSV0 U24436 ( .A1(n28471), .A2(\pe11/got [5]), .ZN(n21947) );
  NAND2HSV0 U24437 ( .A1(\pe11/bq[13] ), .A2(\pe11/aot [2]), .ZN(n21912) );
  NAND2HSV0 U24438 ( .A1(\pe11/bq[14] ), .A2(\pe11/aot [1]), .ZN(n21911) );
  XOR2HSV0 U24439 ( .A1(n21912), .A2(n21911), .Z(n21916) );
  NAND2HSV0 U24440 ( .A1(\pe11/bq[1] ), .A2(n24771), .ZN(n21914) );
  NAND2HSV0 U24441 ( .A1(\pe11/bq[8] ), .A2(\pe11/aot [7]), .ZN(n21913) );
  XOR2HSV0 U24442 ( .A1(n21914), .A2(n21913), .Z(n21915) );
  XOR2HSV0 U24443 ( .A1(n21916), .A2(n21915), .Z(n21924) );
  NAND2HSV0 U24444 ( .A1(\pe11/bq[3] ), .A2(\pe11/aot [12]), .ZN(n21918) );
  NAND2HSV0 U24445 ( .A1(\pe11/bq[11] ), .A2(\pe11/aot [4]), .ZN(n21917) );
  XOR2HSV0 U24446 ( .A1(n21918), .A2(n21917), .Z(n21922) );
  NAND2HSV0 U24447 ( .A1(\pe11/bq[12] ), .A2(\pe11/aot [3]), .ZN(n21920) );
  NAND2HSV0 U24448 ( .A1(\pe11/bq[10] ), .A2(\pe11/aot [5]), .ZN(n21919) );
  XOR2HSV0 U24449 ( .A1(n21920), .A2(n21919), .Z(n21921) );
  XOR2HSV0 U24450 ( .A1(n21922), .A2(n21921), .Z(n21923) );
  XOR2HSV0 U24451 ( .A1(n21924), .A2(n21923), .Z(n21936) );
  NAND2HSV0 U24452 ( .A1(\pe11/bq[6] ), .A2(\pe11/aot [9]), .ZN(n21926) );
  NAND2HSV0 U24453 ( .A1(\pe11/bq[7] ), .A2(\pe11/aot [8]), .ZN(n21925) );
  XOR2HSV0 U24454 ( .A1(n21926), .A2(n21925), .Z(n21930) );
  NAND2HSV0 U24455 ( .A1(\pe11/bq[2] ), .A2(n12011), .ZN(n21928) );
  NAND2HSV0 U24456 ( .A1(\pe11/bq[4] ), .A2(\pe11/aot [11]), .ZN(n21927) );
  XOR2HSV0 U24457 ( .A1(n21928), .A2(n21927), .Z(n21929) );
  XOR2HSV0 U24458 ( .A1(n21930), .A2(n21929), .Z(n21934) );
  NAND2HSV0 U24459 ( .A1(\pe11/bq[9] ), .A2(\pe11/aot [6]), .ZN(n21931) );
  XOR2HSV0 U24460 ( .A1(n21932), .A2(n21931), .Z(n21933) );
  XNOR2HSV1 U24461 ( .A1(n21934), .A2(n21933), .ZN(n21935) );
  XNOR2HSV1 U24462 ( .A1(n21936), .A2(n21935), .ZN(n21938) );
  NAND2HSV0 U24463 ( .A1(n20506), .A2(\pe11/got [1]), .ZN(n21937) );
  XNOR2HSV1 U24464 ( .A1(n21938), .A2(n21937), .ZN(n21940) );
  NAND2HSV0 U24465 ( .A1(\pe11/got [2]), .A2(n25008), .ZN(n21939) );
  XOR2HSV0 U24466 ( .A1(n21940), .A2(n21939), .Z(n21943) );
  CLKNHSV0 U24467 ( .I(n21941), .ZN(n24966) );
  NAND2HSV0 U24468 ( .A1(n11804), .A2(\pe11/got [3]), .ZN(n21942) );
  XOR2HSV0 U24469 ( .A1(n21943), .A2(n21942), .Z(n21945) );
  NAND2HSV0 U24470 ( .A1(n11852), .A2(\pe11/got [4]), .ZN(n21944) );
  XOR2HSV0 U24471 ( .A1(n21945), .A2(n21944), .Z(n21946) );
  XOR2HSV0 U24472 ( .A1(n21947), .A2(n21946), .Z(n21948) );
  XOR2HSV0 U24473 ( .A1(n21949), .A2(n21948), .Z(n21950) );
  XOR2HSV0 U24474 ( .A1(n21951), .A2(n21950), .Z(n21953) );
  NAND2HSV0 U24475 ( .A1(n25169), .A2(\pe11/got [8]), .ZN(n21952) );
  XOR2HSV0 U24476 ( .A1(n21953), .A2(n21952), .Z(n21954) );
  XOR2HSV0 U24477 ( .A1(n21955), .A2(n21954), .Z(n21956) );
  XNOR2HSV1 U24478 ( .A1(n21957), .A2(n21956), .ZN(n21959) );
  XNOR2HSV4 U24479 ( .A1(n21963), .A2(n21962), .ZN(n21965) );
  INHSV1 U24480 ( .I(n21967), .ZN(n21970) );
  NAND2HSV2 U24481 ( .A1(n21988), .A2(n21968), .ZN(n21969) );
  NOR2HSV1 U24482 ( .A1(n21968), .A2(\pe4/ti_7t [13]), .ZN(n22820) );
  NOR2HSV1 U24483 ( .A1(n22820), .A2(n22895), .ZN(n26924) );
  NAND3HSV4 U24484 ( .A1(n13970), .A2(n21975), .A3(n21974), .ZN(n22915) );
  INHSV3 U24485 ( .I(n22915), .ZN(n26930) );
  NOR2HSV2 U24486 ( .A1(n21977), .A2(n21976), .ZN(n21978) );
  NAND2HSV2 U24487 ( .A1(n21978), .A2(n27907), .ZN(n22886) );
  NOR2HSV0 U24488 ( .A1(n21979), .A2(n15813), .ZN(n21982) );
  NAND3HSV1 U24489 ( .A1(n21981), .A2(n21982), .A3(n21980), .ZN(n22884) );
  NAND3HSV2 U24490 ( .A1(n21984), .A2(n21983), .A3(n21982), .ZN(n22883) );
  NOR2HSV0 U24491 ( .A1(n22881), .A2(n26919), .ZN(n21985) );
  NAND3HSV2 U24492 ( .A1(n22884), .A2(n22883), .A3(n21985), .ZN(n21986) );
  INHSV2 U24493 ( .I(n21986), .ZN(n21987) );
  CLKNHSV2 U24494 ( .I(n13963), .ZN(n21991) );
  INHSV4 U24495 ( .I(n21988), .ZN(n21989) );
  INHSV4 U24496 ( .I(n21989), .ZN(n22887) );
  CLKNHSV2 U24497 ( .I(n22887), .ZN(n21990) );
  CLKNAND2HSV2 U24498 ( .A1(n13963), .A2(n22887), .ZN(n22903) );
  CLKNHSV0 U24499 ( .I(n21992), .ZN(n21993) );
  NAND2HSV0 U24500 ( .A1(n21994), .A2(n13994), .ZN(n21995) );
  NAND2HSV0 U24501 ( .A1(n22825), .A2(\pe4/got [9]), .ZN(n22036) );
  NAND2HSV0 U24502 ( .A1(n28671), .A2(\pe4/got [5]), .ZN(n22012) );
  NAND2HSV0 U24503 ( .A1(n26958), .A2(\pe4/aot [4]), .ZN(n21999) );
  NAND2HSV0 U24504 ( .A1(\pe4/got [3]), .A2(n27128), .ZN(n21998) );
  XOR2HSV0 U24505 ( .A1(n21999), .A2(n21998), .Z(n22010) );
  NAND2HSV0 U24506 ( .A1(\pe4/aot [13]), .A2(\pe4/bq[3] ), .ZN(n22960) );
  NAND2HSV0 U24507 ( .A1(\pe4/bq[5] ), .A2(\pe4/aot [14]), .ZN(n22003) );
  NAND2HSV0 U24508 ( .A1(\pe4/aot [6]), .A2(n26961), .ZN(n22002) );
  XOR2HSV0 U24509 ( .A1(n22003), .A2(n22002), .Z(n22007) );
  NAND2HSV0 U24510 ( .A1(\pe4/aot [10]), .A2(\pe4/bq[9] ), .ZN(n22005) );
  NAND2HSV0 U24511 ( .A1(n28433), .A2(\pe4/bq[4] ), .ZN(n22004) );
  XOR2HSV0 U24512 ( .A1(n22005), .A2(n22004), .Z(n22006) );
  XOR2HSV0 U24513 ( .A1(n22007), .A2(n22006), .Z(n22008) );
  XOR3HSV2 U24514 ( .A1(n22010), .A2(n22009), .A3(n22008), .Z(n22011) );
  XOR2HSV0 U24515 ( .A1(n22012), .A2(n22011), .Z(n22029) );
  NAND2HSV0 U24516 ( .A1(\pe4/aot [8]), .A2(\pe4/bq[11] ), .ZN(n22014) );
  NAND2HSV0 U24517 ( .A1(\pe4/aot [11]), .A2(\pe4/bq[8] ), .ZN(n22013) );
  XOR2HSV0 U24518 ( .A1(n22014), .A2(n22013), .Z(n22018) );
  NAND2HSV0 U24519 ( .A1(\pe4/aot [12]), .A2(\pe4/bq[7] ), .ZN(n22016) );
  NAND2HSV0 U24520 ( .A1(\pe4/aot [5]), .A2(n27060), .ZN(n22015) );
  XOR2HSV0 U24521 ( .A1(n22016), .A2(n22015), .Z(n22017) );
  XOR2HSV0 U24522 ( .A1(n22018), .A2(n22017), .Z(n22025) );
  NAND2HSV0 U24523 ( .A1(\pe4/aot [9]), .A2(\pe4/bq[10] ), .ZN(n22020) );
  NAND2HSV0 U24524 ( .A1(\pe4/aot [7]), .A2(\pe4/bq[12] ), .ZN(n22019) );
  XOR2HSV0 U24525 ( .A1(n22020), .A2(n22019), .Z(n22023) );
  CLKNAND2HSV0 U24526 ( .A1(n27089), .A2(\pe4/pvq [14]), .ZN(n22021) );
  XOR2HSV0 U24527 ( .A1(n22021), .A2(\pe4/phq [14]), .Z(n22022) );
  XOR2HSV0 U24528 ( .A1(n22023), .A2(n22022), .Z(n22024) );
  XOR2HSV0 U24529 ( .A1(n22025), .A2(n22024), .Z(n22027) );
  NAND2HSV0 U24530 ( .A1(n28653), .A2(\pe4/got [4]), .ZN(n22026) );
  XNOR2HSV1 U24531 ( .A1(n22027), .A2(n22026), .ZN(n22028) );
  XNOR2HSV1 U24532 ( .A1(n22029), .A2(n22028), .ZN(n22032) );
  NOR2HSV0 U24533 ( .A1(n26981), .A2(n27905), .ZN(n22031) );
  NAND2HSV0 U24534 ( .A1(n27739), .A2(n13996), .ZN(n22030) );
  XOR3HSV2 U24535 ( .A1(n22032), .A2(n22031), .A3(n22030), .Z(n22034) );
  NAND2HSV0 U24536 ( .A1(n27830), .A2(\pe4/got [8]), .ZN(n22033) );
  XOR2HSV0 U24537 ( .A1(n22034), .A2(n22033), .Z(n22035) );
  XNOR2HSV1 U24538 ( .A1(n22036), .A2(n22035), .ZN(n22037) );
  XNOR2HSV1 U24539 ( .A1(n22038), .A2(n22037), .ZN(n22039) );
  XNOR2HSV4 U24540 ( .A1(n22045), .A2(n22044), .ZN(n22904) );
  INHSV2 U24541 ( .I(n22051), .ZN(n22066) );
  NOR3HSV2 U24542 ( .A1(n26825), .A2(n22074), .A3(n22054), .ZN(n22049) );
  INHSV2 U24543 ( .I(n22047), .ZN(n22048) );
  CLKNAND2HSV1 U24544 ( .A1(n22049), .A2(n22048), .ZN(n22065) );
  NAND2HSV2 U24545 ( .A1(n22050), .A2(\pe1/ti_7t [14]), .ZN(n22053) );
  OAI21HSV2 U24546 ( .A1(n22051), .A2(n22050), .B(n22053), .ZN(n22063) );
  BUFHSV3 U24547 ( .I(n22052), .Z(n27137) );
  CLKNHSV0 U24548 ( .I(n22053), .ZN(n22055) );
  NOR2HSV2 U24549 ( .A1(n22055), .A2(n22054), .ZN(n22057) );
  NAND3HSV2 U24550 ( .A1(n27137), .A2(n22057), .A3(n22075), .ZN(n22060) );
  NAND3HSV2 U24551 ( .A1(n22058), .A2(n22057), .A3(n22056), .ZN(n22059) );
  NAND2HSV2 U24552 ( .A1(n22060), .A2(n22059), .ZN(n22061) );
  INHSV2 U24553 ( .I(n22061), .ZN(n22062) );
  INHSV4 U24554 ( .I(n22067), .ZN(n25914) );
  BUFHSV2 U24555 ( .I(n22068), .Z(n22070) );
  NOR2HSV4 U24556 ( .A1(n22070), .A2(n25678), .ZN(n27220) );
  CLKNAND2HSV1 U24557 ( .A1(n22072), .A2(n12277), .ZN(n22073) );
  NOR2HSV4 U24558 ( .A1(n22073), .A2(n25678), .ZN(n27217) );
  OA21HSV2 U24559 ( .A1(n27217), .A2(n22074), .B(n26827), .Z(n22076) );
  MUX2NHSV2 U24560 ( .I0(n22077), .I1(n22076), .S(n22075), .ZN(n26415) );
  CLKNAND2HSV3 U24561 ( .A1(n26415), .A2(n26414), .ZN(n28700) );
  INHSV2 U24562 ( .I(n22081), .ZN(n28616) );
  XNOR2HSV0 U24563 ( .A1(n22083), .A2(n22082), .ZN(n28976) );
  CLKBUFHSV4 U24564 ( .I(n12624), .Z(n27614) );
  NAND2HSV0 U24565 ( .A1(n27614), .A2(n22085), .ZN(n22087) );
  XNOR2HSV0 U24566 ( .A1(n22087), .A2(n21150), .ZN(n22088) );
  XNOR2HSV0 U24567 ( .A1(n22088), .A2(n21218), .ZN(\pov2[10] ) );
  NAND2HSV0 U24568 ( .A1(n14067), .A2(n28610), .ZN(n22090) );
  XOR2HSV0 U24569 ( .A1(n22090), .A2(n22089), .Z(n29014) );
  NAND2HSV0 U24570 ( .A1(n22093), .A2(n14631), .ZN(n22098) );
  CLKNHSV0 U24571 ( .I(n22094), .ZN(n22095) );
  CLKNHSV0 U24572 ( .I(n22095), .ZN(n22096) );
  NAND3HSV0 U24573 ( .A1(n22098), .A2(n22096), .A3(n22097), .ZN(n22101) );
  CLKNHSV0 U24574 ( .I(n22099), .ZN(n22100) );
  XNOR2HSV0 U24575 ( .A1(n22101), .A2(n22100), .ZN(n28992) );
  DELHS4 U24576 ( .I(n22104), .Z(n22105) );
  CLKNHSV0 U24577 ( .I(rst), .ZN(n23791) );
  CLKNHSV0 U24578 ( .I(n23799), .ZN(n28530) );
  MUX2HSV2 U24579 ( .I0(bo11[5]), .I1(n22106), .S(n24980), .Z(n28722) );
  CLKNHSV0 U24580 ( .I(\pe6/bq[10] ), .ZN(n22108) );
  INHSV2 U24581 ( .I(n22108), .ZN(n22110) );
  MUX2HSV2 U24582 ( .I0(bo6[10]), .I1(n22110), .S(n22109), .Z(n28873) );
  MUX2HSV1 U24583 ( .I0(bo10[10]), .I1(\pe10/bq[10] ), .S(n23513), .Z(n28905)
         );
  BUFHSV2 U24584 ( .I(n22111), .Z(n27057) );
  MUX2HSV2 U24585 ( .I0(bo11[12]), .I1(\pe11/bq[12] ), .S(n27057), .Z(n28915)
         );
  CLKNHSV0 U24586 ( .I(\pe2/bq[15] ), .ZN(n22113) );
  INHSV2 U24587 ( .I(n22113), .ZN(n27239) );
  MUX2HSV1 U24588 ( .I0(bo2[15]), .I1(n27239), .S(n23537), .Z(n28823) );
  INHSV2 U24589 ( .I(\pe1/bq[3] ), .ZN(n27157) );
  INHSV2 U24590 ( .I(n24316), .ZN(n27062) );
  MUX2HSV2 U24591 ( .I0(bo1[4]), .I1(\pe1/bq[4] ), .S(n27062), .Z(n28820) );
  INHSV2 U24592 ( .I(n28623), .ZN(n23547) );
  MUX2HSV2 U24593 ( .I0(bo8[7]), .I1(\pe8/bq[7] ), .S(n25625), .Z(n28890) );
  CLKNHSV0 U24594 ( .I(n22115), .ZN(n28660) );
  NAND2HSV2 U24595 ( .A1(n28420), .A2(n25602), .ZN(n22193) );
  NOR2HSV2 U24596 ( .A1(n22126), .A2(n22118), .ZN(n22120) );
  CLKNAND2HSV1 U24597 ( .A1(n22120), .A2(n22119), .ZN(n22123) );
  CLKNHSV0 U24598 ( .I(\pe8/ti_7t [13]), .ZN(n22121) );
  AOI21HSV2 U24599 ( .A1(n22121), .A2(n18767), .B(n28667), .ZN(n22122) );
  NAND2HSV2 U24600 ( .A1(n22123), .A2(n22122), .ZN(n23422) );
  CLKNHSV0 U24601 ( .I(n23422), .ZN(n22124) );
  NAND2HSV2 U24602 ( .A1(n22124), .A2(n23423), .ZN(n22133) );
  CLKAND2HSV1 U24603 ( .A1(n22126), .A2(n22125), .Z(n22127) );
  NAND2HSV2 U24604 ( .A1(n23444), .A2(n22127), .ZN(n23421) );
  CLKNAND2HSV1 U24605 ( .A1(n23421), .A2(n22128), .ZN(n22132) );
  OAI22HSV2 U24606 ( .A1(n23423), .A2(n23421), .B1(n28685), .B2(n22129), .ZN(
        n22130) );
  INHSV2 U24607 ( .I(n22130), .ZN(n22131) );
  OAI21HSV4 U24608 ( .A1(n22133), .A2(n22132), .B(n22131), .ZN(n22135) );
  NOR2HSV2 U24609 ( .A1(n23423), .A2(ctro8), .ZN(n22134) );
  NOR2HSV8 U24610 ( .A1(n22135), .A2(n13961), .ZN(n28692) );
  CLKNHSV1 U24611 ( .I(n28692), .ZN(n22246) );
  CLKNAND2HSV1 U24612 ( .A1(n22246), .A2(n22136), .ZN(n22191) );
  CLKNAND2HSV1 U24613 ( .A1(n23757), .A2(\pe8/got [12]), .ZN(n22189) );
  CLKNAND2HSV4 U24614 ( .A1(pov8[12]), .A2(n22137), .ZN(n22248) );
  NAND2HSV2 U24615 ( .A1(n22138), .A2(\pe8/ti_7t [12]), .ZN(n22247) );
  NAND2HSV0 U24616 ( .A1(n28698), .A2(n23653), .ZN(n22187) );
  INHSV1 U24617 ( .I(n22139), .ZN(n25186) );
  NAND2HSV0 U24618 ( .A1(n25186), .A2(n23605), .ZN(n22181) );
  NAND2HSV0 U24619 ( .A1(n28616), .A2(n14060), .ZN(n22179) );
  INHSV1 U24620 ( .I(n22141), .ZN(n25351) );
  NOR2HSV1 U24621 ( .A1(n25351), .A2(n22142), .ZN(n22177) );
  INAND2HSV2 U24622 ( .A1(n25582), .B1(\pe8/got [3]), .ZN(n22172) );
  NAND2HSV0 U24623 ( .A1(n25578), .A2(\pe8/got [2]), .ZN(n22170) );
  NAND2HSV0 U24624 ( .A1(\pe8/bq[5] ), .A2(\pe8/aot [10]), .ZN(n25559) );
  NAND2HSV0 U24625 ( .A1(\pe8/aot [9]), .A2(\pe8/bq[6] ), .ZN(n22143) );
  XOR2HSV0 U24626 ( .A1(n25559), .A2(n22143), .Z(n22166) );
  NAND2HSV0 U24627 ( .A1(\pe8/aot [3]), .A2(\pe8/bq[12] ), .ZN(n22145) );
  NAND2HSV0 U24628 ( .A1(\pe8/aot [4]), .A2(\pe8/bq[11] ), .ZN(n22144) );
  XOR2HSV0 U24629 ( .A1(n22145), .A2(n22144), .Z(n22149) );
  NAND2HSV0 U24630 ( .A1(\pe8/aot [12]), .A2(\pe8/bq[3] ), .ZN(n22147) );
  NAND2HSV0 U24631 ( .A1(\pe8/aot [11]), .A2(\pe8/bq[4] ), .ZN(n22146) );
  XOR2HSV0 U24632 ( .A1(n22147), .A2(n22146), .Z(n22148) );
  XNOR2HSV1 U24633 ( .A1(n22149), .A2(n22148), .ZN(n22165) );
  CLKNHSV0 U24634 ( .I(\pe8/aot [1]), .ZN(n25543) );
  NAND2HSV0 U24635 ( .A1(\pe8/aot [1]), .A2(\pe8/bq[7] ), .ZN(n23856) );
  NOR2HSV0 U24636 ( .A1(n22150), .A2(n23856), .ZN(n22152) );
  AOI22HSV0 U24637 ( .A1(\pe8/aot [8]), .A2(\pe8/bq[7] ), .B1(n23627), .B2(
        \pe8/aot [1]), .ZN(n22151) );
  NOR2HSV2 U24638 ( .A1(n22152), .A2(n22151), .ZN(n22156) );
  NAND2HSV0 U24639 ( .A1(\pe8/bq[2] ), .A2(\pe8/aot [14]), .ZN(n25558) );
  NAND2HSV0 U24640 ( .A1(\pe8/aot [13]), .A2(\pe8/bq[1] ), .ZN(n23606) );
  NOR2HSV0 U24641 ( .A1(n25558), .A2(n23606), .ZN(n22154) );
  AOI22HSV0 U24642 ( .A1(\pe8/bq[1] ), .A2(\pe8/aot [14]), .B1(\pe8/aot [13]), 
        .B2(\pe8/bq[2] ), .ZN(n22153) );
  NOR2HSV1 U24643 ( .A1(n22154), .A2(n22153), .ZN(n22155) );
  XOR2HSV0 U24644 ( .A1(n22156), .A2(n22155), .Z(n22164) );
  NAND2HSV0 U24645 ( .A1(\pe8/aot [2]), .A2(n25565), .ZN(n22158) );
  NAND2HSV0 U24646 ( .A1(\pe8/aot [5]), .A2(\pe8/bq[10] ), .ZN(n22157) );
  XOR2HSV0 U24647 ( .A1(n22158), .A2(n22157), .Z(n22162) );
  NAND2HSV0 U24648 ( .A1(\pe8/aot [6]), .A2(\pe8/bq[9] ), .ZN(n22160) );
  NAND2HSV0 U24649 ( .A1(\pe8/aot [7]), .A2(\pe8/bq[8] ), .ZN(n22159) );
  XOR2HSV0 U24650 ( .A1(n22160), .A2(n22159), .Z(n22161) );
  XOR2HSV0 U24651 ( .A1(n22162), .A2(n22161), .Z(n22163) );
  XOR4HSV1 U24652 ( .A1(n22166), .A2(n22165), .A3(n22164), .A4(n22163), .Z(
        n22168) );
  NAND2HSV0 U24653 ( .A1(n26230), .A2(n28788), .ZN(n22167) );
  XNOR2HSV1 U24654 ( .A1(n22168), .A2(n22167), .ZN(n22169) );
  XNOR2HSV1 U24655 ( .A1(n22170), .A2(n22169), .ZN(n22171) );
  XOR2HSV0 U24656 ( .A1(n22172), .A2(n22171), .Z(n22175) );
  NOR2HSV0 U24657 ( .A1(n22310), .A2(n22230), .ZN(n22173) );
  XOR3HSV1 U24658 ( .A1(n22175), .A2(n22174), .A3(n22173), .Z(n22176) );
  XNOR2HSV1 U24659 ( .A1(n22177), .A2(n22176), .ZN(n22178) );
  XNOR2HSV1 U24660 ( .A1(n22179), .A2(n22178), .ZN(n22180) );
  XOR2HSV0 U24661 ( .A1(n22181), .A2(n22180), .Z(n22183) );
  NAND2HSV0 U24662 ( .A1(n23721), .A2(n14059), .ZN(n22182) );
  XOR2HSV0 U24663 ( .A1(n22183), .A2(n22182), .Z(n22185) );
  NAND2HSV0 U24664 ( .A1(n25204), .A2(\pe8/got [10]), .ZN(n22184) );
  XNOR2HSV1 U24665 ( .A1(n22185), .A2(n22184), .ZN(n22186) );
  CLKNHSV0 U24666 ( .I(n22194), .ZN(n22192) );
  CLKNAND2HSV1 U24667 ( .A1(n22193), .A2(n22192), .ZN(n22197) );
  CLKNHSV1 U24668 ( .I(n22193), .ZN(n22195) );
  CLKNAND2HSV1 U24669 ( .A1(n22195), .A2(n22194), .ZN(n22196) );
  NAND2HSV0 U24670 ( .A1(\pe8/got [9]), .A2(n26229), .ZN(n22224) );
  NAND2HSV0 U24671 ( .A1(n26231), .A2(\pe8/got [8]), .ZN(n22223) );
  NAND2HSV0 U24672 ( .A1(n25186), .A2(\pe8/got [3]), .ZN(n22219) );
  NAND2HSV0 U24673 ( .A1(n28616), .A2(\pe8/got [2]), .ZN(n22217) );
  INHSV2 U24674 ( .I(\pe8/got [1]), .ZN(n25530) );
  NOR2HSV1 U24675 ( .A1(n25351), .A2(n25530), .ZN(n22215) );
  NAND2HSV0 U24676 ( .A1(\pe8/aot [8]), .A2(\pe8/bq[2] ), .ZN(n25195) );
  NAND2HSV0 U24677 ( .A1(\pe8/aot [6]), .A2(\pe8/bq[6] ), .ZN(n22261) );
  CLKNHSV0 U24678 ( .I(n22261), .ZN(n22201) );
  CLKNHSV0 U24679 ( .I(\pe8/aot [4]), .ZN(n22297) );
  INHSV2 U24680 ( .I(\pe8/bq[4] ), .ZN(n23722) );
  NOR2HSV0 U24681 ( .A1(n22297), .A2(n23722), .ZN(n23851) );
  AOI22HSV0 U24682 ( .A1(\pe8/aot [6]), .A2(\pe8/bq[4] ), .B1(\pe8/bq[6] ), 
        .B2(\pe8/aot [4]), .ZN(n22200) );
  AOI21HSV2 U24683 ( .A1(n22201), .A2(n23851), .B(n22200), .ZN(n22205) );
  NAND2HSV0 U24684 ( .A1(\pe8/aot [2]), .A2(\pe8/bq[8] ), .ZN(n22203) );
  NAND2HSV0 U24685 ( .A1(\pe8/aot [9]), .A2(\pe8/bq[1] ), .ZN(n22202) );
  XOR2HSV0 U24686 ( .A1(n22203), .A2(n22202), .Z(n22204) );
  XOR3HSV2 U24687 ( .A1(n25195), .A2(n22205), .A3(n22204), .Z(n22213) );
  NAND2HSV0 U24688 ( .A1(\pe8/aot [7]), .A2(\pe8/bq[3] ), .ZN(n22207) );
  NAND2HSV0 U24689 ( .A1(\pe8/aot [1]), .A2(\pe8/bq[9] ), .ZN(n22206) );
  XOR2HSV0 U24690 ( .A1(n22207), .A2(n22206), .Z(n22211) );
  NAND2HSV0 U24691 ( .A1(\pe8/aot [5]), .A2(\pe8/bq[5] ), .ZN(n22209) );
  NAND2HSV0 U24692 ( .A1(\pe8/aot [3]), .A2(\pe8/bq[7] ), .ZN(n22208) );
  XOR2HSV0 U24693 ( .A1(n22209), .A2(n22208), .Z(n22210) );
  XOR2HSV0 U24694 ( .A1(n22211), .A2(n22210), .Z(n22212) );
  XOR2HSV0 U24695 ( .A1(n22213), .A2(n22212), .Z(n22214) );
  XNOR2HSV1 U24696 ( .A1(n22215), .A2(n22214), .ZN(n22216) );
  XNOR2HSV1 U24697 ( .A1(n22217), .A2(n22216), .ZN(n22218) );
  XOR2HSV0 U24698 ( .A1(n22219), .A2(n22218), .Z(n22221) );
  NAND2HSV0 U24699 ( .A1(n28457), .A2(n25577), .ZN(n22220) );
  CLKNAND2HSV0 U24700 ( .A1(n22224), .A2(n22225), .ZN(n22229) );
  CLKNHSV0 U24701 ( .I(n22224), .ZN(n22227) );
  CLKNHSV0 U24702 ( .I(n22225), .ZN(n22226) );
  CLKNAND2HSV1 U24703 ( .A1(n22227), .A2(n22226), .ZN(n22228) );
  CLKNAND2HSV1 U24704 ( .A1(n22229), .A2(n22228), .ZN(\pe8/poht [7]) );
  NAND2HSV0 U24705 ( .A1(n23757), .A2(\pe8/got [3]), .ZN(n22243) );
  NAND2HSV0 U24706 ( .A1(n28698), .A2(\pe8/got [2]), .ZN(n22241) );
  NAND2HSV0 U24707 ( .A1(n25204), .A2(n26230), .ZN(n22239) );
  NAND2HSV0 U24708 ( .A1(\pe8/aot [1]), .A2(\pe8/bq[5] ), .ZN(n22232) );
  NAND2HSV0 U24709 ( .A1(\pe8/aot [2]), .A2(\pe8/bq[4] ), .ZN(n22231) );
  XOR2HSV0 U24710 ( .A1(n22232), .A2(n22231), .Z(n22233) );
  NAND2HSV0 U24711 ( .A1(\pe8/aot [4]), .A2(\pe8/bq[2] ), .ZN(n23726) );
  XNOR2HSV1 U24712 ( .A1(n22233), .A2(n23726), .ZN(n22237) );
  NAND2HSV0 U24713 ( .A1(\pe8/aot [3]), .A2(\pe8/bq[3] ), .ZN(n22235) );
  NAND2HSV0 U24714 ( .A1(\pe8/aot [5]), .A2(\pe8/bq[1] ), .ZN(n22234) );
  XOR2HSV0 U24715 ( .A1(n22235), .A2(n22234), .Z(n22236) );
  XNOR2HSV1 U24716 ( .A1(n22237), .A2(n22236), .ZN(n22238) );
  XOR2HSV0 U24717 ( .A1(n22239), .A2(n22238), .Z(n22240) );
  XOR2HSV0 U24718 ( .A1(n22241), .A2(n22240), .Z(n22242) );
  XNOR2HSV1 U24719 ( .A1(n22243), .A2(n22242), .ZN(n22244) );
  NAND2HSV2 U24720 ( .A1(n28420), .A2(n28618), .ZN(n22278) );
  NAND2HSV0 U24721 ( .A1(n22246), .A2(\pe8/got [10]), .ZN(n22276) );
  NAND2HSV4 U24722 ( .A1(n22248), .A2(n22247), .ZN(n25185) );
  NAND2HSV0 U24723 ( .A1(n28631), .A2(\pe8/got [5]), .ZN(n22274) );
  CLKNAND2HSV1 U24724 ( .A1(n22140), .A2(n25577), .ZN(n22272) );
  CLKNHSV0 U24725 ( .I(\pe8/got [3]), .ZN(n22309) );
  NOR2HSV1 U24726 ( .A1(n25528), .A2(n22309), .ZN(n22270) );
  NAND2HSV0 U24727 ( .A1(\pe8/aot [5]), .A2(\pe8/bq[7] ), .ZN(n23563) );
  NAND2HSV0 U24728 ( .A1(\pe8/aot [9]), .A2(\pe8/bq[3] ), .ZN(n22250) );
  NAND2HSV0 U24729 ( .A1(\pe8/aot [7]), .A2(\pe8/bq[5] ), .ZN(n22249) );
  XOR2HSV0 U24730 ( .A1(n22250), .A2(n22249), .Z(n22257) );
  CLKNHSV0 U24731 ( .I(\pe8/aot [10]), .ZN(n22251) );
  NOR2HSV0 U24732 ( .A1(n22251), .A2(n25555), .ZN(n23561) );
  CLKNHSV0 U24733 ( .I(\pe8/aot [2]), .ZN(n23760) );
  CLKNHSV0 U24734 ( .I(\pe8/bq[10] ), .ZN(n23723) );
  CLKNAND2HSV1 U24735 ( .A1(\pe8/bq[2] ), .A2(\pe8/aot [2]), .ZN(n26226) );
  NAND2HSV0 U24736 ( .A1(\pe8/aot [11]), .A2(\pe8/bq[1] ), .ZN(n22254) );
  NAND2HSV0 U24737 ( .A1(\pe8/aot [8]), .A2(\pe8/bq[4] ), .ZN(n22253) );
  XOR2HSV0 U24738 ( .A1(n22254), .A2(n22253), .Z(n22255) );
  XOR4HSV1 U24739 ( .A1(n23563), .A2(n22257), .A3(n22256), .A4(n22255), .Z(
        n22265) );
  NAND2HSV0 U24740 ( .A1(\pe8/aot [1]), .A2(\pe8/bq[11] ), .ZN(n22259) );
  NAND2HSV0 U24741 ( .A1(\pe8/aot [4]), .A2(\pe8/bq[8] ), .ZN(n22258) );
  XOR2HSV0 U24742 ( .A1(n22259), .A2(n22258), .Z(n22263) );
  NAND2HSV0 U24743 ( .A1(\pe8/aot [3]), .A2(\pe8/bq[9] ), .ZN(n22260) );
  XOR2HSV0 U24744 ( .A1(n22261), .A2(n22260), .Z(n22262) );
  XOR2HSV0 U24745 ( .A1(n22263), .A2(n22262), .Z(n22264) );
  XNOR2HSV1 U24746 ( .A1(n22265), .A2(n22264), .ZN(n22268) );
  NAND2HSV0 U24747 ( .A1(n26230), .A2(n28462), .ZN(n22266) );
  XOR3HSV1 U24748 ( .A1(n22268), .A2(n22267), .A3(n22266), .Z(n22269) );
  XNOR2HSV1 U24749 ( .A1(n22270), .A2(n22269), .ZN(n22271) );
  XNOR2HSV1 U24750 ( .A1(n22272), .A2(n22271), .ZN(n22273) );
  CLKNAND2HSV1 U24751 ( .A1(n22278), .A2(n22277), .ZN(n22282) );
  CLKNHSV1 U24752 ( .I(n22278), .ZN(n22280) );
  CLKNAND2HSV1 U24753 ( .A1(n22280), .A2(n22279), .ZN(n22281) );
  CLKNAND2HSV1 U24754 ( .A1(n22282), .A2(n22281), .ZN(\pe8/poht [5]) );
  CLKNAND2HSV0 U24755 ( .A1(\pe8/got [12]), .A2(n26231), .ZN(n22328) );
  CLKNAND2HSV1 U24756 ( .A1(n28426), .A2(n23653), .ZN(n22327) );
  NAND2HSV0 U24757 ( .A1(n25185), .A2(\pe8/got [10]), .ZN(n22325) );
  CLKNAND2HSV0 U24758 ( .A1(n28631), .A2(n14060), .ZN(n22319) );
  CLKNAND2HSV0 U24759 ( .A1(n28616), .A2(\pe8/got [6]), .ZN(n22317) );
  NOR2HSV1 U24760 ( .A1(n25351), .A2(n22283), .ZN(n22315) );
  NAND2HSV0 U24761 ( .A1(\pe8/bq[2] ), .A2(\pe8/aot [5]), .ZN(n23765) );
  NOR2HSV0 U24762 ( .A1(n22284), .A2(n23765), .ZN(n22286) );
  AOI22HSV0 U24763 ( .A1(\pe8/aot [12]), .A2(\pe8/bq[2] ), .B1(\pe8/bq[9] ), 
        .B2(\pe8/aot [5]), .ZN(n22285) );
  NOR2HSV2 U24764 ( .A1(n22286), .A2(n22285), .ZN(n22287) );
  NAND2HSV0 U24765 ( .A1(\pe8/aot [9]), .A2(\pe8/bq[5] ), .ZN(n23614) );
  XOR2HSV0 U24766 ( .A1(n22287), .A2(n23614), .Z(n22289) );
  NAND2HSV0 U24767 ( .A1(\pe8/aot [6]), .A2(\pe8/bq[8] ), .ZN(n23562) );
  XOR2HSV0 U24768 ( .A1(n23606), .A2(n23562), .Z(n22288) );
  XOR2HSV0 U24769 ( .A1(n22289), .A2(n22288), .Z(n22306) );
  NAND2HSV0 U24770 ( .A1(\pe8/aot [7]), .A2(\pe8/bq[7] ), .ZN(n22291) );
  NAND2HSV0 U24771 ( .A1(\pe8/aot [3]), .A2(\pe8/bq[11] ), .ZN(n22290) );
  XOR2HSV0 U24772 ( .A1(n22291), .A2(n22290), .Z(n22295) );
  NAND2HSV0 U24773 ( .A1(\pe8/aot [10]), .A2(\pe8/bq[4] ), .ZN(n22293) );
  NAND2HSV0 U24774 ( .A1(\pe8/aot [1]), .A2(n25565), .ZN(n22292) );
  XOR2HSV0 U24775 ( .A1(n22293), .A2(n22292), .Z(n22294) );
  XOR2HSV0 U24776 ( .A1(n22295), .A2(n22294), .Z(n22303) );
  NAND2HSV0 U24777 ( .A1(\pe8/bq[3] ), .A2(\pe8/aot [11]), .ZN(n23560) );
  NAND2HSV0 U24778 ( .A1(\pe8/aot [2]), .A2(\pe8/bq[12] ), .ZN(n22296) );
  XOR2HSV0 U24779 ( .A1(n23560), .A2(n22296), .Z(n22301) );
  NOR2HSV0 U24780 ( .A1(n22297), .A2(n23723), .ZN(n22299) );
  NAND2HSV0 U24781 ( .A1(\pe8/aot [8]), .A2(\pe8/bq[6] ), .ZN(n22298) );
  XOR2HSV0 U24782 ( .A1(n22299), .A2(n22298), .Z(n22300) );
  XOR2HSV0 U24783 ( .A1(n22301), .A2(n22300), .Z(n22302) );
  XOR2HSV0 U24784 ( .A1(n22303), .A2(n22302), .Z(n22305) );
  NAND2HSV0 U24785 ( .A1(n25578), .A2(n26230), .ZN(n22304) );
  XOR3HSV2 U24786 ( .A1(n22306), .A2(n22305), .A3(n22304), .Z(n22308) );
  INAND2HSV0 U24787 ( .A1(n23642), .B1(\pe8/got [2]), .ZN(n22307) );
  XOR2HSV0 U24788 ( .A1(n22308), .A2(n22307), .Z(n22313) );
  NOR2HSV0 U24789 ( .A1(n22310), .A2(n22309), .ZN(n22311) );
  XOR3HSV1 U24790 ( .A1(n22313), .A2(n22312), .A3(n22311), .Z(n22314) );
  XNOR2HSV1 U24791 ( .A1(n22315), .A2(n22314), .ZN(n22316) );
  XNOR2HSV1 U24792 ( .A1(n22317), .A2(n22316), .ZN(n22318) );
  XOR2HSV0 U24793 ( .A1(n22319), .A2(n22318), .Z(n22321) );
  NAND2HSV0 U24794 ( .A1(\pe8/got [8]), .A2(n28457), .ZN(n22320) );
  XOR2HSV0 U24795 ( .A1(n22321), .A2(n22320), .Z(n22323) );
  NAND2HSV0 U24796 ( .A1(n25204), .A2(n23721), .ZN(n22322) );
  XNOR2HSV1 U24797 ( .A1(n22323), .A2(n22322), .ZN(n22324) );
  XNOR2HSV1 U24798 ( .A1(n22325), .A2(n22324), .ZN(n22326) );
  XNOR2HSV1 U24799 ( .A1(n22327), .A2(n22326), .ZN(n22329) );
  CLKNHSV0 U24800 ( .I(\pe9/got [8]), .ZN(n28124) );
  NOR2HSV2 U24801 ( .A1(n28368), .A2(n28124), .ZN(n22365) );
  CLKNAND2HSV1 U24802 ( .A1(n28231), .A2(\pe9/got [7]), .ZN(n22363) );
  NAND2HSV0 U24803 ( .A1(n28437), .A2(\pe9/got [6]), .ZN(n22361) );
  NAND2HSV0 U24804 ( .A1(n28264), .A2(n28389), .ZN(n22357) );
  CLKNAND2HSV0 U24805 ( .A1(n28059), .A2(n28658), .ZN(n22352) );
  NAND2HSV0 U24806 ( .A1(\pe9/aot [6]), .A2(\pe9/bq[2] ), .ZN(n28326) );
  INHSV2 U24807 ( .I(\pe9/bq[7] ), .ZN(n28240) );
  NAND2HSV0 U24808 ( .A1(\pe9/aot [11]), .A2(\pe9/bq[2] ), .ZN(n28088) );
  OAI21HSV0 U24809 ( .A1(n22330), .A2(n28240), .B(n28088), .ZN(n22331) );
  OAI21HSV0 U24810 ( .A1(n28326), .A2(n22332), .B(n22331), .ZN(n22335) );
  NAND2HSV0 U24811 ( .A1(\pe9/aot [2]), .A2(\pe9/bq[5] ), .ZN(n28363) );
  XOR2HSV0 U24812 ( .A1(n22335), .A2(n22334), .Z(n22350) );
  NAND2HSV0 U24813 ( .A1(\pe9/aot [12]), .A2(\pe9/bq[1] ), .ZN(n22337) );
  NAND2HSV0 U24814 ( .A1(\pe9/aot [5]), .A2(\pe9/bq[8] ), .ZN(n22336) );
  XOR2HSV0 U24815 ( .A1(n22337), .A2(n22336), .Z(n22341) );
  NAND2HSV0 U24816 ( .A1(\pe9/aot [9]), .A2(\pe9/bq[4] ), .ZN(n22339) );
  NAND2HSV0 U24817 ( .A1(\pe9/aot [3]), .A2(\pe9/bq[10] ), .ZN(n22338) );
  XOR2HSV0 U24818 ( .A1(n22339), .A2(n22338), .Z(n22340) );
  XNOR2HSV1 U24819 ( .A1(n22341), .A2(n22340), .ZN(n22349) );
  NAND2HSV0 U24820 ( .A1(\pe9/aot [1]), .A2(\pe9/bq[12] ), .ZN(n22342) );
  XOR2HSV0 U24821 ( .A1(n22343), .A2(n22342), .Z(n22347) );
  NAND2HSV0 U24822 ( .A1(\pe9/aot [4]), .A2(\pe9/bq[9] ), .ZN(n22345) );
  NAND2HSV0 U24823 ( .A1(\pe9/aot [10]), .A2(\pe9/bq[3] ), .ZN(n22344) );
  XOR2HSV0 U24824 ( .A1(n22345), .A2(n22344), .Z(n22346) );
  XOR2HSV0 U24825 ( .A1(n22347), .A2(n22346), .Z(n22348) );
  XOR3HSV2 U24826 ( .A1(n22350), .A2(n22349), .A3(n22348), .Z(n22351) );
  XNOR2HSV1 U24827 ( .A1(n22352), .A2(n22351), .ZN(n22355) );
  CLKNAND2HSV0 U24828 ( .A1(n28189), .A2(\pe9/got [3]), .ZN(n22354) );
  NAND2HSV0 U24829 ( .A1(n28166), .A2(\pe9/got [2]), .ZN(n22353) );
  XOR3HSV2 U24830 ( .A1(n22355), .A2(n22354), .A3(n22353), .Z(n22356) );
  XNOR2HSV1 U24831 ( .A1(n22357), .A2(n22356), .ZN(n22359) );
  INHSV2 U24832 ( .I(n28790), .ZN(n28287) );
  OR2HSV1 U24833 ( .A1(n28287), .A2(n28262), .Z(n22358) );
  XNOR2HSV1 U24834 ( .A1(n22359), .A2(n22358), .ZN(n22360) );
  XNOR2HSV1 U24835 ( .A1(n22361), .A2(n22360), .ZN(n22362) );
  XNOR2HSV1 U24836 ( .A1(n22363), .A2(n22362), .ZN(n22364) );
  XOR2HSV0 U24837 ( .A1(n22365), .A2(n22364), .Z(n22367) );
  NAND2HSV0 U24838 ( .A1(n28580), .A2(n14073), .ZN(n22366) );
  NAND2HSV0 U24839 ( .A1(n28394), .A2(n28227), .ZN(n22368) );
  XOR2HSV0 U24840 ( .A1(n22369), .A2(n22368), .Z(n22372) );
  NAND3HSV2 U24841 ( .A1(n28404), .A2(n28423), .A3(n28412), .ZN(n22371) );
  NAND2HSV2 U24842 ( .A1(n25692), .A2(n25691), .ZN(n28414) );
  NAND2HSV0 U24843 ( .A1(n28414), .A2(n28134), .ZN(n22370) );
  XNOR3HSV1 U24844 ( .A1(n22372), .A2(n22371), .A3(n22370), .ZN(\pe9/poht [4])
         );
  INHSV2 U24845 ( .I(n28419), .ZN(n28316) );
  NOR2HSV2 U24846 ( .A1(n28316), .A2(n22116), .ZN(n22415) );
  CLKNAND2HSV1 U24847 ( .A1(n28317), .A2(n14073), .ZN(n22413) );
  NAND2HSV0 U24848 ( .A1(n28437), .A2(\pe9/got [8]), .ZN(n22411) );
  NAND2HSV0 U24849 ( .A1(n28264), .A2(\pe9/got [6]), .ZN(n22407) );
  NAND2HSV0 U24850 ( .A1(n18399), .A2(n28405), .ZN(n22402) );
  NAND2HSV0 U24851 ( .A1(\pe9/got [2]), .A2(n28804), .ZN(n22400) );
  NAND2HSV0 U24852 ( .A1(\pe9/aot [12]), .A2(\pe9/bq[3] ), .ZN(n22376) );
  XOR2HSV0 U24853 ( .A1(n22377), .A2(n22376), .Z(n22396) );
  NOR2HSV0 U24854 ( .A1(n28398), .A2(n22378), .ZN(n28095) );
  CLKNHSV0 U24855 ( .I(n22379), .ZN(n22381) );
  AOI22HSV0 U24856 ( .A1(\pe9/aot [2]), .A2(\pe9/bq[13] ), .B1(n23822), .B2(
        \pe9/aot [1]), .ZN(n22380) );
  AOI21HSV2 U24857 ( .A1(n28095), .A2(n22381), .B(n22380), .ZN(n22386) );
  NAND2HSV0 U24858 ( .A1(\pe9/aot [10]), .A2(\pe9/bq[2] ), .ZN(n28149) );
  NOR2HSV0 U24859 ( .A1(n22382), .A2(n28149), .ZN(n22384) );
  AOI22HSV0 U24860 ( .A1(\pe9/bq[2] ), .A2(\pe9/aot [13]), .B1(\pe9/aot [10]), 
        .B2(\pe9/bq[5] ), .ZN(n22383) );
  NOR2HSV1 U24861 ( .A1(n22384), .A2(n22383), .ZN(n22385) );
  XOR2HSV0 U24862 ( .A1(n22386), .A2(n22385), .Z(n22394) );
  NAND2HSV0 U24863 ( .A1(\pe9/aot [11]), .A2(\pe9/bq[4] ), .ZN(n22388) );
  NAND2HSV0 U24864 ( .A1(\pe9/aot [3]), .A2(\pe9/bq[12] ), .ZN(n22387) );
  XOR2HSV0 U24865 ( .A1(n22388), .A2(n22387), .Z(n22392) );
  NAND2HSV0 U24866 ( .A1(\pe9/aot [4]), .A2(\pe9/bq[11] ), .ZN(n22390) );
  NAND2HSV0 U24867 ( .A1(\pe9/aot [14]), .A2(\pe9/bq[1] ), .ZN(n22389) );
  XOR2HSV0 U24868 ( .A1(n22390), .A2(n22389), .Z(n22391) );
  XOR2HSV0 U24869 ( .A1(n22392), .A2(n22391), .Z(n22393) );
  XOR4HSV1 U24870 ( .A1(n22396), .A2(n22395), .A3(n22394), .A4(n22393), .Z(
        n22398) );
  NAND2HSV0 U24871 ( .A1(n11863), .A2(\pe9/got [1]), .ZN(n22397) );
  XNOR2HSV1 U24872 ( .A1(n22398), .A2(n22397), .ZN(n22399) );
  XNOR2HSV1 U24873 ( .A1(n22400), .A2(n22399), .ZN(n22401) );
  XNOR2HSV1 U24874 ( .A1(n22402), .A2(n22401), .ZN(n22405) );
  NAND2HSV0 U24875 ( .A1(n28689), .A2(n28643), .ZN(n22404) );
  NAND2HSV0 U24876 ( .A1(n28166), .A2(\pe9/got [4]), .ZN(n22403) );
  XOR3HSV1 U24877 ( .A1(n22405), .A2(n22404), .A3(n22403), .Z(n22406) );
  XNOR2HSV1 U24878 ( .A1(n22407), .A2(n22406), .ZN(n22409) );
  CLKNHSV1 U24879 ( .I(\pe9/got [7]), .ZN(n28348) );
  OR2HSV1 U24880 ( .A1(n28287), .A2(n28348), .Z(n22408) );
  XNOR2HSV1 U24881 ( .A1(n22409), .A2(n22408), .ZN(n22410) );
  XNOR2HSV1 U24882 ( .A1(n22411), .A2(n22410), .ZN(n22412) );
  XNOR2HSV1 U24883 ( .A1(n22413), .A2(n22412), .ZN(n22414) );
  XOR2HSV0 U24884 ( .A1(n22415), .A2(n22414), .Z(n22417) );
  CLKNAND2HSV0 U24885 ( .A1(n28580), .A2(n28423), .ZN(n22416) );
  NAND2HSV2 U24886 ( .A1(n22419), .A2(\pe10/ti_7t [13]), .ZN(n22689) );
  NOR2HSV2 U24887 ( .A1(n24451), .A2(n22637), .ZN(n22438) );
  CLKNAND2HSV1 U24888 ( .A1(n22419), .A2(\pe10/ti_7t [11]), .ZN(n22599) );
  NOR2HSV2 U24889 ( .A1(n26093), .A2(n27194), .ZN(n22429) );
  INHSV2 U24890 ( .I(n28674), .ZN(n26209) );
  BUFHSV2 U24891 ( .I(\pe10/got [1]), .Z(n27196) );
  NAND2HSV0 U24892 ( .A1(n26209), .A2(n27196), .ZN(n22427) );
  NAND2HSV0 U24893 ( .A1(\pe10/aot [4]), .A2(\pe10/bq[4] ), .ZN(n22766) );
  CLKNAND2HSV0 U24894 ( .A1(\pe10/aot [3]), .A2(\pe10/bq[3] ), .ZN(n22703) );
  NAND2HSV0 U24895 ( .A1(\pe10/bq[2] ), .A2(\pe10/aot [5]), .ZN(n22705) );
  NAND2HSV0 U24896 ( .A1(\pe10/aot [6]), .A2(\pe10/bq[1] ), .ZN(n22420) );
  XOR2HSV0 U24897 ( .A1(n22705), .A2(n22420), .Z(n22424) );
  NAND2HSV0 U24898 ( .A1(\pe10/aot [2]), .A2(\pe10/bq[5] ), .ZN(n22422) );
  NAND2HSV0 U24899 ( .A1(\pe10/aot [1]), .A2(\pe10/bq[6] ), .ZN(n22421) );
  XOR2HSV0 U24900 ( .A1(n22422), .A2(n22421), .Z(n22423) );
  XOR3HSV2 U24901 ( .A1(n22425), .A2(n22424), .A3(n22423), .Z(n22426) );
  XOR2HSV0 U24902 ( .A1(n22427), .A2(n22426), .Z(n22428) );
  XOR2HSV0 U24903 ( .A1(n22429), .A2(n22428), .Z(n22436) );
  CLKAND2HSV4 U24904 ( .A1(n22692), .A2(n22691), .Z(n22434) );
  CLKNAND2HSV2 U24905 ( .A1(n22433), .A2(n23716), .ZN(n22696) );
  INHSV2 U24906 ( .I(n22675), .ZN(n22598) );
  NAND2HSV0 U24907 ( .A1(n27197), .A2(\pe10/got [3]), .ZN(n22435) );
  XOR2HSV0 U24908 ( .A1(n22436), .A2(n22435), .Z(n22437) );
  CLKNHSV2 U24909 ( .I(n22440), .ZN(n22441) );
  CLKNAND2HSV0 U24910 ( .A1(n22509), .A2(n28644), .ZN(n22489) );
  INHSV2 U24911 ( .I(\pe10/got [8]), .ZN(n24452) );
  NOR2HSV2 U24912 ( .A1(n26096), .A2(n24452), .ZN(n22485) );
  NAND2HSV0 U24913 ( .A1(n28794), .A2(\pe10/got [6]), .ZN(n22481) );
  NAND2HSV0 U24914 ( .A1(\pe10/bq[4] ), .A2(\pe10/aot [14]), .ZN(n22527) );
  NAND2HSV0 U24915 ( .A1(\pe10/aot [11]), .A2(\pe10/bq[7] ), .ZN(n22443) );
  XOR2HSV0 U24916 ( .A1(n22527), .A2(n22443), .Z(n22457) );
  NAND2HSV0 U24917 ( .A1(\pe10/aot [10]), .A2(\pe10/bq[2] ), .ZN(n25224) );
  NOR2HSV0 U24918 ( .A1(n22444), .A2(n25224), .ZN(n22446) );
  AOI22HSV0 U24919 ( .A1(\pe10/bq[2] ), .A2(n28424), .B1(\pe10/aot [10]), .B2(
        \pe10/bq[8] ), .ZN(n22445) );
  NOR2HSV2 U24920 ( .A1(n22446), .A2(n22445), .ZN(n22447) );
  XNOR2HSV1 U24921 ( .A1(n22448), .A2(n22447), .ZN(n22456) );
  NAND2HSV0 U24922 ( .A1(\pe10/aot [4]), .A2(\pe10/bq[14] ), .ZN(n22450) );
  NAND2HSV0 U24923 ( .A1(\pe10/aot [9]), .A2(\pe10/bq[9] ), .ZN(n22449) );
  XOR2HSV0 U24924 ( .A1(n22450), .A2(n22449), .Z(n22454) );
  NAND2HSV0 U24925 ( .A1(\pe10/aot [8]), .A2(\pe10/bq[10] ), .ZN(n22452) );
  NAND2HSV0 U24926 ( .A1(\pe10/aot [3]), .A2(\pe10/bq[15] ), .ZN(n22451) );
  XOR2HSV0 U24927 ( .A1(n22452), .A2(n22451), .Z(n22453) );
  XOR2HSV0 U24928 ( .A1(n22454), .A2(n22453), .Z(n22455) );
  XOR3HSV2 U24929 ( .A1(n22457), .A2(n22456), .A3(n22455), .Z(n22477) );
  CLKNAND2HSV0 U24930 ( .A1(n28630), .A2(n26132), .ZN(n22476) );
  NAND2HSV0 U24931 ( .A1(n22458), .A2(n28637), .ZN(n22460) );
  NAND2HSV0 U24932 ( .A1(n16973), .A2(\pe10/bq[3] ), .ZN(n22459) );
  XOR2HSV0 U24933 ( .A1(n22460), .A2(n22459), .Z(n22464) );
  NAND2HSV0 U24934 ( .A1(\pe10/aot [13]), .A2(\pe10/bq[5] ), .ZN(n22462) );
  NAND2HSV0 U24935 ( .A1(\pe10/aot [12]), .A2(\pe10/bq[6] ), .ZN(n22461) );
  XOR2HSV0 U24936 ( .A1(n22462), .A2(n22461), .Z(n22463) );
  XOR2HSV0 U24937 ( .A1(n22464), .A2(n22463), .Z(n22472) );
  NAND2HSV0 U24938 ( .A1(\pe10/aot [2]), .A2(\pe10/bq[16] ), .ZN(n22466) );
  NAND2HSV0 U24939 ( .A1(\pe10/aot [5]), .A2(\pe10/bq[13] ), .ZN(n22465) );
  XOR2HSV0 U24940 ( .A1(n22466), .A2(n22465), .Z(n22470) );
  NAND2HSV0 U24941 ( .A1(\pe10/aot [6]), .A2(\pe10/bq[12] ), .ZN(n22468) );
  NAND2HSV0 U24942 ( .A1(\pe10/aot [7]), .A2(\pe10/bq[11] ), .ZN(n22467) );
  XOR2HSV0 U24943 ( .A1(n22468), .A2(n22467), .Z(n22469) );
  XOR2HSV0 U24944 ( .A1(n22470), .A2(n22469), .Z(n22471) );
  XOR2HSV0 U24945 ( .A1(n22472), .A2(n22471), .Z(n22474) );
  NAND2HSV0 U24946 ( .A1(n28666), .A2(\pe10/got [3]), .ZN(n22473) );
  XNOR2HSV1 U24947 ( .A1(n22474), .A2(n22473), .ZN(n22475) );
  XOR3HSV2 U24948 ( .A1(n22477), .A2(n22476), .A3(n22475), .Z(n22479) );
  NAND2HSV0 U24949 ( .A1(n28679), .A2(\pe10/got [5]), .ZN(n22478) );
  XNOR2HSV1 U24950 ( .A1(n22479), .A2(n22478), .ZN(n22480) );
  XNOR2HSV1 U24951 ( .A1(n22481), .A2(n22480), .ZN(n22483) );
  NAND2HSV0 U24952 ( .A1(n26131), .A2(\pe10/got [7]), .ZN(n22482) );
  XNOR2HSV1 U24953 ( .A1(n22483), .A2(n22482), .ZN(n22484) );
  XOR2HSV0 U24954 ( .A1(n22485), .A2(n22484), .Z(n22486) );
  XOR2HSV0 U24955 ( .A1(n22487), .A2(n22486), .Z(n22488) );
  XOR2HSV0 U24956 ( .A1(n22489), .A2(n22488), .Z(n22492) );
  NAND2HSV0 U24957 ( .A1(n21741), .A2(n16759), .ZN(n22491) );
  XNOR2HSV1 U24958 ( .A1(n22492), .A2(n22491), .ZN(n22494) );
  NAND2HSV0 U24959 ( .A1(n25244), .A2(n26212), .ZN(n22493) );
  XOR2HSV0 U24960 ( .A1(n22494), .A2(n22493), .Z(n22495) );
  XNOR2HSV4 U24961 ( .A1(n12278), .A2(n22495), .ZN(n22497) );
  CLKNAND2HSV2 U24962 ( .A1(n22675), .A2(n14070), .ZN(n22496) );
  XNOR2HSV4 U24963 ( .A1(n22497), .A2(n22496), .ZN(n25260) );
  CLKNAND2HSV1 U24964 ( .A1(n26218), .A2(n28988), .ZN(n22500) );
  CLKNHSV0 U24965 ( .I(n22500), .ZN(n22498) );
  CLKNAND2HSV2 U24966 ( .A1(n25260), .A2(n22500), .ZN(n22501) );
  INHSV2 U24967 ( .I(\pe10/ti_7t [15]), .ZN(n22503) );
  NAND2HSV0 U24968 ( .A1(n26221), .A2(\pe10/got [6]), .ZN(n22507) );
  CLKNHSV0 U24969 ( .I(n22507), .ZN(n22505) );
  NAND2HSV0 U24970 ( .A1(n13995), .A2(n23219), .ZN(n22563) );
  CLKNHSV0 U24971 ( .I(n22563), .ZN(n22560) );
  NOR2HSV2 U24972 ( .A1(n24451), .A2(n16729), .ZN(n22557) );
  NOR2HSV2 U24973 ( .A1(n26093), .A2(n22636), .ZN(n22553) );
  INHSV2 U24974 ( .I(n22509), .ZN(n22566) );
  INHSV2 U24975 ( .I(n22566), .ZN(n28620) );
  NAND2HSV0 U24976 ( .A1(n28620), .A2(n28642), .ZN(n22547) );
  NAND2HSV0 U24977 ( .A1(\pe10/got [7]), .A2(n26094), .ZN(n22545) );
  INHSV2 U24978 ( .I(\pe10/got [6]), .ZN(n26199) );
  NOR2HSV0 U24979 ( .A1(n26096), .A2(n26199), .ZN(n22543) );
  NAND2HSV0 U24980 ( .A1(n28794), .A2(n26132), .ZN(n22539) );
  NAND2HSV0 U24981 ( .A1(n26189), .A2(n27196), .ZN(n22535) );
  NAND2HSV0 U24982 ( .A1(n28630), .A2(n14065), .ZN(n22534) );
  NAND2HSV0 U24983 ( .A1(\pe10/aot [10]), .A2(\pe10/bq[6] ), .ZN(n22511) );
  NAND2HSV0 U24984 ( .A1(\pe10/aot [5]), .A2(\pe10/bq[11] ), .ZN(n22510) );
  XOR2HSV0 U24985 ( .A1(n22511), .A2(n22510), .Z(n22515) );
  NAND2HSV0 U24986 ( .A1(\pe10/aot [9]), .A2(\pe10/bq[7] ), .ZN(n22513) );
  NAND2HSV0 U24987 ( .A1(\pe10/aot [7]), .A2(\pe10/bq[9] ), .ZN(n22512) );
  XOR2HSV0 U24988 ( .A1(n22513), .A2(n22512), .Z(n22514) );
  XOR2HSV0 U24989 ( .A1(n22515), .A2(n22514), .Z(n22524) );
  NAND2HSV0 U24990 ( .A1(\pe10/aot [1]), .A2(n16897), .ZN(n22517) );
  NAND2HSV0 U24991 ( .A1(\pe10/aot [6]), .A2(\pe10/bq[10] ), .ZN(n22516) );
  XOR2HSV0 U24992 ( .A1(n22517), .A2(n22516), .Z(n22522) );
  CLKNHSV0 U24993 ( .I(\pe10/aot [8]), .ZN(n22518) );
  NOR2HSV0 U24994 ( .A1(n22518), .A2(n26101), .ZN(n22520) );
  NAND2HSV0 U24995 ( .A1(\pe10/aot [4]), .A2(\pe10/bq[12] ), .ZN(n22519) );
  XOR2HSV0 U24996 ( .A1(n22520), .A2(n22519), .Z(n22521) );
  XOR2HSV0 U24997 ( .A1(n22522), .A2(n22521), .Z(n22523) );
  XOR2HSV0 U24998 ( .A1(n22524), .A2(n22523), .Z(n22532) );
  CLKNHSV0 U24999 ( .I(\pe10/aot [2]), .ZN(n22723) );
  CLKNHSV0 U25000 ( .I(\pe10/bq[13] ), .ZN(n23511) );
  NOR2HSV0 U25001 ( .A1(n22723), .A2(n23511), .ZN(n26106) );
  INHSV2 U25002 ( .I(\pe10/aot [3]), .ZN(n23222) );
  CLKNHSV0 U25003 ( .I(\pe10/bq[14] ), .ZN(n23509) );
  NOR2HSV0 U25004 ( .A1(n23222), .A2(n23509), .ZN(n26164) );
  NAND2HSV0 U25005 ( .A1(n16973), .A2(\pe10/bq[1] ), .ZN(n22526) );
  NAND2HSV0 U25006 ( .A1(\pe10/aot [11]), .A2(\pe10/bq[5] ), .ZN(n22525) );
  XOR2HSV0 U25007 ( .A1(n22526), .A2(n22525), .Z(n22529) );
  NAND2HSV0 U25008 ( .A1(\pe10/bq[2] ), .A2(\pe10/aot [12]), .ZN(n24465) );
  XOR3HSV2 U25009 ( .A1(n22530), .A2(n22529), .A3(n22528), .Z(n22531) );
  XNOR2HSV1 U25010 ( .A1(n22532), .A2(n22531), .ZN(n22533) );
  XOR3HSV2 U25011 ( .A1(n22535), .A2(n22534), .A3(n22533), .Z(n22537) );
  NAND2HSV0 U25012 ( .A1(\pe10/got [3]), .A2(n23474), .ZN(n22536) );
  XNOR2HSV1 U25013 ( .A1(n22537), .A2(n22536), .ZN(n22538) );
  XNOR2HSV1 U25014 ( .A1(n22539), .A2(n22538), .ZN(n22541) );
  NOR2HSV0 U25015 ( .A1(n26200), .A2(n26095), .ZN(n22540) );
  XNOR2HSV1 U25016 ( .A1(n22541), .A2(n22540), .ZN(n22542) );
  XNOR2HSV1 U25017 ( .A1(n22543), .A2(n22542), .ZN(n22544) );
  XNOR2HSV1 U25018 ( .A1(n22545), .A2(n22544), .ZN(n22546) );
  XNOR2HSV1 U25019 ( .A1(n22547), .A2(n22546), .ZN(n22549) );
  NAND2HSV0 U25020 ( .A1(n28585), .A2(\pe10/got [9]), .ZN(n22548) );
  XOR2HSV0 U25021 ( .A1(n22549), .A2(n22548), .Z(n22551) );
  NAND2HSV0 U25022 ( .A1(n26209), .A2(n28644), .ZN(n22550) );
  XNOR2HSV1 U25023 ( .A1(n22551), .A2(n22550), .ZN(n22552) );
  INHSV2 U25024 ( .I(n22598), .ZN(n28469) );
  NAND2HSV0 U25025 ( .A1(n28469), .A2(n26212), .ZN(n22554) );
  XOR2HSV0 U25026 ( .A1(n22555), .A2(n22554), .Z(n22556) );
  CLKNAND2HSV1 U25027 ( .A1(n22560), .A2(n22561), .ZN(n22565) );
  CLKNAND2HSV0 U25028 ( .A1(n22563), .A2(n22562), .ZN(n22564) );
  CLKNAND2HSV1 U25029 ( .A1(n22565), .A2(n22564), .ZN(\pe10/poht [1]) );
  NAND2HSV0 U25030 ( .A1(n27197), .A2(\pe10/got [5]), .ZN(n22588) );
  NAND2HSV0 U25031 ( .A1(\pe10/aot [4]), .A2(\pe10/bq[5] ), .ZN(n22568) );
  NAND2HSV0 U25032 ( .A1(\pe10/aot [3]), .A2(\pe10/bq[6] ), .ZN(n22567) );
  XOR2HSV0 U25033 ( .A1(n22568), .A2(n22567), .Z(n22572) );
  NAND2HSV0 U25034 ( .A1(\pe10/aot [1]), .A2(\pe10/bq[8] ), .ZN(n22570) );
  NAND2HSV0 U25035 ( .A1(\pe10/aot [8]), .A2(\pe10/bq[1] ), .ZN(n22569) );
  XOR2HSV0 U25036 ( .A1(n22570), .A2(n22569), .Z(n22571) );
  XOR2HSV0 U25037 ( .A1(n22572), .A2(n22571), .Z(n22578) );
  NAND2HSV0 U25038 ( .A1(\pe10/aot [7]), .A2(\pe10/bq[2] ), .ZN(n22574) );
  NAND2HSV0 U25039 ( .A1(\pe10/aot [2]), .A2(\pe10/bq[7] ), .ZN(n22573) );
  XOR2HSV0 U25040 ( .A1(n22574), .A2(n22573), .Z(n22576) );
  NAND2HSV0 U25041 ( .A1(\pe10/bq[3] ), .A2(\pe10/aot [5]), .ZN(n22769) );
  NAND2HSV0 U25042 ( .A1(\pe10/bq[4] ), .A2(\pe10/aot [6]), .ZN(n22601) );
  XNOR2HSV1 U25043 ( .A1(n22576), .A2(n22575), .ZN(n22577) );
  XNOR2HSV1 U25044 ( .A1(n22578), .A2(n22577), .ZN(n22579) );
  XNOR2HSV1 U25045 ( .A1(n22580), .A2(n22579), .ZN(n22582) );
  NAND2HSV0 U25046 ( .A1(n28585), .A2(n14065), .ZN(n22581) );
  XOR2HSV0 U25047 ( .A1(n22582), .A2(n22581), .Z(n22584) );
  NAND2HSV0 U25048 ( .A1(n25244), .A2(\pe10/got [3]), .ZN(n22583) );
  XNOR2HSV1 U25049 ( .A1(n22584), .A2(n22583), .ZN(n22585) );
  XOR2HSV0 U25050 ( .A1(n22586), .A2(n22585), .Z(n22587) );
  XOR2HSV0 U25051 ( .A1(n22588), .A2(n22587), .Z(n22591) );
  NOR2HSV2 U25052 ( .A1(n27195), .A2(n26199), .ZN(n22590) );
  INAND2HSV2 U25053 ( .A1(n22680), .B1(\pe10/got [7]), .ZN(n22589) );
  XOR3HSV2 U25054 ( .A1(n22591), .A2(n22590), .A3(n22589), .Z(n22593) );
  NAND2HSV0 U25055 ( .A1(n26221), .A2(n28642), .ZN(n22594) );
  CLKNAND2HSV1 U25056 ( .A1(n22593), .A2(n22592), .ZN(n22597) );
  CLKNHSV1 U25057 ( .I(n22593), .ZN(n22595) );
  CLKNAND2HSV1 U25058 ( .A1(n22595), .A2(n22594), .ZN(n22596) );
  NAND2HSV0 U25059 ( .A1(n26221), .A2(\pe10/got [9]), .ZN(n22631) );
  INAND2HSV2 U25060 ( .A1(n22598), .B1(\pe10/got [6]), .ZN(n22627) );
  INHSV4 U25061 ( .I(n26215), .ZN(n25215) );
  NOR2HSV0 U25062 ( .A1(n25215), .A2(n26095), .ZN(n22623) );
  NAND2HSV0 U25063 ( .A1(n28620), .A2(n14065), .ZN(n22617) );
  NAND2HSV0 U25064 ( .A1(n27196), .A2(n26094), .ZN(n22615) );
  NAND2HSV0 U25065 ( .A1(\pe10/aot [2]), .A2(\pe10/bq[8] ), .ZN(n22600) );
  XOR2HSV0 U25066 ( .A1(n22601), .A2(n22600), .Z(n22613) );
  NAND2HSV0 U25067 ( .A1(\pe10/aot [5]), .A2(\pe10/bq[5] ), .ZN(n22603) );
  NAND2HSV0 U25068 ( .A1(\pe10/aot [3]), .A2(\pe10/bq[7] ), .ZN(n22602) );
  XOR2HSV0 U25069 ( .A1(n22603), .A2(n22602), .Z(n22604) );
  NAND2HSV0 U25070 ( .A1(\pe10/bq[9] ), .A2(\pe10/aot [1]), .ZN(n22724) );
  XNOR2HSV1 U25071 ( .A1(n22604), .A2(n22724), .ZN(n22612) );
  NAND2HSV0 U25072 ( .A1(\pe10/aot [9]), .A2(\pe10/bq[1] ), .ZN(n22606) );
  NAND2HSV0 U25073 ( .A1(\pe10/aot [8]), .A2(\pe10/bq[2] ), .ZN(n22605) );
  XOR2HSV0 U25074 ( .A1(n22606), .A2(n22605), .Z(n22610) );
  NAND2HSV0 U25075 ( .A1(\pe10/aot [4]), .A2(\pe10/bq[6] ), .ZN(n22608) );
  NAND2HSV0 U25076 ( .A1(\pe10/aot [7]), .A2(\pe10/bq[3] ), .ZN(n22607) );
  XOR2HSV0 U25077 ( .A1(n22608), .A2(n22607), .Z(n22609) );
  XOR2HSV0 U25078 ( .A1(n22610), .A2(n22609), .Z(n22611) );
  XOR3HSV2 U25079 ( .A1(n22613), .A2(n22612), .A3(n22611), .Z(n22614) );
  XNOR2HSV1 U25080 ( .A1(n22615), .A2(n22614), .ZN(n22616) );
  XNOR2HSV1 U25081 ( .A1(n22617), .A2(n22616), .ZN(n22619) );
  NAND2HSV0 U25082 ( .A1(n28585), .A2(\pe10/got [3]), .ZN(n22618) );
  XOR2HSV0 U25083 ( .A1(n22619), .A2(n22618), .Z(n22621) );
  CLKNAND2HSV0 U25084 ( .A1(n26209), .A2(n26132), .ZN(n22620) );
  XNOR2HSV1 U25085 ( .A1(n22621), .A2(n22620), .ZN(n22622) );
  XOR2HSV0 U25086 ( .A1(n22623), .A2(n22622), .Z(n22626) );
  CLKNHSV2 U25087 ( .I(\pe10/got [7]), .ZN(n26158) );
  XOR3HSV2 U25088 ( .A1(n22627), .A2(n22626), .A3(n22625), .Z(n22629) );
  NAND2HSV2 U25089 ( .A1(n28642), .A2(n28603), .ZN(n22628) );
  INHSV1 U25090 ( .I(n22633), .ZN(n22630) );
  CLKNAND2HSV1 U25091 ( .A1(n22632), .A2(n22633), .ZN(n22634) );
  NAND2HSV0 U25092 ( .A1(n28479), .A2(n23219), .ZN(n22684) );
  NOR2HSV2 U25093 ( .A1(n24451), .A2(n22636), .ZN(n22679) );
  CLKNAND2HSV0 U25094 ( .A1(n25216), .A2(\pe10/got [6]), .ZN(n22670) );
  NOR2HSV0 U25095 ( .A1(n26096), .A2(n22637), .ZN(n22666) );
  NAND2HSV0 U25096 ( .A1(n28794), .A2(n14065), .ZN(n22662) );
  NAND2HSV0 U25097 ( .A1(n23474), .A2(n27196), .ZN(n22660) );
  NAND2HSV0 U25098 ( .A1(\pe10/aot [6]), .A2(\pe10/bq[8] ), .ZN(n22639) );
  NAND2HSV0 U25099 ( .A1(\pe10/aot [4]), .A2(\pe10/bq[10] ), .ZN(n22638) );
  XOR2HSV0 U25100 ( .A1(n22639), .A2(n22638), .Z(n22658) );
  NAND2HSV0 U25101 ( .A1(\pe10/aot [1]), .A2(\pe10/bq[13] ), .ZN(n22641) );
  NAND2HSV0 U25102 ( .A1(\pe10/aot [11]), .A2(\pe10/bq[3] ), .ZN(n22640) );
  XOR2HSV0 U25103 ( .A1(n22641), .A2(n22640), .Z(n22645) );
  NAND2HSV0 U25104 ( .A1(\pe10/aot [7]), .A2(\pe10/bq[7] ), .ZN(n22643) );
  NAND2HSV0 U25105 ( .A1(\pe10/aot [9]), .A2(\pe10/bq[5] ), .ZN(n22642) );
  XOR2HSV0 U25106 ( .A1(n22643), .A2(n22642), .Z(n22644) );
  XNOR2HSV1 U25107 ( .A1(n22645), .A2(n22644), .ZN(n22657) );
  NAND2HSV0 U25108 ( .A1(\pe10/aot [3]), .A2(\pe10/bq[12] ), .ZN(n26105) );
  NAND2HSV0 U25109 ( .A1(\pe10/aot [2]), .A2(\pe10/bq[11] ), .ZN(n24474) );
  NOR2HSV0 U25110 ( .A1(n26105), .A2(n24474), .ZN(n22647) );
  AOI22HSV0 U25111 ( .A1(\pe10/aot [3]), .A2(\pe10/bq[11] ), .B1(\pe10/bq[12] ), .B2(\pe10/aot [2]), .ZN(n22646) );
  NOR2HSV2 U25112 ( .A1(n22647), .A2(n22646), .ZN(n22648) );
  XOR2HSV0 U25113 ( .A1(n22648), .A2(n24465), .Z(n22656) );
  NAND2HSV0 U25114 ( .A1(\pe10/aot [10]), .A2(\pe10/bq[4] ), .ZN(n22650) );
  NAND2HSV0 U25115 ( .A1(\pe10/aot [13]), .A2(\pe10/bq[1] ), .ZN(n22649) );
  XOR2HSV0 U25116 ( .A1(n22650), .A2(n22649), .Z(n22654) );
  NAND2HSV0 U25117 ( .A1(\pe10/aot [8]), .A2(\pe10/bq[6] ), .ZN(n22652) );
  NAND2HSV0 U25118 ( .A1(\pe10/aot [5]), .A2(\pe10/bq[9] ), .ZN(n22651) );
  XOR2HSV0 U25119 ( .A1(n22652), .A2(n22651), .Z(n22653) );
  XOR2HSV0 U25120 ( .A1(n22654), .A2(n22653), .Z(n22655) );
  XOR4HSV1 U25121 ( .A1(n22658), .A2(n22657), .A3(n22656), .A4(n22655), .Z(
        n22659) );
  XNOR2HSV1 U25122 ( .A1(n22660), .A2(n22659), .ZN(n22661) );
  XNOR2HSV1 U25123 ( .A1(n22662), .A2(n22661), .ZN(n22664) );
  NAND2HSV0 U25124 ( .A1(n26131), .A2(\pe10/got [3]), .ZN(n22663) );
  XNOR2HSV1 U25125 ( .A1(n22664), .A2(n22663), .ZN(n22665) );
  XNOR2HSV1 U25126 ( .A1(n22666), .A2(n22665), .ZN(n22667) );
  XNOR2HSV1 U25127 ( .A1(n22668), .A2(n22667), .ZN(n22669) );
  XNOR2HSV1 U25128 ( .A1(n22670), .A2(n22669), .ZN(n22672) );
  NAND2HSV0 U25129 ( .A1(n28585), .A2(\pe10/got [7]), .ZN(n22671) );
  XOR2HSV0 U25130 ( .A1(n22672), .A2(n22671), .Z(n22674) );
  NAND2HSV0 U25131 ( .A1(n25244), .A2(n28642), .ZN(n22673) );
  XNOR2HSV1 U25132 ( .A1(n22674), .A2(n22673), .ZN(n22678) );
  NOR2HSV2 U25133 ( .A1(n25215), .A2(n25214), .ZN(n22677) );
  NAND2HSV2 U25134 ( .A1(n28469), .A2(n28644), .ZN(n22676) );
  XNOR2HSV1 U25135 ( .A1(n22679), .A2(n13974), .ZN(n22682) );
  NAND2HSV2 U25136 ( .A1(n28603), .A2(\pe10/got [12]), .ZN(n22681) );
  XNOR2HSV4 U25137 ( .A1(n22682), .A2(n22681), .ZN(n22685) );
  INHSV2 U25138 ( .I(n22685), .ZN(n22683) );
  CLKNAND2HSV1 U25139 ( .A1(n22684), .A2(n22683), .ZN(n22688) );
  CLKNHSV0 U25140 ( .I(n22684), .ZN(n22686) );
  CLKNAND2HSV1 U25141 ( .A1(n22686), .A2(n22685), .ZN(n22687) );
  CLKNAND2HSV1 U25142 ( .A1(n22688), .A2(n22687), .ZN(\pe10/poht [3]) );
  INHSV2 U25143 ( .I(\pe10/got [3]), .ZN(n24453) );
  CLKNAND2HSV0 U25144 ( .A1(\pe10/aot [1]), .A2(\pe10/bq[5] ), .ZN(n22693) );
  XNOR2HSV0 U25145 ( .A1(n28637), .A2(n22693), .ZN(n22701) );
  NAND3HSV0 U25146 ( .A1(n22696), .A2(n22691), .A3(n22693), .ZN(n22700) );
  CLKNHSV0 U25147 ( .I(n22693), .ZN(n22698) );
  NOR2HSV0 U25148 ( .A1(n22694), .A2(n22693), .ZN(n22695) );
  NAND3HSV0 U25149 ( .A1(n22696), .A2(n22695), .A3(n22692), .ZN(n22697) );
  AOI21HSV2 U25150 ( .A1(n22701), .A2(n22700), .B(n22699), .ZN(n22711) );
  NOR2HSV2 U25151 ( .A1(n25215), .A2(n26186), .ZN(n22709) );
  NAND2HSV0 U25152 ( .A1(\pe10/aot [2]), .A2(\pe10/bq[4] ), .ZN(n22702) );
  XOR2HSV0 U25153 ( .A1(n22703), .A2(n22702), .Z(n22707) );
  CLKNAND2HSV0 U25154 ( .A1(\pe10/aot [4]), .A2(\pe10/bq[1] ), .ZN(n27198) );
  AO22HSV2 U25155 ( .A1(\pe10/aot [5]), .A2(\pe10/bq[1] ), .B1(\pe10/aot [4]), 
        .B2(\pe10/bq[2] ), .Z(n22704) );
  OAI21HSV1 U25156 ( .A1(n27198), .A2(n22705), .B(n22704), .ZN(n22706) );
  XNOR2HSV1 U25157 ( .A1(n22707), .A2(n22706), .ZN(n22708) );
  NAND2HSV0 U25158 ( .A1(n23219), .A2(\pe10/got [5]), .ZN(n22715) );
  CLKNHSV0 U25159 ( .I(n22715), .ZN(n22712) );
  CLKNAND2HSV1 U25160 ( .A1(n22713), .A2(n22712), .ZN(n22717) );
  CLKNAND2HSV1 U25161 ( .A1(n22715), .A2(n22714), .ZN(n22716) );
  CLKNAND2HSV1 U25162 ( .A1(n22717), .A2(n22716), .ZN(\pe10/poht [11]) );
  INOR2HSV1 U25163 ( .A1(n22718), .B1(n24452), .ZN(n22755) );
  NOR2HSV2 U25164 ( .A1(n25215), .A2(n26199), .ZN(n22751) );
  NAND2HSV0 U25165 ( .A1(n25216), .A2(\pe10/got [3]), .ZN(n22745) );
  NOR2HSV0 U25166 ( .A1(n26159), .A2(n26186), .ZN(n22741) );
  INHSV2 U25167 ( .I(\pe10/bq[1] ), .ZN(n26163) );
  NOR2HSV0 U25168 ( .A1(n22719), .A2(n26163), .ZN(n22721) );
  NAND2HSV0 U25169 ( .A1(\pe10/aot [4]), .A2(\pe10/bq[7] ), .ZN(n22720) );
  XOR2HSV0 U25170 ( .A1(n22721), .A2(n22720), .Z(n22739) );
  NOR2HSV0 U25171 ( .A1(n22723), .A2(n22722), .ZN(n25221) );
  CLKNHSV0 U25172 ( .I(n22724), .ZN(n22726) );
  AOI22HSV0 U25173 ( .A1(\pe10/aot [2]), .A2(\pe10/bq[9] ), .B1(\pe10/bq[10] ), 
        .B2(\pe10/aot [1]), .ZN(n22725) );
  AOI21HSV2 U25174 ( .A1(n25221), .A2(n22726), .B(n22725), .ZN(n22730) );
  CLKNHSV0 U25175 ( .I(n26161), .ZN(n22728) );
  CLKNHSV0 U25176 ( .I(\pe10/bq[2] ), .ZN(n24462) );
  NOR2HSV2 U25177 ( .A1(n23222), .A2(n24462), .ZN(n27199) );
  AOI22HSV0 U25178 ( .A1(\pe10/aot [9]), .A2(\pe10/bq[2] ), .B1(\pe10/bq[8] ), 
        .B2(\pe10/aot [3]), .ZN(n22727) );
  AOI21HSV0 U25179 ( .A1(n22728), .A2(n27199), .B(n22727), .ZN(n22729) );
  XNOR2HSV1 U25180 ( .A1(n22730), .A2(n22729), .ZN(n22738) );
  NAND2HSV0 U25181 ( .A1(\pe10/aot [8]), .A2(\pe10/bq[3] ), .ZN(n22732) );
  NAND2HSV0 U25182 ( .A1(\pe10/aot [7]), .A2(\pe10/bq[4] ), .ZN(n22731) );
  XOR2HSV0 U25183 ( .A1(n22732), .A2(n22731), .Z(n22736) );
  NAND2HSV0 U25184 ( .A1(\pe10/aot [6]), .A2(\pe10/bq[5] ), .ZN(n22734) );
  NAND2HSV0 U25185 ( .A1(\pe10/aot [5]), .A2(\pe10/bq[6] ), .ZN(n22733) );
  XOR2HSV0 U25186 ( .A1(n22734), .A2(n22733), .Z(n22735) );
  XOR2HSV0 U25187 ( .A1(n22736), .A2(n22735), .Z(n22737) );
  XOR3HSV2 U25188 ( .A1(n22739), .A2(n22738), .A3(n22737), .Z(n22740) );
  XOR2HSV0 U25189 ( .A1(n22741), .A2(n22740), .Z(n22742) );
  XNOR2HSV1 U25190 ( .A1(n22743), .A2(n22742), .ZN(n22744) );
  XNOR2HSV1 U25191 ( .A1(n22745), .A2(n22744), .ZN(n22747) );
  NAND2HSV0 U25192 ( .A1(n28585), .A2(\pe10/got [4]), .ZN(n22746) );
  XOR2HSV0 U25193 ( .A1(n22747), .A2(n22746), .Z(n22749) );
  NAND2HSV0 U25194 ( .A1(n26209), .A2(\pe10/got [5]), .ZN(n22748) );
  XNOR2HSV1 U25195 ( .A1(n22749), .A2(n22748), .ZN(n22750) );
  XOR2HSV0 U25196 ( .A1(n22751), .A2(n22750), .Z(n22753) );
  NAND2HSV0 U25197 ( .A1(n27197), .A2(\pe10/got [7]), .ZN(n22752) );
  XOR2HSV0 U25198 ( .A1(n22753), .A2(n22752), .Z(n22754) );
  CLKNHSV0 U25199 ( .I(n22760), .ZN(n22759) );
  NAND2HSV0 U25200 ( .A1(n26221), .A2(n28644), .ZN(n22761) );
  CLKNHSV0 U25201 ( .I(n22761), .ZN(n22758) );
  CLKNAND2HSV1 U25202 ( .A1(n22759), .A2(n22758), .ZN(n22763) );
  CLKNAND2HSV0 U25203 ( .A1(n22761), .A2(n22760), .ZN(n22762) );
  CLKNAND2HSV1 U25204 ( .A1(n22763), .A2(n22762), .ZN(\pe10/poht [6]) );
  NAND2HSV0 U25205 ( .A1(n23219), .A2(\pe10/got [7]), .ZN(n22788) );
  CLKNHSV0 U25206 ( .I(n22788), .ZN(n22786) );
  NOR2HSV2 U25207 ( .A1(n12304), .A2(n26095), .ZN(n22782) );
  NOR2HSV2 U25208 ( .A1(n26093), .A2(n24453), .ZN(n22778) );
  NAND2HSV0 U25209 ( .A1(n28585), .A2(n27196), .ZN(n22774) );
  NAND2HSV0 U25210 ( .A1(\pe10/bq[2] ), .A2(\pe10/aot [6]), .ZN(n26097) );
  CLKNHSV0 U25211 ( .I(\pe10/aot [7]), .ZN(n26102) );
  NAND2HSV0 U25212 ( .A1(\pe10/aot [2]), .A2(\pe10/bq[6] ), .ZN(n22768) );
  NAND2HSV0 U25213 ( .A1(\pe10/aot [1]), .A2(\pe10/bq[7] ), .ZN(n22767) );
  XOR2HSV0 U25214 ( .A1(n22768), .A2(n22767), .Z(n22770) );
  XNOR2HSV1 U25215 ( .A1(n22770), .A2(n22769), .ZN(n22771) );
  XNOR2HSV1 U25216 ( .A1(n22772), .A2(n22771), .ZN(n22773) );
  XNOR2HSV1 U25217 ( .A1(n22774), .A2(n22773), .ZN(n22776) );
  NAND2HSV0 U25218 ( .A1(n26209), .A2(n14065), .ZN(n22775) );
  XOR2HSV0 U25219 ( .A1(n22776), .A2(n22775), .Z(n22777) );
  XOR2HSV0 U25220 ( .A1(n22778), .A2(n22777), .Z(n22780) );
  NAND2HSV0 U25221 ( .A1(n27197), .A2(\pe10/got [4]), .ZN(n22779) );
  XOR2HSV0 U25222 ( .A1(n22780), .A2(n22779), .Z(n22781) );
  NAND2HSV2 U25223 ( .A1(n25060), .A2(\pe10/got [6]), .ZN(n22783) );
  CLKNAND2HSV1 U25224 ( .A1(n22786), .A2(n22785), .ZN(n22790) );
  CLKNAND2HSV0 U25225 ( .A1(n22788), .A2(n22787), .ZN(n22789) );
  CLKNAND2HSV1 U25226 ( .A1(n22790), .A2(n22789), .ZN(\pe10/poht [9]) );
  CLKNAND2HSV2 U25227 ( .A1(n26929), .A2(n22792), .ZN(n22795) );
  INAND2HSV2 U25228 ( .A1(n26923), .B1(n22792), .ZN(n22793) );
  AND2HSV2 U25229 ( .A1(n22915), .A2(n22918), .Z(n22797) );
  NAND2HSV4 U25230 ( .A1(n22799), .A2(n22798), .ZN(n27904) );
  NOR2HSV2 U25231 ( .A1(n27999), .A2(n21997), .ZN(n22926) );
  CLKNAND2HSV0 U25232 ( .A1(n28480), .A2(\pe4/got [4]), .ZN(n22819) );
  MUX2NHSV4 U25233 ( .I0(\pe4/ti_7t [12]), .I1(n29028), .S(n26923), .ZN(n27941) );
  INHSV2 U25234 ( .I(n25079), .ZN(n27979) );
  INHSV2 U25235 ( .I(\pe4/got [3]), .ZN(n27998) );
  NOR2HSV2 U25236 ( .A1(n27979), .A2(n27998), .ZN(n22817) );
  INHSV2 U25237 ( .I(\pe4/got [2]), .ZN(n22848) );
  NAND2HSV0 U25238 ( .A1(n28591), .A2(n14038), .ZN(n22815) );
  INHSV2 U25239 ( .I(\pe4/got [1]), .ZN(n28000) );
  NOR2HSV0 U25240 ( .A1(n27876), .A2(n28000), .ZN(n22813) );
  NAND2HSV0 U25241 ( .A1(\pe4/aot [1]), .A2(\pe4/bq[6] ), .ZN(n22804) );
  NAND2HSV0 U25242 ( .A1(\pe4/aot [3]), .A2(\pe4/bq[4] ), .ZN(n22803) );
  XOR2HSV0 U25243 ( .A1(n22804), .A2(n22803), .Z(n22808) );
  NAND2HSV0 U25244 ( .A1(\pe4/aot [6]), .A2(\pe4/bq[2] ), .ZN(n27886) );
  NAND2HSV0 U25245 ( .A1(\pe4/bq[1] ), .A2(\pe4/aot [5]), .ZN(n27983) );
  NOR2HSV0 U25246 ( .A1(n27886), .A2(n27983), .ZN(n22806) );
  AOI22HSV0 U25247 ( .A1(\pe4/aot [6]), .A2(\pe4/bq[1] ), .B1(\pe4/aot [5]), 
        .B2(\pe4/bq[2] ), .ZN(n22805) );
  NOR2HSV2 U25248 ( .A1(n22806), .A2(n22805), .ZN(n22807) );
  XNOR2HSV1 U25249 ( .A1(n22808), .A2(n22807), .ZN(n22811) );
  NAND2HSV0 U25250 ( .A1(\pe4/aot [2]), .A2(\pe4/bq[5] ), .ZN(n27795) );
  NAND2HSV0 U25251 ( .A1(\pe4/aot [4]), .A2(\pe4/bq[3] ), .ZN(n22809) );
  XOR2HSV0 U25252 ( .A1(n27795), .A2(n22809), .Z(n22810) );
  XNOR2HSV1 U25253 ( .A1(n22811), .A2(n22810), .ZN(n22812) );
  XOR2HSV0 U25254 ( .A1(n22813), .A2(n22812), .Z(n22814) );
  XOR2HSV0 U25255 ( .A1(n22815), .A2(n22814), .Z(n22816) );
  XOR2HSV0 U25256 ( .A1(n22817), .A2(n22816), .Z(n22818) );
  XOR2HSV2 U25257 ( .A1(n22819), .A2(n22818), .Z(n22925) );
  INAND2HSV2 U25258 ( .A1(n22820), .B1(n28592), .ZN(n22821) );
  CLKNAND2HSV1 U25259 ( .A1(n27907), .A2(n25131), .ZN(n22879) );
  INHSV2 U25260 ( .I(n25128), .ZN(n27780) );
  NOR2HSV2 U25261 ( .A1(n27876), .A2(n27780), .ZN(n22877) );
  CLKNAND2HSV2 U25262 ( .A1(n27957), .A2(\pe4/got [10]), .ZN(n22823) );
  XNOR2HSV4 U25263 ( .A1(n22824), .A2(n22823), .ZN(n22875) );
  NAND2HSV0 U25264 ( .A1(\pe4/ti_7[7] ), .A2(\pe4/got [9]), .ZN(n22874) );
  NAND2HSV0 U25265 ( .A1(n22825), .A2(\pe4/got [8]), .ZN(n22872) );
  CLKNAND2HSV0 U25266 ( .A1(n22827), .A2(n22826), .ZN(n22866) );
  NAND2HSV0 U25267 ( .A1(n28671), .A2(\pe4/got [4]), .ZN(n22845) );
  NAND2HSV0 U25268 ( .A1(\pe4/aot [11]), .A2(\pe4/bq[7] ), .ZN(n27748) );
  NAND2HSV0 U25269 ( .A1(\pe4/aot [4]), .A2(n27060), .ZN(n22952) );
  XOR2HSV0 U25270 ( .A1(n27748), .A2(n22952), .Z(n22843) );
  INHSV2 U25271 ( .I(n21332), .ZN(n27066) );
  NAND2HSV0 U25272 ( .A1(n27066), .A2(\pe4/pvq [15]), .ZN(n22828) );
  XNOR2HSV1 U25273 ( .A1(n22828), .A2(\pe4/phq [15]), .ZN(n22833) );
  NAND2HSV0 U25274 ( .A1(\pe4/aot [13]), .A2(\pe4/bq[2] ), .ZN(n25103) );
  NOR2HSV0 U25275 ( .A1(n22829), .A2(n25103), .ZN(n22831) );
  AOI22HSV0 U25276 ( .A1(n28683), .A2(\pe4/bq[2] ), .B1(\pe4/aot [13]), .B2(
        \pe4/bq[5] ), .ZN(n22830) );
  NOR2HSV2 U25277 ( .A1(n22831), .A2(n22830), .ZN(n22832) );
  XNOR2HSV1 U25278 ( .A1(n22833), .A2(n22832), .ZN(n22842) );
  NAND2HSV0 U25279 ( .A1(\pe4/aot [2]), .A2(n22834), .ZN(n22836) );
  NAND2HSV0 U25280 ( .A1(\pe4/aot [12]), .A2(\pe4/bq[6] ), .ZN(n22835) );
  XOR2HSV0 U25281 ( .A1(n22836), .A2(n22835), .Z(n22840) );
  NAND2HSV0 U25282 ( .A1(\pe4/aot [9]), .A2(\pe4/bq[9] ), .ZN(n22837) );
  XOR2HSV0 U25283 ( .A1(n22838), .A2(n22837), .Z(n22839) );
  XOR2HSV0 U25284 ( .A1(n22840), .A2(n22839), .Z(n22841) );
  XOR3HSV2 U25285 ( .A1(n22843), .A2(n22842), .A3(n22841), .Z(n22844) );
  XOR2HSV0 U25286 ( .A1(n22845), .A2(n22844), .Z(n22864) );
  NAND2HSV0 U25287 ( .A1(\pe4/aot [7]), .A2(\pe4/bq[11] ), .ZN(n22847) );
  NAND2HSV0 U25288 ( .A1(\pe4/aot [5]), .A2(n23076), .ZN(n22846) );
  XOR2HSV0 U25289 ( .A1(n22847), .A2(n22846), .Z(n22852) );
  NAND2HSV0 U25290 ( .A1(\pe4/got [2]), .A2(n27128), .ZN(n22850) );
  NAND2HSV0 U25291 ( .A1(n28433), .A2(\pe4/bq[3] ), .ZN(n22849) );
  XOR2HSV0 U25292 ( .A1(n22850), .A2(n22849), .Z(n22851) );
  XOR2HSV0 U25293 ( .A1(n22852), .A2(n22851), .Z(n22860) );
  NAND2HSV0 U25294 ( .A1(n22943), .A2(\pe4/aot [3]), .ZN(n22854) );
  NAND2HSV0 U25295 ( .A1(\pe4/bq[4] ), .A2(\pe4/aot [14]), .ZN(n22853) );
  XOR2HSV0 U25296 ( .A1(n22854), .A2(n22853), .Z(n22858) );
  NAND2HSV0 U25297 ( .A1(\pe4/aot [8]), .A2(\pe4/bq[10] ), .ZN(n22856) );
  NAND2HSV0 U25298 ( .A1(\pe4/aot [6]), .A2(\pe4/bq[12] ), .ZN(n22855) );
  XOR2HSV0 U25299 ( .A1(n22856), .A2(n22855), .Z(n22857) );
  XOR2HSV0 U25300 ( .A1(n22858), .A2(n22857), .Z(n22859) );
  XOR2HSV0 U25301 ( .A1(n22860), .A2(n22859), .Z(n22862) );
  NAND2HSV0 U25302 ( .A1(n23482), .A2(\pe4/got [3]), .ZN(n22861) );
  XNOR2HSV1 U25303 ( .A1(n22862), .A2(n22861), .ZN(n22863) );
  XNOR2HSV1 U25304 ( .A1(n22864), .A2(n22863), .ZN(n22865) );
  XNOR2HSV1 U25305 ( .A1(n22866), .A2(n22865), .ZN(n22868) );
  NAND2HSV0 U25306 ( .A1(n28951), .A2(\pe4/got [5]), .ZN(n22867) );
  XNOR2HSV1 U25307 ( .A1(n22868), .A2(n22867), .ZN(n22870) );
  NAND2HSV0 U25308 ( .A1(n27830), .A2(n13996), .ZN(n22869) );
  XOR2HSV0 U25309 ( .A1(n22870), .A2(n22869), .Z(n22871) );
  XNOR2HSV1 U25310 ( .A1(n22872), .A2(n22871), .ZN(n22873) );
  XNOR2HSV4 U25311 ( .A1(n22875), .A2(n13966), .ZN(n22876) );
  NOR2HSV0 U25312 ( .A1(n22881), .A2(n22880), .ZN(n22882) );
  AND3HSV1 U25313 ( .A1(n22884), .A2(n22883), .A3(n22882), .Z(n22885) );
  NAND3HSV2 U25314 ( .A1(n22887), .A2(n22886), .A3(n22885), .ZN(n22888) );
  INHSV3 U25315 ( .I(n22889), .ZN(n22892) );
  INHSV2 U25316 ( .I(n22890), .ZN(n22891) );
  NAND2HSV4 U25317 ( .A1(n22892), .A2(n22891), .ZN(n22893) );
  CLKNAND2HSV4 U25318 ( .A1(n22893), .A2(n22894), .ZN(n25372) );
  AND2HSV2 U25319 ( .A1(n27976), .A2(\pe4/ti_7t [15]), .Z(n22913) );
  NOR2HSV1 U25320 ( .A1(n15484), .A2(\pe4/ti_7t [14]), .ZN(n27974) );
  NOR2HSV0 U25321 ( .A1(n27974), .A2(n22895), .ZN(n25369) );
  CLKNHSV0 U25322 ( .I(n22913), .ZN(n22896) );
  CLKNAND2HSV1 U25323 ( .A1(n25369), .A2(n22896), .ZN(n22902) );
  CLKNHSV2 U25324 ( .I(n22903), .ZN(n22897) );
  NAND2HSV2 U25325 ( .A1(n26916), .A2(n22897), .ZN(n22898) );
  NAND2HSV2 U25326 ( .A1(n22899), .A2(n22898), .ZN(n22916) );
  NOR2HSV2 U25327 ( .A1(n26930), .A2(n22900), .ZN(n22901) );
  AOI22HSV2 U25328 ( .A1(n22902), .A2(n13991), .B1(n22916), .B2(n22901), .ZN(
        n22911) );
  INHSV2 U25329 ( .I(n22903), .ZN(n22910) );
  CLKNHSV2 U25330 ( .I(n22904), .ZN(n22906) );
  CLKNAND2HSV2 U25331 ( .A1(n22906), .A2(n22905), .ZN(n22907) );
  AOI21HSV4 U25332 ( .A1(n26916), .A2(n22910), .B(n22907), .ZN(n22908) );
  OAI21HSV4 U25333 ( .A1(n22910), .A2(n22909), .B(n22908), .ZN(n25371) );
  OAI21HSV4 U25334 ( .A1(n25372), .A2(n22913), .B(n22912), .ZN(n25074) );
  NAND2HSV0 U25335 ( .A1(n22915), .A2(n22914), .ZN(n22917) );
  AND2HSV2 U25336 ( .A1(n25369), .A2(n22918), .Z(n22919) );
  INHSV3 U25337 ( .I(n25371), .ZN(n22920) );
  INHSV4 U25338 ( .I(n25372), .ZN(n22922) );
  CLKNAND2HSV4 U25339 ( .A1(n22923), .A2(n22922), .ZN(n25075) );
  NAND2HSV4 U25340 ( .A1(n25074), .A2(n25075), .ZN(n23681) );
  INHSV6 U25341 ( .I(n23681), .ZN(n27900) );
  NOR2HSV0 U25342 ( .A1(n27900), .A2(n27905), .ZN(n22924) );
  XOR3HSV1 U25343 ( .A1(n22926), .A2(n22925), .A3(n22924), .Z(\pe4/poht [10])
         );
  AND2HSV2 U25344 ( .A1(n27904), .A2(n25134), .Z(n22990) );
  NOR2HSV2 U25345 ( .A1(n27977), .A2(n26932), .ZN(n22986) );
  NOR2HSV2 U25346 ( .A1(n28001), .A2(n27780), .ZN(n22984) );
  NAND2HSV0 U25347 ( .A1(n13994), .A2(n28523), .ZN(n22982) );
  NOR2HSV0 U25348 ( .A1(n27942), .A2(n27825), .ZN(n22980) );
  NAND2HSV0 U25349 ( .A1(\pe4/got [9]), .A2(n27877), .ZN(n22930) );
  NAND2HSV0 U25350 ( .A1(n27957), .A2(\pe4/got [8]), .ZN(n22929) );
  XNOR2HSV1 U25351 ( .A1(n22930), .A2(n22929), .ZN(n22978) );
  NAND2HSV0 U25352 ( .A1(\pe4/ti_7[7] ), .A2(n13996), .ZN(n22976) );
  NAND2HSV0 U25353 ( .A1(n22825), .A2(n22826), .ZN(n22974) );
  NAND2HSV0 U25354 ( .A1(n28671), .A2(n28591), .ZN(n22934) );
  NOR2HSV0 U25355 ( .A1(n22932), .A2(n28000), .ZN(n22933) );
  XNOR2HSV1 U25356 ( .A1(n22934), .A2(n22933), .ZN(n22967) );
  NAND2HSV0 U25357 ( .A1(\pe4/aot [3]), .A2(n23076), .ZN(n22936) );
  NAND2HSV0 U25358 ( .A1(\pe4/aot [8]), .A2(\pe4/bq[8] ), .ZN(n22935) );
  XOR2HSV0 U25359 ( .A1(n22936), .A2(n22935), .Z(n22940) );
  NAND2HSV0 U25360 ( .A1(\pe4/aot [9]), .A2(\pe4/bq[7] ), .ZN(n22938) );
  NAND2HSV0 U25361 ( .A1(\pe4/aot [12]), .A2(\pe4/bq[4] ), .ZN(n22937) );
  XOR2HSV0 U25362 ( .A1(n22938), .A2(n22937), .Z(n22939) );
  XOR2HSV0 U25363 ( .A1(n22940), .A2(n22939), .Z(n22949) );
  NAND2HSV0 U25364 ( .A1(n28433), .A2(\pe4/bq[1] ), .ZN(n22942) );
  NAND2HSV0 U25365 ( .A1(\pe4/aot [5]), .A2(\pe4/bq[11] ), .ZN(n22941) );
  XOR2HSV0 U25366 ( .A1(n22942), .A2(n22941), .Z(n22947) );
  NAND2HSV0 U25367 ( .A1(\pe4/aot [10]), .A2(\pe4/bq[6] ), .ZN(n22945) );
  NAND2HSV0 U25368 ( .A1(n22943), .A2(\pe4/aot [1]), .ZN(n22944) );
  XOR2HSV0 U25369 ( .A1(n22945), .A2(n22944), .Z(n22946) );
  XNOR2HSV1 U25370 ( .A1(n22947), .A2(n22946), .ZN(n22948) );
  XNOR2HSV1 U25371 ( .A1(n22949), .A2(n22948), .ZN(n22965) );
  NAND2HSV0 U25372 ( .A1(\pe4/aot [11]), .A2(\pe4/bq[5] ), .ZN(n22951) );
  NAND2HSV0 U25373 ( .A1(\pe4/aot [7]), .A2(\pe4/bq[9] ), .ZN(n22950) );
  XOR2HSV0 U25374 ( .A1(n22951), .A2(n22950), .Z(n22956) );
  NAND2HSV0 U25375 ( .A1(\pe4/bq[12] ), .A2(\pe4/aot [2]), .ZN(n23072) );
  NOR2HSV0 U25376 ( .A1(n22952), .A2(n23072), .ZN(n22954) );
  AOI22HSV0 U25377 ( .A1(\pe4/aot [4]), .A2(\pe4/bq[12] ), .B1(n27060), .B2(
        \pe4/aot [2]), .ZN(n22953) );
  NOR2HSV2 U25378 ( .A1(n22954), .A2(n22953), .ZN(n22955) );
  XNOR2HSV1 U25379 ( .A1(n22956), .A2(n22955), .ZN(n22963) );
  NOR2HSV0 U25380 ( .A1(n22957), .A2(n27886), .ZN(n22959) );
  AOI22HSV0 U25381 ( .A1(\pe4/bq[2] ), .A2(\pe4/aot [14]), .B1(\pe4/bq[10] ), 
        .B2(\pe4/aot [6]), .ZN(n22958) );
  NOR2HSV2 U25382 ( .A1(n22959), .A2(n22958), .ZN(n22961) );
  XOR2HSV0 U25383 ( .A1(n22961), .A2(n22960), .Z(n22962) );
  XNOR2HSV1 U25384 ( .A1(n22963), .A2(n22962), .ZN(n22964) );
  XNOR2HSV1 U25385 ( .A1(n22965), .A2(n22964), .ZN(n22966) );
  XNOR2HSV1 U25386 ( .A1(n22967), .A2(n22966), .ZN(n22970) );
  NOR2HSV0 U25387 ( .A1(n26981), .A2(n27998), .ZN(n22969) );
  NAND2HSV0 U25388 ( .A1(n27739), .A2(\pe4/got [4]), .ZN(n22968) );
  XOR3HSV2 U25389 ( .A1(n22970), .A2(n22969), .A3(n22968), .Z(n22972) );
  NAND2HSV0 U25390 ( .A1(\pe4/got [5]), .A2(n27830), .ZN(n22971) );
  XOR2HSV0 U25391 ( .A1(n22972), .A2(n22971), .Z(n22973) );
  XNOR2HSV1 U25392 ( .A1(n22974), .A2(n22973), .ZN(n22975) );
  XNOR2HSV1 U25393 ( .A1(n22976), .A2(n22975), .ZN(n22977) );
  XNOR2HSV1 U25394 ( .A1(n22978), .A2(n22977), .ZN(n22979) );
  XOR2HSV0 U25395 ( .A1(n22980), .A2(n22979), .Z(n22981) );
  XNOR2HSV1 U25396 ( .A1(n22982), .A2(n22981), .ZN(n22983) );
  XNOR2HSV1 U25397 ( .A1(n22986), .A2(n22985), .ZN(n22989) );
  NOR2HSV0 U25398 ( .A1(n27900), .A2(n22987), .ZN(n22988) );
  XOR3HSV1 U25399 ( .A1(n22990), .A2(n22989), .A3(n22988), .Z(\pe4/poht [1])
         );
  INHSV2 U25400 ( .I(n28925), .ZN(n22991) );
  INHSV4 U25401 ( .I(n22991), .ZN(n25980) );
  CLKNAND2HSV1 U25402 ( .A1(n26084), .A2(n22992), .ZN(n23055) );
  NAND2HSV0 U25403 ( .A1(n22078), .A2(n28593), .ZN(n23051) );
  NOR2HSV2 U25404 ( .A1(n25818), .A2(n22994), .ZN(n23049) );
  CLKNAND2HSV0 U25405 ( .A1(n25952), .A2(\pe6/got [10]), .ZN(n23047) );
  NAND2HSV0 U25406 ( .A1(\pe6/ti_7[7] ), .A2(\pe6/got [7]), .ZN(n23040) );
  NAND2HSV0 U25407 ( .A1(n25982), .A2(n26033), .ZN(n23038) );
  INAND2HSV0 U25408 ( .A1(n14029), .B1(n26065), .ZN(n23036) );
  CLKNHSV0 U25409 ( .I(n22996), .ZN(n25849) );
  NAND2HSV0 U25410 ( .A1(n25849), .A2(\pe6/got [3]), .ZN(n23034) );
  NAND2HSV0 U25411 ( .A1(n25846), .A2(\pe6/got [2]), .ZN(n22998) );
  NAND2HSV0 U25412 ( .A1(\pe6/ti_7[1] ), .A2(n28608), .ZN(n22997) );
  XNOR2HSV1 U25413 ( .A1(n22998), .A2(n22997), .ZN(n23031) );
  NAND2HSV0 U25414 ( .A1(\pe6/aot [1]), .A2(\pe6/bq[15] ), .ZN(n23000) );
  NAND2HSV0 U25415 ( .A1(\pe6/aot [7]), .A2(\pe6/bq[9] ), .ZN(n22999) );
  XOR2HSV0 U25416 ( .A1(n23000), .A2(n22999), .Z(n23004) );
  NAND2HSV0 U25417 ( .A1(n28680), .A2(\pe6/bq[1] ), .ZN(n23002) );
  NAND2HSV0 U25418 ( .A1(\pe6/bq[2] ), .A2(\pe6/aot [14]), .ZN(n23001) );
  XOR2HSV0 U25419 ( .A1(n23002), .A2(n23001), .Z(n23003) );
  XOR2HSV0 U25420 ( .A1(n23004), .A2(n23003), .Z(n23012) );
  NAND2HSV0 U25421 ( .A1(\pe6/aot [3]), .A2(\pe6/bq[13] ), .ZN(n23006) );
  NAND2HSV0 U25422 ( .A1(\pe6/aot [9]), .A2(\pe6/bq[7] ), .ZN(n23005) );
  XOR2HSV0 U25423 ( .A1(n23006), .A2(n23005), .Z(n23010) );
  NAND2HSV0 U25424 ( .A1(\pe6/aot [6]), .A2(\pe6/bq[10] ), .ZN(n23008) );
  NAND2HSV0 U25425 ( .A1(\pe6/bq[4] ), .A2(\pe6/aot [12]), .ZN(n23007) );
  XOR2HSV0 U25426 ( .A1(n23008), .A2(n23007), .Z(n23009) );
  XOR2HSV0 U25427 ( .A1(n23010), .A2(n23009), .Z(n23011) );
  XOR2HSV0 U25428 ( .A1(n23012), .A2(n23011), .Z(n23029) );
  NAND2HSV0 U25429 ( .A1(\pe6/bq[6] ), .A2(\pe6/aot [10]), .ZN(n23014) );
  NAND2HSV0 U25430 ( .A1(\pe6/aot [4]), .A2(n25701), .ZN(n23013) );
  XOR2HSV0 U25431 ( .A1(n23014), .A2(n23013), .Z(n23020) );
  NAND2HSV0 U25432 ( .A1(\pe6/bq[8] ), .A2(\pe6/aot [5]), .ZN(n26053) );
  CLKNHSV0 U25433 ( .I(\pe6/aot [5]), .ZN(n23017) );
  CLKNHSV0 U25434 ( .I(\pe6/bq[11] ), .ZN(n23016) );
  OAI21HSV0 U25435 ( .A1(n23017), .A2(n23016), .B(n23015), .ZN(n23018) );
  OAI21HSV0 U25436 ( .A1(n26044), .A2(n26053), .B(n23018), .ZN(n23019) );
  XNOR2HSV1 U25437 ( .A1(n23020), .A2(n23019), .ZN(n23027) );
  NOR2HSV0 U25438 ( .A1(n23021), .A2(n26043), .ZN(n23024) );
  CLKNHSV0 U25439 ( .I(\pe6/bq[14] ), .ZN(n23022) );
  INHSV2 U25440 ( .I(n23022), .ZN(n23485) );
  AOI22HSV0 U25441 ( .A1(\pe6/aot [11]), .A2(\pe6/bq[5] ), .B1(n23485), .B2(
        \pe6/aot [2]), .ZN(n23023) );
  NOR2HSV2 U25442 ( .A1(n23024), .A2(n23023), .ZN(n23025) );
  NAND2HSV0 U25443 ( .A1(\pe6/bq[3] ), .A2(\pe6/aot [13]), .ZN(n25426) );
  XOR2HSV0 U25444 ( .A1(n23025), .A2(n25426), .Z(n23026) );
  XNOR2HSV1 U25445 ( .A1(n23027), .A2(n23026), .ZN(n23028) );
  XNOR2HSV1 U25446 ( .A1(n23029), .A2(n23028), .ZN(n23030) );
  XNOR2HSV1 U25447 ( .A1(n23031), .A2(n23030), .ZN(n23033) );
  NAND2HSV0 U25448 ( .A1(n28792), .A2(\pe6/got [4]), .ZN(n23032) );
  XOR3HSV2 U25449 ( .A1(n23034), .A2(n23033), .A3(n23032), .Z(n23035) );
  XOR2HSV0 U25450 ( .A1(n23036), .A2(n23035), .Z(n23037) );
  XNOR2HSV1 U25451 ( .A1(n23038), .A2(n23037), .ZN(n23039) );
  XNOR2HSV1 U25452 ( .A1(n23040), .A2(n23039), .ZN(n23043) );
  NAND2HSV0 U25453 ( .A1(n23041), .A2(\pe6/got [8]), .ZN(n23042) );
  XOR2HSV0 U25454 ( .A1(n23043), .A2(n23042), .Z(n23045) );
  BUFHSV8 U25455 ( .I(n25767), .Z(n26068) );
  NAND2HSV2 U25456 ( .A1(n26068), .A2(\pe6/got [9]), .ZN(n23044) );
  XNOR2HSV1 U25457 ( .A1(n23045), .A2(n23044), .ZN(n23046) );
  XNOR2HSV1 U25458 ( .A1(n23047), .A2(n23046), .ZN(n23048) );
  XOR2HSV0 U25459 ( .A1(n23049), .A2(n23048), .Z(n23050) );
  XOR2HSV0 U25460 ( .A1(n23051), .A2(n23050), .Z(n23052) );
  XOR2HSV0 U25461 ( .A1(n23053), .A2(n23052), .Z(n23054) );
  XNOR2HSV1 U25462 ( .A1(n23055), .A2(n23054), .ZN(n23056) );
  AND2HSV2 U25463 ( .A1(n27904), .A2(n25128), .Z(n23106) );
  NAND2HSV0 U25464 ( .A1(n13994), .A2(n28480), .ZN(n23103) );
  INHSV2 U25465 ( .I(n25079), .ZN(n27906) );
  NOR2HSV2 U25466 ( .A1(n27906), .A2(n27825), .ZN(n23101) );
  NAND2HSV0 U25467 ( .A1(\pe4/got [9]), .A2(n14038), .ZN(n23099) );
  NOR2HSV0 U25468 ( .A1(n27942), .A2(n27827), .ZN(n23097) );
  NAND2HSV0 U25469 ( .A1(n13996), .A2(n27877), .ZN(n23061) );
  NAND2HSV2 U25470 ( .A1(n23059), .A2(n23058), .ZN(n28578) );
  NAND2HSV0 U25471 ( .A1(n28578), .A2(n22826), .ZN(n23060) );
  XNOR2HSV1 U25472 ( .A1(n23061), .A2(n23060), .ZN(n23095) );
  NAND2HSV0 U25473 ( .A1(\pe4/ti_7[7] ), .A2(\pe4/got [5]), .ZN(n23093) );
  CLKNAND2HSV0 U25474 ( .A1(n22931), .A2(\pe4/got [4]), .ZN(n23091) );
  NAND2HSV0 U25475 ( .A1(n27830), .A2(n28626), .ZN(n23089) );
  NAND2HSV0 U25476 ( .A1(\pe4/aot [7]), .A2(\pe4/bq[7] ), .ZN(n23063) );
  NAND2HSV0 U25477 ( .A1(\pe4/aot [5]), .A2(\pe4/bq[9] ), .ZN(n23062) );
  XOR2HSV0 U25478 ( .A1(n23063), .A2(n23062), .Z(n23084) );
  NAND2HSV0 U25479 ( .A1(\pe4/aot [13]), .A2(\pe4/bq[1] ), .ZN(n23065) );
  NAND2HSV0 U25480 ( .A1(\pe4/aot [4]), .A2(\pe4/bq[10] ), .ZN(n23064) );
  XOR2HSV0 U25481 ( .A1(n23065), .A2(n23064), .Z(n23069) );
  NAND2HSV0 U25482 ( .A1(\pe4/aot [8]), .A2(\pe4/bq[6] ), .ZN(n23067) );
  NAND2HSV0 U25483 ( .A1(\pe4/aot [6]), .A2(\pe4/bq[8] ), .ZN(n23066) );
  XOR2HSV0 U25484 ( .A1(n23067), .A2(n23066), .Z(n23068) );
  XNOR2HSV1 U25485 ( .A1(n23069), .A2(n23068), .ZN(n23083) );
  NAND2HSV0 U25486 ( .A1(\pe4/aot [12]), .A2(\pe4/bq[2] ), .ZN(n26943) );
  NAND2HSV0 U25487 ( .A1(\pe4/aot [9]), .A2(\pe4/bq[5] ), .ZN(n23071) );
  CLKNAND2HSV0 U25488 ( .A1(\pe4/bq[2] ), .A2(\pe4/aot [9]), .ZN(n27841) );
  NOR2HSV0 U25489 ( .A1(n26939), .A2(n27841), .ZN(n23070) );
  AOI21HSV2 U25490 ( .A1(n26943), .A2(n23071), .B(n23070), .ZN(n23073) );
  XOR2HSV0 U25491 ( .A1(n23073), .A2(n23072), .Z(n23082) );
  NAND2HSV0 U25492 ( .A1(\pe4/aot [3]), .A2(\pe4/bq[11] ), .ZN(n23075) );
  NAND2HSV0 U25493 ( .A1(\pe4/aot [10]), .A2(\pe4/bq[4] ), .ZN(n23074) );
  XOR2HSV0 U25494 ( .A1(n23075), .A2(n23074), .Z(n23080) );
  NAND2HSV0 U25495 ( .A1(\pe4/aot [11]), .A2(\pe4/bq[3] ), .ZN(n23078) );
  NAND2HSV0 U25496 ( .A1(\pe4/aot [1]), .A2(n23076), .ZN(n23077) );
  XOR2HSV0 U25497 ( .A1(n23078), .A2(n23077), .Z(n23079) );
  XOR2HSV0 U25498 ( .A1(n23080), .A2(n23079), .Z(n23081) );
  XOR4HSV1 U25499 ( .A1(n23084), .A2(n23083), .A3(n23082), .A4(n23081), .Z(
        n23087) );
  NOR2HSV0 U25500 ( .A1(n26981), .A2(n28000), .ZN(n23086) );
  NAND2HSV0 U25501 ( .A1(n27739), .A2(n28591), .ZN(n23085) );
  XOR3HSV1 U25502 ( .A1(n23087), .A2(n23086), .A3(n23085), .Z(n23088) );
  XOR2HSV0 U25503 ( .A1(n23089), .A2(n23088), .Z(n23090) );
  XOR2HSV0 U25504 ( .A1(n23091), .A2(n23090), .Z(n23092) );
  XNOR2HSV1 U25505 ( .A1(n23093), .A2(n23092), .ZN(n23094) );
  XOR2HSV0 U25506 ( .A1(n23095), .A2(n23094), .Z(n23096) );
  XOR2HSV0 U25507 ( .A1(n23097), .A2(n23096), .Z(n23098) );
  XOR2HSV0 U25508 ( .A1(n23099), .A2(n23098), .Z(n23100) );
  XOR2HSV0 U25509 ( .A1(n23101), .A2(n23100), .Z(n23102) );
  NOR2HSV0 U25510 ( .A1(n27900), .A2(n26932), .ZN(n23104) );
  INAND2HSV2 U25511 ( .A1(n24073), .B1(n28610), .ZN(n23107) );
  INHSV3 U25512 ( .I(n23108), .ZN(n23109) );
  CLKNAND2HSV4 U25513 ( .A1(n23113), .A2(n28610), .ZN(n23114) );
  CLKNHSV3 U25514 ( .I(n23114), .ZN(n23117) );
  NAND2HSV2 U25515 ( .A1(n23120), .A2(n28948), .ZN(n23176) );
  NAND2HSV0 U25516 ( .A1(n25377), .A2(\pe7/got [12]), .ZN(n23166) );
  NAND2HSV2 U25517 ( .A1(n28430), .A2(n14022), .ZN(n23164) );
  NAND2HSV0 U25518 ( .A1(n14066), .A2(\pe7/got [9]), .ZN(n23160) );
  NAND2HSV0 U25519 ( .A1(\pe7/got [8]), .A2(n11935), .ZN(n23158) );
  NAND2HSV0 U25520 ( .A1(n11936), .A2(\pe7/got [6]), .ZN(n23156) );
  NAND2HSV0 U25521 ( .A1(n27083), .A2(\pe7/aot [3]), .ZN(n25277) );
  NAND2HSV0 U25522 ( .A1(\pe7/aot [6]), .A2(\pe7/bq[12] ), .ZN(n23121) );
  XOR2HSV0 U25523 ( .A1(n25277), .A2(n23121), .Z(n23136) );
  NAND2HSV0 U25524 ( .A1(n28876), .A2(\pe7/pvq [15]), .ZN(n23122) );
  XNOR2HSV1 U25525 ( .A1(n23122), .A2(\pe7/phq [15]), .ZN(n23127) );
  NAND2HSV0 U25526 ( .A1(\pe7/aot [14]), .A2(\pe7/bq[2] ), .ZN(n24228) );
  NAND2HSV0 U25527 ( .A1(n14078), .A2(\pe7/bq[2] ), .ZN(n25303) );
  NAND2HSV0 U25528 ( .A1(\pe7/aot [14]), .A2(\pe7/bq[4] ), .ZN(n23123) );
  CLKNAND2HSV1 U25529 ( .A1(n25303), .A2(n23123), .ZN(n23124) );
  OAI21HSV2 U25530 ( .A1(n23125), .A2(n24228), .B(n23124), .ZN(n23126) );
  XNOR2HSV1 U25531 ( .A1(n23127), .A2(n23126), .ZN(n23135) );
  NAND2HSV0 U25532 ( .A1(\pe7/aot [12]), .A2(\pe7/bq[6] ), .ZN(n23129) );
  NAND2HSV0 U25533 ( .A1(\pe7/aot [2]), .A2(n25273), .ZN(n23128) );
  XOR2HSV0 U25534 ( .A1(n23129), .A2(n23128), .Z(n23133) );
  NAND2HSV0 U25535 ( .A1(\pe7/aot [11]), .A2(\pe7/bq[7] ), .ZN(n23131) );
  NAND2HSV0 U25536 ( .A1(\pe7/aot [15]), .A2(\pe7/bq[3] ), .ZN(n23130) );
  XOR2HSV0 U25537 ( .A1(n23131), .A2(n23130), .Z(n23132) );
  XOR2HSV0 U25538 ( .A1(n23133), .A2(n23132), .Z(n23134) );
  XOR3HSV2 U25539 ( .A1(n23136), .A2(n23135), .A3(n23134), .Z(n23151) );
  NAND2HSV0 U25540 ( .A1(n25292), .A2(n25272), .ZN(n23150) );
  NAND2HSV0 U25541 ( .A1(\pe7/aot [9]), .A2(\pe7/bq[9] ), .ZN(n23140) );
  NAND2HSV0 U25542 ( .A1(\pe7/got [2]), .A2(n23138), .ZN(n23139) );
  XOR2HSV0 U25543 ( .A1(n23140), .A2(n23139), .Z(n23144) );
  NAND2HSV0 U25544 ( .A1(\pe7/aot [8]), .A2(\pe7/bq[10] ), .ZN(n23142) );
  NAND2HSV0 U25545 ( .A1(n14050), .A2(\pe7/bq[5] ), .ZN(n23141) );
  XOR2HSV0 U25546 ( .A1(n23142), .A2(n23141), .Z(n23143) );
  XOR2HSV0 U25547 ( .A1(n23144), .A2(n23143), .Z(n23146) );
  XOR2HSV0 U25548 ( .A1(n23146), .A2(n23145), .Z(n23148) );
  CLKNHSV2 U25549 ( .I(\pe7/got [3]), .ZN(n24285) );
  NOR2HSV0 U25550 ( .A1(n25309), .A2(n24285), .ZN(n23147) );
  XOR2HSV0 U25551 ( .A1(n23148), .A2(n23147), .Z(n23149) );
  XOR3HSV2 U25552 ( .A1(n23151), .A2(n23150), .A3(n23149), .Z(n23153) );
  NAND2HSV0 U25553 ( .A1(n24250), .A2(n25375), .ZN(n23152) );
  XOR2HSV0 U25554 ( .A1(n23153), .A2(n23152), .Z(n23155) );
  NAND2HSV0 U25555 ( .A1(n25318), .A2(n25271), .ZN(n23154) );
  XOR3HSV2 U25556 ( .A1(n23156), .A2(n23155), .A3(n23154), .Z(n23157) );
  XOR2HSV0 U25557 ( .A1(n23158), .A2(n23157), .Z(n23159) );
  XOR2HSV0 U25558 ( .A1(n23160), .A2(n23159), .Z(n23162) );
  XOR2HSV0 U25559 ( .A1(n23162), .A2(n23161), .Z(n23163) );
  XNOR2HSV4 U25560 ( .A1(n23164), .A2(n23163), .ZN(n23165) );
  XOR2HSV2 U25561 ( .A1(n23166), .A2(n23165), .Z(n23169) );
  INHSV2 U25562 ( .I(n23169), .ZN(n23167) );
  AOI21HSV2 U25563 ( .A1(n24287), .A2(n24181), .B(n23167), .ZN(n23168) );
  INHSV2 U25564 ( .I(n23168), .ZN(n23172) );
  NOR2HSV2 U25565 ( .A1(n23169), .A2(n19242), .ZN(n23170) );
  NAND2HSV2 U25566 ( .A1(n24287), .A2(n23170), .ZN(n23171) );
  CLKNAND2HSV3 U25567 ( .A1(n23172), .A2(n23171), .ZN(n23174) );
  NAND2HSV2 U25568 ( .A1(n23210), .A2(n24271), .ZN(n23173) );
  XNOR2HSV4 U25569 ( .A1(n23174), .A2(n23173), .ZN(n23430) );
  INHSV2 U25570 ( .I(n23430), .ZN(n23175) );
  NAND2HSV2 U25571 ( .A1(n23176), .A2(n23175), .ZN(n23179) );
  INHSV2 U25572 ( .I(n23176), .ZN(n23177) );
  NAND2HSV4 U25573 ( .A1(n23179), .A2(n23178), .ZN(n23186) );
  INHSV2 U25574 ( .I(\pe7/ti_7t [15]), .ZN(n23182) );
  NOR2HSV2 U25575 ( .A1(n23180), .A2(n23182), .ZN(n23183) );
  OAI21HSV4 U25576 ( .A1(n23187), .A2(n23186), .B(n23185), .ZN(n23549) );
  INHSV4 U25577 ( .I(n23549), .ZN(n24220) );
  NAND2HSV2 U25578 ( .A1(n23188), .A2(\pe7/ti_7t [13]), .ZN(n23189) );
  NAND2HSV4 U25579 ( .A1(n23190), .A2(n23189), .ZN(n23555) );
  INHSV2 U25580 ( .I(n23555), .ZN(n24032) );
  NOR2HSV2 U25581 ( .A1(n24032), .A2(n23191), .ZN(n23214) );
  CLKNAND2HSV0 U25582 ( .A1(n24287), .A2(\pe7/got [3]), .ZN(n23209) );
  NAND2HSV0 U25583 ( .A1(n28656), .A2(\pe7/got [2]), .ZN(n23207) );
  NAND2HSV0 U25584 ( .A1(n28430), .A2(\pe7/got [1]), .ZN(n23205) );
  NAND2HSV0 U25585 ( .A1(\pe7/aot [7]), .A2(\pe7/bq[1] ), .ZN(n23193) );
  NAND2HSV0 U25586 ( .A1(\pe7/aot [2]), .A2(\pe7/bq[6] ), .ZN(n23192) );
  XOR2HSV0 U25587 ( .A1(n23193), .A2(n23192), .Z(n23197) );
  NAND2HSV0 U25588 ( .A1(\pe7/aot [4]), .A2(\pe7/bq[4] ), .ZN(n23195) );
  NAND2HSV0 U25589 ( .A1(\pe7/aot [1]), .A2(\pe7/bq[7] ), .ZN(n23194) );
  XOR2HSV0 U25590 ( .A1(n23195), .A2(n23194), .Z(n23196) );
  XOR2HSV0 U25591 ( .A1(n23197), .A2(n23196), .Z(n23203) );
  NAND2HSV0 U25592 ( .A1(\pe7/aot [6]), .A2(\pe7/bq[2] ), .ZN(n23199) );
  NAND2HSV0 U25593 ( .A1(\pe7/aot [5]), .A2(\pe7/bq[3] ), .ZN(n23198) );
  XOR2HSV0 U25594 ( .A1(n23199), .A2(n23198), .Z(n23201) );
  NAND2HSV0 U25595 ( .A1(\pe7/aot [3]), .A2(\pe7/bq[5] ), .ZN(n23200) );
  XNOR2HSV1 U25596 ( .A1(n23201), .A2(n23200), .ZN(n23202) );
  XNOR2HSV1 U25597 ( .A1(n23203), .A2(n23202), .ZN(n23204) );
  XOR2HSV0 U25598 ( .A1(n23205), .A2(n23204), .Z(n23206) );
  XNOR2HSV1 U25599 ( .A1(n23207), .A2(n23206), .ZN(n23208) );
  XOR2HSV0 U25600 ( .A1(n23209), .A2(n23208), .Z(n23212) );
  BUFHSV4 U25601 ( .I(n23210), .Z(n25335) );
  NAND2HSV0 U25602 ( .A1(n25335), .A2(n25272), .ZN(n23211) );
  XOR2HSV0 U25603 ( .A1(n23212), .A2(n23211), .Z(n23213) );
  NOR2HSV4 U25604 ( .A1(n27195), .A2(n26186), .ZN(n23224) );
  NAND2HSV0 U25605 ( .A1(\pe10/aot [1]), .A2(\pe10/bq[3] ), .ZN(n23221) );
  NAND2HSV0 U25606 ( .A1(\pe10/aot [2]), .A2(\pe10/bq[2] ), .ZN(n23220) );
  XOR2HSV0 U25607 ( .A1(n23221), .A2(n23220), .Z(n23223) );
  NOR2HSV2 U25608 ( .A1(n23222), .A2(n26163), .ZN(n26162) );
  XNOR2HSV1 U25609 ( .A1(n23228), .A2(n23227), .ZN(\pe10/poht [13]) );
  NAND2HSV0 U25610 ( .A1(n14055), .A2(n27736), .ZN(n23231) );
  INHSV2 U25611 ( .I(\pe2/aot [1]), .ZN(n27693) );
  INHSV2 U25612 ( .I(\pe2/bq[1] ), .ZN(n27652) );
  NOR2HSV2 U25613 ( .A1(n27693), .A2(n27652), .ZN(n27672) );
  XNOR2HSV0 U25614 ( .A1(n23231), .A2(n27672), .ZN(\pe2/poht [15]) );
  CLKNHSV0 U25615 ( .I(n23239), .ZN(n23237) );
  NAND2HSV2 U25616 ( .A1(n12517), .A2(n28640), .ZN(n23235) );
  NAND2HSV0 U25617 ( .A1(\pe5/aot [1]), .A2(\pe5/bq[3] ), .ZN(n23232) );
  XOR2HSV0 U25618 ( .A1(n23233), .A2(n23232), .Z(n23234) );
  CLKNHSV0 U25619 ( .I(n23238), .ZN(n23236) );
  CLKNAND2HSV1 U25620 ( .A1(n23237), .A2(n23236), .ZN(n23241) );
  CLKNAND2HSV0 U25621 ( .A1(n23239), .A2(n23238), .ZN(n23240) );
  CLKNAND2HSV0 U25622 ( .A1(n23243), .A2(n23242), .ZN(pov9[14]) );
  NAND2HSV0 U25623 ( .A1(\pe5/ti_7[10] ), .A2(\pe5/got [3]), .ZN(n23265) );
  NAND2HSV0 U25624 ( .A1(\pe5/aot [3]), .A2(\pe5/bq[6] ), .ZN(n23247) );
  NAND2HSV0 U25625 ( .A1(\pe5/aot [2]), .A2(\pe5/bq[7] ), .ZN(n23246) );
  XOR2HSV0 U25626 ( .A1(n23247), .A2(n23246), .Z(n23251) );
  NAND2HSV0 U25627 ( .A1(\pe5/aot [5]), .A2(\pe5/bq[4] ), .ZN(n23249) );
  NAND2HSV0 U25628 ( .A1(\pe5/aot [1]), .A2(\pe5/bq[8] ), .ZN(n23248) );
  XOR2HSV0 U25629 ( .A1(n23249), .A2(n23248), .Z(n23250) );
  XOR2HSV0 U25630 ( .A1(n23251), .A2(n23250), .Z(n23259) );
  NAND2HSV0 U25631 ( .A1(\pe5/aot [8]), .A2(\pe5/bq[1] ), .ZN(n23253) );
  NAND2HSV0 U25632 ( .A1(\pe5/aot [4]), .A2(\pe5/bq[5] ), .ZN(n23252) );
  XOR2HSV0 U25633 ( .A1(n23253), .A2(n23252), .Z(n23257) );
  XNOR2HSV1 U25634 ( .A1(n23257), .A2(n23256), .ZN(n23258) );
  XNOR2HSV1 U25635 ( .A1(n23259), .A2(n23258), .ZN(n23263) );
  NOR2HSV2 U25636 ( .A1(n24684), .A2(n24638), .ZN(n23262) );
  OR2HSV1 U25637 ( .A1(n24686), .A2(n23260), .Z(n23261) );
  XOR3HSV2 U25638 ( .A1(n23263), .A2(n23262), .A3(n23261), .Z(n23264) );
  XNOR2HSV1 U25639 ( .A1(n23265), .A2(n23264), .ZN(n23268) );
  BUFHSV2 U25640 ( .I(n23266), .Z(n28803) );
  XNOR2HSV1 U25641 ( .A1(n23268), .A2(n23267), .ZN(n23269) );
  AOI21HSV0 U25642 ( .A1(n23275), .A2(n20870), .B(n24683), .ZN(n23276) );
  NAND2HSV0 U25643 ( .A1(n25137), .A2(\pe11/got [6]), .ZN(n23306) );
  NAND2HSV0 U25644 ( .A1(n14063), .A2(\pe11/got [5]), .ZN(n23304) );
  NAND2HSV0 U25645 ( .A1(n25138), .A2(\pe11/got [3]), .ZN(n23299) );
  NAND2HSV0 U25646 ( .A1(n25139), .A2(\pe11/got [2]), .ZN(n23297) );
  NAND2HSV0 U25647 ( .A1(n28471), .A2(\pe11/got [1]), .ZN(n23295) );
  NAND2HSV0 U25648 ( .A1(\pe11/bq[9] ), .A2(\pe11/aot [2]), .ZN(n24766) );
  NAND2HSV0 U25649 ( .A1(\pe11/bq[6] ), .A2(\pe11/aot [5]), .ZN(n23278) );
  XOR2HSV0 U25650 ( .A1(n24766), .A2(n23278), .Z(n23293) );
  NAND2HSV0 U25651 ( .A1(\pe11/bq[8] ), .A2(\pe11/aot [3]), .ZN(n23280) );
  NAND2HSV0 U25652 ( .A1(\pe11/bq[4] ), .A2(\pe11/aot [7]), .ZN(n23279) );
  XOR2HSV0 U25653 ( .A1(n23280), .A2(n23279), .Z(n23284) );
  NAND2HSV0 U25654 ( .A1(\pe11/bq[10] ), .A2(\pe11/aot [1]), .ZN(n23282) );
  NAND2HSV0 U25655 ( .A1(\pe11/bq[5] ), .A2(\pe11/aot [6]), .ZN(n23281) );
  XOR2HSV0 U25656 ( .A1(n23282), .A2(n23281), .Z(n23283) );
  XNOR2HSV1 U25657 ( .A1(n23284), .A2(n23283), .ZN(n23292) );
  NAND2HSV0 U25658 ( .A1(\pe11/bq[3] ), .A2(\pe11/aot [8]), .ZN(n23286) );
  NAND2HSV0 U25659 ( .A1(\pe11/bq[1] ), .A2(\pe11/aot [10]), .ZN(n23285) );
  XOR2HSV0 U25660 ( .A1(n23286), .A2(n23285), .Z(n23290) );
  NAND2HSV0 U25661 ( .A1(\pe11/bq[2] ), .A2(\pe11/aot [9]), .ZN(n23288) );
  NAND2HSV0 U25662 ( .A1(\pe11/bq[7] ), .A2(\pe11/aot [4]), .ZN(n23287) );
  XOR2HSV0 U25663 ( .A1(n23288), .A2(n23287), .Z(n23289) );
  XOR2HSV0 U25664 ( .A1(n23290), .A2(n23289), .Z(n23291) );
  XOR3HSV2 U25665 ( .A1(n23293), .A2(n23292), .A3(n23291), .Z(n23294) );
  XNOR2HSV1 U25666 ( .A1(n23295), .A2(n23294), .ZN(n23296) );
  XNOR2HSV1 U25667 ( .A1(n23297), .A2(n23296), .ZN(n23298) );
  XNOR2HSV1 U25668 ( .A1(n23299), .A2(n23298), .ZN(n23302) );
  INHSV2 U25669 ( .I(n23300), .ZN(n28464) );
  NAND2HSV0 U25670 ( .A1(n28464), .A2(\pe11/got [4]), .ZN(n23301) );
  XOR2HSV0 U25671 ( .A1(n23302), .A2(n23301), .Z(n23303) );
  XOR2HSV0 U25672 ( .A1(n23304), .A2(n23303), .Z(n23305) );
  XNOR2HSV1 U25673 ( .A1(n23306), .A2(n23305), .ZN(n23308) );
  NAND2HSV0 U25674 ( .A1(n28919), .A2(\pe11/got [7]), .ZN(n23307) );
  NAND2HSV2 U25675 ( .A1(n24902), .A2(\pe11/got [4]), .ZN(n23318) );
  NAND2HSV0 U25676 ( .A1(\pe11/bq[1] ), .A2(\pe11/aot [5]), .ZN(n23315) );
  NAND2HSV0 U25677 ( .A1(\pe11/bq[5] ), .A2(\pe11/aot [1]), .ZN(n23310) );
  NAND2HSV0 U25678 ( .A1(\pe11/bq[2] ), .A2(\pe11/aot [4]), .ZN(n23309) );
  XNOR2HSV1 U25679 ( .A1(n23310), .A2(n23309), .ZN(n23314) );
  NAND2HSV0 U25680 ( .A1(\pe11/bq[4] ), .A2(\pe11/aot [2]), .ZN(n23312) );
  NAND2HSV0 U25681 ( .A1(\pe11/bq[3] ), .A2(\pe11/aot [3]), .ZN(n23311) );
  XOR2HSV0 U25682 ( .A1(n23312), .A2(n23311), .Z(n23313) );
  XOR3HSV2 U25683 ( .A1(n23315), .A2(n23314), .A3(n23313), .Z(n23316) );
  XNOR2HSV4 U25684 ( .A1(n23318), .A2(n23317), .ZN(n23322) );
  CLKNAND2HSV1 U25685 ( .A1(n28927), .A2(\pe11/got [5]), .ZN(n23321) );
  NAND2HSV0 U25686 ( .A1(\pe11/bq[2] ), .A2(\pe11/aot [2]), .ZN(n23324) );
  NAND2HSV0 U25687 ( .A1(\pe11/bq[3] ), .A2(\pe11/aot [1]), .ZN(n23323) );
  XOR2HSV0 U25688 ( .A1(n23324), .A2(n23323), .Z(n23326) );
  NAND2HSV0 U25689 ( .A1(\pe11/bq[1] ), .A2(\pe11/aot [3]), .ZN(n23325) );
  CLKBUFHSV4 U25690 ( .I(n28945), .Z(n26634) );
  NAND2HSV0 U25691 ( .A1(n23327), .A2(\pe3/got [10]), .ZN(n23371) );
  NAND2HSV0 U25692 ( .A1(n26682), .A2(n28648), .ZN(n23365) );
  NAND2HSV0 U25693 ( .A1(n15240), .A2(\pe3/got [6]), .ZN(n23363) );
  NAND2HSV0 U25694 ( .A1(n26350), .A2(\pe3/got [4]), .ZN(n23361) );
  NAND2HSV0 U25695 ( .A1(n26242), .A2(\pe3/got [5]), .ZN(n23360) );
  NAND2HSV0 U25696 ( .A1(\pe3/aot [4]), .A2(n14026), .ZN(n23331) );
  NAND2HSV0 U25697 ( .A1(\pe3/aot [12]), .A2(\pe3/bq[6] ), .ZN(n23330) );
  XOR2HSV0 U25698 ( .A1(n23331), .A2(n23330), .Z(n23335) );
  NAND2HSV0 U25699 ( .A1(\pe3/aot [11]), .A2(\pe3/bq[7] ), .ZN(n23333) );
  NAND2HSV0 U25700 ( .A1(\pe3/got [2]), .A2(n15044), .ZN(n23332) );
  XOR2HSV0 U25701 ( .A1(n23333), .A2(n23332), .Z(n23334) );
  XOR2HSV0 U25702 ( .A1(n23335), .A2(n23334), .Z(n23338) );
  CLKNHSV0 U25703 ( .I(\pe3/bq[12] ), .ZN(n24535) );
  XOR2HSV0 U25704 ( .A1(n23338), .A2(n23337), .Z(n23341) );
  NAND2HSV0 U25705 ( .A1(n26367), .A2(\pe3/got [3]), .ZN(n23340) );
  XNOR2HSV1 U25706 ( .A1(n23341), .A2(n23340), .ZN(n23358) );
  CLKNHSV0 U25707 ( .I(\pe3/bq[10] ), .ZN(n23342) );
  INHSV2 U25708 ( .I(n23342), .ZN(n23490) );
  NAND2HSV0 U25709 ( .A1(\pe3/aot [8]), .A2(n23490), .ZN(n23686) );
  NAND2HSV0 U25710 ( .A1(\pe3/aot [7]), .A2(\pe3/bq[11] ), .ZN(n26688) );
  XOR2HSV0 U25711 ( .A1(n23686), .A2(n26688), .Z(n23356) );
  NAND2HSV0 U25712 ( .A1(\pe3/aot [10]), .A2(\pe3/bq[8] ), .ZN(n23344) );
  NAND2HSV0 U25713 ( .A1(\pe3/aot [5]), .A2(\pe3/bq[13] ), .ZN(n23343) );
  XOR2HSV0 U25714 ( .A1(n23344), .A2(n23343), .Z(n23347) );
  XNOR2HSV1 U25715 ( .A1(n23347), .A2(n23346), .ZN(n23355) );
  NAND2HSV0 U25716 ( .A1(\pe3/aot [9]), .A2(\pe3/bq[9] ), .ZN(n24532) );
  XOR2HSV0 U25717 ( .A1(n23348), .A2(n24532), .Z(n23353) );
  NAND2HSV0 U25718 ( .A1(\pe3/aot [14]), .A2(\pe3/bq[4] ), .ZN(n23351) );
  NAND2HSV0 U25719 ( .A1(\pe3/aot [3]), .A2(n26373), .ZN(n23350) );
  XOR2HSV0 U25720 ( .A1(n23351), .A2(n23350), .Z(n23352) );
  XOR2HSV0 U25721 ( .A1(n23353), .A2(n23352), .Z(n23354) );
  XOR3HSV2 U25722 ( .A1(n23356), .A2(n23355), .A3(n23354), .Z(n23357) );
  XNOR2HSV1 U25723 ( .A1(n23358), .A2(n23357), .ZN(n23359) );
  XOR3HSV1 U25724 ( .A1(n23361), .A2(n23360), .A3(n23359), .Z(n23362) );
  XNOR2HSV1 U25725 ( .A1(n23363), .A2(n23362), .ZN(n23364) );
  XNOR2HSV1 U25726 ( .A1(n23365), .A2(n23364), .ZN(n23367) );
  CLKNHSV1 U25727 ( .I(\pe3/got [7]), .ZN(n23682) );
  NOR2HSV0 U25728 ( .A1(n26625), .A2(n23682), .ZN(n23366) );
  XNOR2HSV1 U25729 ( .A1(n23367), .A2(n23366), .ZN(n23368) );
  INHSV2 U25730 ( .I(n23374), .ZN(n24499) );
  NAND2HSV0 U25731 ( .A1(n26291), .A2(\pe3/got [13]), .ZN(n23380) );
  XNOR2HSV4 U25732 ( .A1(n23381), .A2(n23380), .ZN(n23389) );
  INHSV2 U25733 ( .I(n23389), .ZN(n23388) );
  AND2HSV2 U25734 ( .A1(n23382), .A2(n15086), .Z(n23386) );
  NOR2HSV0 U25735 ( .A1(n23384), .A2(n23383), .ZN(n23385) );
  AOI21HSV2 U25736 ( .A1(n21312), .A2(n23386), .B(n23385), .ZN(n23387) );
  NAND2HSV2 U25737 ( .A1(n23409), .A2(n23408), .ZN(n23413) );
  CLKNHSV1 U25738 ( .I(n23390), .ZN(n23391) );
  NOR2HSV2 U25739 ( .A1(n23391), .A2(n21732), .ZN(n23407) );
  CLKNHSV1 U25740 ( .I(n23392), .ZN(n23394) );
  CLKNHSV0 U25741 ( .I(n23396), .ZN(n23393) );
  NOR2HSV2 U25742 ( .A1(n23394), .A2(n23393), .ZN(n23406) );
  CLKNHSV0 U25743 ( .I(n23395), .ZN(n23399) );
  NAND2HSV0 U25744 ( .A1(n23397), .A2(n23396), .ZN(n23398) );
  NOR2HSV2 U25745 ( .A1(n23399), .A2(n23398), .ZN(n23401) );
  CLKNAND2HSV1 U25746 ( .A1(n23401), .A2(n23400), .ZN(n23404) );
  AOI21HSV4 U25747 ( .A1(n23407), .A2(n23406), .B(n23405), .ZN(n23412) );
  CLKNAND2HSV2 U25748 ( .A1(n23410), .A2(n23412), .ZN(n23411) );
  OAI21HSV4 U25749 ( .A1(n23413), .A2(n12301), .B(n23411), .ZN(n23668) );
  OAI21HSV2 U25750 ( .A1(n23417), .A2(n23416), .B(n23415), .ZN(n23418) );
  INHSV3 U25751 ( .I(n24628), .ZN(n23670) );
  INHSV4 U25752 ( .I(n23670), .ZN(n24522) );
  BUFHSV2 U25753 ( .I(n23423), .Z(n23424) );
  NOR2HSV2 U25754 ( .A1(n24032), .A2(n25339), .ZN(n23429) );
  CLKNHSV0 U25755 ( .I(n23425), .ZN(n23426) );
  INHSV2 U25756 ( .I(n23426), .ZN(n23427) );
  XOR3HSV1 U25757 ( .A1(n23430), .A2(n23429), .A3(n23428), .Z(n28978) );
  INHSV2 U25758 ( .I(n14972), .ZN(n27218) );
  INHSV2 U25759 ( .I(n25914), .ZN(n27185) );
  XNOR2HSV0 U25760 ( .A1(n23444), .A2(n23443), .ZN(n28994) );
  CLKNAND2HSV1 U25761 ( .A1(n23446), .A2(n23445), .ZN(n27283) );
  CLKNHSV0 U25762 ( .I(n23453), .ZN(n28474) );
  INHSV4 U25763 ( .I(n23455), .ZN(n25981) );
  INHSV2 U25764 ( .I(n25981), .ZN(n28937) );
  INHSV2 U25765 ( .I(n23456), .ZN(n26416) );
  INHSV2 U25766 ( .I(n27876), .ZN(n28583) );
  CLKNHSV0 U25767 ( .I(n28508), .ZN(n23801) );
  BUFHSV2 U25768 ( .I(n23801), .Z(n23795) );
  CLKNHSV0 U25769 ( .I(n23796), .ZN(n28597) );
  CLKNHSV0 U25770 ( .I(n28597), .ZN(n23800) );
  BUFHSV2 U25771 ( .I(n23800), .Z(n23797) );
  CLKNHSV0 U25772 ( .I(n23798), .ZN(n28553) );
  CLKNHSV0 U25773 ( .I(n28553), .ZN(n23799) );
  CLKNHSV0 U25774 ( .I(n26094), .ZN(n28675) );
  CLKNHSV0 U25775 ( .I(n28547), .ZN(n24308) );
  CLKNHSV0 U25776 ( .I(n23462), .ZN(n28672) );
  CLKNHSV0 U25777 ( .I(n23467), .ZN(pov5[6]) );
  BUFHSV2 U25778 ( .I(n23468), .Z(n23469) );
  NAND2HSV0 U25779 ( .A1(n28427), .A2(n28693), .ZN(n23472) );
  XNOR2HSV0 U25780 ( .A1(n23472), .A2(n23471), .ZN(n29042) );
  CLKNHSV0 U25781 ( .I(n28487), .ZN(n24309) );
  CLKNHSV0 U25782 ( .I(n23801), .ZN(n28524) );
  INHSV1 U25783 ( .I(n27423), .ZN(n28953) );
  CLKNHSV0 U25784 ( .I(n23801), .ZN(n28452) );
  CLKNHSV0 U25785 ( .I(n24308), .ZN(n28602) );
  CLKNHSV0 U25786 ( .I(n23795), .ZN(n28542) );
  MUX2HSV2 U25787 ( .I0(bo6[14]), .I1(n23485), .S(n23486), .Z(n28869) );
  MUX2HSV1 U25788 ( .I0(bo6[9]), .I1(n14012), .S(n23486), .Z(n28874) );
  CLKNHSV0 U25789 ( .I(\pe4/bq[5] ), .ZN(n27793) );
  MUX2HSV2 U25790 ( .I0(bo4[5]), .I1(\pe4/bq[5] ), .S(n27066), .Z(n28858) );
  MUX2HSV2 U25791 ( .I0(bo4[9]), .I1(\pe4/bq[9] ), .S(n27129), .Z(n28857) );
  MUX2HSV2 U25792 ( .I0(bo11[6]), .I1(\pe11/bq[6] ), .S(n20650), .Z(n28724) );
  INHSV2 U25793 ( .I(n28682), .ZN(n23487) );
  MUX2HSV2 U25794 ( .I0(n23909), .I1(bo5[12]), .S(n23487), .Z(n28861) );
  MUX2HSV2 U25795 ( .I0(n24647), .I1(bo5[15]), .S(n23487), .Z(n28860) );
  CLKNHSV0 U25796 ( .I(\pe7/bq[9] ), .ZN(n23488) );
  INHSV2 U25797 ( .I(n23488), .ZN(n23489) );
  MUX2HSV2 U25798 ( .I0(bo7[9]), .I1(n23489), .S(n27094), .Z(n28879) );
  MUX2HSV2 U25799 ( .I0(bo3[7]), .I1(\pe3/bq[7] ), .S(n23543), .Z(n28847) );
  MUX2HSV1 U25800 ( .I0(bo3[3]), .I1(\pe3/bq[3] ), .S(n23524), .Z(n28850) );
  MUX2HSV2 U25801 ( .I0(bo3[10]), .I1(n23490), .S(n23520), .Z(n28844) );
  CLKNHSV0 U25802 ( .I(\pe3/bq[9] ), .ZN(n23491) );
  INHSV2 U25803 ( .I(n23491), .ZN(n23492) );
  MUX2HSV2 U25804 ( .I0(bo3[9]), .I1(n23492), .S(n23524), .Z(n28843) );
  CLKNHSV0 U25805 ( .I(\pe3/bq[8] ), .ZN(n23493) );
  INHSV2 U25806 ( .I(n23493), .ZN(n23494) );
  MUX2HSV2 U25807 ( .I0(bo3[8]), .I1(n23494), .S(n23517), .Z(n28846) );
  CLKNHSV0 U25808 ( .I(\pe7/bq[6] ), .ZN(n23495) );
  INHSV2 U25809 ( .I(n23495), .ZN(n23496) );
  MUX2HSV2 U25810 ( .I0(bo7[6]), .I1(n23496), .S(n27102), .Z(n28880) );
  MUX2HSV1 U25811 ( .I0(bo6[11]), .I1(\pe6/bq[11] ), .S(n23498), .Z(n28872) );
  CLKNHSV0 U25812 ( .I(\pe11/bq[1] ), .ZN(n25413) );
  MUX2HSV2 U25813 ( .I0(bo11[2]), .I1(\pe11/bq[2] ), .S(n23499), .Z(n28721) );
  BUFHSV2 U25814 ( .I(n27074), .Z(n24305) );
  MUX2HSV2 U25815 ( .I0(\pe6/bq[4] ), .I1(bo6[4]), .S(n24305), .Z(n28875) );
  BUFHSV2 U25816 ( .I(n28639), .Z(n24320) );
  MUX2HSV1 U25817 ( .I0(bo11[8]), .I1(\pe11/bq[8] ), .S(n24320), .Z(n28718) );
  MUX2HSV2 U25818 ( .I0(bo11[9]), .I1(\pe11/bq[9] ), .S(n27055), .Z(n28917) );
  MUX2HSV2 U25819 ( .I0(bo11[10]), .I1(\pe11/bq[10] ), .S(n22111), .Z(n28916)
         );
  MUX2HSV2 U25820 ( .I0(bo8[13]), .I1(n25565), .S(n23545), .Z(n28886) );
  MUX2HSV2 U25821 ( .I0(bo8[15]), .I1(n18720), .S(n23547), .Z(n28881) );
  MUX2HSV1 U25822 ( .I0(bo10[8]), .I1(\pe10/bq[8] ), .S(n14035), .Z(n28907) );
  MUX2HSV1 U25823 ( .I0(bo10[6]), .I1(\pe10/bq[6] ), .S(n14035), .Z(n28909) );
  MUX2HSV1 U25824 ( .I0(bo10[4]), .I1(\pe10/bq[4] ), .S(n14035), .Z(n28911) );
  BUFHSV2 U25825 ( .I(n27311), .Z(n25623) );
  MUX2HSV2 U25826 ( .I0(bo2[14]), .I1(n27312), .S(n25623), .Z(n28824) );
  BUFHSV2 U25827 ( .I(n27311), .Z(n27059) );
  MUX2HSV1 U25828 ( .I0(bo2[12]), .I1(n14016), .S(n27059), .Z(n28829) );
  CLKNHSV0 U25829 ( .I(\pe2/bq[11] ), .ZN(n23500) );
  INHSV2 U25830 ( .I(n23500), .ZN(n23501) );
  MUX2HSV2 U25831 ( .I0(bo2[11]), .I1(n23501), .S(n23503), .Z(n28828) );
  MUX2HSV1 U25832 ( .I0(bo2[8]), .I1(\pe2/bq[8] ), .S(n27059), .Z(n28831) );
  INHSV2 U25833 ( .I(n23505), .ZN(n23506) );
  MUX2HSV2 U25834 ( .I0(\pe5/bq[8] ), .I1(bo5[8]), .S(n23506), .Z(n28862) );
  INHSV2 U25835 ( .I(n23505), .ZN(n27051) );
  INHSV2 U25836 ( .I(n27050), .ZN(n27048) );
  MUX2HSV2 U25837 ( .I0(\pe5/bq[5] ), .I1(bo5[5]), .S(n27048), .Z(n28864) );
  MUX2HSV2 U25838 ( .I0(\pe5/bq[4] ), .I1(bo5[4]), .S(n23506), .Z(n28865) );
  MUX2HSV2 U25839 ( .I0(n23507), .I1(bo5[14]), .S(n23506), .Z(n28859) );
  BUFHSV2 U25840 ( .I(n28811), .Z(n23510) );
  MUX2HSV1 U25841 ( .I0(bo10[7]), .I1(n14010), .S(n23510), .Z(n28908) );
  BUFHSV2 U25842 ( .I(n28811), .Z(n23512) );
  MUX2HSV2 U25843 ( .I0(bo10[5]), .I1(\pe10/bq[5] ), .S(n23512), .Z(n28910) );
  MUX2HSV2 U25844 ( .I0(bo10[3]), .I1(\pe10/bq[3] ), .S(n23512), .Z(n28914) );
  BUFHSV2 U25845 ( .I(n28811), .Z(n23514) );
  MUX2HSV1 U25846 ( .I0(bo10[2]), .I1(\pe10/bq[2] ), .S(n23514), .Z(n28913) );
  BUFHSV2 U25847 ( .I(n23537), .Z(n28835) );
  INHSV2 U25848 ( .I(n27652), .ZN(n27723) );
  MUX2HSV2 U25849 ( .I0(bo2[1]), .I1(n27723), .S(n28835), .Z(n28836) );
  CLKNHSV0 U25850 ( .I(\pe2/bq[2] ), .ZN(n27554) );
  MUX2HSV1 U25851 ( .I0(bo4[11]), .I1(\pe4/bq[11] ), .S(n23508), .Z(n28774) );
  MUX2HSV2 U25852 ( .I0(bo2[3]), .I1(\pe2/bq[3] ), .S(n25623), .Z(n28837) );
  MUX2HSV2 U25853 ( .I0(bo10[15]), .I1(n16897), .S(n23514), .Z(n28899) );
  MUX2HSV2 U25854 ( .I0(bo10[11]), .I1(\pe10/bq[11] ), .S(n23513), .Z(n28904)
         );
  MUX2HSV2 U25855 ( .I0(bo10[9]), .I1(n23515), .S(n23514), .Z(n28906) );
  INHSV2 U25856 ( .I(n24316), .ZN(n23534) );
  MUX2HSV2 U25857 ( .I0(bo1[15]), .I1(n26548), .S(n23534), .Z(n28817) );
  MUX2HSV2 U25858 ( .I0(bo3[15]), .I1(n26373), .S(n23518), .Z(n28842) );
  MUX2HSV2 U25859 ( .I0(bo3[14]), .I1(n14026), .S(n23517), .Z(n28841) );
  MUX2HSV2 U25860 ( .I0(bo8[1]), .I1(\pe8/bq[1] ), .S(n23519), .Z(n28895) );
  MUX2HSV2 U25861 ( .I0(bo3[1]), .I1(\pe3/bq[1] ), .S(n23520), .Z(n28853) );
  CLKNHSV0 U25862 ( .I(\pe7/bq[12] ), .ZN(n23521) );
  INHSV2 U25863 ( .I(n23521), .ZN(n23523) );
  MUX2HSV2 U25864 ( .I0(bo7[12]), .I1(n23523), .S(n27102), .Z(n28877) );
  MUX2HSV1 U25865 ( .I0(bo3[2]), .I1(\pe3/bq[2] ), .S(n15937), .Z(n28852) );
  MUX2HSV2 U25866 ( .I0(bo3[4]), .I1(\pe3/bq[4] ), .S(n15937), .Z(n28851) );
  INHSV2 U25867 ( .I(n28623), .ZN(n23545) );
  MUX2HSV2 U25868 ( .I0(bo8[9]), .I1(\pe8/bq[9] ), .S(n14036), .Z(n28888) );
  MUX2HSV1 U25869 ( .I0(bo6[2]), .I1(\pe6/bq[2] ), .S(n23525), .Z(n28783) );
  MUX2HSV2 U25870 ( .I0(bo8[8]), .I1(\pe8/bq[8] ), .S(n23545), .Z(n28889) );
  CLKNHSV0 U25871 ( .I(\pe8/bq[6] ), .ZN(n23526) );
  INHSV2 U25872 ( .I(n23526), .ZN(n23527) );
  MUX2HSV2 U25873 ( .I0(bo8[6]), .I1(n23527), .S(n23545), .Z(n28894) );
  MUX2HSV2 U25874 ( .I0(bo8[5]), .I1(n23529), .S(n14036), .Z(n28892) );
  INHSV2 U25875 ( .I(n28623), .ZN(n25625) );
  MUX2HSV1 U25876 ( .I0(bo8[4]), .I1(\pe8/bq[4] ), .S(n23547), .Z(n28893) );
  MUX2HSV1 U25877 ( .I0(bo8[3]), .I1(\pe8/bq[3] ), .S(n18673), .Z(n28891) );
  MUX2HSV1 U25878 ( .I0(bo9[1]), .I1(\pe9/bq[1] ), .S(n23530), .Z(n28755) );
  MUX2HSV1 U25879 ( .I0(bo9[9]), .I1(\pe9/bq[9] ), .S(n23530), .Z(n28771) );
  CLKNHSV0 U25880 ( .I(\pe8/bq[12] ), .ZN(n23532) );
  INHSV1 U25881 ( .I(n23532), .ZN(n23533) );
  MUX2HSV1 U25882 ( .I0(bo8[12]), .I1(n23533), .S(n25625), .Z(n28885) );
  INHSV2 U25883 ( .I(n24316), .ZN(n28598) );
  MUX2HSV2 U25884 ( .I0(bo1[9]), .I1(\pe1/bq[9] ), .S(n28598), .Z(n28819) );
  MUX2HSV2 U25885 ( .I0(bo1[11]), .I1(\pe1/bq[11] ), .S(n23534), .Z(n28818) );
  MUX2HSV2 U25886 ( .I0(bo4[15]), .I1(n26958), .S(n23508), .Z(n28855) );
  MUX2HSV1 U25887 ( .I0(bo2[13]), .I1(n14014), .S(n23537), .Z(n28825) );
  MUX2HSV2 U25888 ( .I0(bo10[12]), .I1(\pe10/bq[12] ), .S(n23536), .Z(n28903)
         );
  MUX2HSV1 U25889 ( .I0(bo2[10]), .I1(n14018), .S(n23537), .Z(n28826) );
  INHSV2 U25890 ( .I(\pe2/bq[6] ), .ZN(n27654) );
  INHSV2 U25891 ( .I(n27654), .ZN(n27668) );
  MUX2HSV2 U25892 ( .I0(bo2[6]), .I1(n27668), .S(n23539), .Z(n28833) );
  MUX2HSV2 U25893 ( .I0(bo2[5]), .I1(\pe2/bq[5] ), .S(n23539), .Z(n28832) );
  CLKNHSV0 U25894 ( .I(\pe3/bq[5] ), .ZN(n23540) );
  INHSV2 U25895 ( .I(n23540), .ZN(n23542) );
  MUX2HSV2 U25896 ( .I0(bo3[5]), .I1(n23542), .S(n23543), .Z(n28849) );
  MUX2HSV1 U25897 ( .I0(bo3[6]), .I1(n14076), .S(n23543), .Z(n28848) );
  MUX2HSV1 U25898 ( .I0(bo10[16]), .I1(\pe10/bq[16] ), .S(n23544), .Z(n28901)
         );
  MUX2HSV1 U25899 ( .I0(bo8[16]), .I1(n25539), .S(n23545), .Z(n28884) );
  MUX2HSV1 U25900 ( .I0(bo8[14]), .I1(n23627), .S(n25625), .Z(n28882) );
  MUX2HSV1 U25901 ( .I0(bo8[11]), .I1(\pe8/bq[11] ), .S(n23547), .Z(n28883) );
  NAND2HSV2 U25902 ( .A1(n24500), .A2(n24499), .ZN(n28438) );
  CLKNHSV0 U25903 ( .I(n24309), .ZN(n28439) );
  CLKNHSV0 U25904 ( .I(n24310), .ZN(n28440) );
  CLKNHSV0 U25905 ( .I(n23791), .ZN(n28441) );
  CLKNHSV0 U25906 ( .I(n23791), .ZN(n28442) );
  CLKNHSV0 U25907 ( .I(n23790), .ZN(n28443) );
  CLKNHSV0 U25908 ( .I(n23791), .ZN(n28444) );
  CLKNHSV0 U25909 ( .I(n23791), .ZN(n28445) );
  CLKNHSV0 U25910 ( .I(n24309), .ZN(n28446) );
  CLKNHSV0 U25911 ( .I(n23793), .ZN(n28447) );
  CLKNHSV0 U25912 ( .I(n23791), .ZN(n28565) );
  CLKNHSV0 U25913 ( .I(n24310), .ZN(n28448) );
  CLKNHSV0 U25914 ( .I(n24310), .ZN(n28449) );
  CLKNHSV0 U25915 ( .I(n14021), .ZN(n23796) );
  CLKNHSV0 U25916 ( .I(n23796), .ZN(n28450) );
  CLKNHSV0 U25917 ( .I(n23796), .ZN(n28451) );
  CLKNHSV0 U25918 ( .I(n23791), .ZN(n28453) );
  NAND2HSV0 U25919 ( .A1(\pe7/aot [2]), .A2(\pe7/bq[2] ), .ZN(n23552) );
  NAND2HSV0 U25920 ( .A1(\pe7/aot [1]), .A2(\pe7/bq[3] ), .ZN(n23551) );
  XOR2HSV0 U25921 ( .A1(n23552), .A2(n23551), .Z(n23554) );
  NAND2HSV0 U25922 ( .A1(\pe7/aot [3]), .A2(\pe7/bq[1] ), .ZN(n23553) );
  XNOR2HSV1 U25923 ( .A1(n23554), .A2(n23553), .ZN(n23558) );
  INHSV2 U25924 ( .I(n23555), .ZN(n24045) );
  CLKNHSV2 U25925 ( .I(\pe7/got [1]), .ZN(n24221) );
  NOR2HSV2 U25926 ( .A1(n24045), .A2(n24221), .ZN(n23557) );
  INHSV2 U25927 ( .I(\pe7/got [2]), .ZN(n25308) );
  NOR2HSV2 U25928 ( .A1(n25340), .A2(n25308), .ZN(n23556) );
  XNOR3HSV2 U25929 ( .A1(n23558), .A2(n23557), .A3(n23556), .ZN(n23559) );
  NAND2HSV2 U25930 ( .A1(n28420), .A2(\pe8/got [12]), .ZN(n23604) );
  NAND2HSV2 U25931 ( .A1(n25525), .A2(n28618), .ZN(n23602) );
  CLKNAND2HSV1 U25932 ( .A1(n23757), .A2(\pe8/got [10]), .ZN(n23600) );
  NAND2HSV2 U25933 ( .A1(n25185), .A2(\pe8/got [9]), .ZN(n23598) );
  NAND2HSV0 U25934 ( .A1(n25186), .A2(\pe8/got [6]), .ZN(n23592) );
  CLKNAND2HSV0 U25935 ( .A1(n28616), .A2(\pe8/got [5]), .ZN(n23590) );
  NOR2HSV1 U25936 ( .A1(n25351), .A2(n22230), .ZN(n23588) );
  NAND2HSV0 U25937 ( .A1(n28462), .A2(\pe8/got [2]), .ZN(n23584) );
  INAND2HSV0 U25938 ( .A1(n23642), .B1(n26230), .ZN(n23582) );
  XOR2HSV0 U25939 ( .A1(n23565), .A2(n23564), .Z(n23580) );
  NAND2HSV0 U25940 ( .A1(\pe8/aot [9]), .A2(\pe8/bq[4] ), .ZN(n23567) );
  NAND2HSV0 U25941 ( .A1(\pe8/aot [8]), .A2(\pe8/bq[5] ), .ZN(n23566) );
  XOR2HSV0 U25942 ( .A1(n23567), .A2(n23566), .Z(n23571) );
  NAND2HSV0 U25943 ( .A1(\pe8/aot [1]), .A2(\pe8/bq[12] ), .ZN(n23569) );
  NAND2HSV0 U25944 ( .A1(\pe8/aot [2]), .A2(\pe8/bq[11] ), .ZN(n23568) );
  XOR2HSV0 U25945 ( .A1(n23569), .A2(n23568), .Z(n23570) );
  XNOR2HSV1 U25946 ( .A1(n23571), .A2(n23570), .ZN(n23579) );
  NAND2HSV0 U25947 ( .A1(\pe8/aot [3]), .A2(\pe8/bq[10] ), .ZN(n23573) );
  NAND2HSV0 U25948 ( .A1(\pe8/aot [4]), .A2(\pe8/bq[9] ), .ZN(n23572) );
  XOR2HSV0 U25949 ( .A1(n23573), .A2(n23572), .Z(n23577) );
  NAND2HSV0 U25950 ( .A1(\pe8/aot [7]), .A2(\pe8/bq[6] ), .ZN(n23575) );
  NAND2HSV0 U25951 ( .A1(\pe8/aot [12]), .A2(\pe8/bq[1] ), .ZN(n23574) );
  XOR2HSV0 U25952 ( .A1(n23575), .A2(n23574), .Z(n23576) );
  XOR2HSV0 U25953 ( .A1(n23577), .A2(n23576), .Z(n23578) );
  XOR3HSV2 U25954 ( .A1(n23580), .A2(n23579), .A3(n23578), .Z(n23581) );
  XNOR2HSV1 U25955 ( .A1(n23582), .A2(n23581), .ZN(n23583) );
  XNOR2HSV1 U25956 ( .A1(n23584), .A2(n23583), .ZN(n23586) );
  XNOR2HSV1 U25957 ( .A1(n23586), .A2(n23585), .ZN(n23587) );
  XNOR2HSV1 U25958 ( .A1(n23588), .A2(n23587), .ZN(n23589) );
  XNOR2HSV1 U25959 ( .A1(n23590), .A2(n23589), .ZN(n23591) );
  XOR2HSV0 U25960 ( .A1(n23592), .A2(n23591), .Z(n23594) );
  NAND2HSV0 U25961 ( .A1(n14060), .A2(n28457), .ZN(n23593) );
  XOR2HSV0 U25962 ( .A1(n23594), .A2(n23593), .Z(n23596) );
  NAND2HSV0 U25963 ( .A1(n25204), .A2(\pe8/got [8]), .ZN(n23595) );
  XNOR2HSV1 U25964 ( .A1(n23604), .A2(n23603), .ZN(\pe8/poht [4]) );
  CLKNAND2HSV1 U25965 ( .A1(n28420), .A2(n28695), .ZN(n23663) );
  NAND2HSV2 U25966 ( .A1(n25525), .A2(n25602), .ZN(n23661) );
  CLKNAND2HSV1 U25967 ( .A1(n23757), .A2(n22136), .ZN(n23659) );
  NAND2HSV2 U25968 ( .A1(n25185), .A2(\pe8/got [12]), .ZN(n23657) );
  CLKNAND2HSV0 U25969 ( .A1(n25186), .A2(n23721), .ZN(n23650) );
  CLKNAND2HSV0 U25970 ( .A1(n22140), .A2(n23605), .ZN(n23649) );
  NOR2HSV1 U25971 ( .A1(n25528), .A2(n23869), .ZN(n23648) );
  NAND2HSV0 U25972 ( .A1(\pe8/got [2]), .A2(n28788), .ZN(n23641) );
  NOR2HSV0 U25973 ( .A1(n25557), .A2(n23606), .ZN(n23608) );
  AOI22HSV0 U25974 ( .A1(\pe8/bq[1] ), .A2(n28641), .B1(\pe8/aot [13]), .B2(
        \pe8/bq[3] ), .ZN(n23607) );
  NOR2HSV2 U25975 ( .A1(n23608), .A2(n23607), .ZN(n23613) );
  NAND2HSV0 U25976 ( .A1(\pe8/aot [3]), .A2(\pe8/bq[8] ), .ZN(n23730) );
  NOR2HSV0 U25977 ( .A1(n23609), .A2(n23730), .ZN(n23611) );
  AOI22HSV0 U25978 ( .A1(\pe8/aot [8]), .A2(\pe8/bq[8] ), .B1(n25565), .B2(
        \pe8/aot [3]), .ZN(n23610) );
  NOR2HSV2 U25979 ( .A1(n23611), .A2(n23610), .ZN(n23612) );
  XNOR2HSV1 U25980 ( .A1(n23613), .A2(n23612), .ZN(n23620) );
  NAND2HSV0 U25981 ( .A1(\pe8/aot [11]), .A2(\pe8/bq[5] ), .ZN(n23617) );
  NOR2HSV0 U25982 ( .A1(n23615), .A2(n23614), .ZN(n23616) );
  AOI21HSV0 U25983 ( .A1(n23727), .A2(n23617), .B(n23616), .ZN(n23618) );
  XNOR2HSV1 U25984 ( .A1(n23618), .A2(n25558), .ZN(n23619) );
  XNOR2HSV1 U25985 ( .A1(n23620), .A2(n23619), .ZN(n23638) );
  NOR2HSV1 U25986 ( .A1(n27225), .A2(n25530), .ZN(n23637) );
  NAND2HSV0 U25987 ( .A1(\pe8/aot [5]), .A2(\pe8/bq[11] ), .ZN(n23622) );
  NAND2HSV0 U25988 ( .A1(\pe8/aot [7]), .A2(\pe8/bq[9] ), .ZN(n23621) );
  XOR2HSV0 U25989 ( .A1(n23622), .A2(n23621), .Z(n23626) );
  NAND2HSV0 U25990 ( .A1(\pe8/aot [4]), .A2(\pe8/bq[12] ), .ZN(n23624) );
  NAND2HSV0 U25991 ( .A1(\pe8/aot [6]), .A2(\pe8/bq[10] ), .ZN(n23623) );
  XOR2HSV0 U25992 ( .A1(n23624), .A2(n23623), .Z(n23625) );
  XOR2HSV0 U25993 ( .A1(n23626), .A2(n23625), .Z(n23635) );
  NAND2HSV0 U25994 ( .A1(\pe8/aot [1]), .A2(n25532), .ZN(n23629) );
  NAND2HSV0 U25995 ( .A1(n23627), .A2(\pe8/aot [2]), .ZN(n23628) );
  XOR2HSV0 U25996 ( .A1(n23629), .A2(n23628), .Z(n23633) );
  NAND2HSV0 U25997 ( .A1(\pe8/aot [12]), .A2(\pe8/bq[4] ), .ZN(n23631) );
  NAND2HSV0 U25998 ( .A1(\pe8/aot [10]), .A2(\pe8/bq[6] ), .ZN(n23630) );
  XOR2HSV0 U25999 ( .A1(n23631), .A2(n23630), .Z(n23632) );
  XOR2HSV0 U26000 ( .A1(n23633), .A2(n23632), .Z(n23634) );
  XOR2HSV0 U26001 ( .A1(n23635), .A2(n23634), .Z(n23636) );
  XOR3HSV2 U26002 ( .A1(n23638), .A2(n23637), .A3(n23636), .Z(n23640) );
  NAND2HSV0 U26003 ( .A1(n25578), .A2(\pe8/got [3]), .ZN(n23639) );
  XOR3HSV2 U26004 ( .A1(n23641), .A2(n23640), .A3(n23639), .Z(n23644) );
  INAND2HSV2 U26005 ( .A1(n23642), .B1(n25203), .ZN(n23643) );
  XOR2HSV0 U26006 ( .A1(n23644), .A2(n23643), .Z(n23647) );
  NAND2HSV0 U26007 ( .A1(n12007), .A2(\pe8/got [5]), .ZN(n23645) );
  NAND2HSV0 U26008 ( .A1(\pe8/got [10]), .A2(n14059), .ZN(n23651) );
  XOR2HSV0 U26009 ( .A1(n23652), .A2(n23651), .Z(n23655) );
  NAND2HSV0 U26010 ( .A1(n25204), .A2(n23653), .ZN(n23654) );
  XNOR2HSV1 U26011 ( .A1(n23655), .A2(n23654), .ZN(n23656) );
  XNOR2HSV1 U26012 ( .A1(n23663), .A2(n23662), .ZN(\pe8/poht [1]) );
  CLKNAND2HSV3 U26013 ( .A1(n23665), .A2(n23668), .ZN(n23803) );
  NOR2HSV4 U26014 ( .A1(n23668), .A2(n23667), .ZN(n23805) );
  INHSV4 U26015 ( .I(n23669), .ZN(n23804) );
  CLKNAND2HSV2 U26016 ( .A1(n23805), .A2(n23804), .ZN(n23677) );
  NAND2HSV4 U26017 ( .A1(n23676), .A2(n23677), .ZN(n28661) );
  INHSV4 U26018 ( .I(n23670), .ZN(n26760) );
  INHSV2 U26019 ( .I(n26349), .ZN(n26681) );
  CLKNHSV1 U26020 ( .I(\pe3/got [2]), .ZN(n26713) );
  NOR2HSV2 U26021 ( .A1(n26681), .A2(n26713), .ZN(n23675) );
  INHSV2 U26022 ( .I(n24516), .ZN(n28584) );
  NAND2HSV0 U26023 ( .A1(\pe3/aot [1]), .A2(\pe3/bq[5] ), .ZN(n23672) );
  NAND2HSV0 U26024 ( .A1(\pe3/aot [3]), .A2(\pe3/bq[3] ), .ZN(n23671) );
  XOR2HSV0 U26025 ( .A1(n23672), .A2(n23671), .Z(n23673) );
  CLKNAND2HSV0 U26026 ( .A1(\pe3/bq[2] ), .A2(\pe3/aot [4]), .ZN(n26683) );
  CLKNAND2HSV1 U26027 ( .A1(n28652), .A2(\pe3/got [1]), .ZN(n23680) );
  CLKNAND2HSV0 U26028 ( .A1(\pe3/aot [3]), .A2(\pe3/bq[1] ), .ZN(n24584) );
  NAND2HSV0 U26029 ( .A1(\pe3/aot [2]), .A2(\pe3/bq[2] ), .ZN(n23678) );
  XOR2HSV0 U26030 ( .A1(n24584), .A2(n23678), .Z(n23679) );
  CLKNAND2HSV1 U26031 ( .A1(\pe3/bq[3] ), .A2(\pe3/aot [1]), .ZN(n26309) );
  INHSV2 U26032 ( .I(n23681), .ZN(n23993) );
  INHSV4 U26033 ( .I(n23993), .ZN(n28461) );
  INHSV2 U26034 ( .I(n26349), .ZN(n26602) );
  NOR2HSV2 U26035 ( .A1(n26602), .A2(n23682), .ZN(n23700) );
  NAND2HSV0 U26036 ( .A1(n28438), .A2(\pe3/got [4]), .ZN(n23694) );
  NAND2HSV0 U26037 ( .A1(n23327), .A2(n26751), .ZN(n23692) );
  NAND2HSV0 U26038 ( .A1(\pe3/bq[7] ), .A2(\pe3/aot [4]), .ZN(n26610) );
  NAND2HSV0 U26039 ( .A1(\pe3/aot [10]), .A2(\pe3/bq[1] ), .ZN(n23685) );
  NAND2HSV0 U26040 ( .A1(\pe3/aot [7]), .A2(\pe3/bq[4] ), .ZN(n23684) );
  NOR2HSV0 U26041 ( .A1(n23686), .A2(n26309), .ZN(n23688) );
  AOI22HSV0 U26042 ( .A1(\pe3/aot [8]), .A2(\pe3/bq[3] ), .B1(\pe3/bq[10] ), 
        .B2(\pe3/aot [1]), .ZN(n23687) );
  NAND2HSV0 U26043 ( .A1(\pe3/aot [2]), .A2(\pe3/bq[9] ), .ZN(n23690) );
  NAND2HSV0 U26044 ( .A1(\pe3/aot [5]), .A2(\pe3/bq[6] ), .ZN(n23689) );
  XNOR2HSV1 U26045 ( .A1(n23692), .A2(n23691), .ZN(n23693) );
  XOR2HSV0 U26046 ( .A1(n23694), .A2(n23693), .Z(n23696) );
  NAND2HSV0 U26047 ( .A1(n26752), .A2(\pe3/got [5]), .ZN(n23695) );
  XOR2HSV0 U26048 ( .A1(n23696), .A2(n23695), .Z(n23698) );
  NAND2HSV0 U26049 ( .A1(\pe3/got [6]), .A2(n28584), .ZN(n23697) );
  XOR2HSV0 U26050 ( .A1(n23698), .A2(n23697), .Z(n23699) );
  NAND2HSV2 U26051 ( .A1(n28467), .A2(n28608), .ZN(n23708) );
  NAND2HSV0 U26052 ( .A1(\pe6/aot [3]), .A2(\pe6/bq[2] ), .ZN(n23702) );
  NAND2HSV0 U26053 ( .A1(\pe6/aot [1]), .A2(\pe6/bq[4] ), .ZN(n23701) );
  XOR2HSV0 U26054 ( .A1(n23702), .A2(n23701), .Z(n23706) );
  NAND2HSV0 U26055 ( .A1(\pe6/aot [2]), .A2(\pe6/bq[3] ), .ZN(n23703) );
  XOR2HSV0 U26056 ( .A1(n23704), .A2(n23703), .Z(n23705) );
  XOR2HSV0 U26057 ( .A1(n23706), .A2(n23705), .Z(n23707) );
  XNOR2HSV1 U26058 ( .A1(n23708), .A2(n23707), .ZN(n23709) );
  XOR2HSV0 U26059 ( .A1(n23709), .A2(n23710), .Z(n23711) );
  BUFHSV4 U26060 ( .I(n23720), .Z(n28347) );
  NAND2HSV0 U26061 ( .A1(n28698), .A2(n14060), .ZN(n23755) );
  CLKNAND2HSV0 U26062 ( .A1(n28631), .A2(n25577), .ZN(n23749) );
  NAND2HSV0 U26063 ( .A1(n28616), .A2(\pe8/got [3]), .ZN(n23747) );
  NOR2HSV1 U26064 ( .A1(n25528), .A2(n28650), .ZN(n23745) );
  NOR2HSV2 U26065 ( .A1(n25543), .A2(n23722), .ZN(n23776) );
  CLKNHSV0 U26066 ( .I(\pe8/aot [7]), .ZN(n23724) );
  NOR2HSV0 U26067 ( .A1(n23724), .A2(n23723), .ZN(n25553) );
  AOI22HSV0 U26068 ( .A1(\pe8/aot [7]), .A2(\pe8/bq[4] ), .B1(\pe8/bq[10] ), 
        .B2(\pe8/aot [1]), .ZN(n23725) );
  AOI21HSV0 U26069 ( .A1(n23776), .A2(n25553), .B(n23725), .ZN(n23729) );
  XOR2HSV0 U26070 ( .A1(n23729), .A2(n23728), .Z(n23733) );
  XOR2HSV0 U26071 ( .A1(n23731), .A2(n23730), .Z(n23732) );
  XNOR2HSV1 U26072 ( .A1(n23733), .A2(n23732), .ZN(n23741) );
  NAND2HSV0 U26073 ( .A1(\pe8/aot [10]), .A2(\pe8/bq[1] ), .ZN(n23735) );
  NAND2HSV0 U26074 ( .A1(\pe8/aot [2]), .A2(\pe8/bq[9] ), .ZN(n23734) );
  XOR2HSV0 U26075 ( .A1(n23735), .A2(n23734), .Z(n23739) );
  NAND2HSV0 U26076 ( .A1(\pe8/aot [5]), .A2(\pe8/bq[6] ), .ZN(n23737) );
  NAND2HSV0 U26077 ( .A1(\pe8/aot [8]), .A2(\pe8/bq[3] ), .ZN(n23736) );
  XOR2HSV0 U26078 ( .A1(n23737), .A2(n23736), .Z(n23738) );
  XOR2HSV0 U26079 ( .A1(n23739), .A2(n23738), .Z(n23740) );
  XOR2HSV0 U26080 ( .A1(n23741), .A2(n23740), .Z(n23742) );
  XNOR2HSV1 U26081 ( .A1(n23743), .A2(n23742), .ZN(n23744) );
  XOR2HSV0 U26082 ( .A1(n23745), .A2(n23744), .Z(n23746) );
  XNOR2HSV1 U26083 ( .A1(n23747), .A2(n23746), .ZN(n23748) );
  XOR2HSV0 U26084 ( .A1(n23749), .A2(n23748), .Z(n23751) );
  NAND2HSV0 U26085 ( .A1(n14059), .A2(\pe8/got [5]), .ZN(n23750) );
  XOR2HSV0 U26086 ( .A1(n23751), .A2(n23750), .Z(n23753) );
  NAND2HSV0 U26087 ( .A1(n25204), .A2(\pe8/got [6]), .ZN(n23752) );
  XOR2HSV0 U26088 ( .A1(n23753), .A2(n23752), .Z(n23754) );
  XNOR2HSV1 U26089 ( .A1(n23755), .A2(n23754), .ZN(n23756) );
  NAND2HSV0 U26090 ( .A1(n25185), .A2(\pe8/got [3]), .ZN(n23773) );
  NAND2HSV0 U26091 ( .A1(n28457), .A2(n26230), .ZN(n23769) );
  NAND2HSV0 U26092 ( .A1(\pe8/aot [1]), .A2(\pe8/bq[6] ), .ZN(n23759) );
  NAND2HSV0 U26093 ( .A1(\pe8/aot [6]), .A2(\pe8/bq[1] ), .ZN(n23758) );
  XOR2HSV0 U26094 ( .A1(n23759), .A2(n23758), .Z(n23764) );
  NOR2HSV0 U26095 ( .A1(n23760), .A2(n23847), .ZN(n23762) );
  NAND2HSV0 U26096 ( .A1(\pe8/aot [4]), .A2(\pe8/bq[3] ), .ZN(n23761) );
  XOR2HSV0 U26097 ( .A1(n23762), .A2(n23761), .Z(n23763) );
  XNOR2HSV1 U26098 ( .A1(n23764), .A2(n23763), .ZN(n23767) );
  NAND2HSV0 U26099 ( .A1(\pe8/aot [3]), .A2(\pe8/bq[4] ), .ZN(n23849) );
  XOR2HSV0 U26100 ( .A1(n23849), .A2(n23765), .Z(n23766) );
  XNOR2HSV1 U26101 ( .A1(n23767), .A2(n23766), .ZN(n23768) );
  XNOR2HSV1 U26102 ( .A1(n23769), .A2(n23768), .ZN(n23771) );
  NAND2HSV0 U26103 ( .A1(n28706), .A2(\pe8/got [2]), .ZN(n23770) );
  XOR2HSV0 U26104 ( .A1(n23771), .A2(n23770), .Z(n23772) );
  NAND2HSV0 U26105 ( .A1(n26229), .A2(n25577), .ZN(n23788) );
  NAND2HSV0 U26106 ( .A1(n28698), .A2(n26230), .ZN(n23782) );
  NAND2HSV0 U26107 ( .A1(\pe8/aot [4]), .A2(\pe8/bq[1] ), .ZN(n23775) );
  XOR2HSV0 U26108 ( .A1(n23776), .A2(n23775), .Z(n23780) );
  CLKNHSV0 U26109 ( .I(\pe8/aot [3]), .ZN(n23848) );
  NOR2HSV1 U26110 ( .A1(n23848), .A2(n25555), .ZN(n23778) );
  NAND2HSV0 U26111 ( .A1(\pe8/aot [2]), .A2(\pe8/bq[3] ), .ZN(n23777) );
  XOR2HSV0 U26112 ( .A1(n23778), .A2(n23777), .Z(n23779) );
  XOR2HSV0 U26113 ( .A1(n23780), .A2(n23779), .Z(n23781) );
  XOR2HSV0 U26114 ( .A1(n23782), .A2(n23781), .Z(n23784) );
  NAND2HSV0 U26115 ( .A1(n23846), .A2(\pe8/got [2]), .ZN(n23783) );
  XNOR2HSV1 U26116 ( .A1(n23784), .A2(n23783), .ZN(n23785) );
  XNOR2HSV1 U26117 ( .A1(n23786), .A2(n23785), .ZN(n23787) );
  XOR2HSV0 U26118 ( .A1(n23788), .A2(n23787), .Z(\pe8/poht [12]) );
  CLKNHSV0 U26119 ( .I(n28547), .ZN(n23790) );
  CLKNHSV0 U26120 ( .I(n23790), .ZN(n28561) );
  CLKNHSV0 U26121 ( .I(n23799), .ZN(n28458) );
  CLKNHSV0 U26122 ( .I(n23798), .ZN(n28459) );
  CLKNHSV0 U26123 ( .I(n23790), .ZN(n28476) );
  CLKNHSV0 U26124 ( .I(n23798), .ZN(n28477) );
  CLKNHSV0 U26125 ( .I(n23796), .ZN(n28552) );
  CLKNHSV0 U26126 ( .I(n28552), .ZN(n23793) );
  CLKNHSV0 U26127 ( .I(n28921), .ZN(n28522) );
  CLKNHSV0 U26128 ( .I(n28522), .ZN(n24310) );
  CLKNHSV0 U26129 ( .I(n24310), .ZN(n28482) );
  CLKNHSV0 U26130 ( .I(n24310), .ZN(n28483) );
  CLKNHSV0 U26131 ( .I(n28921), .ZN(n28484) );
  CLKNHSV0 U26132 ( .I(n23799), .ZN(n28486) );
  CLKNHSV0 U26133 ( .I(n24308), .ZN(n28487) );
  CLKNHSV0 U26134 ( .I(n23790), .ZN(n28488) );
  CLKNHSV0 U26135 ( .I(n23790), .ZN(n28489) );
  CLKNHSV0 U26136 ( .I(n24308), .ZN(n28490) );
  CLKNHSV0 U26137 ( .I(n23790), .ZN(n28491) );
  CLKNHSV0 U26138 ( .I(n24308), .ZN(n28492) );
  CLKNHSV0 U26139 ( .I(n23793), .ZN(n28493) );
  CLKNHSV0 U26140 ( .I(n24310), .ZN(n28511) );
  CLKNHSV0 U26141 ( .I(n23795), .ZN(n28494) );
  CLKNHSV0 U26142 ( .I(n23799), .ZN(n28495) );
  CLKNHSV0 U26143 ( .I(n23790), .ZN(n28496) );
  CLKNHSV0 U26144 ( .I(n23790), .ZN(n28497) );
  CLKNHSV0 U26145 ( .I(n24308), .ZN(n28498) );
  CLKNHSV0 U26146 ( .I(n23796), .ZN(n28499) );
  CLKNHSV0 U26147 ( .I(n23790), .ZN(n28500) );
  CLKNHSV0 U26148 ( .I(n28595), .ZN(n23792) );
  CLKNHSV0 U26149 ( .I(n23790), .ZN(n28501) );
  CLKNHSV0 U26150 ( .I(n23796), .ZN(n28502) );
  CLKNHSV0 U26151 ( .I(n23801), .ZN(n28503) );
  CLKNHSV0 U26152 ( .I(n28921), .ZN(n28504) );
  CLKNHSV0 U26153 ( .I(n23801), .ZN(n28505) );
  CLKNHSV0 U26154 ( .I(n24309), .ZN(n28506) );
  CLKNHSV0 U26155 ( .I(n23797), .ZN(n28507) );
  CLKNHSV0 U26156 ( .I(n23800), .ZN(n28508) );
  CLKNHSV0 U26157 ( .I(n23800), .ZN(n28509) );
  CLKNHSV0 U26158 ( .I(n23795), .ZN(n28510) );
  CLKNHSV0 U26159 ( .I(n23791), .ZN(n28528) );
  CLKNHSV0 U26160 ( .I(n28564), .ZN(n23794) );
  CLKNHSV0 U26161 ( .I(n23796), .ZN(n28512) );
  CLKNHSV0 U26162 ( .I(n23794), .ZN(n28513) );
  CLKNHSV0 U26163 ( .I(n23795), .ZN(n28514) );
  CLKNHSV0 U26164 ( .I(n23795), .ZN(n28515) );
  CLKNHSV0 U26165 ( .I(n28921), .ZN(n28516) );
  CLKNHSV0 U26166 ( .I(n28921), .ZN(n28517) );
  CLKNHSV0 U26167 ( .I(n24308), .ZN(n28518) );
  CLKNHSV0 U26168 ( .I(n23799), .ZN(n28519) );
  CLKNHSV0 U26169 ( .I(n28500), .ZN(n23798) );
  CLKNHSV0 U26170 ( .I(n23798), .ZN(n28520) );
  CLKNHSV0 U26171 ( .I(n23800), .ZN(n28521) );
  CLKNHSV0 U26172 ( .I(n28921), .ZN(n28525) );
  CLKNHSV0 U26173 ( .I(n23798), .ZN(n28527) );
  CLKNHSV0 U26174 ( .I(n23791), .ZN(n28529) );
  CLKNHSV0 U26175 ( .I(n24310), .ZN(n28531) );
  CLKNHSV0 U26176 ( .I(n23795), .ZN(n28532) );
  CLKNHSV0 U26177 ( .I(n23795), .ZN(n28533) );
  CLKNHSV0 U26178 ( .I(n23796), .ZN(n28534) );
  CLKNHSV0 U26179 ( .I(n24308), .ZN(n28535) );
  CLKNHSV0 U26180 ( .I(n28921), .ZN(n28536) );
  CLKNHSV0 U26181 ( .I(n23799), .ZN(n28537) );
  CLKNHSV0 U26182 ( .I(n23795), .ZN(n28538) );
  CLKNHSV0 U26183 ( .I(n23801), .ZN(n28539) );
  CLKNHSV0 U26184 ( .I(n23798), .ZN(n28540) );
  CLKNHSV0 U26185 ( .I(n23798), .ZN(n28541) );
  CLKNHSV0 U26186 ( .I(n23798), .ZN(n28543) );
  CLKNHSV0 U26187 ( .I(n23800), .ZN(n28544) );
  CLKNHSV0 U26188 ( .I(n23800), .ZN(n28545) );
  CLKNHSV0 U26189 ( .I(n23791), .ZN(n28546) );
  CLKNHSV0 U26190 ( .I(n23791), .ZN(n28547) );
  CLKNHSV0 U26191 ( .I(n24310), .ZN(n28548) );
  CLKNHSV0 U26192 ( .I(n23793), .ZN(n28549) );
  CLKNHSV0 U26193 ( .I(n23796), .ZN(n28550) );
  CLKNHSV0 U26194 ( .I(n23793), .ZN(n28551) );
  CLKNHSV0 U26195 ( .I(n23801), .ZN(n28554) );
  CLKNHSV0 U26196 ( .I(n23801), .ZN(n28555) );
  CLKNHSV0 U26197 ( .I(n23795), .ZN(n28556) );
  CLKNHSV0 U26198 ( .I(n23795), .ZN(n28557) );
  CLKNHSV0 U26199 ( .I(n23796), .ZN(n28558) );
  CLKNHSV0 U26200 ( .I(n23795), .ZN(n28559) );
  CLKNHSV0 U26201 ( .I(n23799), .ZN(n28560) );
  CLKNHSV0 U26202 ( .I(n24308), .ZN(n28562) );
  CLKNHSV0 U26203 ( .I(n23796), .ZN(n28563) );
  CLKNHSV0 U26204 ( .I(n28921), .ZN(n28564) );
  CLKNHSV0 U26205 ( .I(n23792), .ZN(n28566) );
  CLKNHSV0 U26206 ( .I(n24310), .ZN(n28567) );
  CLKNHSV0 U26207 ( .I(n23799), .ZN(n28568) );
  CLKNHSV0 U26208 ( .I(n23800), .ZN(n28569) );
  CLKNHSV0 U26209 ( .I(n23798), .ZN(n28570) );
  CLKNHSV0 U26210 ( .I(n23800), .ZN(n28571) );
  CLKNHSV0 U26211 ( .I(n23800), .ZN(n28572) );
  CLKNHSV0 U26212 ( .I(n24310), .ZN(n28573) );
  CLKNHSV0 U26213 ( .I(n23801), .ZN(n28574) );
  CLKNHSV0 U26214 ( .I(n23791), .ZN(n28575) );
  CLKNHSV0 U26215 ( .I(n23790), .ZN(n28576) );
  CLKNHSV0 U26216 ( .I(n28921), .ZN(n28577) );
  NAND2HSV0 U26217 ( .A1(n26600), .A2(\pe3/got [4]), .ZN(n23821) );
  NAND2HSV2 U26218 ( .A1(n24522), .A2(n26751), .ZN(n23819) );
  CLKNHSV1 U26219 ( .I(\pe3/got [1]), .ZN(n26624) );
  NAND2HSV0 U26220 ( .A1(\pe3/aot [1]), .A2(\pe3/bq[4] ), .ZN(n23807) );
  NAND2HSV0 U26221 ( .A1(\pe3/aot [4]), .A2(\pe3/bq[1] ), .ZN(n23806) );
  XOR2HSV0 U26222 ( .A1(n23807), .A2(n23806), .Z(n23811) );
  NAND2HSV0 U26223 ( .A1(\pe3/aot [3]), .A2(\pe3/bq[2] ), .ZN(n23809) );
  NAND2HSV0 U26224 ( .A1(\pe3/aot [2]), .A2(\pe3/bq[3] ), .ZN(n23808) );
  XOR2HSV0 U26225 ( .A1(n23809), .A2(n23808), .Z(n23810) );
  XOR2HSV0 U26226 ( .A1(n23811), .A2(n23810), .Z(n23812) );
  CLKXOR2HSV4 U26227 ( .A1(n23813), .A2(n23812), .Z(n23817) );
  CLKNAND2HSV3 U26228 ( .A1(n23815), .A2(n23814), .ZN(n26759) );
  NAND2HSV0 U26229 ( .A1(n26759), .A2(\pe3/got [2]), .ZN(n23816) );
  XOR2HSV2 U26230 ( .A1(n23817), .A2(n23816), .Z(n23818) );
  XNOR2HSV2 U26231 ( .A1(n23819), .A2(n23818), .ZN(n23820) );
  XOR2HSV0 U26232 ( .A1(n23821), .A2(n23820), .Z(\pe3/poht [12]) );
  MUX2HSV2 U26233 ( .I0(bo9[14]), .I1(n23822), .S(n27093), .Z(n28780) );
  INHSV4 U26234 ( .I(n24220), .ZN(n24277) );
  CLKNAND2HSV0 U26235 ( .A1(n28665), .A2(\pe7/got [2]), .ZN(n23836) );
  NAND2HSV0 U26236 ( .A1(n28656), .A2(\pe7/got [1]), .ZN(n23834) );
  NAND2HSV0 U26237 ( .A1(\pe7/aot [3]), .A2(\pe7/bq[4] ), .ZN(n23824) );
  NAND2HSV0 U26238 ( .A1(\pe7/aot [5]), .A2(\pe7/bq[2] ), .ZN(n23823) );
  XOR2HSV0 U26239 ( .A1(n23824), .A2(n23823), .Z(n23828) );
  NAND2HSV0 U26240 ( .A1(\pe7/aot [2]), .A2(\pe7/bq[5] ), .ZN(n23826) );
  NAND2HSV0 U26241 ( .A1(\pe7/aot [1]), .A2(\pe7/bq[6] ), .ZN(n23825) );
  XOR2HSV0 U26242 ( .A1(n23826), .A2(n23825), .Z(n23827) );
  XOR2HSV0 U26243 ( .A1(n23828), .A2(n23827), .Z(n23832) );
  NAND2HSV0 U26244 ( .A1(\pe7/aot [6]), .A2(\pe7/bq[1] ), .ZN(n23830) );
  NAND2HSV0 U26245 ( .A1(\pe7/aot [4]), .A2(\pe7/bq[3] ), .ZN(n23829) );
  XOR2HSV0 U26246 ( .A1(n23830), .A2(n23829), .Z(n23831) );
  XNOR2HSV1 U26247 ( .A1(n23832), .A2(n23831), .ZN(n23833) );
  XNOR2HSV1 U26248 ( .A1(n23834), .A2(n23833), .ZN(n23835) );
  XOR2HSV0 U26249 ( .A1(n23836), .A2(n23835), .Z(n23838) );
  NAND2HSV0 U26250 ( .A1(n25335), .A2(\pe7/got [3]), .ZN(n23837) );
  XOR2HSV0 U26251 ( .A1(n23838), .A2(n23837), .Z(n23842) );
  NOR2HSV2 U26252 ( .A1(n24045), .A2(n23839), .ZN(n23841) );
  NAND2HSV0 U26253 ( .A1(n25408), .A2(n25375), .ZN(n23840) );
  XNOR3HSV2 U26254 ( .A1(n23842), .A2(n23841), .A3(n23840), .ZN(n23843) );
  NAND2HSV0 U26255 ( .A1(n28621), .A2(n28610), .ZN(n23845) );
  XOR2HSV0 U26256 ( .A1(n23845), .A2(n23844), .Z(n28960) );
  NAND2HSV0 U26257 ( .A1(n28631), .A2(n26230), .ZN(n23860) );
  NOR2HSV0 U26258 ( .A1(n23848), .A2(n23847), .ZN(n23850) );
  NAND2HSV0 U26259 ( .A1(\pe8/aot [4]), .A2(\pe8/bq[5] ), .ZN(n25190) );
  OAI22HSV1 U26260 ( .A1(n23851), .A2(n23850), .B1(n23849), .B2(n25190), .ZN(
        n23858) );
  NAND2HSV0 U26261 ( .A1(\pe8/aot [5]), .A2(\pe8/bq[3] ), .ZN(n23853) );
  NAND2HSV0 U26262 ( .A1(\pe8/aot [2]), .A2(\pe8/bq[6] ), .ZN(n23852) );
  XOR2HSV0 U26263 ( .A1(n23853), .A2(n23852), .Z(n23857) );
  NAND2HSV0 U26264 ( .A1(\pe8/aot [7]), .A2(\pe8/bq[1] ), .ZN(n25196) );
  NAND2HSV0 U26265 ( .A1(\pe8/aot [6]), .A2(\pe8/bq[2] ), .ZN(n23854) );
  XOR2HSV0 U26266 ( .A1(n25196), .A2(n23854), .Z(n23855) );
  XOR4HSV1 U26267 ( .A1(n23858), .A2(n23857), .A3(n23856), .A4(n23855), .Z(
        n23859) );
  XOR2HSV0 U26268 ( .A1(n23860), .A2(n23859), .Z(n23862) );
  NAND2HSV0 U26269 ( .A1(n28457), .A2(\pe8/got [2]), .ZN(n23861) );
  XOR2HSV0 U26270 ( .A1(n23862), .A2(n23861), .Z(n23864) );
  NAND2HSV0 U26271 ( .A1(n25204), .A2(\pe8/got [3]), .ZN(n23863) );
  NAND2HSV0 U26272 ( .A1(n28698), .A2(n25203), .ZN(n23865) );
  XNOR2HSV0 U26273 ( .A1(n23867), .A2(n23866), .ZN(n23868) );
  INHSV2 U26274 ( .I(n23871), .ZN(n25376) );
  NAND2HSV0 U26275 ( .A1(n14067), .A2(n25272), .ZN(n23900) );
  NAND2HSV0 U26276 ( .A1(\pe7/got [3]), .A2(n28466), .ZN(n23899) );
  NAND2HSV0 U26277 ( .A1(n25318), .A2(\pe7/got [2]), .ZN(n23897) );
  NAND2HSV0 U26278 ( .A1(n11936), .A2(\pe7/got [1]), .ZN(n23895) );
  NAND2HSV0 U26279 ( .A1(\pe7/aot [6]), .A2(\pe7/bq[7] ), .ZN(n23873) );
  NAND2HSV0 U26280 ( .A1(\pe7/aot [4]), .A2(\pe7/bq[9] ), .ZN(n23872) );
  XOR2HSV0 U26281 ( .A1(n23873), .A2(n23872), .Z(n23877) );
  NAND2HSV0 U26282 ( .A1(\pe7/aot [3]), .A2(\pe7/bq[10] ), .ZN(n23875) );
  NAND2HSV0 U26283 ( .A1(\pe7/aot [7]), .A2(\pe7/bq[6] ), .ZN(n23874) );
  XOR2HSV0 U26284 ( .A1(n23875), .A2(n23874), .Z(n23876) );
  XOR2HSV0 U26285 ( .A1(n23877), .A2(n23876), .Z(n23885) );
  NAND2HSV0 U26286 ( .A1(\pe7/aot [1]), .A2(\pe7/bq[12] ), .ZN(n23879) );
  NAND2HSV0 U26287 ( .A1(\pe7/aot [2]), .A2(\pe7/bq[11] ), .ZN(n23878) );
  XOR2HSV0 U26288 ( .A1(n23879), .A2(n23878), .Z(n23883) );
  NAND2HSV0 U26289 ( .A1(\pe7/aot [11]), .A2(\pe7/bq[2] ), .ZN(n23881) );
  NAND2HSV0 U26290 ( .A1(\pe7/aot [12]), .A2(\pe7/bq[1] ), .ZN(n23880) );
  XOR2HSV0 U26291 ( .A1(n23881), .A2(n23880), .Z(n23882) );
  XOR2HSV0 U26292 ( .A1(n23883), .A2(n23882), .Z(n23884) );
  XOR2HSV0 U26293 ( .A1(n23885), .A2(n23884), .Z(n23893) );
  NAND2HSV0 U26294 ( .A1(\pe7/aot [8]), .A2(\pe7/bq[5] ), .ZN(n23887) );
  NAND2HSV0 U26295 ( .A1(\pe7/aot [9]), .A2(\pe7/bq[4] ), .ZN(n23886) );
  XOR2HSV0 U26296 ( .A1(n23887), .A2(n23886), .Z(n23891) );
  CLKNHSV0 U26297 ( .I(\pe7/bq[3] ), .ZN(n27098) );
  NOR2HSV0 U26298 ( .A1(n24105), .A2(n27098), .ZN(n23889) );
  NAND2HSV0 U26299 ( .A1(\pe7/aot [5]), .A2(\pe7/bq[8] ), .ZN(n23888) );
  XOR2HSV0 U26300 ( .A1(n23889), .A2(n23888), .Z(n23890) );
  XOR2HSV0 U26301 ( .A1(n23891), .A2(n23890), .Z(n23892) );
  XNOR2HSV1 U26302 ( .A1(n23893), .A2(n23892), .ZN(n23894) );
  XNOR2HSV1 U26303 ( .A1(n23895), .A2(n23894), .ZN(n23896) );
  XOR2HSV0 U26304 ( .A1(n23897), .A2(n23896), .Z(n23898) );
  CLKNHSV3 U26305 ( .I(n23901), .ZN(n25397) );
  NAND2HSV0 U26306 ( .A1(n25335), .A2(\pe7/got [9]), .ZN(n23902) );
  INHSV4 U26307 ( .I(n23555), .ZN(n24286) );
  NOR2HSV2 U26308 ( .A1(n24286), .A2(n24084), .ZN(n23905) );
  XOR2HSV0 U26309 ( .A1(n23908), .A2(n23907), .Z(\pe7/poht [4]) );
  NAND2HSV0 U26310 ( .A1(n21718), .A2(n20977), .ZN(n23950) );
  NAND2HSV0 U26311 ( .A1(n24341), .A2(n24637), .ZN(n23949) );
  NAND2HSV0 U26312 ( .A1(\pe5/ti_7[10] ), .A2(n24340), .ZN(n23945) );
  CLKNAND2HSV0 U26313 ( .A1(n21523), .A2(\pe5/got [5]), .ZN(n23939) );
  NAND2HSV0 U26314 ( .A1(n28614), .A2(n28640), .ZN(n23932) );
  NAND2HSV0 U26315 ( .A1(\pe5/aot [3]), .A2(\pe5/bq[11] ), .ZN(n23911) );
  NAND2HSV0 U26316 ( .A1(\pe5/aot [2]), .A2(n23909), .ZN(n23910) );
  XOR2HSV0 U26317 ( .A1(n23911), .A2(n23910), .Z(n23930) );
  NAND2HSV0 U26318 ( .A1(\pe5/aot [4]), .A2(\pe5/bq[10] ), .ZN(n23913) );
  NAND2HSV0 U26319 ( .A1(\pe5/aot [9]), .A2(\pe5/bq[5] ), .ZN(n23912) );
  XOR2HSV0 U26320 ( .A1(n23913), .A2(n23912), .Z(n23915) );
  XNOR2HSV1 U26321 ( .A1(n23915), .A2(n23914), .ZN(n23929) );
  NAND2HSV0 U26322 ( .A1(\pe5/aot [13]), .A2(\pe5/bq[3] ), .ZN(n24664) );
  NOR2HSV0 U26323 ( .A1(n24664), .A2(n23916), .ZN(n23918) );
  AOI22HSV0 U26324 ( .A1(n14019), .A2(\pe5/bq[1] ), .B1(\pe5/aot [11]), .B2(
        \pe5/bq[3] ), .ZN(n23917) );
  NOR2HSV2 U26325 ( .A1(n23918), .A2(n23917), .ZN(n23920) );
  XOR2HSV0 U26326 ( .A1(n23920), .A2(n23919), .Z(n23928) );
  NAND2HSV0 U26327 ( .A1(\pe5/aot [1]), .A2(\pe5/bq[13] ), .ZN(n23922) );
  NAND2HSV0 U26328 ( .A1(\pe5/aot [10]), .A2(\pe5/bq[4] ), .ZN(n23921) );
  XOR2HSV0 U26329 ( .A1(n23922), .A2(n23921), .Z(n23926) );
  XOR2HSV0 U26330 ( .A1(n23926), .A2(n23925), .Z(n23927) );
  XOR4HSV1 U26331 ( .A1(n23930), .A2(n23929), .A3(n23928), .A4(n23927), .Z(
        n23931) );
  XNOR2HSV1 U26332 ( .A1(n23932), .A2(n23931), .ZN(n23934) );
  NAND2HSV0 U26333 ( .A1(n24411), .A2(\pe5/got [2]), .ZN(n23933) );
  XOR2HSV0 U26334 ( .A1(n23934), .A2(n23933), .Z(n23937) );
  NOR2HSV0 U26335 ( .A1(n25350), .A2(n24364), .ZN(n23936) );
  NAND2HSV0 U26336 ( .A1(n28478), .A2(n13993), .ZN(n23935) );
  XOR3HSV1 U26337 ( .A1(n23937), .A2(n23936), .A3(n23935), .Z(n23938) );
  XNOR2HSV1 U26338 ( .A1(n23939), .A2(n23938), .ZN(n23943) );
  NOR2HSV2 U26339 ( .A1(n24684), .A2(n23940), .ZN(n23942) );
  OR2HSV1 U26340 ( .A1(n24686), .A2(n24420), .Z(n23941) );
  XOR3HSV2 U26341 ( .A1(n23943), .A2(n23942), .A3(n23941), .Z(n23944) );
  XNOR2HSV1 U26342 ( .A1(n23945), .A2(n23944), .ZN(n23947) );
  NAND2HSV0 U26343 ( .A1(n28803), .A2(n14071), .ZN(n23946) );
  XNOR2HSV1 U26344 ( .A1(n23947), .A2(n23946), .ZN(n23948) );
  NAND2HSV0 U26345 ( .A1(n28700), .A2(\pe1/got [7]), .ZN(n23980) );
  CLKNAND2HSV0 U26346 ( .A1(n27137), .A2(n28434), .ZN(n23978) );
  CLKNHSV0 U26347 ( .I(\pe1/got [5]), .ZN(n25878) );
  NOR2HSV2 U26348 ( .A1(n27002), .A2(n25878), .ZN(n23976) );
  NOR2HSV2 U26349 ( .A1(n26830), .A2(n26852), .ZN(n23974) );
  NAND2HSV0 U26350 ( .A1(n26854), .A2(\pe1/got [3]), .ZN(n23972) );
  NAND2HSV0 U26351 ( .A1(n26541), .A2(\pe1/got [1]), .ZN(n23968) );
  NAND2HSV0 U26352 ( .A1(\pe1/aot [8]), .A2(\pe1/bq[2] ), .ZN(n26863) );
  NAND2HSV2 U26353 ( .A1(\pe1/bq[1] ), .A2(\pe1/aot [1]), .ZN(n26805) );
  INHSV2 U26354 ( .I(\pe1/bq[1] ), .ZN(n27064) );
  NAND2HSV0 U26355 ( .A1(\pe1/bq[9] ), .A2(\pe1/aot [1]), .ZN(n27020) );
  OAI21HSV0 U26356 ( .A1(n27064), .A2(n27158), .B(n27020), .ZN(n23955) );
  OAI21HSV0 U26357 ( .A1(n26487), .A2(n26805), .B(n23955), .ZN(n23958) );
  NAND2HSV0 U26358 ( .A1(\pe1/bq[7] ), .A2(\pe1/aot [3]), .ZN(n26769) );
  NAND2HSV0 U26359 ( .A1(\pe1/aot [6]), .A2(\pe1/bq[4] ), .ZN(n23956) );
  XOR2HSV0 U26360 ( .A1(n26769), .A2(n23956), .Z(n23957) );
  XOR3HSV2 U26361 ( .A1(n26863), .A2(n23958), .A3(n23957), .Z(n23966) );
  NAND2HSV0 U26362 ( .A1(\pe1/aot [2]), .A2(\pe1/bq[8] ), .ZN(n23960) );
  NAND2HSV0 U26363 ( .A1(\pe1/aot [4]), .A2(\pe1/bq[6] ), .ZN(n23959) );
  XOR2HSV0 U26364 ( .A1(n23960), .A2(n23959), .Z(n23964) );
  NOR2HSV0 U26365 ( .A1(n26764), .A2(n27157), .ZN(n23962) );
  NAND2HSV0 U26366 ( .A1(\pe1/aot [5]), .A2(\pe1/bq[5] ), .ZN(n23961) );
  XOR2HSV0 U26367 ( .A1(n23962), .A2(n23961), .Z(n23963) );
  XOR2HSV0 U26368 ( .A1(n23964), .A2(n23963), .Z(n23965) );
  XNOR2HSV1 U26369 ( .A1(n23966), .A2(n23965), .ZN(n23967) );
  XNOR2HSV1 U26370 ( .A1(n23968), .A2(n23967), .ZN(n23970) );
  NAND2HSV0 U26371 ( .A1(n28589), .A2(\pe1/got [2]), .ZN(n23969) );
  XNOR2HSV1 U26372 ( .A1(n23970), .A2(n23969), .ZN(n23971) );
  XNOR2HSV1 U26373 ( .A1(n23972), .A2(n23971), .ZN(n23973) );
  XOR2HSV0 U26374 ( .A1(n23974), .A2(n23973), .Z(n23975) );
  XOR2HSV0 U26375 ( .A1(n23976), .A2(n23975), .Z(n23977) );
  XNOR2HSV1 U26376 ( .A1(n23978), .A2(n23977), .ZN(n23979) );
  XNOR2HSV1 U26377 ( .A1(n23980), .A2(n23979), .ZN(n23982) );
  NAND2HSV0 U26378 ( .A1(n26909), .A2(\pe1/got [8]), .ZN(n23981) );
  XOR2HSV0 U26379 ( .A1(n23982), .A2(n23981), .Z(n23984) );
  XOR2HSV0 U26380 ( .A1(n23984), .A2(n23983), .Z(\pe1/poht [7]) );
  CLKNHSV0 U26381 ( .I(n23985), .ZN(n28581) );
  INHSV2 U26382 ( .I(\pe4/got [2]), .ZN(n27978) );
  NOR2HSV2 U26383 ( .A1(n27999), .A2(n27978), .ZN(n23996) );
  CLKAND2HSV2 U26384 ( .A1(n28480), .A2(\pe4/got [1]), .Z(n23992) );
  NAND2HSV0 U26385 ( .A1(\pe4/aot [1]), .A2(\pe4/bq[3] ), .ZN(n23988) );
  NAND2HSV0 U26386 ( .A1(\pe4/aot [2]), .A2(\pe4/bq[2] ), .ZN(n23987) );
  XOR2HSV0 U26387 ( .A1(n23988), .A2(n23987), .Z(n23990) );
  NAND2HSV0 U26388 ( .A1(\pe4/aot [3]), .A2(\pe4/bq[1] ), .ZN(n23989) );
  XNOR2HSV1 U26389 ( .A1(n23990), .A2(n23989), .ZN(n23991) );
  XOR2HSV2 U26390 ( .A1(n23992), .A2(n23991), .Z(n23995) );
  NOR2HSV2 U26391 ( .A1(n23993), .A2(n27998), .ZN(n23994) );
  XOR3HSV2 U26392 ( .A1(n23996), .A2(n23995), .A3(n23994), .Z(\pe4/poht [13])
         );
  CLKNHSV6 U26393 ( .I(n23997), .ZN(n26082) );
  NAND2HSV0 U26394 ( .A1(n26084), .A2(\pe6/got [2]), .ZN(n24005) );
  CLKNAND2HSV1 U26395 ( .A1(n28699), .A2(n28608), .ZN(n24003) );
  NAND2HSV0 U26396 ( .A1(\pe6/aot [2]), .A2(\pe6/bq[2] ), .ZN(n23999) );
  NAND2HSV0 U26397 ( .A1(\pe6/aot [1]), .A2(\pe6/bq[3] ), .ZN(n23998) );
  XOR2HSV0 U26398 ( .A1(n23999), .A2(n23998), .Z(n24001) );
  XNOR2HSV1 U26399 ( .A1(n24001), .A2(n24000), .ZN(n24002) );
  XOR2HSV0 U26400 ( .A1(n24003), .A2(n24002), .Z(n24004) );
  NAND2HSV2 U26401 ( .A1(n24277), .A2(\pe7/got [8]), .ZN(n24036) );
  CLKNAND2HSV0 U26402 ( .A1(n28665), .A2(\pe7/got [4]), .ZN(n24029) );
  NAND2HSV0 U26403 ( .A1(n28656), .A2(\pe7/got [3]), .ZN(n24027) );
  NAND2HSV0 U26404 ( .A1(n11978), .A2(\pe7/got [1]), .ZN(n24023) );
  NAND2HSV0 U26405 ( .A1(\pe7/aot [2]), .A2(\pe7/bq[7] ), .ZN(n24009) );
  NAND2HSV0 U26406 ( .A1(\pe7/aot [1]), .A2(\pe7/bq[8] ), .ZN(n24008) );
  XOR2HSV0 U26407 ( .A1(n24009), .A2(n24008), .Z(n24013) );
  NAND2HSV0 U26408 ( .A1(\pe7/aot [5]), .A2(\pe7/bq[4] ), .ZN(n24011) );
  NAND2HSV0 U26409 ( .A1(\pe7/aot [6]), .A2(\pe7/bq[3] ), .ZN(n24010) );
  XOR2HSV0 U26410 ( .A1(n24011), .A2(n24010), .Z(n24012) );
  XOR2HSV0 U26411 ( .A1(n24013), .A2(n24012), .Z(n24021) );
  NAND2HSV0 U26412 ( .A1(\pe7/aot [7]), .A2(\pe7/bq[2] ), .ZN(n24015) );
  NAND2HSV0 U26413 ( .A1(\pe7/aot [8]), .A2(\pe7/bq[1] ), .ZN(n24014) );
  XOR2HSV0 U26414 ( .A1(n24015), .A2(n24014), .Z(n24019) );
  NAND2HSV0 U26415 ( .A1(\pe7/aot [3]), .A2(\pe7/bq[6] ), .ZN(n24017) );
  NAND2HSV0 U26416 ( .A1(\pe7/aot [4]), .A2(\pe7/bq[5] ), .ZN(n24016) );
  XOR2HSV0 U26417 ( .A1(n24017), .A2(n24016), .Z(n24018) );
  XOR2HSV0 U26418 ( .A1(n24019), .A2(n24018), .Z(n24020) );
  XOR2HSV0 U26419 ( .A1(n24021), .A2(n24020), .Z(n24022) );
  XNOR2HSV1 U26420 ( .A1(n24023), .A2(n24022), .ZN(n24025) );
  NAND2HSV0 U26421 ( .A1(n25397), .A2(\pe7/got [2]), .ZN(n24024) );
  XOR2HSV0 U26422 ( .A1(n24025), .A2(n24024), .Z(n24026) );
  XNOR2HSV1 U26423 ( .A1(n24027), .A2(n24026), .ZN(n24028) );
  XOR2HSV0 U26424 ( .A1(n24029), .A2(n24028), .Z(n24031) );
  NAND2HSV0 U26425 ( .A1(n28926), .A2(\pe7/got [5]), .ZN(n24030) );
  XOR2HSV0 U26426 ( .A1(n24031), .A2(n24030), .Z(n24034) );
  NOR2HSV2 U26427 ( .A1(n24032), .A2(n19532), .ZN(n24033) );
  NAND2HSV0 U26428 ( .A1(n14030), .A2(\pe7/got [1]), .ZN(n24044) );
  NAND2HSV0 U26429 ( .A1(\pe7/aot [2]), .A2(\pe7/bq[3] ), .ZN(n24038) );
  NAND2HSV0 U26430 ( .A1(\pe7/aot [1]), .A2(\pe7/bq[4] ), .ZN(n24037) );
  XOR2HSV0 U26431 ( .A1(n24038), .A2(n24037), .Z(n24042) );
  NAND2HSV0 U26432 ( .A1(\pe7/aot [3]), .A2(\pe7/bq[2] ), .ZN(n24040) );
  NAND2HSV0 U26433 ( .A1(\pe7/aot [4]), .A2(\pe7/bq[1] ), .ZN(n24039) );
  XOR2HSV0 U26434 ( .A1(n24040), .A2(n24039), .Z(n24041) );
  XOR2HSV0 U26435 ( .A1(n24042), .A2(n24041), .Z(n24043) );
  XNOR2HSV1 U26436 ( .A1(n24044), .A2(n24043), .ZN(n24048) );
  NOR2HSV2 U26437 ( .A1(n24045), .A2(n25308), .ZN(n24047) );
  AND2HSV2 U26438 ( .A1(n28703), .A2(\pe7/got [3]), .Z(n24046) );
  XNOR3HSV2 U26439 ( .A1(n24048), .A2(n24047), .A3(n24046), .ZN(n24049) );
  NAND2HSV2 U26440 ( .A1(n24277), .A2(n24214), .ZN(n24080) );
  NAND2HSV0 U26441 ( .A1(n14066), .A2(\pe7/got [2]), .ZN(n24070) );
  NAND2HSV0 U26442 ( .A1(\pe7/got [1]), .A2(n11935), .ZN(n24068) );
  NAND2HSV0 U26443 ( .A1(\pe7/aot [1]), .A2(\pe7/bq[10] ), .ZN(n24051) );
  NAND2HSV0 U26444 ( .A1(\pe7/aot [9]), .A2(\pe7/bq[2] ), .ZN(n24050) );
  XOR2HSV0 U26445 ( .A1(n24051), .A2(n24050), .Z(n24066) );
  NAND2HSV0 U26446 ( .A1(\pe7/aot [2]), .A2(\pe7/bq[9] ), .ZN(n24053) );
  NAND2HSV0 U26447 ( .A1(\pe7/aot [3]), .A2(\pe7/bq[8] ), .ZN(n24052) );
  XOR2HSV0 U26448 ( .A1(n24053), .A2(n24052), .Z(n24057) );
  INHSV2 U26449 ( .I(\pe7/bq[1] ), .ZN(n27095) );
  NOR2HSV0 U26450 ( .A1(n24105), .A2(n27095), .ZN(n24055) );
  NAND2HSV0 U26451 ( .A1(\pe7/aot [4]), .A2(\pe7/bq[7] ), .ZN(n24054) );
  XOR2HSV0 U26452 ( .A1(n24055), .A2(n24054), .Z(n24056) );
  XNOR2HSV1 U26453 ( .A1(n24057), .A2(n24056), .ZN(n24065) );
  NAND2HSV0 U26454 ( .A1(\pe7/aot [5]), .A2(\pe7/bq[6] ), .ZN(n24059) );
  NAND2HSV0 U26455 ( .A1(\pe7/aot [6]), .A2(\pe7/bq[5] ), .ZN(n24058) );
  XOR2HSV0 U26456 ( .A1(n24059), .A2(n24058), .Z(n24063) );
  NAND2HSV0 U26457 ( .A1(\pe7/aot [7]), .A2(\pe7/bq[4] ), .ZN(n24061) );
  NAND2HSV0 U26458 ( .A1(\pe7/aot [8]), .A2(\pe7/bq[3] ), .ZN(n24060) );
  XOR2HSV0 U26459 ( .A1(n24061), .A2(n24060), .Z(n24062) );
  XOR2HSV0 U26460 ( .A1(n24063), .A2(n24062), .Z(n24064) );
  XOR3HSV2 U26461 ( .A1(n24066), .A2(n24065), .A3(n24064), .Z(n24067) );
  XNOR2HSV1 U26462 ( .A1(n24068), .A2(n24067), .ZN(n24069) );
  NAND2HSV0 U26463 ( .A1(\pe7/got [7]), .A2(n28926), .ZN(n24071) );
  XOR2HSV0 U26464 ( .A1(n24072), .A2(n24071), .Z(n24078) );
  AOI31HSV0 U26465 ( .A1(n24075), .A2(n24074), .A3(n24073), .B(n24213), .ZN(
        n24076) );
  XOR3HSV2 U26466 ( .A1(n24078), .A2(n24077), .A3(n24076), .Z(n24079) );
  NAND2HSV2 U26467 ( .A1(n28659), .A2(n25334), .ZN(n24132) );
  NAND2HSV0 U26468 ( .A1(n25377), .A2(\pe7/got [8]), .ZN(n24083) );
  NAND2HSV0 U26469 ( .A1(n25397), .A2(\pe7/got [7]), .ZN(n24081) );
  INHSV1 U26470 ( .I(n24081), .ZN(n24082) );
  XNOR2HSV1 U26471 ( .A1(n24083), .A2(n24082), .ZN(n24086) );
  CLKNHSV0 U26472 ( .I(n24086), .ZN(n24085) );
  NOR2HSV1 U26473 ( .A1(n24085), .A2(n24084), .ZN(n24088) );
  AOI21HSV0 U26474 ( .A1(n28926), .A2(n24214), .B(n24086), .ZN(n24087) );
  AOI21HSV2 U26475 ( .A1(n24088), .A2(n25335), .B(n24087), .ZN(n24127) );
  CLKNAND2HSV0 U26476 ( .A1(n24287), .A2(\pe7/got [9]), .ZN(n24125) );
  NAND2HSV0 U26477 ( .A1(n14067), .A2(\pe7/got [5]), .ZN(n24121) );
  NAND2HSV0 U26478 ( .A1(n25272), .A2(n19579), .ZN(n24119) );
  NAND2HSV0 U26479 ( .A1(n25318), .A2(\pe7/got [3]), .ZN(n24117) );
  NAND2HSV0 U26480 ( .A1(n11936), .A2(\pe7/got [2]), .ZN(n24115) );
  NAND2HSV0 U26481 ( .A1(n28621), .A2(\pe7/got [1]), .ZN(n24113) );
  NAND2HSV0 U26482 ( .A1(n14050), .A2(\pe7/bq[1] ), .ZN(n24090) );
  NAND2HSV0 U26483 ( .A1(\pe7/aot [7]), .A2(\pe7/bq[7] ), .ZN(n24089) );
  XOR2HSV0 U26484 ( .A1(n24090), .A2(n24089), .Z(n24094) );
  NAND2HSV0 U26485 ( .A1(\pe7/aot [2]), .A2(\pe7/bq[12] ), .ZN(n24092) );
  NAND2HSV0 U26486 ( .A1(\pe7/aot [5]), .A2(\pe7/bq[9] ), .ZN(n24091) );
  XOR2HSV0 U26487 ( .A1(n24092), .A2(n24091), .Z(n24093) );
  XOR2HSV0 U26488 ( .A1(n24094), .A2(n24093), .Z(n24102) );
  NAND2HSV0 U26489 ( .A1(\pe7/aot [3]), .A2(\pe7/bq[11] ), .ZN(n24096) );
  NAND2HSV0 U26490 ( .A1(\pe7/aot [1]), .A2(\pe7/bq[13] ), .ZN(n24095) );
  XOR2HSV0 U26491 ( .A1(n24096), .A2(n24095), .Z(n24100) );
  NAND2HSV0 U26492 ( .A1(\pe7/aot [9]), .A2(\pe7/bq[5] ), .ZN(n24098) );
  NAND2HSV0 U26493 ( .A1(\pe7/aot [6]), .A2(\pe7/bq[8] ), .ZN(n24097) );
  XOR2HSV0 U26494 ( .A1(n24098), .A2(n24097), .Z(n24099) );
  XOR2HSV0 U26495 ( .A1(n24100), .A2(n24099), .Z(n24101) );
  XOR2HSV0 U26496 ( .A1(n24102), .A2(n24101), .Z(n24111) );
  NAND2HSV0 U26497 ( .A1(\pe7/aot [11]), .A2(\pe7/bq[3] ), .ZN(n25279) );
  NAND2HSV0 U26498 ( .A1(\pe7/aot [8]), .A2(\pe7/bq[6] ), .ZN(n24104) );
  NAND2HSV0 U26499 ( .A1(\pe7/aot [4]), .A2(\pe7/bq[10] ), .ZN(n24103) );
  XOR2HSV0 U26500 ( .A1(n24104), .A2(n24103), .Z(n24109) );
  NOR2HSV0 U26501 ( .A1(n24105), .A2(n19649), .ZN(n24107) );
  NAND2HSV0 U26502 ( .A1(\pe7/aot [12]), .A2(\pe7/bq[2] ), .ZN(n24106) );
  XOR2HSV0 U26503 ( .A1(n24107), .A2(n24106), .Z(n24108) );
  XOR3HSV2 U26504 ( .A1(n25279), .A2(n24109), .A3(n24108), .Z(n24110) );
  XNOR2HSV1 U26505 ( .A1(n24111), .A2(n24110), .ZN(n24112) );
  XNOR2HSV1 U26506 ( .A1(n24113), .A2(n24112), .ZN(n24114) );
  XNOR2HSV1 U26507 ( .A1(n24115), .A2(n24114), .ZN(n24116) );
  XNOR2HSV1 U26508 ( .A1(n24117), .A2(n24116), .ZN(n24118) );
  XOR2HSV0 U26509 ( .A1(n24119), .A2(n24118), .Z(n24120) );
  XNOR2HSV1 U26510 ( .A1(n24121), .A2(n24120), .ZN(n24123) );
  NAND2HSV0 U26511 ( .A1(n28587), .A2(\pe7/got [6]), .ZN(n24122) );
  XOR2HSV0 U26512 ( .A1(n24123), .A2(n24122), .Z(n24124) );
  XOR2HSV0 U26513 ( .A1(n24125), .A2(n24124), .Z(n24126) );
  XOR2HSV0 U26514 ( .A1(n24127), .A2(n24126), .Z(n24130) );
  AND2HSV2 U26515 ( .A1(n25408), .A2(\pe7/got [12]), .Z(n24129) );
  XOR2HSV0 U26516 ( .A1(n24131), .A2(n24132), .Z(\pe7/poht [3]) );
  NAND2HSV2 U26517 ( .A1(n24277), .A2(n24271), .ZN(n24186) );
  CLKNAND2HSV1 U26518 ( .A1(n25376), .A2(n24214), .ZN(n24178) );
  NAND2HSV0 U26519 ( .A1(n25377), .A2(\pe7/got [9]), .ZN(n24176) );
  NAND2HSV0 U26520 ( .A1(n11978), .A2(n25271), .ZN(n24172) );
  NAND2HSV0 U26521 ( .A1(n14067), .A2(\pe7/got [6]), .ZN(n24170) );
  NAND2HSV0 U26522 ( .A1(n25375), .A2(n28466), .ZN(n24168) );
  NAND2HSV0 U26523 ( .A1(n11936), .A2(\pe7/got [3]), .ZN(n24164) );
  NAND2HSV0 U26524 ( .A1(n14050), .A2(\pe7/bq[2] ), .ZN(n24134) );
  NAND2HSV0 U26525 ( .A1(\pe7/aot [10]), .A2(\pe7/bq[5] ), .ZN(n24133) );
  XOR2HSV0 U26526 ( .A1(n24134), .A2(n24133), .Z(n24138) );
  NAND2HSV0 U26527 ( .A1(\pe7/aot [12]), .A2(\pe7/bq[3] ), .ZN(n24136) );
  NAND2HSV0 U26528 ( .A1(\pe7/aot [14]), .A2(\pe7/bq[1] ), .ZN(n24135) );
  XOR2HSV0 U26529 ( .A1(n24136), .A2(n24135), .Z(n24137) );
  XOR2HSV0 U26530 ( .A1(n24138), .A2(n24137), .Z(n24146) );
  NAND2HSV0 U26531 ( .A1(\pe7/aot [7]), .A2(\pe7/bq[8] ), .ZN(n24140) );
  NAND2HSV0 U26532 ( .A1(\pe7/aot [11]), .A2(\pe7/bq[4] ), .ZN(n24139) );
  XOR2HSV0 U26533 ( .A1(n24140), .A2(n24139), .Z(n24144) );
  NAND2HSV0 U26534 ( .A1(\pe7/aot [3]), .A2(\pe7/bq[12] ), .ZN(n24142) );
  NAND2HSV0 U26535 ( .A1(\pe7/aot [4]), .A2(\pe7/bq[11] ), .ZN(n24141) );
  XOR2HSV0 U26536 ( .A1(n24142), .A2(n24141), .Z(n24143) );
  XOR2HSV0 U26537 ( .A1(n24144), .A2(n24143), .Z(n24145) );
  XOR2HSV0 U26538 ( .A1(n24146), .A2(n24145), .Z(n24158) );
  NAND2HSV0 U26539 ( .A1(\pe7/aot [2]), .A2(\pe7/bq[13] ), .ZN(n24148) );
  NAND2HSV0 U26540 ( .A1(\pe7/aot [1]), .A2(\pe7/bq[14] ), .ZN(n24147) );
  XOR2HSV0 U26541 ( .A1(n24148), .A2(n24147), .Z(n24152) );
  NAND2HSV0 U26542 ( .A1(\pe7/aot [8]), .A2(\pe7/bq[7] ), .ZN(n24150) );
  NAND2HSV0 U26543 ( .A1(\pe7/aot [9]), .A2(\pe7/bq[6] ), .ZN(n24149) );
  XOR2HSV0 U26544 ( .A1(n24150), .A2(n24149), .Z(n24151) );
  XOR2HSV0 U26545 ( .A1(n24152), .A2(n24151), .Z(n24156) );
  NAND2HSV0 U26546 ( .A1(\pe7/aot [5]), .A2(\pe7/bq[10] ), .ZN(n24154) );
  NAND2HSV0 U26547 ( .A1(\pe7/aot [6]), .A2(\pe7/bq[9] ), .ZN(n24153) );
  XOR2HSV0 U26548 ( .A1(n24154), .A2(n24153), .Z(n24155) );
  XNOR2HSV1 U26549 ( .A1(n24156), .A2(n24155), .ZN(n24157) );
  XNOR2HSV1 U26550 ( .A1(n24158), .A2(n24157), .ZN(n24160) );
  NAND2HSV0 U26551 ( .A1(n25292), .A2(\pe7/got [1]), .ZN(n24159) );
  XNOR2HSV1 U26552 ( .A1(n24160), .A2(n24159), .ZN(n24162) );
  NAND2HSV0 U26553 ( .A1(n24250), .A2(\pe7/got [2]), .ZN(n24161) );
  XOR2HSV0 U26554 ( .A1(n24162), .A2(n24161), .Z(n24163) );
  XOR2HSV0 U26555 ( .A1(n24164), .A2(n24163), .Z(n24166) );
  NAND2HSV0 U26556 ( .A1(n25318), .A2(n25272), .ZN(n24165) );
  XOR2HSV0 U26557 ( .A1(n24166), .A2(n24165), .Z(n24167) );
  XOR2HSV0 U26558 ( .A1(n24168), .A2(n24167), .Z(n24169) );
  XNOR2HSV1 U26559 ( .A1(n24170), .A2(n24169), .ZN(n24171) );
  XNOR2HSV1 U26560 ( .A1(n24172), .A2(n24171), .ZN(n24174) );
  NAND2HSV0 U26561 ( .A1(n25397), .A2(\pe7/got [8]), .ZN(n24173) );
  XNOR2HSV1 U26562 ( .A1(n24174), .A2(n24173), .ZN(n24175) );
  XNOR2HSV1 U26563 ( .A1(n24176), .A2(n24175), .ZN(n24177) );
  XOR2HSV0 U26564 ( .A1(n24178), .A2(n24177), .Z(n24180) );
  NAND2HSV0 U26565 ( .A1(n25335), .A2(n14022), .ZN(n24179) );
  NOR2HSV2 U26566 ( .A1(n24286), .A2(n24321), .ZN(n24183) );
  AND2HSV2 U26567 ( .A1(n25408), .A2(n24181), .Z(n24182) );
  XOR3HSV2 U26568 ( .A1(n24184), .A2(n24183), .A3(n24182), .Z(n24185) );
  XOR2HSV0 U26569 ( .A1(n24186), .A2(n24185), .Z(\pe7/poht [2]) );
  NAND2HSV2 U26570 ( .A1(n28659), .A2(n14022), .ZN(n24219) );
  NAND2HSV0 U26571 ( .A1(\pe7/got [2]), .A2(n11935), .ZN(n24210) );
  NAND2HSV0 U26572 ( .A1(n25318), .A2(\pe7/got [1]), .ZN(n24208) );
  NAND2HSV0 U26573 ( .A1(\pe7/aot [8]), .A2(\pe7/bq[4] ), .ZN(n24188) );
  NAND2HSV0 U26574 ( .A1(\pe7/aot [11]), .A2(\pe7/bq[1] ), .ZN(n24187) );
  XOR2HSV0 U26575 ( .A1(n24188), .A2(n24187), .Z(n24192) );
  NAND2HSV0 U26576 ( .A1(\pe7/aot [1]), .A2(\pe7/bq[11] ), .ZN(n24190) );
  NAND2HSV0 U26577 ( .A1(\pe7/aot [7]), .A2(\pe7/bq[5] ), .ZN(n24189) );
  XOR2HSV0 U26578 ( .A1(n24190), .A2(n24189), .Z(n24191) );
  XOR2HSV0 U26579 ( .A1(n24192), .A2(n24191), .Z(n24198) );
  NAND2HSV0 U26580 ( .A1(\pe7/aot [2]), .A2(\pe7/bq[10] ), .ZN(n24194) );
  NAND2HSV0 U26581 ( .A1(\pe7/aot [6]), .A2(\pe7/bq[6] ), .ZN(n24193) );
  XOR2HSV0 U26582 ( .A1(n24194), .A2(n24193), .Z(n24196) );
  NAND2HSV0 U26583 ( .A1(\pe7/aot [5]), .A2(\pe7/bq[7] ), .ZN(n24195) );
  XNOR2HSV1 U26584 ( .A1(n24196), .A2(n24195), .ZN(n24197) );
  XNOR2HSV1 U26585 ( .A1(n24198), .A2(n24197), .ZN(n24206) );
  NAND2HSV0 U26586 ( .A1(\pe7/aot [4]), .A2(\pe7/bq[8] ), .ZN(n24200) );
  NAND2HSV0 U26587 ( .A1(\pe7/aot [9]), .A2(\pe7/bq[3] ), .ZN(n24199) );
  XOR2HSV0 U26588 ( .A1(n24200), .A2(n24199), .Z(n24204) );
  NAND2HSV0 U26589 ( .A1(\pe7/aot [3]), .A2(\pe7/bq[9] ), .ZN(n24202) );
  NAND2HSV0 U26590 ( .A1(\pe7/aot [10]), .A2(\pe7/bq[2] ), .ZN(n24201) );
  XOR2HSV0 U26591 ( .A1(n24202), .A2(n24201), .Z(n24203) );
  XOR2HSV0 U26592 ( .A1(n24204), .A2(n24203), .Z(n24205) );
  XNOR2HSV1 U26593 ( .A1(n24206), .A2(n24205), .ZN(n24207) );
  XOR2HSV0 U26594 ( .A1(n24208), .A2(n24207), .Z(n24209) );
  NAND2HSV0 U26595 ( .A1(\pe7/got [8]), .A2(n14030), .ZN(n24211) );
  XNOR2HSV1 U26596 ( .A1(n24212), .A2(n24211), .ZN(n24217) );
  NOR2HSV2 U26597 ( .A1(n24286), .A2(n24213), .ZN(n24216) );
  XOR3HSV2 U26598 ( .A1(n24217), .A2(n24216), .A3(n24215), .Z(n24218) );
  XOR2HSV0 U26599 ( .A1(n24219), .A2(n24218), .Z(\pe7/poht [5]) );
  CLKNAND2HSV0 U26600 ( .A1(n28665), .A2(n14022), .ZN(n24268) );
  NAND2HSV0 U26601 ( .A1(n25377), .A2(n24214), .ZN(n24266) );
  NAND2HSV0 U26602 ( .A1(n14067), .A2(n25271), .ZN(n24260) );
  NAND2HSV0 U26603 ( .A1(\pe7/got [6]), .A2(n28466), .ZN(n24258) );
  NOR2HSV0 U26604 ( .A1(n25309), .A2(n24221), .ZN(n24249) );
  NAND2HSV0 U26605 ( .A1(n25292), .A2(\pe7/got [2]), .ZN(n24248) );
  NAND2HSV0 U26606 ( .A1(\pe7/aot [6]), .A2(\pe7/bq[10] ), .ZN(n24223) );
  NAND2HSV0 U26607 ( .A1(\pe7/aot [10]), .A2(\pe7/bq[6] ), .ZN(n24222) );
  XOR2HSV0 U26608 ( .A1(n24223), .A2(n24222), .Z(n24227) );
  NAND2HSV0 U26609 ( .A1(\pe7/aot [9]), .A2(\pe7/bq[7] ), .ZN(n24225) );
  NAND2HSV0 U26610 ( .A1(\pe7/aot [12]), .A2(\pe7/bq[4] ), .ZN(n24224) );
  XOR2HSV0 U26611 ( .A1(n24225), .A2(n24224), .Z(n24226) );
  XOR2HSV0 U26612 ( .A1(n24227), .A2(n24226), .Z(n24234) );
  NAND2HSV0 U26613 ( .A1(\pe7/bq[1] ), .A2(\pe7/aot [15]), .ZN(n25302) );
  XOR2HSV0 U26614 ( .A1(n24228), .A2(n25302), .Z(n24232) );
  NAND2HSV0 U26615 ( .A1(n14050), .A2(\pe7/bq[3] ), .ZN(n24230) );
  NAND2HSV0 U26616 ( .A1(\pe7/aot [8]), .A2(\pe7/bq[8] ), .ZN(n24229) );
  XOR2HSV0 U26617 ( .A1(n24230), .A2(n24229), .Z(n24231) );
  XOR2HSV0 U26618 ( .A1(n24232), .A2(n24231), .Z(n24233) );
  XOR2HSV0 U26619 ( .A1(n24234), .A2(n24233), .Z(n24246) );
  NAND2HSV0 U26620 ( .A1(\pe7/aot [7]), .A2(\pe7/bq[9] ), .ZN(n24236) );
  NAND2HSV0 U26621 ( .A1(\pe7/aot [3]), .A2(\pe7/bq[13] ), .ZN(n24235) );
  XOR2HSV0 U26622 ( .A1(n24236), .A2(n24235), .Z(n24240) );
  NAND2HSV0 U26623 ( .A1(\pe7/aot [4]), .A2(\pe7/bq[12] ), .ZN(n24238) );
  NAND2HSV0 U26624 ( .A1(\pe7/aot [1]), .A2(\pe7/bq[15] ), .ZN(n24237) );
  XOR2HSV0 U26625 ( .A1(n24238), .A2(n24237), .Z(n24239) );
  XOR2HSV0 U26626 ( .A1(n24240), .A2(n24239), .Z(n24244) );
  NAND2HSV0 U26627 ( .A1(\pe7/aot [5]), .A2(\pe7/bq[5] ), .ZN(n25382) );
  NAND2HSV0 U26628 ( .A1(\pe7/aot [2]), .A2(\pe7/bq[14] ), .ZN(n25276) );
  XOR2HSV0 U26629 ( .A1(n24242), .A2(n25276), .Z(n24243) );
  XNOR2HSV1 U26630 ( .A1(n24244), .A2(n24243), .ZN(n24245) );
  XNOR2HSV1 U26631 ( .A1(n24246), .A2(n24245), .ZN(n24247) );
  XOR3HSV2 U26632 ( .A1(n24249), .A2(n24248), .A3(n24247), .Z(n24252) );
  NAND2HSV0 U26633 ( .A1(n24250), .A2(\pe7/got [3]), .ZN(n24251) );
  XNOR2HSV1 U26634 ( .A1(n24252), .A2(n24251), .ZN(n24254) );
  NAND2HSV0 U26635 ( .A1(n11936), .A2(n25272), .ZN(n24253) );
  XOR2HSV0 U26636 ( .A1(n24254), .A2(n24253), .Z(n24256) );
  NAND2HSV0 U26637 ( .A1(n25318), .A2(n25375), .ZN(n24255) );
  XOR2HSV0 U26638 ( .A1(n24256), .A2(n24255), .Z(n24257) );
  XOR2HSV0 U26639 ( .A1(n24258), .A2(n24257), .Z(n24259) );
  XOR2HSV0 U26640 ( .A1(n24260), .A2(n24259), .Z(n24262) );
  NAND2HSV0 U26641 ( .A1(n11978), .A2(\pe7/got [8]), .ZN(n24261) );
  XOR2HSV0 U26642 ( .A1(n24262), .A2(n24261), .Z(n24264) );
  NAND2HSV0 U26643 ( .A1(n25397), .A2(\pe7/got [9]), .ZN(n24263) );
  XNOR2HSV1 U26644 ( .A1(n24264), .A2(n24263), .ZN(n24265) );
  XNOR2HSV1 U26645 ( .A1(n24266), .A2(n24265), .ZN(n24267) );
  XOR2HSV0 U26646 ( .A1(n24268), .A2(n24267), .Z(n24270) );
  NAND2HSV0 U26647 ( .A1(n28926), .A2(\pe7/got [12]), .ZN(n24269) );
  XNOR2HSV1 U26648 ( .A1(n24270), .A2(n24269), .ZN(n24274) );
  NAND2HSV0 U26649 ( .A1(n28703), .A2(\pe7/got [1]), .ZN(n24281) );
  NAND2HSV0 U26650 ( .A1(\pe7/aot [2]), .A2(\pe7/bq[1] ), .ZN(n24279) );
  NAND2HSV0 U26651 ( .A1(\pe7/aot [1]), .A2(\pe7/bq[2] ), .ZN(n24278) );
  XOR2HSV0 U26652 ( .A1(n24279), .A2(n24278), .Z(n24280) );
  XOR2HSV0 U26653 ( .A1(n24281), .A2(n24280), .Z(n24282) );
  XOR2HSV0 U26654 ( .A1(n24283), .A2(n24282), .Z(\pe7/poht [14]) );
  CLKNAND2HSV2 U26655 ( .A1(n24284), .A2(\pe7/got [5]), .ZN(n24304) );
  NOR2HSV2 U26656 ( .A1(n25374), .A2(n24285), .ZN(n24301) );
  CLKNAND2HSV1 U26657 ( .A1(n25335), .A2(\pe7/got [2]), .ZN(n24299) );
  CLKNAND2HSV1 U26658 ( .A1(n24287), .A2(\pe7/got [1]), .ZN(n24297) );
  NAND2HSV0 U26659 ( .A1(\pe7/aot [5]), .A2(\pe7/bq[1] ), .ZN(n24289) );
  NAND2HSV0 U26660 ( .A1(\pe7/aot [3]), .A2(\pe7/bq[3] ), .ZN(n24288) );
  XOR2HSV0 U26661 ( .A1(n24289), .A2(n24288), .Z(n24291) );
  NAND2HSV0 U26662 ( .A1(\pe7/aot [4]), .A2(\pe7/bq[2] ), .ZN(n24290) );
  XNOR2HSV1 U26663 ( .A1(n24291), .A2(n24290), .ZN(n24295) );
  NAND2HSV0 U26664 ( .A1(\pe7/aot [2]), .A2(\pe7/bq[4] ), .ZN(n24293) );
  NAND2HSV0 U26665 ( .A1(\pe7/aot [1]), .A2(\pe7/bq[5] ), .ZN(n24292) );
  XOR2HSV0 U26666 ( .A1(n24293), .A2(n24292), .Z(n24294) );
  XNOR2HSV1 U26667 ( .A1(n24295), .A2(n24294), .ZN(n24296) );
  XOR2HSV0 U26668 ( .A1(n24297), .A2(n24296), .Z(n24298) );
  XNOR2HSV1 U26669 ( .A1(n24299), .A2(n24298), .ZN(n24300) );
  XNOR2HSV4 U26670 ( .A1(n24301), .A2(n24300), .ZN(n24302) );
  XNOR2HSV4 U26671 ( .A1(n24302), .A2(n13960), .ZN(n24303) );
  CLKNHSV0 U26672 ( .I(bo6[8]), .ZN(n24306) );
  MUX2NHSV1 U26673 ( .I0(n24307), .I1(n24306), .S(n24305), .ZN(n28748) );
  MUX2HSV2 U26674 ( .I0(bo6[16]), .I1(n14028), .S(n27072), .Z(n28732) );
  CLKNHSV0 U26675 ( .I(n23793), .ZN(n28596) );
  CLKNHSV0 U26676 ( .I(n24310), .ZN(n28605) );
  INHSV2 U26677 ( .I(n24312), .ZN(n28619) );
  CLKNHSV0 U26678 ( .I(\pe1/bq[8] ), .ZN(n24315) );
  INHSV2 U26679 ( .I(n24315), .ZN(n24317) );
  INHSV2 U26680 ( .I(n24316), .ZN(n27065) );
  MUX2HSV2 U26681 ( .I0(bo1[8]), .I1(n24317), .S(n27065), .Z(n28736) );
  CLKNHSV0 U26682 ( .I(\pe1/bq[14] ), .ZN(n24318) );
  INHSV2 U26683 ( .I(n24318), .ZN(n24319) );
  MUX2HSV2 U26684 ( .I0(bo1[14]), .I1(n24319), .S(n28598), .Z(n28734) );
  MUX2HSV2 U26685 ( .I0(bo11[4]), .I1(\pe11/bq[4] ), .S(n27057), .Z(n28723) );
  MUX2HSV2 U26686 ( .I0(bo11[3]), .I1(\pe11/bq[3] ), .S(n24320), .Z(n28720) );
  MUX2HSV2 U26687 ( .I0(bo11[7]), .I1(\pe11/bq[7] ), .S(n24320), .Z(n28719) );
  CLKNHSV0 U26688 ( .I(n25374), .ZN(n28934) );
  INHSV2 U26689 ( .I(go7[16]), .ZN(n28670) );
  NAND2HSV0 U26690 ( .A1(n28473), .A2(\pe5/got [2]), .ZN(n24336) );
  NAND2HSV0 U26691 ( .A1(n21452), .A2(n28640), .ZN(n24334) );
  NAND2HSV0 U26692 ( .A1(\pe5/aot [4]), .A2(\pe5/bq[2] ), .ZN(n24332) );
  NOR2HSV0 U26693 ( .A1(n24443), .A2(n24323), .ZN(n24325) );
  AOI22HSV0 U26694 ( .A1(\pe5/aot [2]), .A2(\pe5/bq[4] ), .B1(\pe5/bq[5] ), 
        .B2(\pe5/aot [1]), .ZN(n24324) );
  NOR2HSV2 U26695 ( .A1(n24325), .A2(n24324), .ZN(n24331) );
  IOA22HSV1 U26696 ( .B1(n24440), .B2(n24326), .A1(\pe5/aot [3]), .A2(
        \pe5/bq[3] ), .ZN(n24327) );
  OAI21HSV1 U26697 ( .A1(n24329), .A2(n24328), .B(n24327), .ZN(n24330) );
  XOR3HSV2 U26698 ( .A1(n24332), .A2(n24331), .A3(n24330), .Z(n24333) );
  XOR2HSV0 U26699 ( .A1(n24334), .A2(n24333), .Z(n24335) );
  XOR2HSV0 U26700 ( .A1(n24336), .A2(n24335), .Z(n24337) );
  NAND2HSV0 U26701 ( .A1(n12517), .A2(n24340), .ZN(n24375) );
  NAND2HSV0 U26702 ( .A1(n24341), .A2(n28645), .ZN(n24373) );
  NAND2HSV0 U26703 ( .A1(n21523), .A2(\pe5/got [2]), .ZN(n24363) );
  NAND2HSV0 U26704 ( .A1(n28478), .A2(n28640), .ZN(n24361) );
  NAND2HSV0 U26705 ( .A1(\pe5/aot [10]), .A2(\pe5/bq[1] ), .ZN(n24343) );
  NAND2HSV0 U26706 ( .A1(\pe5/aot [6]), .A2(\pe5/bq[5] ), .ZN(n24342) );
  XOR2HSV0 U26707 ( .A1(n24343), .A2(n24342), .Z(n24359) );
  NAND2HSV0 U26708 ( .A1(\pe5/aot [9]), .A2(\pe5/bq[2] ), .ZN(n24345) );
  NAND2HSV0 U26709 ( .A1(\pe5/aot [4]), .A2(\pe5/bq[7] ), .ZN(n24344) );
  XOR2HSV0 U26710 ( .A1(n24345), .A2(n24344), .Z(n24350) );
  NOR2HSV0 U26711 ( .A1(n24440), .A2(n24346), .ZN(n24348) );
  NAND2HSV0 U26712 ( .A1(\pe5/aot [2]), .A2(\pe5/bq[9] ), .ZN(n24347) );
  XOR2HSV0 U26713 ( .A1(n24348), .A2(n24347), .Z(n24349) );
  XNOR2HSV1 U26714 ( .A1(n24350), .A2(n24349), .ZN(n24358) );
  NAND2HSV0 U26715 ( .A1(\pe5/aot [7]), .A2(\pe5/bq[4] ), .ZN(n24352) );
  NAND2HSV0 U26716 ( .A1(\pe5/aot [3]), .A2(\pe5/bq[8] ), .ZN(n24351) );
  XOR2HSV0 U26717 ( .A1(n24352), .A2(n24351), .Z(n24356) );
  NAND2HSV0 U26718 ( .A1(\pe5/aot [8]), .A2(\pe5/bq[3] ), .ZN(n24354) );
  NAND2HSV0 U26719 ( .A1(\pe5/aot [1]), .A2(\pe5/bq[10] ), .ZN(n24353) );
  XOR2HSV0 U26720 ( .A1(n24354), .A2(n24353), .Z(n24355) );
  XOR2HSV0 U26721 ( .A1(n24356), .A2(n24355), .Z(n24357) );
  XOR3HSV2 U26722 ( .A1(n24359), .A2(n24358), .A3(n24357), .Z(n24360) );
  XNOR2HSV1 U26723 ( .A1(n24361), .A2(n24360), .ZN(n24362) );
  XNOR2HSV1 U26724 ( .A1(n24363), .A2(n24362), .ZN(n24367) );
  NOR2HSV2 U26725 ( .A1(n24684), .A2(n24364), .ZN(n24366) );
  OR2HSV1 U26726 ( .A1(n24686), .A2(n24414), .Z(n24365) );
  XOR3HSV2 U26727 ( .A1(n24367), .A2(n24366), .A3(n24365), .Z(n24368) );
  XNOR2HSV1 U26728 ( .A1(n24371), .A2(n24370), .ZN(n24372) );
  XOR2HSV0 U26729 ( .A1(n24373), .A2(n24372), .Z(n24374) );
  NAND2HSV0 U26730 ( .A1(n21718), .A2(n24636), .ZN(n24432) );
  NAND2HSV0 U26731 ( .A1(\pe5/ti_7[10] ), .A2(n14069), .ZN(n24426) );
  NAND2HSV0 U26732 ( .A1(n11931), .A2(n28647), .ZN(n24419) );
  NAND2HSV0 U26733 ( .A1(n28614), .A2(\pe5/got [2]), .ZN(n24410) );
  NAND2HSV0 U26734 ( .A1(\pe5/aot [10]), .A2(\pe5/bq[5] ), .ZN(n24380) );
  NAND2HSV0 U26735 ( .A1(\pe5/aot [12]), .A2(\pe5/bq[3] ), .ZN(n24379) );
  XOR2HSV0 U26736 ( .A1(n24380), .A2(n24379), .Z(n24405) );
  NAND2HSV0 U26737 ( .A1(\pe5/aot [9]), .A2(\pe5/bq[6] ), .ZN(n24382) );
  NAND2HSV0 U26738 ( .A1(\pe5/aot [8]), .A2(\pe5/bq[7] ), .ZN(n24381) );
  XOR2HSV0 U26739 ( .A1(n24382), .A2(n24381), .Z(n24386) );
  NAND2HSV0 U26740 ( .A1(\pe5/aot [5]), .A2(\pe5/bq[10] ), .ZN(n24384) );
  INAND2HSV0 U26741 ( .A1(n14766), .B1(\pe5/aot [3]), .ZN(n24383) );
  XOR2HSV0 U26742 ( .A1(n24384), .A2(n24383), .Z(n24385) );
  XNOR2HSV1 U26743 ( .A1(n24386), .A2(n24385), .ZN(n24404) );
  AOI22HSV0 U26744 ( .A1(\pe5/aot [13]), .A2(\pe5/bq[2] ), .B1(\pe5/bq[9] ), 
        .B2(\pe5/aot [6]), .ZN(n24387) );
  AOI21HSV0 U26745 ( .A1(n24389), .A2(n24388), .B(n24387), .ZN(n24395) );
  NOR2HSV0 U26746 ( .A1(n24391), .A2(n24390), .ZN(n24393) );
  AOI22HSV0 U26747 ( .A1(\pe5/bq[1] ), .A2(\pe5/aot [14]), .B1(\pe5/bq[11] ), 
        .B2(\pe5/aot [4]), .ZN(n24392) );
  NOR2HSV1 U26748 ( .A1(n24393), .A2(n24392), .ZN(n24394) );
  XOR2HSV0 U26749 ( .A1(n24395), .A2(n24394), .Z(n24403) );
  NAND2HSV0 U26750 ( .A1(\pe5/aot [2]), .A2(\pe5/bq[13] ), .ZN(n24397) );
  NAND2HSV0 U26751 ( .A1(\pe5/aot [1]), .A2(\pe5/bq[14] ), .ZN(n24396) );
  XOR2HSV0 U26752 ( .A1(n24397), .A2(n24396), .Z(n24401) );
  NAND2HSV0 U26753 ( .A1(\pe5/aot [11]), .A2(\pe5/bq[4] ), .ZN(n24399) );
  NAND2HSV0 U26754 ( .A1(\pe5/aot [7]), .A2(\pe5/bq[8] ), .ZN(n24398) );
  XOR2HSV0 U26755 ( .A1(n24399), .A2(n24398), .Z(n24400) );
  XOR2HSV0 U26756 ( .A1(n24401), .A2(n24400), .Z(n24402) );
  XOR4HSV1 U26757 ( .A1(n24405), .A2(n24404), .A3(n24403), .A4(n24402), .Z(
        n24408) );
  NAND2HSV0 U26758 ( .A1(n28594), .A2(n28640), .ZN(n24407) );
  XNOR2HSV1 U26759 ( .A1(n24408), .A2(n24407), .ZN(n24409) );
  XOR2HSV0 U26760 ( .A1(n24410), .A2(n24409), .Z(n24413) );
  NAND2HSV0 U26761 ( .A1(n24411), .A2(\pe5/got [3]), .ZN(n24412) );
  XOR2HSV0 U26762 ( .A1(n24413), .A2(n24412), .Z(n24417) );
  NOR2HSV0 U26763 ( .A1(n25350), .A2(n24414), .ZN(n24416) );
  NAND2HSV0 U26764 ( .A1(n28478), .A2(n14072), .ZN(n24415) );
  XOR3HSV1 U26765 ( .A1(n24417), .A2(n24416), .A3(n24415), .Z(n24418) );
  XNOR2HSV1 U26766 ( .A1(n24419), .A2(n24418), .ZN(n24424) );
  NOR2HSV0 U26767 ( .A1(n24684), .A2(n24420), .ZN(n24423) );
  OR2HSV1 U26768 ( .A1(n24686), .A2(n24421), .Z(n24422) );
  XOR3HSV1 U26769 ( .A1(n24424), .A2(n24423), .A3(n24422), .Z(n24425) );
  XNOR2HSV1 U26770 ( .A1(n24426), .A2(n24425), .ZN(n24428) );
  NAND2HSV0 U26771 ( .A1(n28473), .A2(\pe5/got [3]), .ZN(n24447) );
  NAND2HSV0 U26772 ( .A1(\pe5/aot [1]), .A2(\pe5/bq[6] ), .ZN(n24438) );
  NAND2HSV0 U26773 ( .A1(\pe5/aot [6]), .A2(\pe5/bq[1] ), .ZN(n24437) );
  NOR2HSV0 U26774 ( .A1(n24440), .A2(n24439), .ZN(n24442) );
  NAND2HSV0 U26775 ( .A1(\pe5/aot [4]), .A2(\pe5/bq[3] ), .ZN(n24441) );
  CLKNAND2HSV0 U26776 ( .A1(n28803), .A2(\pe5/got [2]), .ZN(n24444) );
  XNOR2HSV1 U26777 ( .A1(n24445), .A2(n24444), .ZN(n24446) );
  XOR2HSV0 U26778 ( .A1(n24447), .A2(n24446), .Z(n24448) );
  NOR2HSV2 U26779 ( .A1(n24451), .A2(n26092), .ZN(n24498) );
  NOR2HSV2 U26780 ( .A1(n26093), .A2(n24452), .ZN(n24494) );
  NAND2HSV0 U26781 ( .A1(n28620), .A2(\pe10/got [5]), .ZN(n24488) );
  NOR2HSV0 U26782 ( .A1(n26159), .A2(n24453), .ZN(n24484) );
  NAND2HSV0 U26783 ( .A1(n28794), .A2(n27196), .ZN(n24480) );
  NAND2HSV0 U26784 ( .A1(\pe10/aot [3]), .A2(\pe10/bq[10] ), .ZN(n24455) );
  NAND2HSV0 U26785 ( .A1(\pe10/aot [1]), .A2(\pe10/bq[12] ), .ZN(n24454) );
  XOR2HSV0 U26786 ( .A1(n24455), .A2(n24454), .Z(n24459) );
  NAND2HSV0 U26787 ( .A1(\pe10/aot [10]), .A2(\pe10/bq[3] ), .ZN(n24457) );
  NAND2HSV0 U26788 ( .A1(\pe10/aot [4]), .A2(\pe10/bq[9] ), .ZN(n24456) );
  XOR2HSV0 U26789 ( .A1(n24457), .A2(n24456), .Z(n24458) );
  XOR2HSV0 U26790 ( .A1(n24459), .A2(n24458), .Z(n24470) );
  NAND2HSV0 U26791 ( .A1(\pe10/aot [8]), .A2(\pe10/bq[5] ), .ZN(n24461) );
  NAND2HSV0 U26792 ( .A1(\pe10/aot [9]), .A2(\pe10/bq[4] ), .ZN(n24460) );
  XOR2HSV0 U26793 ( .A1(n24461), .A2(n24460), .Z(n24468) );
  NOR2HSV0 U26794 ( .A1(n24463), .A2(n24462), .ZN(n26167) );
  CLKNHSV0 U26795 ( .I(\pe10/aot [12]), .ZN(n24464) );
  NOR2HSV0 U26796 ( .A1(n24464), .A2(n26163), .ZN(n24466) );
  NAND2HSV0 U26797 ( .A1(\pe10/aot [11]), .A2(\pe10/bq[1] ), .ZN(n25220) );
  OAI22HSV2 U26798 ( .A1(n26167), .A2(n24466), .B1(n25220), .B2(n24465), .ZN(
        n24467) );
  XNOR2HSV1 U26799 ( .A1(n24468), .A2(n24467), .ZN(n24469) );
  XNOR2HSV1 U26800 ( .A1(n24470), .A2(n24469), .ZN(n24478) );
  NAND2HSV0 U26801 ( .A1(\pe10/aot [6]), .A2(\pe10/bq[7] ), .ZN(n24472) );
  NAND2HSV0 U26802 ( .A1(\pe10/aot [5]), .A2(\pe10/bq[8] ), .ZN(n24471) );
  XOR2HSV0 U26803 ( .A1(n24472), .A2(n24471), .Z(n24476) );
  NAND2HSV0 U26804 ( .A1(\pe10/aot [7]), .A2(\pe10/bq[6] ), .ZN(n24473) );
  XOR2HSV0 U26805 ( .A1(n24474), .A2(n24473), .Z(n24475) );
  XOR2HSV0 U26806 ( .A1(n24476), .A2(n24475), .Z(n24477) );
  XNOR2HSV1 U26807 ( .A1(n24478), .A2(n24477), .ZN(n24479) );
  XNOR2HSV1 U26808 ( .A1(n24480), .A2(n24479), .ZN(n24482) );
  NOR2HSV0 U26809 ( .A1(n26200), .A2(n27194), .ZN(n24481) );
  XNOR2HSV1 U26810 ( .A1(n24482), .A2(n24481), .ZN(n24483) );
  XNOR2HSV1 U26811 ( .A1(n24484), .A2(n24483), .ZN(n24485) );
  XNOR2HSV1 U26812 ( .A1(n24486), .A2(n24485), .ZN(n24487) );
  XNOR2HSV1 U26813 ( .A1(n24488), .A2(n24487), .ZN(n24490) );
  NAND2HSV0 U26814 ( .A1(n28585), .A2(\pe10/got [6]), .ZN(n24489) );
  XOR2HSV0 U26815 ( .A1(n24490), .A2(n24489), .Z(n24492) );
  NAND2HSV0 U26816 ( .A1(n26209), .A2(\pe10/got [7]), .ZN(n24491) );
  XNOR2HSV1 U26817 ( .A1(n24492), .A2(n24491), .ZN(n24493) );
  XOR2HSV0 U26818 ( .A1(n24494), .A2(n24493), .Z(n24496) );
  NAND2HSV0 U26819 ( .A1(n27197), .A2(\pe10/got [9]), .ZN(n24495) );
  XOR2HSV0 U26820 ( .A1(n24496), .A2(n24495), .Z(n24497) );
  CLKNHSV1 U26821 ( .I(\pe3/got [4]), .ZN(n26333) );
  NOR2HSV2 U26822 ( .A1(n26681), .A2(n26333), .ZN(n24520) );
  NAND2HSV2 U26823 ( .A1(n24500), .A2(n24499), .ZN(n26297) );
  NAND2HSV0 U26824 ( .A1(n26297), .A2(\pe3/got [1]), .ZN(n24513) );
  NAND2HSV0 U26825 ( .A1(\pe3/aot [6]), .A2(\pe3/bq[2] ), .ZN(n24502) );
  NAND2HSV0 U26826 ( .A1(\pe3/aot [4]), .A2(\pe3/bq[4] ), .ZN(n24501) );
  XOR2HSV0 U26827 ( .A1(n24502), .A2(n24501), .Z(n24506) );
  NAND2HSV0 U26828 ( .A1(\pe3/aot [3]), .A2(\pe3/bq[5] ), .ZN(n24504) );
  NAND2HSV0 U26829 ( .A1(\pe3/aot [5]), .A2(\pe3/bq[3] ), .ZN(n24503) );
  XOR2HSV0 U26830 ( .A1(n24504), .A2(n24503), .Z(n24505) );
  XOR2HSV0 U26831 ( .A1(n24506), .A2(n24505), .Z(n24511) );
  NAND2HSV0 U26832 ( .A1(\pe3/aot [1]), .A2(\pe3/bq[7] ), .ZN(n24508) );
  NAND2HSV0 U26833 ( .A1(\pe3/aot [7]), .A2(\pe3/bq[1] ), .ZN(n24507) );
  XOR2HSV0 U26834 ( .A1(n24508), .A2(n24507), .Z(n24509) );
  NAND2HSV0 U26835 ( .A1(\pe3/aot [2]), .A2(\pe3/bq[6] ), .ZN(n26687) );
  XNOR2HSV1 U26836 ( .A1(n24509), .A2(n26687), .ZN(n24510) );
  XNOR2HSV1 U26837 ( .A1(n24511), .A2(n24510), .ZN(n24512) );
  XOR2HSV0 U26838 ( .A1(n24513), .A2(n24512), .Z(n24515) );
  NAND2HSV0 U26839 ( .A1(n26634), .A2(\pe3/got [2]), .ZN(n24514) );
  XOR2HSV0 U26840 ( .A1(n24515), .A2(n24514), .Z(n24518) );
  CLKNHSV0 U26841 ( .I(n24516), .ZN(n26637) );
  NAND2HSV0 U26842 ( .A1(n26637), .A2(n26751), .ZN(n24517) );
  XOR2HSV0 U26843 ( .A1(n24518), .A2(n24517), .Z(n24519) );
  CLKXOR2HSV4 U26844 ( .A1(n24520), .A2(n24519), .Z(n24521) );
  NAND2HSV2 U26845 ( .A1(n28661), .A2(n28628), .ZN(n24573) );
  NAND2HSV2 U26846 ( .A1(n24522), .A2(n11891), .ZN(n24571) );
  NOR2HSV2 U26847 ( .A1(n26681), .A2(n26645), .ZN(n24567) );
  NAND2HSV0 U26848 ( .A1(n26297), .A2(\pe3/got [7]), .ZN(n24561) );
  NAND2HSV0 U26849 ( .A1(n23327), .A2(\pe3/got [6]), .ZN(n24559) );
  NAND2HSV0 U26850 ( .A1(n28588), .A2(n26603), .ZN(n24557) );
  NAND2HSV0 U26851 ( .A1(n26682), .A2(\pe3/got [4]), .ZN(n24553) );
  NAND2HSV0 U26852 ( .A1(n15240), .A2(\pe3/got [2]), .ZN(n24551) );
  NAND2HSV0 U26853 ( .A1(n26242), .A2(\pe3/got [1]), .ZN(n24549) );
  NAND2HSV0 U26854 ( .A1(\pe3/aot [1]), .A2(\pe3/bq[13] ), .ZN(n24523) );
  XOR2HSV0 U26855 ( .A1(n24524), .A2(n24523), .Z(n24547) );
  NAND2HSV0 U26856 ( .A1(\pe3/aot [4]), .A2(\pe3/bq[10] ), .ZN(n24526) );
  NAND2HSV0 U26857 ( .A1(\pe3/aot [10]), .A2(\pe3/bq[4] ), .ZN(n24525) );
  XOR2HSV0 U26858 ( .A1(n24526), .A2(n24525), .Z(n24531) );
  CLKNHSV0 U26859 ( .I(\pe3/aot [3]), .ZN(n26247) );
  NOR2HSV0 U26860 ( .A1(n26247), .A2(n24527), .ZN(n24529) );
  NAND2HSV0 U26861 ( .A1(n11932), .A2(\pe3/bq[1] ), .ZN(n24528) );
  XOR2HSV0 U26862 ( .A1(n24529), .A2(n24528), .Z(n24530) );
  XNOR2HSV1 U26863 ( .A1(n24531), .A2(n24530), .ZN(n24546) );
  NAND2HSV0 U26864 ( .A1(\pe3/aot [5]), .A2(\pe3/bq[5] ), .ZN(n24587) );
  NOR2HSV0 U26865 ( .A1(n24532), .A2(n24587), .ZN(n24534) );
  AOI22HSV0 U26866 ( .A1(\pe3/aot [9]), .A2(\pe3/bq[5] ), .B1(\pe3/bq[9] ), 
        .B2(\pe3/aot [5]), .ZN(n24533) );
  NOR2HSV2 U26867 ( .A1(n24534), .A2(n24533), .ZN(n24537) );
  CLKNHSV0 U26868 ( .I(\pe3/aot [2]), .ZN(n24536) );
  NOR2HSV0 U26869 ( .A1(n24536), .A2(n24535), .ZN(n26307) );
  XOR2HSV0 U26870 ( .A1(n24537), .A2(n26307), .Z(n24545) );
  NAND2HSV0 U26871 ( .A1(\pe3/aot [8]), .A2(\pe3/bq[6] ), .ZN(n24539) );
  NAND2HSV0 U26872 ( .A1(\pe3/aot [6]), .A2(\pe3/bq[8] ), .ZN(n24538) );
  XOR2HSV0 U26873 ( .A1(n24539), .A2(n24538), .Z(n24543) );
  NAND2HSV0 U26874 ( .A1(\pe3/aot [11]), .A2(\pe3/bq[3] ), .ZN(n24541) );
  NAND2HSV0 U26875 ( .A1(\pe3/aot [12]), .A2(\pe3/bq[2] ), .ZN(n24540) );
  XOR2HSV0 U26876 ( .A1(n24541), .A2(n24540), .Z(n24542) );
  XOR2HSV0 U26877 ( .A1(n24543), .A2(n24542), .Z(n24544) );
  XOR4HSV1 U26878 ( .A1(n24547), .A2(n24546), .A3(n24545), .A4(n24544), .Z(
        n24548) );
  XNOR2HSV1 U26879 ( .A1(n24549), .A2(n24548), .ZN(n24550) );
  XNOR2HSV1 U26880 ( .A1(n24551), .A2(n24550), .ZN(n24552) );
  XNOR2HSV1 U26881 ( .A1(n24553), .A2(n24552), .ZN(n24555) );
  CLKNHSV1 U26882 ( .I(\pe3/got [3]), .ZN(n24610) );
  NOR2HSV0 U26883 ( .A1(n26714), .A2(n24610), .ZN(n24554) );
  XNOR2HSV1 U26884 ( .A1(n24555), .A2(n24554), .ZN(n24556) );
  XNOR2HSV1 U26885 ( .A1(n24557), .A2(n24556), .ZN(n24558) );
  XNOR2HSV1 U26886 ( .A1(n24559), .A2(n24558), .ZN(n24560) );
  XOR2HSV0 U26887 ( .A1(n24561), .A2(n24560), .Z(n24563) );
  NAND2HSV0 U26888 ( .A1(n26752), .A2(n28648), .ZN(n24562) );
  XOR2HSV0 U26889 ( .A1(n24563), .A2(n24562), .Z(n24565) );
  NAND2HSV0 U26890 ( .A1(n28584), .A2(n26642), .ZN(n24564) );
  XOR2HSV0 U26891 ( .A1(n24565), .A2(n24564), .Z(n24566) );
  CLKXOR2HSV4 U26892 ( .A1(n24567), .A2(n24566), .Z(n24570) );
  NAND2HSV0 U26893 ( .A1(n26759), .A2(\pe3/got [11]), .ZN(n24568) );
  INHSV2 U26894 ( .I(n24568), .ZN(n24569) );
  XOR2HSV0 U26895 ( .A1(n24573), .A2(n24572), .Z(\pe3/poht [3]) );
  NAND2HSV2 U26896 ( .A1(n26679), .A2(\pe3/got [2]), .ZN(n24579) );
  NAND2HSV2 U26897 ( .A1(n26760), .A2(\pe3/got [1]), .ZN(n24577) );
  NAND2HSV0 U26898 ( .A1(\pe3/aot [2]), .A2(\pe3/bq[1] ), .ZN(n24575) );
  NAND2HSV0 U26899 ( .A1(\pe3/aot [1]), .A2(\pe3/bq[2] ), .ZN(n24574) );
  XOR2HSV0 U26900 ( .A1(n24575), .A2(n24574), .Z(n24576) );
  XOR2HSV0 U26901 ( .A1(n24577), .A2(n24576), .Z(n24578) );
  XOR2HSV0 U26902 ( .A1(n24579), .A2(n24578), .Z(\pe3/poht [14]) );
  NAND2HSV2 U26903 ( .A1(n28661), .A2(\pe3/got [1]), .ZN(n24580) );
  NAND2HSV2 U26904 ( .A1(\pe3/bq[1] ), .A2(\pe3/aot [1]), .ZN(n26739) );
  XOR2HSV0 U26905 ( .A1(n24580), .A2(n26739), .Z(\pe3/poht [15]) );
  CLKNHSV0 U26906 ( .I(\pe3/got [6]), .ZN(n26397) );
  NOR2HSV2 U26907 ( .A1(n26730), .A2(n26397), .ZN(n24609) );
  NAND2HSV0 U26908 ( .A1(n26297), .A2(n26751), .ZN(n24603) );
  NAND2HSV0 U26909 ( .A1(n23327), .A2(\pe3/got [2]), .ZN(n24601) );
  CLKNAND2HSV0 U26910 ( .A1(n23328), .A2(\pe3/got [1]), .ZN(n24599) );
  NOR2HSV1 U26911 ( .A1(n24581), .A2(n23349), .ZN(n24583) );
  NAND2HSV0 U26912 ( .A1(\pe3/aot [1]), .A2(\pe3/bq[9] ), .ZN(n24582) );
  XOR2HSV0 U26913 ( .A1(n24583), .A2(n24582), .Z(n24597) );
  NAND2HSV0 U26914 ( .A1(\pe3/aot [9]), .A2(\pe3/bq[7] ), .ZN(n26265) );
  NOR2HSV0 U26915 ( .A1(n26265), .A2(n24584), .ZN(n24586) );
  AOI22HSV0 U26916 ( .A1(\pe3/aot [9]), .A2(\pe3/bq[1] ), .B1(\pe3/bq[7] ), 
        .B2(\pe3/aot [3]), .ZN(n24585) );
  NOR2HSV2 U26917 ( .A1(n24586), .A2(n24585), .ZN(n24588) );
  XOR2HSV0 U26918 ( .A1(n24588), .A2(n24587), .Z(n24596) );
  NAND2HSV0 U26919 ( .A1(\pe3/aot [7]), .A2(\pe3/bq[3] ), .ZN(n24590) );
  NAND2HSV0 U26920 ( .A1(\pe3/aot [2]), .A2(\pe3/bq[8] ), .ZN(n24589) );
  XOR2HSV0 U26921 ( .A1(n24590), .A2(n24589), .Z(n24594) );
  NAND2HSV0 U26922 ( .A1(\pe3/aot [8]), .A2(\pe3/bq[2] ), .ZN(n24592) );
  NAND2HSV0 U26923 ( .A1(\pe3/aot [4]), .A2(\pe3/bq[6] ), .ZN(n24591) );
  XOR2HSV0 U26924 ( .A1(n24592), .A2(n24591), .Z(n24593) );
  XOR2HSV0 U26925 ( .A1(n24594), .A2(n24593), .Z(n24595) );
  XOR3HSV2 U26926 ( .A1(n24597), .A2(n24596), .A3(n24595), .Z(n24598) );
  XNOR2HSV1 U26927 ( .A1(n24599), .A2(n24598), .ZN(n24600) );
  XNOR2HSV1 U26928 ( .A1(n24601), .A2(n24600), .ZN(n24602) );
  XOR2HSV0 U26929 ( .A1(n24603), .A2(n24602), .Z(n24605) );
  NAND2HSV0 U26930 ( .A1(n26752), .A2(\pe3/got [4]), .ZN(n24604) );
  XOR2HSV0 U26931 ( .A1(n24605), .A2(n24604), .Z(n24607) );
  XNOR2HSV1 U26932 ( .A1(n24607), .A2(n24606), .ZN(n24608) );
  NAND2HSV2 U26933 ( .A1(n26679), .A2(\pe3/got [6]), .ZN(n24633) );
  NOR2HSV2 U26934 ( .A1(n26730), .A2(n24610), .ZN(n24625) );
  NAND2HSV0 U26935 ( .A1(n26752), .A2(\pe3/got [1]), .ZN(n24621) );
  NAND2HSV0 U26936 ( .A1(\pe3/aot [1]), .A2(\pe3/bq[6] ), .ZN(n24612) );
  NAND2HSV0 U26937 ( .A1(\pe3/aot [6]), .A2(\pe3/bq[1] ), .ZN(n24611) );
  XOR2HSV0 U26938 ( .A1(n24612), .A2(n24611), .Z(n24616) );
  NAND2HSV0 U26939 ( .A1(\pe3/aot [5]), .A2(\pe3/bq[2] ), .ZN(n24614) );
  NAND2HSV0 U26940 ( .A1(\pe3/aot [3]), .A2(\pe3/bq[4] ), .ZN(n24613) );
  XOR2HSV0 U26941 ( .A1(n24614), .A2(n24613), .Z(n24615) );
  XOR2HSV0 U26942 ( .A1(n24616), .A2(n24615), .Z(n24619) );
  NAND2HSV0 U26943 ( .A1(\pe3/aot [2]), .A2(\pe3/bq[5] ), .ZN(n26604) );
  NAND2HSV0 U26944 ( .A1(\pe3/aot [4]), .A2(\pe3/bq[3] ), .ZN(n24617) );
  XOR2HSV0 U26945 ( .A1(n26604), .A2(n24617), .Z(n24618) );
  XNOR2HSV1 U26946 ( .A1(n24619), .A2(n24618), .ZN(n24620) );
  XOR2HSV0 U26947 ( .A1(n24621), .A2(n24620), .Z(n24623) );
  NAND2HSV0 U26948 ( .A1(\pe3/got [2]), .A2(n28584), .ZN(n24622) );
  XOR2HSV0 U26949 ( .A1(n24623), .A2(n24622), .Z(n24624) );
  NAND2HSV0 U26950 ( .A1(n28652), .A2(\pe3/got [4]), .ZN(n24626) );
  INHSV2 U26951 ( .I(n24628), .ZN(n24629) );
  INHSV4 U26952 ( .I(n24629), .ZN(n26729) );
  NAND2HSV2 U26953 ( .A1(n26603), .A2(n26729), .ZN(n24630) );
  XNOR2HSV4 U26954 ( .A1(n24631), .A2(n24630), .ZN(n24632) );
  XNOR2HSV4 U26955 ( .A1(n24633), .A2(n24632), .ZN(\pe3/poht [10]) );
  NAND2HSV2 U26956 ( .A1(n27112), .A2(n24634), .ZN(n24699) );
  NAND2HSV2 U26957 ( .A1(n12517), .A2(n14503), .ZN(n24696) );
  CLKNAND2HSV0 U26958 ( .A1(n21523), .A2(n28645), .ZN(n24682) );
  NAND2HSV0 U26959 ( .A1(n28594), .A2(\pe5/got [2]), .ZN(n24640) );
  NOR2HSV0 U26960 ( .A1(n27191), .A2(n24638), .ZN(n24639) );
  XNOR2HSV1 U26961 ( .A1(n24640), .A2(n24639), .ZN(n24671) );
  NAND2HSV0 U26962 ( .A1(\pe5/aot [5]), .A2(\pe5/bq[11] ), .ZN(n24642) );
  NAND2HSV0 U26963 ( .A1(\pe5/bq[2] ), .A2(\pe5/aot [14]), .ZN(n24641) );
  XOR2HSV0 U26964 ( .A1(n24642), .A2(n24641), .Z(n24646) );
  NAND2HSV0 U26965 ( .A1(\pe5/aot [11]), .A2(\pe5/bq[5] ), .ZN(n24644) );
  NAND2HSV0 U26966 ( .A1(\pe5/aot [12]), .A2(\pe5/bq[4] ), .ZN(n24643) );
  XOR2HSV0 U26967 ( .A1(n24644), .A2(n24643), .Z(n24645) );
  XOR2HSV0 U26968 ( .A1(n24646), .A2(n24645), .Z(n24655) );
  NAND2HSV0 U26969 ( .A1(\pe5/aot [6]), .A2(\pe5/bq[10] ), .ZN(n24649) );
  NAND2HSV0 U26970 ( .A1(\pe5/aot [1]), .A2(n24647), .ZN(n24648) );
  XOR2HSV0 U26971 ( .A1(n24649), .A2(n24648), .Z(n24653) );
  NAND2HSV0 U26972 ( .A1(\pe5/aot [3]), .A2(\pe5/bq[13] ), .ZN(n24650) );
  XOR2HSV0 U26973 ( .A1(n24651), .A2(n24650), .Z(n24652) );
  XOR2HSV0 U26974 ( .A1(n24653), .A2(n24652), .Z(n24654) );
  XOR2HSV0 U26975 ( .A1(n24655), .A2(n24654), .Z(n24669) );
  NAND2HSV0 U26976 ( .A1(\pe5/aot [7]), .A2(\pe5/bq[9] ), .ZN(n24657) );
  NAND2HSV0 U26977 ( .A1(n14031), .A2(\pe5/bq[1] ), .ZN(n24656) );
  XOR2HSV0 U26978 ( .A1(n24657), .A2(n24656), .Z(n24661) );
  NAND2HSV0 U26979 ( .A1(\pe5/aot [8]), .A2(\pe5/bq[8] ), .ZN(n24659) );
  INAND2HSV0 U26980 ( .A1(n14766), .B1(\pe5/aot [4]), .ZN(n24658) );
  XOR2HSV0 U26981 ( .A1(n24659), .A2(n24658), .Z(n24660) );
  XOR2HSV0 U26982 ( .A1(n24661), .A2(n24660), .Z(n24667) );
  NAND2HSV0 U26983 ( .A1(\pe5/aot [10]), .A2(\pe5/bq[6] ), .ZN(n24663) );
  NAND2HSV0 U26984 ( .A1(\pe5/aot [2]), .A2(\pe5/bq[14] ), .ZN(n24662) );
  XOR2HSV0 U26985 ( .A1(n24663), .A2(n24662), .Z(n24665) );
  XNOR2HSV1 U26986 ( .A1(n24665), .A2(n24664), .ZN(n24666) );
  XNOR2HSV1 U26987 ( .A1(n24667), .A2(n24666), .ZN(n24668) );
  XNOR2HSV1 U26988 ( .A1(n24669), .A2(n24668), .ZN(n24670) );
  XNOR2HSV1 U26989 ( .A1(n24671), .A2(n24670), .ZN(n24673) );
  NAND2HSV0 U26990 ( .A1(n28614), .A2(\pe5/got [3]), .ZN(n24672) );
  XNOR2HSV1 U26991 ( .A1(n24673), .A2(n24672), .ZN(n24676) );
  NAND2HSV0 U26992 ( .A1(n24674), .A2(n13993), .ZN(n24675) );
  XNOR2HSV1 U26993 ( .A1(n24676), .A2(n24675), .ZN(n24680) );
  NOR2HSV0 U26994 ( .A1(n25350), .A2(n24677), .ZN(n24679) );
  NAND2HSV0 U26995 ( .A1(n28478), .A2(n28647), .ZN(n24678) );
  XOR3HSV1 U26996 ( .A1(n24680), .A2(n24679), .A3(n24678), .Z(n24681) );
  XNOR2HSV1 U26997 ( .A1(n24682), .A2(n24681), .ZN(n24689) );
  NOR2HSV2 U26998 ( .A1(n24684), .A2(n24683), .ZN(n24688) );
  OR2HSV1 U26999 ( .A1(n24686), .A2(n24685), .Z(n24687) );
  XOR3HSV2 U27000 ( .A1(n24689), .A2(n24688), .A3(n24687), .Z(n24690) );
  NAND2HSV0 U27001 ( .A1(n28803), .A2(\pe5/got [11]), .ZN(n24691) );
  XNOR2HSV1 U27002 ( .A1(n24692), .A2(n24691), .ZN(n24693) );
  XOR2HSV0 U27003 ( .A1(n24694), .A2(n24693), .Z(n24695) );
  NAND2HSV0 U27004 ( .A1(n14063), .A2(\pe11/got [8]), .ZN(n24738) );
  NAND2HSV0 U27005 ( .A1(n25138), .A2(\pe11/got [6]), .ZN(n24734) );
  NAND2HSV0 U27006 ( .A1(n25139), .A2(\pe11/got [5]), .ZN(n24732) );
  NAND2HSV0 U27007 ( .A1(n28471), .A2(\pe11/got [4]), .ZN(n24730) );
  NAND2HSV0 U27008 ( .A1(n14043), .A2(\pe11/got [3]), .ZN(n24728) );
  NAND2HSV0 U27009 ( .A1(\pe11/got [2]), .A2(n11804), .ZN(n24726) );
  NAND2HSV0 U27010 ( .A1(n25008), .A2(\pe11/got [1]), .ZN(n24724) );
  NAND2HSV0 U27011 ( .A1(\pe11/bq[12] ), .A2(\pe11/aot [2]), .ZN(n24701) );
  NAND2HSV0 U27012 ( .A1(\pe11/bq[1] ), .A2(n12011), .ZN(n24700) );
  XOR2HSV0 U27013 ( .A1(n24701), .A2(n24700), .Z(n24705) );
  NAND2HSV0 U27014 ( .A1(\pe11/bq[13] ), .A2(\pe11/aot [1]), .ZN(n24703) );
  NAND2HSV0 U27015 ( .A1(\pe11/bq[2] ), .A2(\pe11/aot [12]), .ZN(n24702) );
  XOR2HSV0 U27016 ( .A1(n24703), .A2(n24702), .Z(n24704) );
  XOR2HSV0 U27017 ( .A1(n24705), .A2(n24704), .Z(n24713) );
  NAND2HSV0 U27018 ( .A1(\pe11/bq[11] ), .A2(\pe11/aot [3]), .ZN(n24707) );
  NAND2HSV0 U27019 ( .A1(\pe11/bq[9] ), .A2(\pe11/aot [5]), .ZN(n24706) );
  XOR2HSV0 U27020 ( .A1(n24707), .A2(n24706), .Z(n24711) );
  NAND2HSV0 U27021 ( .A1(\pe11/bq[5] ), .A2(\pe11/aot [9]), .ZN(n24709) );
  NAND2HSV0 U27022 ( .A1(\pe11/bq[4] ), .A2(\pe11/aot [10]), .ZN(n24708) );
  XOR2HSV0 U27023 ( .A1(n24709), .A2(n24708), .Z(n24710) );
  XOR2HSV0 U27024 ( .A1(n24711), .A2(n24710), .Z(n24712) );
  XOR2HSV0 U27025 ( .A1(n24713), .A2(n24712), .Z(n24722) );
  NAND2HSV0 U27026 ( .A1(\pe11/bq[6] ), .A2(\pe11/aot [8]), .ZN(n24714) );
  XOR2HSV0 U27027 ( .A1(n24715), .A2(n24714), .Z(n24719) );
  NAND2HSV0 U27028 ( .A1(\pe11/bq[10] ), .A2(\pe11/aot [4]), .ZN(n24717) );
  NAND2HSV0 U27029 ( .A1(\pe11/bq[8] ), .A2(\pe11/aot [6]), .ZN(n24716) );
  XOR2HSV0 U27030 ( .A1(n24717), .A2(n24716), .Z(n24718) );
  XOR3HSV1 U27031 ( .A1(n24720), .A2(n24719), .A3(n24718), .Z(n24721) );
  XNOR2HSV1 U27032 ( .A1(n24722), .A2(n24721), .ZN(n24723) );
  XNOR2HSV1 U27033 ( .A1(n24724), .A2(n24723), .ZN(n24725) );
  XNOR2HSV1 U27034 ( .A1(n24726), .A2(n24725), .ZN(n24727) );
  XOR2HSV0 U27035 ( .A1(n24728), .A2(n24727), .Z(n24729) );
  XOR2HSV0 U27036 ( .A1(n24730), .A2(n24729), .Z(n24731) );
  XOR2HSV0 U27037 ( .A1(n24732), .A2(n24731), .Z(n24733) );
  XOR2HSV0 U27038 ( .A1(n24734), .A2(n24733), .Z(n24736) );
  NAND2HSV0 U27039 ( .A1(n28464), .A2(\pe11/got [7]), .ZN(n24735) );
  XOR2HSV0 U27040 ( .A1(n24736), .A2(n24735), .Z(n24737) );
  XOR2HSV0 U27041 ( .A1(n24738), .A2(n24737), .Z(n24739) );
  NAND2HSV0 U27042 ( .A1(n28919), .A2(\pe11/got [10]), .ZN(n24741) );
  NAND2HSV2 U27043 ( .A1(n25414), .A2(n14049), .ZN(n24746) );
  CLKNAND2HSV1 U27044 ( .A1(n25182), .A2(n20292), .ZN(n24745) );
  XOR3HSV2 U27045 ( .A1(n24747), .A2(n24746), .A3(n24745), .Z(\pe11/poht [3])
         );
  NAND2HSV0 U27046 ( .A1(n28918), .A2(\pe11/got [11]), .ZN(n24799) );
  NAND2HSV0 U27047 ( .A1(n14063), .A2(\pe11/got [10]), .ZN(n24797) );
  NAND2HSV0 U27048 ( .A1(n25138), .A2(\pe11/got [8]), .ZN(n24793) );
  NAND2HSV0 U27049 ( .A1(n25139), .A2(\pe11/got [7]), .ZN(n24791) );
  NAND2HSV0 U27050 ( .A1(n28471), .A2(\pe11/got [6]), .ZN(n24789) );
  NAND2HSV0 U27051 ( .A1(n25008), .A2(\pe11/got [3]), .ZN(n24785) );
  NAND2HSV0 U27052 ( .A1(n20506), .A2(\pe11/got [2]), .ZN(n24749) );
  NAND2HSV0 U27053 ( .A1(n28629), .A2(\pe11/got [1]), .ZN(n24748) );
  XOR2HSV0 U27054 ( .A1(n24749), .A2(n24748), .Z(n24782) );
  NAND2HSV0 U27055 ( .A1(\pe11/bq[5] ), .A2(\pe11/aot [11]), .ZN(n24751) );
  NAND2HSV0 U27056 ( .A1(\pe11/bq[3] ), .A2(n12011), .ZN(n24750) );
  XOR2HSV0 U27057 ( .A1(n24751), .A2(n24750), .Z(n24755) );
  NAND2HSV0 U27058 ( .A1(\pe11/bq[6] ), .A2(\pe11/aot [10]), .ZN(n24753) );
  NAND2HSV0 U27059 ( .A1(\pe11/bq[12] ), .A2(\pe11/aot [4]), .ZN(n24752) );
  XOR2HSV0 U27060 ( .A1(n24753), .A2(n24752), .Z(n24754) );
  XOR2HSV0 U27061 ( .A1(n24755), .A2(n24754), .Z(n24763) );
  NAND2HSV0 U27062 ( .A1(\pe11/bq[11] ), .A2(\pe11/aot [5]), .ZN(n24757) );
  NAND2HSV0 U27063 ( .A1(\pe11/bq[8] ), .A2(\pe11/aot [8]), .ZN(n24756) );
  XOR2HSV0 U27064 ( .A1(n24757), .A2(n24756), .Z(n24761) );
  NAND2HSV0 U27065 ( .A1(\pe11/bq[4] ), .A2(\pe11/aot [12]), .ZN(n24759) );
  NAND2HSV0 U27066 ( .A1(\pe11/bq[13] ), .A2(\pe11/aot [3]), .ZN(n24758) );
  XOR2HSV0 U27067 ( .A1(n24759), .A2(n24758), .Z(n24760) );
  XOR2HSV0 U27068 ( .A1(n24761), .A2(n24760), .Z(n24762) );
  XOR2HSV0 U27069 ( .A1(n24763), .A2(n24762), .Z(n24780) );
  AO22HSV2 U27070 ( .A1(\pe11/bq[14] ), .A2(\pe11/aot [2]), .B1(\pe11/bq[9] ), 
        .B2(\pe11/aot [7]), .Z(n24764) );
  OAI21HSV0 U27071 ( .A1(n24766), .A2(n24765), .B(n24764), .ZN(n24778) );
  NAND2HSV0 U27072 ( .A1(n24994), .A2(\pe11/bq[1] ), .ZN(n24768) );
  NAND2HSV0 U27073 ( .A1(\pe11/bq[7] ), .A2(\pe11/aot [9]), .ZN(n24767) );
  XOR2HSV0 U27074 ( .A1(n24768), .A2(n24767), .Z(n24777) );
  NOR2HSV0 U27075 ( .A1(n24770), .A2(n24769), .ZN(n24773) );
  AOI22HSV0 U27076 ( .A1(\pe11/bq[10] ), .A2(\pe11/aot [6]), .B1(n24771), .B2(
        \pe11/bq[2] ), .ZN(n24772) );
  NOR2HSV2 U27077 ( .A1(n24773), .A2(n24772), .ZN(n24775) );
  NAND2HSV0 U27078 ( .A1(n24997), .A2(\pe11/aot [1]), .ZN(n24774) );
  XNOR2HSV1 U27079 ( .A1(n24775), .A2(n24774), .ZN(n24776) );
  XOR3HSV2 U27080 ( .A1(n24778), .A2(n24777), .A3(n24776), .Z(n24779) );
  XNOR2HSV1 U27081 ( .A1(n24780), .A2(n24779), .ZN(n24781) );
  XOR2HSV0 U27082 ( .A1(n24782), .A2(n24781), .Z(n24784) );
  NAND2HSV0 U27083 ( .A1(n11804), .A2(\pe11/got [4]), .ZN(n24783) );
  XOR3HSV2 U27084 ( .A1(n24785), .A2(n24784), .A3(n24783), .Z(n24787) );
  NAND2HSV0 U27085 ( .A1(n14043), .A2(\pe11/got [5]), .ZN(n24786) );
  XOR2HSV0 U27086 ( .A1(n24787), .A2(n24786), .Z(n24788) );
  XNOR2HSV1 U27087 ( .A1(n24789), .A2(n24788), .ZN(n24790) );
  XNOR2HSV1 U27088 ( .A1(n24791), .A2(n24790), .ZN(n24792) );
  XNOR2HSV1 U27089 ( .A1(n24793), .A2(n24792), .ZN(n24795) );
  NAND2HSV0 U27090 ( .A1(n28464), .A2(\pe11/got [9]), .ZN(n24794) );
  XOR2HSV0 U27091 ( .A1(n24795), .A2(n24794), .Z(n24796) );
  XOR2HSV0 U27092 ( .A1(n24797), .A2(n24796), .Z(n24798) );
  XNOR2HSV1 U27093 ( .A1(n24799), .A2(n24798), .ZN(n24802) );
  XNOR2HSV1 U27094 ( .A1(n24802), .A2(n24801), .ZN(n24803) );
  NAND2HSV2 U27095 ( .A1(n24902), .A2(n25030), .ZN(n24806) );
  CLKNAND2HSV1 U27096 ( .A1(n28927), .A2(n25504), .ZN(n24805) );
  XOR3HSV2 U27097 ( .A1(n24807), .A2(n24806), .A3(n24805), .Z(\pe11/poht [1])
         );
  NAND2HSV0 U27098 ( .A1(n25137), .A2(\pe11/got [8]), .ZN(n24845) );
  NAND2HSV0 U27099 ( .A1(n14063), .A2(\pe11/got [7]), .ZN(n24843) );
  NAND2HSV0 U27100 ( .A1(n28935), .A2(\pe11/got [5]), .ZN(n24839) );
  NAND2HSV0 U27101 ( .A1(n25139), .A2(\pe11/got [4]), .ZN(n24837) );
  NAND2HSV0 U27102 ( .A1(n28471), .A2(\pe11/got [3]), .ZN(n24835) );
  NAND2HSV0 U27103 ( .A1(\pe11/bq[6] ), .A2(\pe11/aot [7]), .ZN(n24809) );
  NAND2HSV0 U27104 ( .A1(\pe11/bq[11] ), .A2(\pe11/aot [2]), .ZN(n24808) );
  XOR2HSV0 U27105 ( .A1(n24809), .A2(n24808), .Z(n24813) );
  NAND2HSV0 U27106 ( .A1(\pe11/bq[3] ), .A2(\pe11/aot [10]), .ZN(n24811) );
  NAND2HSV0 U27107 ( .A1(\pe11/bq[9] ), .A2(\pe11/aot [4]), .ZN(n24810) );
  XOR2HSV0 U27108 ( .A1(n24811), .A2(n24810), .Z(n24812) );
  XOR2HSV0 U27109 ( .A1(n24813), .A2(n24812), .Z(n24830) );
  NAND2HSV0 U27110 ( .A1(\pe11/bq[8] ), .A2(\pe11/aot [5]), .ZN(n24815) );
  NAND2HSV0 U27111 ( .A1(\pe11/bq[7] ), .A2(\pe11/aot [6]), .ZN(n24814) );
  XOR2HSV0 U27112 ( .A1(n24815), .A2(n24814), .Z(n24819) );
  NAND2HSV0 U27113 ( .A1(\pe11/aot [1]), .A2(\pe11/bq[12] ), .ZN(n24817) );
  NAND2HSV0 U27114 ( .A1(\pe11/bq[10] ), .A2(\pe11/aot [3]), .ZN(n24816) );
  XOR2HSV0 U27115 ( .A1(n24817), .A2(n24816), .Z(n24818) );
  XOR2HSV0 U27116 ( .A1(n24819), .A2(n24818), .Z(n24827) );
  NAND2HSV0 U27117 ( .A1(\pe11/bq[4] ), .A2(\pe11/aot [9]), .ZN(n24821) );
  NAND2HSV0 U27118 ( .A1(\pe11/bq[5] ), .A2(\pe11/aot [8]), .ZN(n24820) );
  XOR2HSV0 U27119 ( .A1(n24821), .A2(n24820), .Z(n24825) );
  NAND2HSV0 U27120 ( .A1(\pe11/bq[1] ), .A2(\pe11/aot [12]), .ZN(n24823) );
  NAND2HSV0 U27121 ( .A1(\pe11/bq[2] ), .A2(\pe11/aot [11]), .ZN(n24822) );
  XOR2HSV0 U27122 ( .A1(n24823), .A2(n24822), .Z(n24824) );
  XOR2HSV0 U27123 ( .A1(n24825), .A2(n24824), .Z(n24826) );
  XOR2HSV0 U27124 ( .A1(n24827), .A2(n24826), .Z(n24829) );
  NAND2HSV0 U27125 ( .A1(n20467), .A2(\pe11/got [1]), .ZN(n24828) );
  XOR3HSV2 U27126 ( .A1(n24830), .A2(n24829), .A3(n24828), .Z(n24833) );
  CLKNHSV0 U27127 ( .I(n24831), .ZN(n25140) );
  NAND2HSV0 U27128 ( .A1(n25140), .A2(\pe11/got [2]), .ZN(n24832) );
  XOR2HSV0 U27129 ( .A1(n24833), .A2(n24832), .Z(n24834) );
  XNOR2HSV1 U27130 ( .A1(n24835), .A2(n24834), .ZN(n24836) );
  XNOR2HSV1 U27131 ( .A1(n24837), .A2(n24836), .ZN(n24838) );
  XNOR2HSV1 U27132 ( .A1(n24839), .A2(n24838), .ZN(n24841) );
  NAND2HSV0 U27133 ( .A1(n28464), .A2(\pe11/got [6]), .ZN(n24840) );
  XOR2HSV0 U27134 ( .A1(n24841), .A2(n24840), .Z(n24842) );
  XNOR2HSV1 U27135 ( .A1(n24843), .A2(n24842), .ZN(n24844) );
  XNOR2HSV1 U27136 ( .A1(n24845), .A2(n24844), .ZN(n24847) );
  NAND2HSV2 U27137 ( .A1(n28936), .A2(\pe11/got [11]), .ZN(n24851) );
  CLKNAND2HSV1 U27138 ( .A1(n24957), .A2(\pe11/got [12]), .ZN(n24850) );
  XOR3HSV2 U27139 ( .A1(n24852), .A2(n24851), .A3(n24850), .Z(\pe11/poht [4])
         );
  NAND2HSV2 U27140 ( .A1(n24902), .A2(\pe11/got [7]), .ZN(n24880) );
  NAND2HSV0 U27141 ( .A1(n14064), .A2(\pe11/got [3]), .ZN(n24872) );
  NAND2HSV0 U27142 ( .A1(n25138), .A2(\pe11/got [1]), .ZN(n24868) );
  NAND2HSV0 U27143 ( .A1(\pe11/bq[3] ), .A2(\pe11/aot [6]), .ZN(n24854) );
  NAND2HSV0 U27144 ( .A1(\pe11/bq[6] ), .A2(\pe11/aot [3]), .ZN(n24853) );
  XOR2HSV0 U27145 ( .A1(n24854), .A2(n24853), .Z(n24858) );
  NAND2HSV0 U27146 ( .A1(\pe11/bq[2] ), .A2(\pe11/aot [7]), .ZN(n24856) );
  NAND2HSV0 U27147 ( .A1(\pe11/bq[8] ), .A2(\pe11/aot [1]), .ZN(n24855) );
  XOR2HSV0 U27148 ( .A1(n24856), .A2(n24855), .Z(n24857) );
  XOR2HSV0 U27149 ( .A1(n24858), .A2(n24857), .Z(n24866) );
  NAND2HSV0 U27150 ( .A1(\pe11/bq[7] ), .A2(\pe11/aot [2]), .ZN(n24860) );
  NAND2HSV0 U27151 ( .A1(\pe11/bq[1] ), .A2(\pe11/aot [8]), .ZN(n24859) );
  XOR2HSV0 U27152 ( .A1(n24860), .A2(n24859), .Z(n24864) );
  NAND2HSV0 U27153 ( .A1(\pe11/bq[5] ), .A2(\pe11/aot [4]), .ZN(n24862) );
  NAND2HSV0 U27154 ( .A1(\pe11/bq[4] ), .A2(\pe11/aot [5]), .ZN(n24861) );
  XOR2HSV0 U27155 ( .A1(n24862), .A2(n24861), .Z(n24863) );
  XOR2HSV0 U27156 ( .A1(n24864), .A2(n24863), .Z(n24865) );
  XOR2HSV0 U27157 ( .A1(n24866), .A2(n24865), .Z(n24867) );
  XNOR2HSV1 U27158 ( .A1(n24868), .A2(n24867), .ZN(n24870) );
  CLKNAND2HSV0 U27159 ( .A1(n28464), .A2(\pe11/got [2]), .ZN(n24869) );
  XOR2HSV0 U27160 ( .A1(n24870), .A2(n24869), .Z(n24871) );
  XOR2HSV0 U27161 ( .A1(n24872), .A2(n24871), .Z(n24873) );
  XNOR2HSV1 U27162 ( .A1(n24874), .A2(n24873), .ZN(n24876) );
  XNOR2HSV4 U27163 ( .A1(n24880), .A2(n24879), .ZN(n24892) );
  AND2HSV2 U27164 ( .A1(n24881), .A2(n20561), .Z(n24882) );
  NOR2HSV1 U27165 ( .A1(n24882), .A2(n25415), .ZN(n24890) );
  NAND2HSV0 U27166 ( .A1(n24883), .A2(\pe11/got [8]), .ZN(n24886) );
  CLKNHSV0 U27167 ( .I(\pe11/got [8]), .ZN(n24885) );
  OAI22HSV1 U27168 ( .A1(n24887), .A2(n24886), .B1(n24885), .B2(n24884), .ZN(
        n24888) );
  AOI31HSV2 U27169 ( .A1(\pe11/got [8]), .A2(n24890), .A3(n24889), .B(n24888), 
        .ZN(n24891) );
  XNOR2HSV4 U27170 ( .A1(n24892), .A2(n24891), .ZN(\pe11/poht [8]) );
  NAND2HSV0 U27171 ( .A1(n28919), .A2(\pe11/got [1]), .ZN(n24901) );
  NAND2HSV0 U27172 ( .A1(\pe11/bq[4] ), .A2(\pe11/aot [1]), .ZN(n24895) );
  NAND2HSV0 U27173 ( .A1(\pe11/bq[1] ), .A2(\pe11/aot [4]), .ZN(n24894) );
  XOR2HSV0 U27174 ( .A1(n24895), .A2(n24894), .Z(n24899) );
  NAND2HSV0 U27175 ( .A1(\pe11/bq[2] ), .A2(\pe11/aot [3]), .ZN(n24897) );
  NAND2HSV0 U27176 ( .A1(\pe11/bq[3] ), .A2(\pe11/aot [2]), .ZN(n24896) );
  XOR2HSV0 U27177 ( .A1(n24897), .A2(n24896), .Z(n24898) );
  XOR2HSV0 U27178 ( .A1(n24899), .A2(n24898), .Z(n24900) );
  NAND2HSV2 U27179 ( .A1(n24902), .A2(\pe11/got [5]), .ZN(n24923) );
  NAND2HSV2 U27180 ( .A1(n24903), .A2(\pe11/got [4]), .ZN(n24921) );
  NAND2HSV0 U27181 ( .A1(n25137), .A2(\pe11/got [2]), .ZN(n24917) );
  NAND2HSV0 U27182 ( .A1(n14064), .A2(\pe11/got [1]), .ZN(n24915) );
  NAND2HSV0 U27183 ( .A1(\pe11/bq[6] ), .A2(\pe11/aot [1]), .ZN(n24905) );
  NAND2HSV0 U27184 ( .A1(\pe11/bq[5] ), .A2(\pe11/aot [2]), .ZN(n24904) );
  XOR2HSV0 U27185 ( .A1(n24905), .A2(n24904), .Z(n24909) );
  NAND2HSV0 U27186 ( .A1(\pe11/bq[4] ), .A2(\pe11/aot [3]), .ZN(n24907) );
  NAND2HSV0 U27187 ( .A1(\pe11/bq[3] ), .A2(\pe11/aot [4]), .ZN(n24906) );
  XOR2HSV0 U27188 ( .A1(n24907), .A2(n24906), .Z(n24908) );
  XOR2HSV0 U27189 ( .A1(n24909), .A2(n24908), .Z(n24913) );
  NAND2HSV0 U27190 ( .A1(\pe11/bq[2] ), .A2(\pe11/aot [5]), .ZN(n24911) );
  NAND2HSV0 U27191 ( .A1(\pe11/bq[1] ), .A2(\pe11/aot [6]), .ZN(n24910) );
  XOR2HSV0 U27192 ( .A1(n24911), .A2(n24910), .Z(n24912) );
  XNOR2HSV1 U27193 ( .A1(n24913), .A2(n24912), .ZN(n24914) );
  XOR2HSV0 U27194 ( .A1(n24915), .A2(n24914), .Z(n24916) );
  XNOR2HSV1 U27195 ( .A1(n24917), .A2(n24916), .ZN(n24919) );
  NAND2HSV0 U27196 ( .A1(n28919), .A2(\pe11/got [3]), .ZN(n24918) );
  XNOR2HSV4 U27197 ( .A1(n24923), .A2(n24922), .ZN(n24925) );
  CLKNAND2HSV1 U27198 ( .A1(n28927), .A2(\pe11/got [6]), .ZN(n24924) );
  XNOR2HSV4 U27199 ( .A1(n24925), .A2(n24924), .ZN(\pe11/poht [10]) );
  NAND2HSV2 U27200 ( .A1(n25414), .A2(\pe11/got [8]), .ZN(n24956) );
  CLKNAND2HSV1 U27201 ( .A1(n24965), .A2(\pe11/got [5]), .ZN(n24950) );
  NAND2HSV0 U27202 ( .A1(n14064), .A2(\pe11/got [4]), .ZN(n24948) );
  NAND2HSV0 U27203 ( .A1(\pe11/got [2]), .A2(n25138), .ZN(n24944) );
  NAND2HSV0 U27204 ( .A1(n25139), .A2(\pe11/got [1]), .ZN(n24942) );
  NAND2HSV0 U27205 ( .A1(\pe11/bq[2] ), .A2(\pe11/aot [8]), .ZN(n24927) );
  NAND2HSV0 U27206 ( .A1(\pe11/bq[4] ), .A2(\pe11/aot [6]), .ZN(n24926) );
  XOR2HSV0 U27207 ( .A1(n24927), .A2(n24926), .Z(n24940) );
  NAND2HSV0 U27208 ( .A1(\pe11/bq[6] ), .A2(\pe11/aot [4]), .ZN(n24929) );
  NAND2HSV0 U27209 ( .A1(\pe11/bq[5] ), .A2(\pe11/aot [5]), .ZN(n24928) );
  XOR2HSV0 U27210 ( .A1(n24929), .A2(n24928), .Z(n24931) );
  NAND2HSV0 U27211 ( .A1(\pe11/bq[7] ), .A2(\pe11/aot [3]), .ZN(n24930) );
  XNOR2HSV1 U27212 ( .A1(n24931), .A2(n24930), .ZN(n24939) );
  NAND2HSV0 U27213 ( .A1(\pe11/bq[9] ), .A2(\pe11/aot [1]), .ZN(n24933) );
  NAND2HSV0 U27214 ( .A1(\pe11/bq[3] ), .A2(\pe11/aot [7]), .ZN(n24932) );
  XOR2HSV0 U27215 ( .A1(n24933), .A2(n24932), .Z(n24937) );
  NAND2HSV0 U27216 ( .A1(\pe11/bq[8] ), .A2(\pe11/aot [2]), .ZN(n24935) );
  NAND2HSV0 U27217 ( .A1(\pe11/bq[1] ), .A2(\pe11/aot [9]), .ZN(n24934) );
  XOR2HSV0 U27218 ( .A1(n24935), .A2(n24934), .Z(n24936) );
  XOR2HSV0 U27219 ( .A1(n24937), .A2(n24936), .Z(n24938) );
  XOR3HSV2 U27220 ( .A1(n24940), .A2(n24939), .A3(n24938), .Z(n24941) );
  XNOR2HSV1 U27221 ( .A1(n24942), .A2(n24941), .ZN(n24943) );
  XNOR2HSV1 U27222 ( .A1(n24944), .A2(n24943), .ZN(n24946) );
  NAND2HSV0 U27223 ( .A1(n25169), .A2(\pe11/got [3]), .ZN(n24945) );
  XOR2HSV0 U27224 ( .A1(n24946), .A2(n24945), .Z(n24947) );
  XOR2HSV0 U27225 ( .A1(n24948), .A2(n24947), .Z(n24949) );
  XNOR2HSV1 U27226 ( .A1(n24950), .A2(n24949), .ZN(n24952) );
  NAND2HSV0 U27227 ( .A1(n28919), .A2(\pe11/got [6]), .ZN(n24951) );
  XOR2HSV0 U27228 ( .A1(n24952), .A2(n24951), .Z(n24953) );
  XNOR2HSV4 U27229 ( .A1(n24956), .A2(n24955), .ZN(n24959) );
  XNOR2HSV4 U27230 ( .A1(n24959), .A2(n24958), .ZN(\pe11/poht [7]) );
  XNOR2HSV1 U27231 ( .A1(n12298), .A2(n24960), .ZN(n29015) );
  CLKNAND2HSV1 U27232 ( .A1(n24965), .A2(\pe11/got [12]), .ZN(n25025) );
  NAND2HSV0 U27233 ( .A1(n14064), .A2(\pe11/got [11]), .ZN(n25023) );
  NAND2HSV0 U27234 ( .A1(n25138), .A2(\pe11/got [9]), .ZN(n25019) );
  NAND2HSV0 U27235 ( .A1(n25139), .A2(\pe11/got [8]), .ZN(n25017) );
  NAND2HSV0 U27236 ( .A1(n28471), .A2(\pe11/got [7]), .ZN(n25015) );
  NAND2HSV0 U27237 ( .A1(n11804), .A2(\pe11/got [5]), .ZN(n25013) );
  NAND2HSV0 U27238 ( .A1(\pe11/bq[3] ), .A2(\pe11/aot [14]), .ZN(n24968) );
  NAND2HSV0 U27239 ( .A1(\pe11/bq[6] ), .A2(\pe11/aot [11]), .ZN(n24967) );
  XOR2HSV0 U27240 ( .A1(n24968), .A2(n24967), .Z(n24972) );
  NAND2HSV0 U27241 ( .A1(\pe11/bq[7] ), .A2(\pe11/aot [10]), .ZN(n24970) );
  NAND2HSV0 U27242 ( .A1(\pe11/bq[11] ), .A2(\pe11/aot [6]), .ZN(n24969) );
  XOR2HSV0 U27243 ( .A1(n24970), .A2(n24969), .Z(n24971) );
  XOR2HSV0 U27244 ( .A1(n24972), .A2(n24971), .Z(n24987) );
  NAND2HSV0 U27245 ( .A1(\pe11/bq[9] ), .A2(\pe11/aot [8]), .ZN(n24974) );
  NAND2HSV0 U27246 ( .A1(\pe11/bq[14] ), .A2(\pe11/aot [3]), .ZN(n24973) );
  XOR2HSV0 U27247 ( .A1(n24974), .A2(n24973), .Z(n24979) );
  NAND2HSV0 U27248 ( .A1(\pe11/bq[12] ), .A2(\pe11/aot [5]), .ZN(n24977) );
  NAND2HSV0 U27249 ( .A1(n24975), .A2(\pe11/got [1]), .ZN(n24976) );
  XOR2HSV0 U27250 ( .A1(n24977), .A2(n24976), .Z(n24978) );
  XNOR2HSV1 U27251 ( .A1(n24979), .A2(n24978), .ZN(n24984) );
  NAND2HSV0 U27252 ( .A1(n24980), .A2(\pe11/pq ), .ZN(n24982) );
  NAND2HSV0 U27253 ( .A1(n27058), .A2(\pe11/aot [1]), .ZN(n24981) );
  XOR2HSV0 U27254 ( .A1(n24982), .A2(n24981), .Z(n24983) );
  XNOR2HSV1 U27255 ( .A1(n24984), .A2(n24983), .ZN(n24986) );
  NAND2HSV0 U27256 ( .A1(n20506), .A2(\pe11/got [3]), .ZN(n24985) );
  XOR3HSV2 U27257 ( .A1(n24987), .A2(n24986), .A3(n24985), .Z(n25007) );
  NAND2HSV0 U27258 ( .A1(\pe11/aot [16]), .A2(\pe11/bq[1] ), .ZN(n24989) );
  NAND2HSV0 U27259 ( .A1(\pe11/bq[5] ), .A2(\pe11/aot [12]), .ZN(n24988) );
  XOR2HSV0 U27260 ( .A1(n24989), .A2(n24988), .Z(n24993) );
  NAND2HSV0 U27261 ( .A1(\pe11/bq[8] ), .A2(\pe11/aot [9]), .ZN(n24991) );
  NAND2HSV0 U27262 ( .A1(\pe11/bq[10] ), .A2(\pe11/aot [7]), .ZN(n24990) );
  XOR2HSV0 U27263 ( .A1(n24991), .A2(n24990), .Z(n24992) );
  XOR2HSV0 U27264 ( .A1(n24993), .A2(n24992), .Z(n25003) );
  NAND2HSV0 U27265 ( .A1(\pe11/bq[2] ), .A2(n24994), .ZN(n24996) );
  NAND2HSV0 U27266 ( .A1(\pe11/bq[13] ), .A2(\pe11/aot [4]), .ZN(n24995) );
  XOR2HSV0 U27267 ( .A1(n24996), .A2(n24995), .Z(n25001) );
  NAND2HSV0 U27268 ( .A1(n24997), .A2(\pe11/aot [2]), .ZN(n24999) );
  NAND2HSV0 U27269 ( .A1(\pe11/bq[4] ), .A2(n12011), .ZN(n24998) );
  XOR2HSV0 U27270 ( .A1(n24999), .A2(n24998), .Z(n25000) );
  XOR2HSV0 U27271 ( .A1(n25001), .A2(n25000), .Z(n25002) );
  XOR2HSV0 U27272 ( .A1(n25003), .A2(n25002), .Z(n25005) );
  NAND2HSV0 U27273 ( .A1(n25489), .A2(\pe11/got [2]), .ZN(n25004) );
  XNOR2HSV1 U27274 ( .A1(n25005), .A2(n25004), .ZN(n25006) );
  XNOR2HSV1 U27275 ( .A1(n25007), .A2(n25006), .ZN(n25010) );
  NAND2HSV0 U27276 ( .A1(n25008), .A2(\pe11/got [4]), .ZN(n25009) );
  XNOR2HSV1 U27277 ( .A1(n25010), .A2(n25009), .ZN(n25012) );
  NAND2HSV0 U27278 ( .A1(n11852), .A2(\pe11/got [6]), .ZN(n25011) );
  XOR3HSV2 U27279 ( .A1(n25013), .A2(n25012), .A3(n25011), .Z(n25014) );
  XNOR2HSV1 U27280 ( .A1(n25015), .A2(n25014), .ZN(n25016) );
  XNOR2HSV1 U27281 ( .A1(n25017), .A2(n25016), .ZN(n25018) );
  XNOR2HSV1 U27282 ( .A1(n25019), .A2(n25018), .ZN(n25021) );
  NAND2HSV0 U27283 ( .A1(n28464), .A2(\pe11/got [10]), .ZN(n25020) );
  XOR2HSV0 U27284 ( .A1(n25021), .A2(n25020), .Z(n25022) );
  XOR2HSV0 U27285 ( .A1(n25023), .A2(n25022), .Z(n25024) );
  XNOR2HSV1 U27286 ( .A1(n25025), .A2(n25024), .ZN(n25056) );
  INAND2HSV4 U27287 ( .A1(n25027), .B1(n25026), .ZN(n25042) );
  NAND3HSV0 U27288 ( .A1(n25030), .A2(\pe11/ti_7t [13]), .A3(n20770), .ZN(
        n25031) );
  CLKAND2HSV1 U27289 ( .A1(n25042), .A2(n25031), .Z(n25038) );
  NOR2HSV0 U27290 ( .A1(n25028), .A2(n25032), .ZN(n25041) );
  CLKNHSV0 U27291 ( .I(n25041), .ZN(n25033) );
  NOR2HSV0 U27292 ( .A1(n25034), .A2(n25033), .ZN(n25035) );
  INHSV1 U27293 ( .I(n25035), .ZN(n25037) );
  CLKNHSV1 U27294 ( .I(n25045), .ZN(n25047) );
  NAND2HSV2 U27295 ( .A1(n25042), .A2(n25047), .ZN(n25036) );
  NOR2HSV2 U27296 ( .A1(n25042), .A2(n20620), .ZN(n25048) );
  CLKNAND2HSV0 U27297 ( .A1(n25040), .A2(n25048), .ZN(n25044) );
  CLKNHSV1 U27298 ( .I(n25040), .ZN(n25046) );
  NAND3HSV2 U27299 ( .A1(n25046), .A2(n25042), .A3(n25041), .ZN(n25043) );
  NAND3HSV2 U27300 ( .A1(n25048), .A2(n25047), .A3(n25046), .ZN(n25049) );
  NOR2HSV0 U27301 ( .A1(n25053), .A2(n25052), .ZN(n25051) );
  NAND2HSV0 U27302 ( .A1(\pe10/aot [2]), .A2(\pe10/bq[1] ), .ZN(n25062) );
  NAND2HSV0 U27303 ( .A1(\pe10/aot [1]), .A2(\pe10/bq[2] ), .ZN(n25061) );
  XOR2HSV0 U27304 ( .A1(n25062), .A2(n25061), .Z(n25063) );
  XOR2HSV0 U27305 ( .A1(n25064), .A2(n25063), .Z(n25065) );
  XOR2HSV0 U27306 ( .A1(n25065), .A2(n25066), .Z(\pe10/poht [14]) );
  NAND2HSV2 U27307 ( .A1(n25414), .A2(\pe11/got [1]), .ZN(n25070) );
  NAND2HSV0 U27308 ( .A1(\pe11/bq[1] ), .A2(\pe11/aot [2]), .ZN(n25068) );
  NAND2HSV0 U27309 ( .A1(\pe11/bq[2] ), .A2(\pe11/aot [1]), .ZN(n25067) );
  XOR2HSV0 U27310 ( .A1(n25068), .A2(n25067), .Z(n25069) );
  XNOR2HSV4 U27311 ( .A1(n25070), .A2(n25069), .ZN(n25072) );
  CLKNAND2HSV1 U27312 ( .A1(n25182), .A2(\pe11/got [2]), .ZN(n25071) );
  XNOR2HSV4 U27313 ( .A1(n25072), .A2(n25071), .ZN(\pe11/poht [14]) );
  NAND2HSV2 U27314 ( .A1(\pe4/bq[1] ), .A2(\pe4/aot [2]), .ZN(n27831) );
  NAND2HSV0 U27315 ( .A1(\pe4/aot [1]), .A2(\pe4/bq[2] ), .ZN(n25073) );
  XOR2HSV0 U27316 ( .A1(n27831), .A2(n25073), .Z(n25078) );
  NAND2HSV2 U27317 ( .A1(n25075), .A2(n25074), .ZN(n28012) );
  NAND2HSV0 U27318 ( .A1(n28012), .A2(\pe4/got [2]), .ZN(n25076) );
  XOR3HSV2 U27319 ( .A1(n25078), .A2(n25077), .A3(n25076), .Z(\pe4/poht [14])
         );
  CLKNHSV1 U27320 ( .I(n25079), .ZN(n25080) );
  NOR2HSV2 U27321 ( .A1(n25080), .A2(n27871), .ZN(n25127) );
  NAND2HSV0 U27322 ( .A1(\pe4/got [10]), .A2(n27907), .ZN(n25125) );
  NOR2HSV0 U27323 ( .A1(n27942), .A2(n27826), .ZN(n25123) );
  NAND2HSV0 U27324 ( .A1(\pe4/got [8]), .A2(n27877), .ZN(n25082) );
  NAND2HSV0 U27325 ( .A1(n27957), .A2(n13996), .ZN(n25081) );
  XNOR2HSV1 U27326 ( .A1(n25082), .A2(n25081), .ZN(n25121) );
  NAND2HSV0 U27327 ( .A1(\pe4/ti_7[7] ), .A2(n22826), .ZN(n25119) );
  NAND2HSV0 U27328 ( .A1(n22825), .A2(\pe4/got [5]), .ZN(n25117) );
  NAND2HSV0 U27329 ( .A1(n27830), .A2(\pe4/got [4]), .ZN(n25115) );
  NAND2HSV0 U27330 ( .A1(\pe4/bq[1] ), .A2(\pe4/aot [14]), .ZN(n25084) );
  NAND2HSV0 U27331 ( .A1(\pe4/aot [7]), .A2(\pe4/bq[8] ), .ZN(n25083) );
  XOR2HSV0 U27332 ( .A1(n25084), .A2(n25083), .Z(n25088) );
  NAND2HSV0 U27333 ( .A1(\pe4/aot [11]), .A2(\pe4/bq[4] ), .ZN(n25086) );
  NAND2HSV0 U27334 ( .A1(\pe4/aot [9]), .A2(\pe4/bq[6] ), .ZN(n25085) );
  XOR2HSV0 U27335 ( .A1(n25086), .A2(n25085), .Z(n25087) );
  XOR2HSV0 U27336 ( .A1(n25088), .A2(n25087), .Z(n25096) );
  NAND2HSV0 U27337 ( .A1(\pe4/aot [2]), .A2(n26961), .ZN(n25090) );
  NAND2HSV0 U27338 ( .A1(\pe4/aot [12]), .A2(\pe4/bq[3] ), .ZN(n25089) );
  XOR2HSV0 U27339 ( .A1(n25090), .A2(n25089), .Z(n25094) );
  NAND2HSV0 U27340 ( .A1(\pe4/aot [10]), .A2(\pe4/bq[5] ), .ZN(n25092) );
  NAND2HSV0 U27341 ( .A1(\pe4/aot [8]), .A2(\pe4/bq[7] ), .ZN(n25091) );
  XOR2HSV0 U27342 ( .A1(n25092), .A2(n25091), .Z(n25093) );
  XOR2HSV0 U27343 ( .A1(n25094), .A2(n25093), .Z(n25095) );
  XOR2HSV0 U27344 ( .A1(n25096), .A2(n25095), .Z(n25107) );
  NAND2HSV0 U27345 ( .A1(\pe4/aot [4]), .A2(\pe4/bq[11] ), .ZN(n25098) );
  NAND2HSV0 U27346 ( .A1(\pe4/aot [3]), .A2(\pe4/bq[12] ), .ZN(n25097) );
  XOR2HSV0 U27347 ( .A1(n25098), .A2(n25097), .Z(n25102) );
  NAND2HSV0 U27348 ( .A1(\pe4/aot [5]), .A2(\pe4/bq[10] ), .ZN(n25100) );
  NAND2HSV0 U27349 ( .A1(\pe4/aot [1]), .A2(n27060), .ZN(n25099) );
  XOR2HSV0 U27350 ( .A1(n25100), .A2(n25099), .Z(n25101) );
  XOR2HSV0 U27351 ( .A1(n25102), .A2(n25101), .Z(n25105) );
  NAND2HSV0 U27352 ( .A1(\pe4/aot [6]), .A2(\pe4/bq[9] ), .ZN(n27796) );
  XOR2HSV0 U27353 ( .A1(n25103), .A2(n27796), .Z(n25104) );
  XNOR2HSV1 U27354 ( .A1(n25105), .A2(n25104), .ZN(n25106) );
  XNOR2HSV1 U27355 ( .A1(n25107), .A2(n25106), .ZN(n25110) );
  NOR2HSV0 U27356 ( .A1(n25108), .A2(n28000), .ZN(n25109) );
  XNOR2HSV1 U27357 ( .A1(n25110), .A2(n25109), .ZN(n25113) );
  NOR2HSV0 U27358 ( .A1(n26981), .A2(n27978), .ZN(n25112) );
  NAND2HSV0 U27359 ( .A1(n27739), .A2(n28626), .ZN(n25111) );
  XOR3HSV1 U27360 ( .A1(n25113), .A2(n25112), .A3(n25111), .Z(n25114) );
  XOR2HSV0 U27361 ( .A1(n25115), .A2(n25114), .Z(n25116) );
  XNOR2HSV1 U27362 ( .A1(n25117), .A2(n25116), .ZN(n25118) );
  XNOR2HSV1 U27363 ( .A1(n25119), .A2(n25118), .ZN(n25120) );
  XNOR2HSV1 U27364 ( .A1(n25121), .A2(n25120), .ZN(n25122) );
  XOR2HSV0 U27365 ( .A1(n25123), .A2(n25122), .Z(n25124) );
  XNOR2HSV1 U27366 ( .A1(n25125), .A2(n25124), .ZN(n25126) );
  CLKNAND2HSV1 U27367 ( .A1(n27940), .A2(n25128), .ZN(n25129) );
  XNOR2HSV4 U27368 ( .A1(n25130), .A2(n25129), .ZN(n25133) );
  NAND2HSV0 U27369 ( .A1(n27904), .A2(n25131), .ZN(n25132) );
  XNOR2HSV1 U27370 ( .A1(n25136), .A2(n25135), .ZN(\pe4/poht [2]) );
  NAND2HSV2 U27371 ( .A1(n28936), .A2(\pe11/got [10]), .ZN(n25181) );
  NAND2HSV0 U27372 ( .A1(n28918), .A2(\pe11/got [7]), .ZN(n25175) );
  NAND2HSV0 U27373 ( .A1(n14064), .A2(\pe11/got [6]), .ZN(n25173) );
  NAND2HSV0 U27374 ( .A1(n25138), .A2(\pe11/got [4]), .ZN(n25168) );
  NAND2HSV0 U27375 ( .A1(n25139), .A2(\pe11/got [3]), .ZN(n25166) );
  NAND2HSV0 U27376 ( .A1(n28471), .A2(\pe11/got [2]), .ZN(n25164) );
  NAND2HSV0 U27377 ( .A1(n25140), .A2(\pe11/got [1]), .ZN(n25162) );
  NAND2HSV0 U27378 ( .A1(\pe11/bq[5] ), .A2(\pe11/aot [7]), .ZN(n25142) );
  NAND2HSV0 U27379 ( .A1(\pe11/bq[8] ), .A2(\pe11/aot [4]), .ZN(n25141) );
  XOR2HSV0 U27380 ( .A1(n25142), .A2(n25141), .Z(n25146) );
  NAND2HSV0 U27381 ( .A1(\pe11/bq[11] ), .A2(\pe11/aot [1]), .ZN(n25144) );
  NAND2HSV0 U27382 ( .A1(\pe11/bq[7] ), .A2(\pe11/aot [5]), .ZN(n25143) );
  XOR2HSV0 U27383 ( .A1(n25144), .A2(n25143), .Z(n25145) );
  XOR2HSV0 U27384 ( .A1(n25146), .A2(n25145), .Z(n25152) );
  NAND2HSV0 U27385 ( .A1(\pe11/bq[1] ), .A2(\pe11/aot [11]), .ZN(n25148) );
  NAND2HSV0 U27386 ( .A1(\pe11/bq[2] ), .A2(\pe11/aot [10]), .ZN(n25147) );
  XOR2HSV0 U27387 ( .A1(n25148), .A2(n25147), .Z(n25150) );
  NAND2HSV0 U27388 ( .A1(\pe11/bq[3] ), .A2(\pe11/aot [9]), .ZN(n25149) );
  XNOR2HSV1 U27389 ( .A1(n25150), .A2(n25149), .ZN(n25151) );
  XNOR2HSV1 U27390 ( .A1(n25152), .A2(n25151), .ZN(n25160) );
  NAND2HSV0 U27391 ( .A1(\pe11/bq[6] ), .A2(\pe11/aot [6]), .ZN(n25154) );
  NAND2HSV0 U27392 ( .A1(\pe11/bq[10] ), .A2(\pe11/aot [2]), .ZN(n25153) );
  XOR2HSV0 U27393 ( .A1(n25154), .A2(n25153), .Z(n25158) );
  NAND2HSV0 U27394 ( .A1(\pe11/bq[9] ), .A2(\pe11/aot [3]), .ZN(n25156) );
  NAND2HSV0 U27395 ( .A1(\pe11/bq[4] ), .A2(\pe11/aot [8]), .ZN(n25155) );
  XOR2HSV0 U27396 ( .A1(n25156), .A2(n25155), .Z(n25157) );
  XOR2HSV0 U27397 ( .A1(n25158), .A2(n25157), .Z(n25159) );
  XNOR2HSV1 U27398 ( .A1(n25160), .A2(n25159), .ZN(n25161) );
  XOR2HSV0 U27399 ( .A1(n25162), .A2(n25161), .Z(n25163) );
  XOR2HSV0 U27400 ( .A1(n25164), .A2(n25163), .Z(n25165) );
  XOR2HSV0 U27401 ( .A1(n25166), .A2(n25165), .Z(n25167) );
  XOR2HSV0 U27402 ( .A1(n25168), .A2(n25167), .Z(n25171) );
  NAND2HSV0 U27403 ( .A1(n25169), .A2(\pe11/got [5]), .ZN(n25170) );
  XOR2HSV0 U27404 ( .A1(n25171), .A2(n25170), .Z(n25172) );
  XOR2HSV0 U27405 ( .A1(n25173), .A2(n25172), .Z(n25174) );
  XNOR2HSV1 U27406 ( .A1(n25175), .A2(n25174), .ZN(n25177) );
  XNOR2HSV4 U27407 ( .A1(n25181), .A2(n25180), .ZN(n25184) );
  CLKNAND2HSV1 U27408 ( .A1(n25182), .A2(\pe11/got [11]), .ZN(n25183) );
  XNOR2HSV4 U27409 ( .A1(n25184), .A2(n25183), .ZN(\pe11/poht [5]) );
  NAND2HSV0 U27410 ( .A1(n26231), .A2(n14060), .ZN(n25211) );
  CLKNAND2HSV1 U27411 ( .A1(n25185), .A2(\pe8/got [5]), .ZN(n25206) );
  NAND2HSV0 U27412 ( .A1(\pe8/aot [5]), .A2(\pe8/bq[4] ), .ZN(n25188) );
  NAND2HSV0 U27413 ( .A1(\pe8/aot [6]), .A2(\pe8/bq[3] ), .ZN(n25187) );
  XOR2HSV0 U27414 ( .A1(n25188), .A2(n25187), .Z(n25192) );
  NAND2HSV0 U27415 ( .A1(\pe8/aot [1]), .A2(\pe8/bq[8] ), .ZN(n25189) );
  XOR2HSV0 U27416 ( .A1(n25190), .A2(n25189), .Z(n25191) );
  XOR2HSV0 U27417 ( .A1(n25192), .A2(n25191), .Z(n25202) );
  NAND2HSV0 U27418 ( .A1(\pe8/aot [2]), .A2(\pe8/bq[7] ), .ZN(n25194) );
  NAND2HSV0 U27419 ( .A1(\pe8/aot [3]), .A2(\pe8/bq[6] ), .ZN(n25193) );
  XOR2HSV0 U27420 ( .A1(n25194), .A2(n25193), .Z(n25200) );
  NOR2HSV0 U27421 ( .A1(n25196), .A2(n25195), .ZN(n25198) );
  AOI22HSV0 U27422 ( .A1(\pe8/aot [7]), .A2(\pe8/bq[2] ), .B1(\pe8/aot [8]), 
        .B2(\pe8/bq[1] ), .ZN(n25197) );
  NOR2HSV2 U27423 ( .A1(n25198), .A2(n25197), .ZN(n25199) );
  XNOR2HSV1 U27424 ( .A1(n25200), .A2(n25199), .ZN(n25201) );
  XNOR2HSV1 U27425 ( .A1(n25206), .A2(n25205), .ZN(n25209) );
  INHSV1 U27426 ( .I(n25207), .ZN(n25208) );
  XOR2HSV0 U27427 ( .A1(n25209), .A2(n25208), .Z(n25210) );
  XOR2HSV0 U27428 ( .A1(n25211), .A2(n25210), .Z(n25212) );
  XOR2HSV0 U27429 ( .A1(n25212), .A2(n25213), .Z(\pe8/poht [8]) );
  NOR2HSV2 U27430 ( .A1(n12304), .A2(n25214), .ZN(n25252) );
  NOR2HSV2 U27431 ( .A1(n25215), .A2(n26158), .ZN(n25248) );
  NAND2HSV0 U27432 ( .A1(n25216), .A2(n26132), .ZN(n25241) );
  NAND2HSV0 U27433 ( .A1(n26094), .A2(\pe10/got [3]), .ZN(n25239) );
  NOR2HSV0 U27434 ( .A1(n26096), .A2(n27194), .ZN(n25237) );
  NAND2HSV0 U27435 ( .A1(n26131), .A2(n27196), .ZN(n25235) );
  NAND2HSV0 U27436 ( .A1(\pe10/aot [1]), .A2(\pe10/bq[11] ), .ZN(n25219) );
  NAND2HSV2 U27437 ( .A1(\pe10/aot [1]), .A2(\pe10/bq[1] ), .ZN(n25694) );
  NOR2HSV0 U27438 ( .A1(n25217), .A2(n25694), .ZN(n25218) );
  AOI21HSV2 U27439 ( .A1(n25220), .A2(n25219), .B(n25218), .ZN(n25222) );
  XNOR2HSV1 U27440 ( .A1(n25222), .A2(n25221), .ZN(n25233) );
  NAND2HSV0 U27441 ( .A1(\pe10/aot [4]), .A2(\pe10/bq[8] ), .ZN(n25226) );
  NAND2HSV0 U27442 ( .A1(\pe10/aot [5]), .A2(\pe10/bq[7] ), .ZN(n25225) );
  XOR2HSV0 U27443 ( .A1(n25226), .A2(n25225), .Z(n25230) );
  NAND2HSV0 U27444 ( .A1(\pe10/aot [8]), .A2(\pe10/bq[4] ), .ZN(n25228) );
  NAND2HSV0 U27445 ( .A1(\pe10/aot [7]), .A2(\pe10/bq[5] ), .ZN(n25227) );
  XOR2HSV0 U27446 ( .A1(n25228), .A2(n25227), .Z(n25229) );
  XOR2HSV0 U27447 ( .A1(n25230), .A2(n25229), .Z(n25231) );
  XOR3HSV2 U27448 ( .A1(n25233), .A2(n25232), .A3(n25231), .Z(n25234) );
  XNOR2HSV1 U27449 ( .A1(n25235), .A2(n25234), .ZN(n25236) );
  XNOR2HSV1 U27450 ( .A1(n25237), .A2(n25236), .ZN(n25238) );
  XNOR2HSV1 U27451 ( .A1(n25239), .A2(n25238), .ZN(n25240) );
  XNOR2HSV1 U27452 ( .A1(n25241), .A2(n25240), .ZN(n25243) );
  NAND2HSV0 U27453 ( .A1(n28585), .A2(\pe10/got [5]), .ZN(n25242) );
  XOR2HSV0 U27454 ( .A1(n25243), .A2(n25242), .Z(n25246) );
  NAND2HSV0 U27455 ( .A1(n25244), .A2(\pe10/got [6]), .ZN(n25245) );
  XNOR2HSV1 U27456 ( .A1(n25246), .A2(n25245), .ZN(n25247) );
  XOR2HSV0 U27457 ( .A1(n25248), .A2(n25247), .Z(n25250) );
  NAND2HSV0 U27458 ( .A1(n27197), .A2(n28642), .ZN(n25249) );
  XOR2HSV0 U27459 ( .A1(n25250), .A2(n25249), .Z(n25251) );
  CLKXOR2HSV4 U27460 ( .A1(n25252), .A2(n25251), .Z(n25254) );
  NAND2HSV2 U27461 ( .A1(n28644), .A2(n25060), .ZN(n25253) );
  NOR2HSV2 U27462 ( .A1(n25260), .A2(n25256), .ZN(n25264) );
  NOR2HSV2 U27463 ( .A1(n28603), .A2(n25259), .ZN(n25268) );
  OAI21HSV0 U27464 ( .A1(n16998), .A2(\pe10/ti_7t [15]), .B(\pe10/got [11]), 
        .ZN(n25267) );
  NOR2HSV0 U27465 ( .A1(n12304), .A2(n25267), .ZN(n25265) );
  OAI21HSV0 U27466 ( .A1(n27195), .A2(n25261), .B(n25260), .ZN(n25262) );
  NOR2HSV1 U27467 ( .A1(n25262), .A2(n25267), .ZN(n25263) );
  AOI21HSV2 U27468 ( .A1(n25265), .A2(n25264), .B(n25263), .ZN(n25266) );
  OAI21HSV2 U27469 ( .A1(n25268), .A2(n25267), .B(n25266), .ZN(n25269) );
  NAND2HSV2 U27470 ( .A1(n28659), .A2(\pe7/got [16]), .ZN(n25343) );
  CLKNAND2HSV0 U27471 ( .A1(n25376), .A2(\pe7/got [12]), .ZN(n25333) );
  NAND2HSV0 U27472 ( .A1(n28656), .A2(n14022), .ZN(n25331) );
  NAND2HSV0 U27473 ( .A1(n14067), .A2(\pe7/got [8]), .ZN(n25324) );
  NAND2HSV0 U27474 ( .A1(n25271), .A2(n11935), .ZN(n25322) );
  NAND2HSV0 U27475 ( .A1(n28621), .A2(n25272), .ZN(n25317) );
  NAND2HSV0 U27476 ( .A1(\pe7/aot [9]), .A2(\pe7/bq[8] ), .ZN(n25275) );
  NAND2HSV0 U27477 ( .A1(\pe7/aot [1]), .A2(n25273), .ZN(n25274) );
  XOR2HSV0 U27478 ( .A1(n25275), .A2(n25274), .Z(n25291) );
  CLKNHSV0 U27479 ( .I(n25278), .ZN(n27103) );
  XOR2HSV0 U27480 ( .A1(n25282), .A2(n25281), .Z(n25290) );
  NAND2HSV0 U27481 ( .A1(\pe7/aot [8]), .A2(\pe7/bq[9] ), .ZN(n25284) );
  NAND2HSV0 U27482 ( .A1(\pe7/aot [5]), .A2(\pe7/bq[12] ), .ZN(n25283) );
  XOR2HSV0 U27483 ( .A1(n25284), .A2(n25283), .Z(n25288) );
  NAND2HSV0 U27484 ( .A1(\pe7/aot [6]), .A2(\pe7/bq[11] ), .ZN(n25286) );
  NAND2HSV0 U27485 ( .A1(\pe7/aot [7]), .A2(\pe7/bq[10] ), .ZN(n25285) );
  XOR2HSV0 U27486 ( .A1(n25286), .A2(n25285), .Z(n25287) );
  XOR2HSV0 U27487 ( .A1(n25288), .A2(n25287), .Z(n25289) );
  XOR3HSV2 U27488 ( .A1(n25291), .A2(n25290), .A3(n25289), .Z(n25314) );
  NAND2HSV0 U27489 ( .A1(n25292), .A2(\pe7/got [3]), .ZN(n25313) );
  NAND2HSV0 U27490 ( .A1(n14050), .A2(\pe7/bq[4] ), .ZN(n25294) );
  NAND2HSV0 U27491 ( .A1(\pe7/aot [10]), .A2(\pe7/bq[7] ), .ZN(n25293) );
  XOR2HSV0 U27492 ( .A1(n25294), .A2(n25293), .Z(n25298) );
  NAND2HSV0 U27493 ( .A1(\pe7/aot [4]), .A2(\pe7/bq[13] ), .ZN(n25296) );
  NAND2HSV0 U27494 ( .A1(\pe7/aot [12]), .A2(\pe7/bq[5] ), .ZN(n25295) );
  XOR2HSV0 U27495 ( .A1(n25296), .A2(n25295), .Z(n25297) );
  XOR2HSV0 U27496 ( .A1(n25298), .A2(n25297), .Z(n25307) );
  NAND2HSV0 U27497 ( .A1(n28876), .A2(\pe7/pq ), .ZN(n25301) );
  NAND2HSV0 U27498 ( .A1(\pe7/got [1]), .A2(n25299), .ZN(n25300) );
  XOR2HSV0 U27499 ( .A1(n25301), .A2(n25300), .Z(n25305) );
  XNOR2HSV1 U27500 ( .A1(n25305), .A2(n25304), .ZN(n25306) );
  XNOR2HSV1 U27501 ( .A1(n25307), .A2(n25306), .ZN(n25311) );
  NOR2HSV0 U27502 ( .A1(n25309), .A2(n25308), .ZN(n25310) );
  XNOR2HSV1 U27503 ( .A1(n25311), .A2(n25310), .ZN(n25312) );
  XOR3HSV2 U27504 ( .A1(n25314), .A2(n25313), .A3(n25312), .Z(n25316) );
  NAND2HSV0 U27505 ( .A1(n11936), .A2(n25375), .ZN(n25315) );
  XOR3HSV2 U27506 ( .A1(n25317), .A2(n25316), .A3(n25315), .Z(n25320) );
  NAND2HSV0 U27507 ( .A1(\pe7/got [6]), .A2(n25318), .ZN(n25319) );
  XOR2HSV0 U27508 ( .A1(n25320), .A2(n25319), .Z(n25321) );
  XOR2HSV0 U27509 ( .A1(n25322), .A2(n25321), .Z(n25323) );
  XOR2HSV0 U27510 ( .A1(n25324), .A2(n25323), .Z(n25327) );
  NAND2HSV0 U27511 ( .A1(n11978), .A2(\pe7/got [9]), .ZN(n25326) );
  XOR2HSV0 U27512 ( .A1(n25327), .A2(n25326), .Z(n25329) );
  NAND2HSV0 U27513 ( .A1(n25397), .A2(n24214), .ZN(n25328) );
  XNOR2HSV1 U27514 ( .A1(n25329), .A2(n25328), .ZN(n25330) );
  XNOR2HSV1 U27515 ( .A1(n25331), .A2(n25330), .ZN(n25332) );
  XOR2HSV0 U27516 ( .A1(n25333), .A2(n25332), .Z(n25337) );
  CLKNAND2HSV0 U27517 ( .A1(n25335), .A2(n25334), .ZN(n25336) );
  XOR2HSV0 U27518 ( .A1(n25337), .A2(n25336), .Z(n25342) );
  DELHS4 U27519 ( .I(n25347), .Z(n25348) );
  MUX2HSV2 U27520 ( .I0(bo1[6]), .I1(\pe1/bq[6] ), .S(n27065), .Z(n28744) );
  MUX2HSV2 U27521 ( .I0(n25349), .I1(bo5[16]), .S(n27048), .Z(n28709) );
  INHSV2 U27522 ( .I(n25350), .ZN(n28955) );
  INHSV2 U27523 ( .I(n25351), .ZN(n28947) );
  CLKNAND2HSV0 U27524 ( .A1(n26297), .A2(n26240), .ZN(n25354) );
  XOR2HSV0 U27525 ( .A1(n25354), .A2(n25353), .Z(n25356) );
  NAND2HSV0 U27526 ( .A1(n26752), .A2(n26413), .ZN(n25355) );
  XOR2HSV0 U27527 ( .A1(n25356), .A2(n25355), .Z(pov3[11]) );
  CLKNAND2HSV0 U27528 ( .A1(n27657), .A2(n28693), .ZN(n25359) );
  CLKNHSV0 U27529 ( .I(n25357), .ZN(n25358) );
  XNOR2HSV1 U27530 ( .A1(n25359), .A2(n25358), .ZN(n28972) );
  CLKNAND2HSV0 U27531 ( .A1(n27667), .A2(n28421), .ZN(n25360) );
  XNOR2HSV1 U27532 ( .A1(n25360), .A2(n25361), .ZN(n25368) );
  NAND2HSV2 U27533 ( .A1(n25362), .A2(n28693), .ZN(n25363) );
  NAND2HSV0 U27534 ( .A1(n25364), .A2(n25363), .ZN(n25365) );
  NOR2HSV1 U27535 ( .A1(n25366), .A2(n25365), .ZN(n25367) );
  XNOR2HSV1 U27536 ( .A1(n25368), .A2(n25367), .ZN(n28986) );
  NAND2HSV2 U27537 ( .A1(n28659), .A2(\pe7/got [9]), .ZN(n25412) );
  NOR2HSV2 U27538 ( .A1(n25374), .A2(n25373), .ZN(n25407) );
  CLKNAND2HSV1 U27539 ( .A1(n25376), .A2(n25375), .ZN(n25403) );
  NAND2HSV0 U27540 ( .A1(n25377), .A2(\pe7/got [4]), .ZN(n25401) );
  NAND2HSV0 U27541 ( .A1(n14067), .A2(\pe7/got [1]), .ZN(n25394) );
  NAND2HSV0 U27542 ( .A1(\pe7/aot [4]), .A2(\pe7/bq[6] ), .ZN(n25379) );
  NAND2HSV0 U27543 ( .A1(\pe7/aot [9]), .A2(\pe7/bq[1] ), .ZN(n25378) );
  XOR2HSV0 U27544 ( .A1(n25379), .A2(n25378), .Z(n25392) );
  NAND2HSV0 U27545 ( .A1(\pe7/aot [8]), .A2(\pe7/bq[2] ), .ZN(n25381) );
  NAND2HSV0 U27546 ( .A1(\pe7/aot [6]), .A2(\pe7/bq[4] ), .ZN(n25380) );
  XOR2HSV0 U27547 ( .A1(n25381), .A2(n25380), .Z(n25383) );
  XNOR2HSV1 U27548 ( .A1(n25383), .A2(n25382), .ZN(n25391) );
  NAND2HSV0 U27549 ( .A1(\pe7/aot [7]), .A2(\pe7/bq[3] ), .ZN(n25385) );
  NAND2HSV0 U27550 ( .A1(\pe7/aot [3]), .A2(\pe7/bq[7] ), .ZN(n25384) );
  XOR2HSV0 U27551 ( .A1(n25385), .A2(n25384), .Z(n25389) );
  NAND2HSV0 U27552 ( .A1(\pe7/aot [2]), .A2(\pe7/bq[8] ), .ZN(n25387) );
  NAND2HSV0 U27553 ( .A1(\pe7/aot [1]), .A2(\pe7/bq[9] ), .ZN(n25386) );
  XOR2HSV0 U27554 ( .A1(n25387), .A2(n25386), .Z(n25388) );
  XOR2HSV0 U27555 ( .A1(n25389), .A2(n25388), .Z(n25390) );
  XOR3HSV2 U27556 ( .A1(n25392), .A2(n25391), .A3(n25390), .Z(n25393) );
  XNOR2HSV1 U27557 ( .A1(n25394), .A2(n25393), .ZN(n25396) );
  NAND2HSV0 U27558 ( .A1(n28587), .A2(\pe7/got [2]), .ZN(n25395) );
  XOR2HSV0 U27559 ( .A1(n25396), .A2(n25395), .Z(n25399) );
  NAND2HSV0 U27560 ( .A1(n25397), .A2(\pe7/got [3]), .ZN(n25398) );
  XNOR2HSV1 U27561 ( .A1(n25399), .A2(n25398), .ZN(n25400) );
  XOR2HSV0 U27562 ( .A1(n25401), .A2(n25400), .Z(n25402) );
  XOR2HSV0 U27563 ( .A1(n25403), .A2(n25402), .Z(n25405) );
  NAND2HSV0 U27564 ( .A1(n14030), .A2(\pe7/got [6]), .ZN(n25404) );
  XNOR2HSV1 U27565 ( .A1(n25405), .A2(n25404), .ZN(n25406) );
  XNOR2HSV4 U27566 ( .A1(n25407), .A2(n25406), .ZN(n25410) );
  NAND2HSV0 U27567 ( .A1(n25408), .A2(\pe7/got [8]), .ZN(n25409) );
  XNOR2HSV4 U27568 ( .A1(n25410), .A2(n25409), .ZN(n25411) );
  NAND2HSV2 U27569 ( .A1(n25414), .A2(n20182), .ZN(n25416) );
  NOR2HSV4 U27570 ( .A1(n25417), .A2(n24889), .ZN(n25418) );
  CLKXOR2HSV4 U27571 ( .A1(n25418), .A2(poh11[15]), .Z(po[16]) );
  NAND2HSV0 U27572 ( .A1(n25950), .A2(n25420), .ZN(n25486) );
  CLKNAND2HSV1 U27573 ( .A1(n28699), .A2(n28686), .ZN(n25480) );
  NAND2HSV0 U27574 ( .A1(n26031), .A2(n14236), .ZN(n25478) );
  CLKNAND2HSV0 U27575 ( .A1(n25952), .A2(n28586), .ZN(n25474) );
  NAND2HSV0 U27576 ( .A1(\pe6/ti_7[7] ), .A2(\pe6/got [8]), .ZN(n25468) );
  NAND2HSV0 U27577 ( .A1(n28526), .A2(\pe6/got [7]), .ZN(n25466) );
  INAND2HSV0 U27578 ( .A1(n14029), .B1(n25982), .ZN(n25464) );
  NAND2HSV0 U27579 ( .A1(n25849), .A2(\pe6/got [4]), .ZN(n25462) );
  NAND2HSV0 U27580 ( .A1(n25846), .A2(n14008), .ZN(n25440) );
  NAND2HSV0 U27581 ( .A1(n19021), .A2(n28608), .ZN(n25422) );
  NAND2HSV0 U27582 ( .A1(\pe6/aot [4]), .A2(\pe6/bq[13] ), .ZN(n25421) );
  XOR2HSV0 U27583 ( .A1(n25422), .A2(n25421), .Z(n25438) );
  NAND2HSV0 U27584 ( .A1(\pe6/aot [12]), .A2(\pe6/bq[1] ), .ZN(n26054) );
  NOR2HSV0 U27585 ( .A1(n25423), .A2(n26054), .ZN(n25425) );
  AOI22HSV0 U27586 ( .A1(n28681), .A2(\pe6/bq[1] ), .B1(\pe6/aot [12]), .B2(
        \pe6/bq[5] ), .ZN(n25424) );
  NOR2HSV2 U27587 ( .A1(n25425), .A2(n25424), .ZN(n25429) );
  XOR2HSV0 U27588 ( .A1(n25429), .A2(n25428), .Z(n25437) );
  NAND2HSV0 U27589 ( .A1(\pe6/aot [1]), .A2(n14028), .ZN(n25431) );
  NAND2HSV0 U27590 ( .A1(\pe6/aot [8]), .A2(\pe6/bq[9] ), .ZN(n25430) );
  XOR2HSV0 U27591 ( .A1(n25431), .A2(n25430), .Z(n25435) );
  NAND2HSV0 U27592 ( .A1(\pe6/aot [6]), .A2(\pe6/bq[11] ), .ZN(n25433) );
  NAND2HSV0 U27593 ( .A1(\pe6/aot [9]), .A2(\pe6/bq[8] ), .ZN(n25432) );
  XOR2HSV0 U27594 ( .A1(n25433), .A2(n25432), .Z(n25434) );
  XNOR2HSV1 U27595 ( .A1(n25435), .A2(n25434), .ZN(n25436) );
  XOR3HSV2 U27596 ( .A1(n25438), .A2(n25437), .A3(n25436), .Z(n25439) );
  XNOR2HSV1 U27597 ( .A1(n25440), .A2(n25439), .ZN(n25459) );
  NAND2HSV0 U27598 ( .A1(n28867), .A2(\pe6/pq ), .ZN(n25442) );
  NAND2HSV0 U27599 ( .A1(\pe6/aot [11]), .A2(\pe6/bq[6] ), .ZN(n25441) );
  XOR2HSV0 U27600 ( .A1(n25442), .A2(n25441), .Z(n25446) );
  NAND2HSV0 U27601 ( .A1(\pe6/aot [5]), .A2(\pe6/bq[12] ), .ZN(n25444) );
  NAND2HSV0 U27602 ( .A1(\pe6/bq[7] ), .A2(\pe6/aot [10]), .ZN(n25443) );
  XOR2HSV0 U27603 ( .A1(n25444), .A2(n25443), .Z(n25445) );
  XOR2HSV0 U27604 ( .A1(n25446), .A2(n25445), .Z(n25454) );
  NAND2HSV0 U27605 ( .A1(\pe6/bq[15] ), .A2(\pe6/aot [2]), .ZN(n25448) );
  NAND2HSV0 U27606 ( .A1(\pe6/aot [7]), .A2(\pe6/bq[10] ), .ZN(n25447) );
  XOR2HSV0 U27607 ( .A1(n25448), .A2(n25447), .Z(n25452) );
  NAND2HSV0 U27608 ( .A1(n28680), .A2(\pe6/bq[2] ), .ZN(n25450) );
  NAND2HSV0 U27609 ( .A1(\pe6/aot [3]), .A2(\pe6/bq[14] ), .ZN(n25449) );
  XOR2HSV0 U27610 ( .A1(n25450), .A2(n25449), .Z(n25451) );
  XOR2HSV0 U27611 ( .A1(n25452), .A2(n25451), .Z(n25453) );
  XOR2HSV0 U27612 ( .A1(n25454), .A2(n25453), .Z(n25457) );
  NOR2HSV0 U27613 ( .A1(n25455), .A2(n28651), .ZN(n25456) );
  XNOR2HSV1 U27614 ( .A1(n25457), .A2(n25456), .ZN(n25458) );
  XNOR2HSV1 U27615 ( .A1(n25459), .A2(n25458), .ZN(n25461) );
  NAND2HSV0 U27616 ( .A1(n28792), .A2(n26065), .ZN(n25460) );
  XOR3HSV2 U27617 ( .A1(n25462), .A2(n25461), .A3(n25460), .Z(n25463) );
  XOR2HSV0 U27618 ( .A1(n25464), .A2(n25463), .Z(n25465) );
  XNOR2HSV1 U27619 ( .A1(n25466), .A2(n25465), .ZN(n25467) );
  XNOR2HSV1 U27620 ( .A1(n25468), .A2(n25467), .ZN(n25470) );
  NAND2HSV0 U27621 ( .A1(n25764), .A2(\pe6/got [9]), .ZN(n25469) );
  XOR2HSV0 U27622 ( .A1(n25470), .A2(n25469), .Z(n25472) );
  NAND2HSV0 U27623 ( .A1(n26068), .A2(\pe6/got [10]), .ZN(n25471) );
  XNOR2HSV1 U27624 ( .A1(n25472), .A2(n25471), .ZN(n25473) );
  XNOR2HSV1 U27625 ( .A1(n25474), .A2(n25473), .ZN(n25475) );
  XOR2HSV0 U27626 ( .A1(n25476), .A2(n25475), .Z(n25477) );
  XOR2HSV2 U27627 ( .A1(n25478), .A2(n25477), .Z(n25481) );
  INHSV1 U27628 ( .I(n25481), .ZN(n25479) );
  CLKNAND2HSV1 U27629 ( .A1(n25480), .A2(n25479), .ZN(n25484) );
  CLKNHSV0 U27630 ( .I(n25480), .ZN(n25482) );
  CLKNAND2HSV1 U27631 ( .A1(n25482), .A2(n25481), .ZN(n25483) );
  CLKNAND2HSV1 U27632 ( .A1(n25484), .A2(n25483), .ZN(n25485) );
  NAND2HSV0 U27633 ( .A1(n25489), .A2(n25488), .ZN(n25491) );
  XNOR2HSV0 U27634 ( .A1(n25491), .A2(n25490), .ZN(n25492) );
  NOR2HSV1 U27635 ( .A1(n25492), .A2(n25515), .ZN(n25493) );
  XOR2HSV0 U27636 ( .A1(n25493), .A2(poh11[2]), .Z(po[3]) );
  NAND3HSV0 U27637 ( .A1(n23116), .A2(n25495), .A3(n25494), .ZN(n25497) );
  OAI211HSV1 U27638 ( .A1(n25499), .A2(n25498), .B(n25497), .C(n25496), .ZN(
        n25501) );
  XNOR2HSV1 U27639 ( .A1(n25501), .A2(n25500), .ZN(n29013) );
  NOR2HSV0 U27640 ( .A1(n12010), .A2(n25512), .ZN(n25503) );
  XOR2HSV0 U27641 ( .A1(n25503), .A2(poh11[1]), .Z(po[2]) );
  NAND2HSV0 U27642 ( .A1(n28629), .A2(n25504), .ZN(n25507) );
  CLKNHSV0 U27643 ( .I(n25505), .ZN(n25506) );
  XNOR2HSV1 U27644 ( .A1(n25507), .A2(n25506), .ZN(n25509) );
  XNOR2HSV1 U27645 ( .A1(n25509), .A2(n25508), .ZN(n25510) );
  NOR2HSV1 U27646 ( .A1(n25510), .A2(n20463), .ZN(n25511) );
  XOR2HSV0 U27647 ( .A1(n25511), .A2(poh11[3]), .Z(po[4]) );
  NOR2HSV0 U27648 ( .A1(n25513), .A2(n25512), .ZN(n25514) );
  XOR2HSV0 U27649 ( .A1(n25514), .A2(poh11[4]), .Z(po[5]) );
  INHSV2 U27650 ( .I(n27904), .ZN(n27875) );
  CLKNHSV0 U27651 ( .I(n27999), .ZN(n28941) );
  AND2HSV2 U27652 ( .A1(n25524), .A2(n25523), .Z(n25610) );
  NAND2HSV2 U27653 ( .A1(n25525), .A2(n28695), .ZN(n25614) );
  INHSV2 U27654 ( .I(n25614), .ZN(n25526) );
  OAI21HSV2 U27655 ( .A1(n20063), .A2(n25610), .B(n25526), .ZN(n25618) );
  CLKNAND2HSV0 U27656 ( .A1(n28698), .A2(n22136), .ZN(n25601) );
  NAND2HSV0 U27657 ( .A1(n28631), .A2(\pe8/got [10]), .ZN(n25594) );
  NAND2HSV0 U27658 ( .A1(n28616), .A2(\pe8/got [9]), .ZN(n25592) );
  NOR2HSV0 U27659 ( .A1(n25528), .A2(n25527), .ZN(n25590) );
  NAND2HSV0 U27660 ( .A1(n12007), .A2(\pe8/got [6]), .ZN(n25586) );
  NAND2HSV0 U27661 ( .A1(\pe8/aot [11]), .A2(\pe8/bq[6] ), .ZN(n25534) );
  NAND2HSV0 U27662 ( .A1(\pe8/aot [2]), .A2(n25532), .ZN(n25533) );
  XOR2HSV0 U27663 ( .A1(n25534), .A2(n25533), .Z(n25535) );
  XOR2HSV0 U27664 ( .A1(n25536), .A2(n25535), .Z(n25549) );
  NAND2HSV0 U27665 ( .A1(n23547), .A2(\pe8/pq ), .ZN(n25538) );
  NAND2HSV0 U27666 ( .A1(\pe8/aot [9]), .A2(\pe8/bq[8] ), .ZN(n25537) );
  XOR2HSV0 U27667 ( .A1(n25538), .A2(n25537), .Z(n25547) );
  NAND2HSV2 U27668 ( .A1(\pe8/bq[1] ), .A2(\pe8/aot [1]), .ZN(n26222) );
  CLKNHSV0 U27669 ( .I(n25539), .ZN(n25542) );
  CLKNHSV0 U27670 ( .I(n28627), .ZN(n25540) );
  OR2HSV0 U27671 ( .A1(n25542), .A2(n25540), .Z(n25545) );
  NAND2HSV0 U27672 ( .A1(n28627), .A2(\pe8/bq[1] ), .ZN(n25541) );
  OAI21HSV0 U27673 ( .A1(n25543), .A2(n25542), .B(n25541), .ZN(n25544) );
  OAI21HSV0 U27674 ( .A1(n26222), .A2(n25545), .B(n25544), .ZN(n25546) );
  XNOR2HSV1 U27675 ( .A1(n25547), .A2(n25546), .ZN(n25548) );
  XNOR2HSV1 U27676 ( .A1(n25549), .A2(n25548), .ZN(n25551) );
  NOR2HSV0 U27677 ( .A1(n27225), .A2(n28650), .ZN(n25550) );
  XNOR2HSV1 U27678 ( .A1(n25551), .A2(n25550), .ZN(n25581) );
  NAND2HSV0 U27679 ( .A1(n28788), .A2(\pe8/got [3]), .ZN(n25576) );
  NAND2HSV0 U27680 ( .A1(\pe8/aot [8]), .A2(\pe8/bq[9] ), .ZN(n25552) );
  XOR2HSV0 U27681 ( .A1(n25553), .A2(n25552), .Z(n25574) );
  OAI21HSV0 U27682 ( .A1(n19995), .A2(n25555), .B(n25554), .ZN(n25556) );
  OAI21HSV0 U27683 ( .A1(n25558), .A2(n25557), .B(n25556), .ZN(n25564) );
  NOR2HSV0 U27684 ( .A1(n25560), .A2(n25559), .ZN(n25562) );
  AOI22HSV0 U27685 ( .A1(\pe8/aot [12]), .A2(\pe8/bq[5] ), .B1(\pe8/aot [10]), 
        .B2(\pe8/bq[7] ), .ZN(n25561) );
  NOR2HSV1 U27686 ( .A1(n25562), .A2(n25561), .ZN(n25563) );
  XOR2HSV0 U27687 ( .A1(n25564), .A2(n25563), .Z(n25573) );
  NAND2HSV0 U27688 ( .A1(\pe8/aot [4]), .A2(n25565), .ZN(n25567) );
  NAND2HSV0 U27689 ( .A1(\pe8/aot [5]), .A2(\pe8/bq[12] ), .ZN(n25566) );
  XOR2HSV0 U27690 ( .A1(n25567), .A2(n25566), .Z(n25571) );
  NAND2HSV0 U27691 ( .A1(\pe8/aot [6]), .A2(\pe8/bq[11] ), .ZN(n25569) );
  NAND2HSV0 U27692 ( .A1(\pe8/aot [13]), .A2(\pe8/bq[4] ), .ZN(n25568) );
  XOR2HSV0 U27693 ( .A1(n25569), .A2(n25568), .Z(n25570) );
  XOR2HSV0 U27694 ( .A1(n25571), .A2(n25570), .Z(n25572) );
  XOR3HSV2 U27695 ( .A1(n25574), .A2(n25573), .A3(n25572), .Z(n25575) );
  XOR2HSV0 U27696 ( .A1(n25576), .A2(n25575), .Z(n25580) );
  NAND2HSV0 U27697 ( .A1(n25578), .A2(n25577), .ZN(n25579) );
  XOR3HSV2 U27698 ( .A1(n25581), .A2(n25580), .A3(n25579), .Z(n25584) );
  INAND2HSV2 U27699 ( .A1(n25582), .B1(\pe8/got [5]), .ZN(n25583) );
  XOR2HSV0 U27700 ( .A1(n25584), .A2(n25583), .Z(n25585) );
  XNOR2HSV1 U27701 ( .A1(n25586), .A2(n25585), .ZN(n25588) );
  XNOR2HSV1 U27702 ( .A1(n25588), .A2(n25587), .ZN(n25589) );
  XOR2HSV0 U27703 ( .A1(n25590), .A2(n25589), .Z(n25591) );
  XOR2HSV0 U27704 ( .A1(n25592), .A2(n25591), .Z(n25593) );
  XOR2HSV0 U27705 ( .A1(n25594), .A2(n25593), .Z(n25596) );
  NAND2HSV0 U27706 ( .A1(n28618), .A2(n14059), .ZN(n25595) );
  XOR2HSV0 U27707 ( .A1(n25596), .A2(n25595), .Z(n25599) );
  NAND2HSV0 U27708 ( .A1(n28706), .A2(\pe8/got [12]), .ZN(n25598) );
  XOR2HSV0 U27709 ( .A1(n25599), .A2(n25598), .Z(n25600) );
  XNOR2HSV1 U27710 ( .A1(n25601), .A2(n25600), .ZN(n25604) );
  CLKNAND2HSV0 U27711 ( .A1(n28426), .A2(n25602), .ZN(n25603) );
  XNOR2HSV1 U27712 ( .A1(n25604), .A2(n25603), .ZN(n25617) );
  CLKAND2HSV1 U27713 ( .A1(n25618), .A2(n25617), .Z(n25621) );
  INHSV1 U27714 ( .I(n20063), .ZN(n25616) );
  CLKNHSV0 U27715 ( .I(n25605), .ZN(n25612) );
  CLKNAND2HSV0 U27716 ( .A1(n25606), .A2(\pe8/got [16]), .ZN(n25609) );
  CLKNHSV0 U27717 ( .I(n25607), .ZN(n25608) );
  NOR2HSV1 U27718 ( .A1(n25609), .A2(n25608), .ZN(n25611) );
  AOI31HSV0 U27719 ( .A1(n25613), .A2(n25612), .A3(n25611), .B(n25610), .ZN(
        n25615) );
  NAND3HSV2 U27720 ( .A1(n25616), .A2(n25615), .A3(n25614), .ZN(n25620) );
  AOI21HSV2 U27721 ( .A1(n25620), .A2(n25618), .B(n25617), .ZN(n25619) );
  AOI21HSV2 U27722 ( .A1(n25621), .A2(n25620), .B(n25619), .ZN(po8) );
  CLKNHSV0 U27723 ( .I(n28610), .ZN(n25628) );
  NAND2HSV0 U27724 ( .A1(n28697), .A2(n28693), .ZN(n25632) );
  CLKNHSV0 U27725 ( .I(n25630), .ZN(n25631) );
  XNOR2HSV1 U27726 ( .A1(n25632), .A2(n25631), .ZN(n29045) );
  XOR2HSV0 U27727 ( .A1(n25636), .A2(n25635), .Z(n28981) );
  XOR2HSV0 U27728 ( .A1(n25641), .A2(n25640), .Z(n25643) );
  XNOR2HSV1 U27729 ( .A1(n25643), .A2(n25642), .ZN(n29016) );
  XOR2HSV0 U27730 ( .A1(n14496), .A2(n12294), .Z(n25646) );
  XOR2HSV0 U27731 ( .A1(n25646), .A2(n25645), .Z(n29026) );
  CLKNAND2HSV1 U27732 ( .A1(n28649), .A2(n27218), .ZN(n25655) );
  CLKNHSV0 U27733 ( .I(n25653), .ZN(n25654) );
  XNOR2HSV1 U27734 ( .A1(n25655), .A2(n25654), .ZN(pov1[6]) );
  XNOR2HSV1 U27735 ( .A1(n25661), .A2(n25662), .ZN(n28999) );
  BUFHSV2 U27736 ( .I(n25666), .Z(n25671) );
  CLKNHSV0 U27737 ( .I(n25667), .ZN(n25670) );
  CLKNHSV0 U27738 ( .I(n25668), .ZN(n25669) );
  MUX2NHSV1 U27739 ( .I0(n25671), .I1(n25670), .S(n25669), .ZN(n29029) );
  XOR2HSV0 U27740 ( .A1(n25672), .A2(n25673), .Z(n25675) );
  XOR2HSV0 U27741 ( .A1(n25675), .A2(n25674), .Z(n28977) );
  INHSV2 U27742 ( .I(n26416), .ZN(n27139) );
  BUFHSV2 U27743 ( .I(n25683), .Z(n25684) );
  NOR2HSV2 U27744 ( .A1(n12304), .A2(n25688), .ZN(n25686) );
  XOR2HSV0 U27745 ( .A1(n25686), .A2(n25685), .Z(pov10[14]) );
  NAND2HSV2 U27746 ( .A1(\pe9/aot [1]), .A2(\pe9/bq[1] ), .ZN(n28269) );
  XOR2HSV0 U27747 ( .A1(n25693), .A2(n28269), .Z(\pe9/poht [15]) );
  XOR2HSV0 U27748 ( .A1(n25695), .A2(n25694), .Z(\pe10/poht [15]) );
  NAND2HSV0 U27749 ( .A1(n26082), .A2(\pe6/got [13]), .ZN(n25748) );
  CLKNAND2HSV1 U27750 ( .A1(n28787), .A2(n28593), .ZN(n25746) );
  CLKNAND2HSV0 U27751 ( .A1(n28467), .A2(\pe6/got [10]), .ZN(n25743) );
  NOR2HSV2 U27752 ( .A1(n25981), .A2(n25698), .ZN(n25741) );
  NAND2HSV0 U27753 ( .A1(\pe6/ti_7[7] ), .A2(n26065), .ZN(n25733) );
  NAND2HSV0 U27754 ( .A1(\pe6/got [4]), .A2(n28526), .ZN(n25731) );
  INAND2HSV0 U27755 ( .A1(n14029), .B1(\pe6/got [3]), .ZN(n25729) );
  NAND2HSV0 U27756 ( .A1(n28792), .A2(\pe6/got [2]), .ZN(n25727) );
  NAND2HSV0 U27757 ( .A1(n25849), .A2(n26083), .ZN(n25725) );
  NAND2HSV0 U27758 ( .A1(\pe6/bq[4] ), .A2(\pe6/aot [10]), .ZN(n25700) );
  NAND2HSV0 U27759 ( .A1(\pe6/aot [6]), .A2(\pe6/bq[8] ), .ZN(n25699) );
  XOR2HSV0 U27760 ( .A1(n25700), .A2(n25699), .Z(n25705) );
  NAND2HSV0 U27761 ( .A1(\pe6/bq[2] ), .A2(\pe6/aot [12]), .ZN(n25703) );
  NAND2HSV0 U27762 ( .A1(\pe6/aot [2]), .A2(n25701), .ZN(n25702) );
  XOR2HSV0 U27763 ( .A1(n25703), .A2(n25702), .Z(n25704) );
  XOR2HSV0 U27764 ( .A1(n25705), .A2(n25704), .Z(n25715) );
  NOR2HSV0 U27765 ( .A1(n25963), .A2(n25706), .ZN(n25708) );
  NAND2HSV0 U27766 ( .A1(\pe6/aot [3]), .A2(\pe6/bq[11] ), .ZN(n25707) );
  XOR2HSV0 U27767 ( .A1(n25708), .A2(n25707), .Z(n25713) );
  NAND2HSV0 U27768 ( .A1(\pe6/aot [7]), .A2(\pe6/bq[3] ), .ZN(n25755) );
  NOR2HSV0 U27769 ( .A1(n25709), .A2(n25755), .ZN(n25711) );
  AOI22HSV0 U27770 ( .A1(\pe6/aot [11]), .A2(\pe6/bq[3] ), .B1(\pe6/bq[7] ), 
        .B2(\pe6/aot [7]), .ZN(n25710) );
  NOR2HSV2 U27771 ( .A1(n25711), .A2(n25710), .ZN(n25712) );
  XNOR2HSV1 U27772 ( .A1(n25713), .A2(n25712), .ZN(n25714) );
  XNOR2HSV1 U27773 ( .A1(n25715), .A2(n25714), .ZN(n25723) );
  NAND2HSV0 U27774 ( .A1(\pe6/aot [1]), .A2(\pe6/bq[13] ), .ZN(n25721) );
  NAND2HSV0 U27775 ( .A1(\pe6/aot [9]), .A2(\pe6/bq[1] ), .ZN(n25756) );
  NAND2HSV0 U27776 ( .A1(\pe6/aot [4]), .A2(\pe6/bq[10] ), .ZN(n25718) );
  NAND2HSV0 U27777 ( .A1(\pe6/aot [5]), .A2(\pe6/bq[9] ), .ZN(n25717) );
  XOR2HSV0 U27778 ( .A1(n25718), .A2(n25717), .Z(n25719) );
  XOR3HSV2 U27779 ( .A1(n25721), .A2(n25720), .A3(n25719), .Z(n25722) );
  XNOR2HSV1 U27780 ( .A1(n25723), .A2(n25722), .ZN(n25724) );
  XNOR2HSV1 U27781 ( .A1(n25725), .A2(n25724), .ZN(n25726) );
  XNOR2HSV1 U27782 ( .A1(n25727), .A2(n25726), .ZN(n25728) );
  XNOR2HSV1 U27783 ( .A1(n25729), .A2(n25728), .ZN(n25730) );
  XNOR2HSV1 U27784 ( .A1(n25731), .A2(n25730), .ZN(n25732) );
  XNOR2HSV1 U27785 ( .A1(n25733), .A2(n25732), .ZN(n25735) );
  NAND2HSV0 U27786 ( .A1(n23041), .A2(n25982), .ZN(n25734) );
  XOR2HSV0 U27787 ( .A1(n25735), .A2(n25734), .Z(n25737) );
  INHSV2 U27788 ( .I(n25767), .ZN(n26015) );
  NOR2HSV2 U27789 ( .A1(n26015), .A2(n14418), .ZN(n25736) );
  XNOR2HSV1 U27790 ( .A1(n25737), .A2(n25736), .ZN(n25738) );
  XNOR2HSV1 U27791 ( .A1(n25739), .A2(n25738), .ZN(n25740) );
  XOR2HSV0 U27792 ( .A1(n25741), .A2(n25740), .Z(n25742) );
  NAND2HSV2 U27793 ( .A1(n25784), .A2(\pe6/got [9]), .ZN(n25783) );
  CLKNAND2HSV1 U27794 ( .A1(\pe6/got [8]), .A2(n26084), .ZN(n25782) );
  NAND2HSV0 U27795 ( .A1(\pe6/aot [2]), .A2(\pe6/bq[8] ), .ZN(n25750) );
  NAND2HSV0 U27796 ( .A1(\pe6/aot [4]), .A2(\pe6/bq[6] ), .ZN(n25749) );
  XOR2HSV0 U27797 ( .A1(n25750), .A2(n25749), .Z(n25754) );
  NAND2HSV0 U27798 ( .A1(\pe6/aot [6]), .A2(\pe6/bq[4] ), .ZN(n25752) );
  NAND2HSV0 U27799 ( .A1(\pe6/aot [3]), .A2(\pe6/bq[7] ), .ZN(n25751) );
  XOR2HSV0 U27800 ( .A1(n25752), .A2(n25751), .Z(n25753) );
  XNOR2HSV1 U27801 ( .A1(n25754), .A2(n25753), .ZN(n25758) );
  XOR2HSV0 U27802 ( .A1(n25756), .A2(n25755), .Z(n25757) );
  XNOR2HSV1 U27803 ( .A1(n25758), .A2(n25757), .ZN(n25776) );
  NAND2HSV0 U27804 ( .A1(\pe6/ti_7[7] ), .A2(n26083), .ZN(n25763) );
  NAND2HSV0 U27805 ( .A1(\pe6/aot [1]), .A2(\pe6/bq[9] ), .ZN(n25760) );
  NAND2HSV0 U27806 ( .A1(\pe6/aot [5]), .A2(\pe6/bq[5] ), .ZN(n25759) );
  XOR2HSV0 U27807 ( .A1(n25760), .A2(n25759), .Z(n25761) );
  NOR2HSV2 U27808 ( .A1(n25963), .A2(n25990), .ZN(n25961) );
  XNOR2HSV1 U27809 ( .A1(n25761), .A2(n25961), .ZN(n25762) );
  XNOR2HSV1 U27810 ( .A1(n25763), .A2(n25762), .ZN(n25766) );
  NAND2HSV0 U27811 ( .A1(n25764), .A2(\pe6/got [2]), .ZN(n25765) );
  XOR2HSV0 U27812 ( .A1(n25766), .A2(n25765), .Z(n25769) );
  XNOR2HSV1 U27813 ( .A1(n25769), .A2(n25768), .ZN(n25771) );
  CLKNHSV0 U27814 ( .I(n25771), .ZN(n25770) );
  INHSV2 U27815 ( .I(\pe6/got [4]), .ZN(n25951) );
  NOR2HSV2 U27816 ( .A1(n25770), .A2(n25951), .ZN(n25773) );
  AOI21HSV2 U27817 ( .A1(n25773), .A2(n28662), .B(n25772), .ZN(n25775) );
  NOR2HSV2 U27818 ( .A1(n25818), .A2(n26014), .ZN(n25774) );
  XOR3HSV2 U27819 ( .A1(n25776), .A2(n25775), .A3(n25774), .Z(n25778) );
  CLKNAND2HSV0 U27820 ( .A1(n28467), .A2(\pe6/got [6]), .ZN(n25777) );
  XOR2HSV0 U27821 ( .A1(n25778), .A2(n25777), .Z(n25779) );
  XOR2HSV0 U27822 ( .A1(n25780), .A2(n25779), .Z(n25781) );
  NAND2HSV0 U27823 ( .A1(n26031), .A2(\pe6/got [7]), .ZN(n25815) );
  NOR2HSV2 U27824 ( .A1(n25981), .A2(n25785), .ZN(n25813) );
  NAND2HSV0 U27825 ( .A1(n25952), .A2(n26065), .ZN(n25811) );
  NAND2HSV0 U27826 ( .A1(\pe6/ti_7[7] ), .A2(\pe6/got [2]), .ZN(n25805) );
  NAND2HSV0 U27827 ( .A1(n26083), .A2(n26033), .ZN(n25803) );
  NAND2HSV0 U27828 ( .A1(\pe6/aot [6]), .A2(\pe6/bq[5] ), .ZN(n25983) );
  NAND2HSV0 U27829 ( .A1(\pe6/bq[1] ), .A2(\pe6/aot [10]), .ZN(n25786) );
  XOR2HSV0 U27830 ( .A1(n25983), .A2(n25786), .Z(n25801) );
  NAND2HSV0 U27831 ( .A1(\pe6/aot [7]), .A2(\pe6/bq[4] ), .ZN(n25788) );
  NAND2HSV0 U27832 ( .A1(\pe6/aot [4]), .A2(\pe6/bq[7] ), .ZN(n25787) );
  XOR2HSV0 U27833 ( .A1(n25788), .A2(n25787), .Z(n25792) );
  NAND2HSV0 U27834 ( .A1(\pe6/aot [9]), .A2(\pe6/bq[2] ), .ZN(n25992) );
  NOR2HSV0 U27835 ( .A1(n25790), .A2(n25789), .ZN(n25994) );
  XNOR2HSV1 U27836 ( .A1(n25792), .A2(n25791), .ZN(n25800) );
  NAND2HSV0 U27837 ( .A1(\pe6/aot [3]), .A2(\pe6/bq[8] ), .ZN(n25794) );
  NAND2HSV0 U27838 ( .A1(\pe6/aot [1]), .A2(\pe6/bq[10] ), .ZN(n25793) );
  XOR2HSV0 U27839 ( .A1(n25794), .A2(n25793), .Z(n25798) );
  NAND2HSV0 U27840 ( .A1(\pe6/aot [2]), .A2(\pe6/bq[9] ), .ZN(n25796) );
  NAND2HSV0 U27841 ( .A1(\pe6/aot [5]), .A2(\pe6/bq[6] ), .ZN(n25795) );
  XOR2HSV0 U27842 ( .A1(n25796), .A2(n25795), .Z(n25797) );
  XOR2HSV0 U27843 ( .A1(n25798), .A2(n25797), .Z(n25799) );
  XOR3HSV2 U27844 ( .A1(n25801), .A2(n25800), .A3(n25799), .Z(n25802) );
  XNOR2HSV1 U27845 ( .A1(n25803), .A2(n25802), .ZN(n25804) );
  XNOR2HSV1 U27846 ( .A1(n25805), .A2(n25804), .ZN(n25807) );
  NAND2HSV0 U27847 ( .A1(n23041), .A2(n14008), .ZN(n25806) );
  XOR2HSV0 U27848 ( .A1(n25807), .A2(n25806), .Z(n25809) );
  NOR2HSV2 U27849 ( .A1(n26015), .A2(n25951), .ZN(n25808) );
  XNOR2HSV1 U27850 ( .A1(n25809), .A2(n25808), .ZN(n25810) );
  XNOR2HSV1 U27851 ( .A1(n25811), .A2(n25810), .ZN(n25812) );
  XOR2HSV0 U27852 ( .A1(n25813), .A2(n25812), .Z(n25814) );
  NAND2HSV0 U27853 ( .A1(n25980), .A2(n28686), .ZN(n25873) );
  NAND2HSV0 U27854 ( .A1(n26031), .A2(n14061), .ZN(n25869) );
  NOR2HSV2 U27855 ( .A1(n25818), .A2(n18860), .ZN(n25867) );
  CLKNAND2HSV0 U27856 ( .A1(n25952), .A2(\pe6/got [9]), .ZN(n25865) );
  NAND2HSV0 U27857 ( .A1(\pe6/ti_7[7] ), .A2(n25982), .ZN(n25859) );
  NAND2HSV0 U27858 ( .A1(n26033), .A2(n26065), .ZN(n25857) );
  INAND2HSV0 U27859 ( .A1(n14029), .B1(\pe6/got [4]), .ZN(n25855) );
  NAND2HSV0 U27860 ( .A1(\pe6/aot [11]), .A2(\pe6/bq[4] ), .ZN(n25820) );
  NAND2HSV0 U27861 ( .A1(\pe6/bq[3] ), .A2(\pe6/aot [12]), .ZN(n25819) );
  XOR2HSV0 U27862 ( .A1(n25820), .A2(n25819), .Z(n25824) );
  NAND2HSV0 U27863 ( .A1(\pe6/aot [5]), .A2(\pe6/bq[10] ), .ZN(n25822) );
  NAND2HSV0 U27864 ( .A1(\pe6/aot [1]), .A2(\pe6/bq[14] ), .ZN(n25821) );
  XOR2HSV0 U27865 ( .A1(n25822), .A2(n25821), .Z(n25823) );
  XOR2HSV0 U27866 ( .A1(n25824), .A2(n25823), .Z(n25832) );
  NAND2HSV0 U27867 ( .A1(\pe6/aot [4]), .A2(\pe6/bq[11] ), .ZN(n25826) );
  NAND2HSV0 U27868 ( .A1(\pe6/aot [7]), .A2(\pe6/bq[8] ), .ZN(n25825) );
  XOR2HSV0 U27869 ( .A1(n25826), .A2(n25825), .Z(n25830) );
  NAND2HSV0 U27870 ( .A1(\pe6/aot [6]), .A2(\pe6/bq[9] ), .ZN(n25828) );
  NAND2HSV0 U27871 ( .A1(\pe6/aot [14]), .A2(\pe6/bq[1] ), .ZN(n25827) );
  XOR2HSV0 U27872 ( .A1(n25828), .A2(n25827), .Z(n25829) );
  XOR2HSV0 U27873 ( .A1(n25830), .A2(n25829), .Z(n25831) );
  XOR2HSV0 U27874 ( .A1(n25832), .A2(n25831), .Z(n25845) );
  NAND2HSV0 U27875 ( .A1(\pe6/aot [8]), .A2(\pe6/bq[7] ), .ZN(n25834) );
  NAND2HSV0 U27876 ( .A1(\pe6/aot [9]), .A2(\pe6/bq[6] ), .ZN(n25833) );
  XOR2HSV0 U27877 ( .A1(n25834), .A2(n25833), .Z(n25839) );
  NOR2HSV0 U27878 ( .A1(n25835), .A2(n26043), .ZN(n25837) );
  AOI22HSV0 U27879 ( .A1(\pe6/aot [10]), .A2(\pe6/bq[5] ), .B1(\pe6/bq[13] ), 
        .B2(\pe6/aot [2]), .ZN(n25836) );
  NOR2HSV2 U27880 ( .A1(n25837), .A2(n25836), .ZN(n25838) );
  XNOR2HSV1 U27881 ( .A1(n25839), .A2(n25838), .ZN(n25843) );
  NAND2HSV0 U27882 ( .A1(\pe6/aot [3]), .A2(\pe6/bq[12] ), .ZN(n25840) );
  XOR2HSV0 U27883 ( .A1(n25841), .A2(n25840), .Z(n25842) );
  XNOR2HSV1 U27884 ( .A1(n25843), .A2(n25842), .ZN(n25844) );
  XNOR2HSV1 U27885 ( .A1(n25845), .A2(n25844), .ZN(n25848) );
  NAND2HSV0 U27886 ( .A1(n25846), .A2(n26083), .ZN(n25847) );
  XOR2HSV0 U27887 ( .A1(n25848), .A2(n25847), .Z(n25851) );
  NAND2HSV0 U27888 ( .A1(n25849), .A2(\pe6/got [2]), .ZN(n25850) );
  XOR2HSV0 U27889 ( .A1(n25851), .A2(n25850), .Z(n25853) );
  NAND2HSV0 U27890 ( .A1(n28792), .A2(\pe6/got [3]), .ZN(n25852) );
  XOR2HSV0 U27891 ( .A1(n25853), .A2(n25852), .Z(n25854) );
  XNOR2HSV1 U27892 ( .A1(n25855), .A2(n25854), .ZN(n25856) );
  XNOR2HSV1 U27893 ( .A1(n25857), .A2(n25856), .ZN(n25858) );
  XNOR2HSV1 U27894 ( .A1(n25859), .A2(n25858), .ZN(n25861) );
  NAND2HSV0 U27895 ( .A1(n23041), .A2(\pe6/got [7]), .ZN(n25860) );
  XOR2HSV0 U27896 ( .A1(n25861), .A2(n25860), .Z(n25863) );
  NAND2HSV0 U27897 ( .A1(n26068), .A2(\pe6/got [8]), .ZN(n25862) );
  XNOR2HSV1 U27898 ( .A1(n25863), .A2(n25862), .ZN(n25864) );
  XNOR2HSV1 U27899 ( .A1(n25865), .A2(n25864), .ZN(n25866) );
  XOR2HSV0 U27900 ( .A1(n25867), .A2(n25866), .Z(n25868) );
  XOR2HSV0 U27901 ( .A1(n25869), .A2(n25868), .Z(n25870) );
  NAND2HSV0 U27902 ( .A1(n25874), .A2(n28615), .ZN(n25877) );
  NAND2HSV0 U27903 ( .A1(n25875), .A2(n27184), .ZN(n25876) );
  OAI211HSV1 U27904 ( .A1(n26539), .A2(n26482), .B(n25877), .C(n25876), .ZN(
        n25918) );
  NAND2HSV0 U27905 ( .A1(n28700), .A2(\pe1/got [8]), .ZN(n25913) );
  NAND2HSV0 U27906 ( .A1(\pe1/got [7]), .A2(n28460), .ZN(n25911) );
  NOR2HSV2 U27907 ( .A1(n27139), .A2(n27140), .ZN(n25909) );
  INHSV2 U27908 ( .I(n26418), .ZN(n27004) );
  NOR2HSV2 U27909 ( .A1(n27004), .A2(n25878), .ZN(n25907) );
  CLKNAND2HSV0 U27910 ( .A1(n26854), .A2(n28435), .ZN(n25905) );
  NAND2HSV0 U27911 ( .A1(n25880), .A2(\pe1/got [2]), .ZN(n25900) );
  NAND2HSV0 U27912 ( .A1(n27166), .A2(\pe1/got [1]), .ZN(n25898) );
  NAND2HSV0 U27913 ( .A1(\pe1/aot [7]), .A2(\pe1/bq[4] ), .ZN(n27143) );
  NAND2HSV0 U27914 ( .A1(\pe1/aot [5]), .A2(\pe1/bq[6] ), .ZN(n25881) );
  XOR2HSV0 U27915 ( .A1(n27143), .A2(n25881), .Z(n25896) );
  NAND2HSV0 U27916 ( .A1(\pe1/aot [4]), .A2(\pe1/bq[7] ), .ZN(n25883) );
  NAND2HSV0 U27917 ( .A1(\pe1/aot [8]), .A2(\pe1/bq[3] ), .ZN(n25882) );
  XOR2HSV0 U27918 ( .A1(n25883), .A2(n25882), .Z(n25887) );
  NOR2HSV0 U27919 ( .A1(n27158), .A2(n26652), .ZN(n25885) );
  NAND2HSV0 U27920 ( .A1(\pe1/aot [3]), .A2(\pe1/bq[8] ), .ZN(n25884) );
  XOR2HSV0 U27921 ( .A1(n25885), .A2(n25884), .Z(n25886) );
  XNOR2HSV1 U27922 ( .A1(n25887), .A2(n25886), .ZN(n25895) );
  NAND2HSV0 U27923 ( .A1(\pe1/aot [1]), .A2(\pe1/bq[10] ), .ZN(n25889) );
  NAND2HSV0 U27924 ( .A1(\pe1/aot [10]), .A2(\pe1/bq[1] ), .ZN(n25888) );
  XOR2HSV0 U27925 ( .A1(n25889), .A2(n25888), .Z(n25893) );
  NOR2HSV0 U27926 ( .A1(n26653), .A2(n26659), .ZN(n25891) );
  NAND2HSV0 U27927 ( .A1(\pe1/aot [2]), .A2(\pe1/bq[9] ), .ZN(n25890) );
  XOR2HSV0 U27928 ( .A1(n25891), .A2(n25890), .Z(n25892) );
  XOR2HSV0 U27929 ( .A1(n25893), .A2(n25892), .Z(n25894) );
  XOR3HSV2 U27930 ( .A1(n25896), .A2(n25895), .A3(n25894), .Z(n25897) );
  XNOR2HSV1 U27931 ( .A1(n25898), .A2(n25897), .ZN(n25899) );
  XNOR2HSV1 U27932 ( .A1(n25900), .A2(n25899), .ZN(n25903) );
  NAND2HSV0 U27933 ( .A1(n25901), .A2(\pe1/got [3]), .ZN(n25902) );
  XNOR2HSV1 U27934 ( .A1(n25903), .A2(n25902), .ZN(n25904) );
  XNOR2HSV1 U27935 ( .A1(n25905), .A2(n25904), .ZN(n25906) );
  XOR2HSV0 U27936 ( .A1(n25907), .A2(n25906), .Z(n25908) );
  XOR2HSV0 U27937 ( .A1(n25909), .A2(n25908), .Z(n25910) );
  XNOR2HSV1 U27938 ( .A1(n25911), .A2(n25910), .ZN(n25912) );
  XNOR2HSV1 U27939 ( .A1(n25913), .A2(n25912), .ZN(n25916) );
  CLKNAND2HSV0 U27940 ( .A1(n26909), .A2(\pe1/got [9]), .ZN(n25915) );
  XOR2HSV0 U27941 ( .A1(n25916), .A2(n25915), .Z(n25917) );
  XOR2HSV0 U27942 ( .A1(n25917), .A2(n25918), .Z(\pe1/poht [6]) );
  NAND2HSV0 U27943 ( .A1(n25980), .A2(n28608), .ZN(n25920) );
  NAND2HSV0 U27944 ( .A1(\pe6/aot [1]), .A2(\pe6/bq[1] ), .ZN(n25919) );
  XOR2HSV0 U27945 ( .A1(n25920), .A2(n25919), .Z(\pe6/poht [15]) );
  NAND2HSV0 U27946 ( .A1(\pe6/got [7]), .A2(n26082), .ZN(n25949) );
  NAND2HSV0 U27947 ( .A1(\pe6/bq[2] ), .A2(\pe6/aot [7]), .ZN(n25962) );
  NAND2HSV0 U27948 ( .A1(\pe6/aot [7]), .A2(\pe6/bq[1] ), .ZN(n25966) );
  NAND2HSV0 U27949 ( .A1(\pe6/aot [6]), .A2(\pe6/bq[2] ), .ZN(n25921) );
  CLKNAND2HSV1 U27950 ( .A1(n25966), .A2(n25921), .ZN(n25922) );
  OAI21HSV2 U27951 ( .A1(n25923), .A2(n25962), .B(n25922), .ZN(n25925) );
  XNOR2HSV1 U27952 ( .A1(n25925), .A2(n25924), .ZN(n25929) );
  NAND2HSV0 U27953 ( .A1(\pe6/aot [1]), .A2(\pe6/bq[7] ), .ZN(n25927) );
  NAND2HSV0 U27954 ( .A1(\pe6/aot [2]), .A2(\pe6/bq[6] ), .ZN(n25926) );
  XNOR2HSV1 U27955 ( .A1(n25927), .A2(n25926), .ZN(n25928) );
  XNOR2HSV1 U27956 ( .A1(n25929), .A2(n25928), .ZN(n25931) );
  OAI21HSV2 U27957 ( .A1(n25818), .A2(n25932), .B(n25931), .ZN(n25930) );
  OAI31HSV2 U27958 ( .A1(n25818), .A2(n25932), .A3(n25931), .B(n25930), .ZN(
        n25940) );
  NAND2HSV0 U27959 ( .A1(n25952), .A2(\pe6/got [2]), .ZN(n25938) );
  CLKNAND2HSV1 U27960 ( .A1(n26068), .A2(n28608), .ZN(n25936) );
  NAND2HSV0 U27961 ( .A1(\pe6/aot [4]), .A2(\pe6/bq[4] ), .ZN(n25934) );
  NAND2HSV0 U27962 ( .A1(\pe6/aot [3]), .A2(\pe6/bq[5] ), .ZN(n25933) );
  XOR2HSV0 U27963 ( .A1(n25934), .A2(n25933), .Z(n25935) );
  XNOR2HSV1 U27964 ( .A1(n25936), .A2(n25935), .ZN(n25937) );
  XNOR2HSV1 U27965 ( .A1(n25938), .A2(n25937), .ZN(n25939) );
  XOR2HSV0 U27966 ( .A1(n25940), .A2(n25939), .Z(n25942) );
  NAND2HSV0 U27967 ( .A1(n28467), .A2(\pe6/got [4]), .ZN(n25941) );
  XNOR2HSV1 U27968 ( .A1(n25944), .A2(n25943), .ZN(n25947) );
  NAND2HSV0 U27969 ( .A1(n25945), .A2(n25982), .ZN(n25946) );
  XOR2HSV0 U27970 ( .A1(n25949), .A2(n25948), .Z(\pe6/poht [9]) );
  NAND2HSV0 U27971 ( .A1(n25980), .A2(\pe6/got [8]), .ZN(n25979) );
  NAND2HSV0 U27972 ( .A1(n25950), .A2(\pe6/got [7]), .ZN(n25977) );
  NAND2HSV0 U27973 ( .A1(n26031), .A2(n26065), .ZN(n25973) );
  NAND2HSV0 U27974 ( .A1(\pe6/aot [2]), .A2(\pe6/bq[7] ), .ZN(n25954) );
  NAND2HSV0 U27975 ( .A1(\pe6/aot [5]), .A2(\pe6/bq[4] ), .ZN(n25953) );
  XOR2HSV0 U27976 ( .A1(n25954), .A2(n25953), .Z(n25958) );
  NAND2HSV0 U27977 ( .A1(\pe6/aot [3]), .A2(\pe6/bq[6] ), .ZN(n25955) );
  XOR2HSV0 U27978 ( .A1(n25956), .A2(n25955), .Z(n25957) );
  XOR2HSV0 U27979 ( .A1(n25958), .A2(n25957), .Z(n25971) );
  NAND2HSV0 U27980 ( .A1(\pe6/aot [4]), .A2(\pe6/bq[5] ), .ZN(n25960) );
  NAND2HSV0 U27981 ( .A1(\pe6/aot [1]), .A2(\pe6/bq[8] ), .ZN(n25959) );
  XOR2HSV0 U27982 ( .A1(n25960), .A2(n25959), .Z(n25969) );
  CLKNHSV0 U27983 ( .I(n25961), .ZN(n25967) );
  OAI21HSV0 U27984 ( .A1(n25964), .A2(n25963), .B(n25962), .ZN(n25965) );
  OAI21HSV1 U27985 ( .A1(n25967), .A2(n25966), .B(n25965), .ZN(n25968) );
  XNOR2HSV1 U27986 ( .A1(n25969), .A2(n25968), .ZN(n25970) );
  XOR2HSV0 U27987 ( .A1(n25973), .A2(n25972), .Z(n25974) );
  NAND2HSV0 U27988 ( .A1(n25980), .A2(n28586), .ZN(n26029) );
  CLKNAND2HSV1 U27989 ( .A1(n26084), .A2(\pe6/got [10]), .ZN(n26027) );
  CLKNAND2HSV0 U27990 ( .A1(n28467), .A2(\pe6/got [8]), .ZN(n26023) );
  NOR2HSV2 U27991 ( .A1(n25981), .A2(n14418), .ZN(n26021) );
  NAND2HSV0 U27992 ( .A1(n28662), .A2(n25982), .ZN(n26019) );
  NAND2HSV0 U27993 ( .A1(\pe6/ti_7[7] ), .A2(n14008), .ZN(n26011) );
  NAND2HSV0 U27994 ( .A1(\pe6/got [2]), .A2(n28526), .ZN(n26009) );
  INAND2HSV0 U27995 ( .A1(n22995), .B1(n26083), .ZN(n26007) );
  NAND2HSV0 U27996 ( .A1(\pe6/aot [7]), .A2(\pe6/bq[6] ), .ZN(n26052) );
  NOR2HSV0 U27997 ( .A1(n26052), .A2(n25983), .ZN(n25985) );
  AOI22HSV0 U27998 ( .A1(\pe6/aot [7]), .A2(\pe6/bq[5] ), .B1(\pe6/bq[6] ), 
        .B2(\pe6/aot [6]), .ZN(n25984) );
  NOR2HSV2 U27999 ( .A1(n25985), .A2(n25984), .ZN(n25987) );
  NAND2HSV0 U28000 ( .A1(\pe6/aot [11]), .A2(\pe6/bq[1] ), .ZN(n25986) );
  XNOR2HSV1 U28001 ( .A1(n25987), .A2(n25986), .ZN(n26005) );
  NAND2HSV0 U28002 ( .A1(\pe6/aot [4]), .A2(\pe6/bq[8] ), .ZN(n25989) );
  NAND2HSV0 U28003 ( .A1(\pe6/aot [3]), .A2(\pe6/bq[9] ), .ZN(n25988) );
  XOR2HSV0 U28004 ( .A1(n25989), .A2(n25988), .Z(n25996) );
  CLKNHSV0 U28005 ( .I(\pe6/aot [10]), .ZN(n25991) );
  NOR2HSV0 U28006 ( .A1(n25991), .A2(n25990), .ZN(n25993) );
  NAND2HSV0 U28007 ( .A1(\pe6/bq[3] ), .A2(\pe6/aot [10]), .ZN(n26051) );
  OAI22HSV1 U28008 ( .A1(n25994), .A2(n25993), .B1(n26051), .B2(n25992), .ZN(
        n25995) );
  XNOR2HSV1 U28009 ( .A1(n25996), .A2(n25995), .ZN(n26004) );
  NAND2HSV0 U28010 ( .A1(\pe6/aot [5]), .A2(\pe6/bq[7] ), .ZN(n25998) );
  NAND2HSV0 U28011 ( .A1(\pe6/aot [8]), .A2(\pe6/bq[4] ), .ZN(n25997) );
  XOR2HSV0 U28012 ( .A1(n25998), .A2(n25997), .Z(n26002) );
  NAND2HSV0 U28013 ( .A1(\pe6/aot [1]), .A2(\pe6/bq[11] ), .ZN(n26000) );
  NAND2HSV0 U28014 ( .A1(\pe6/aot [2]), .A2(\pe6/bq[10] ), .ZN(n25999) );
  XOR2HSV0 U28015 ( .A1(n26000), .A2(n25999), .Z(n26001) );
  XOR2HSV0 U28016 ( .A1(n26002), .A2(n26001), .Z(n26003) );
  XOR3HSV2 U28017 ( .A1(n26005), .A2(n26004), .A3(n26003), .Z(n26006) );
  XNOR2HSV1 U28018 ( .A1(n26007), .A2(n26006), .ZN(n26008) );
  XNOR2HSV1 U28019 ( .A1(n26009), .A2(n26008), .ZN(n26010) );
  XNOR2HSV1 U28020 ( .A1(n26011), .A2(n26010), .ZN(n26013) );
  NAND2HSV0 U28021 ( .A1(n23041), .A2(\pe6/got [4]), .ZN(n26012) );
  XOR2HSV0 U28022 ( .A1(n26013), .A2(n26012), .Z(n26017) );
  NOR2HSV1 U28023 ( .A1(n26015), .A2(n26014), .ZN(n26016) );
  XNOR2HSV1 U28024 ( .A1(n26017), .A2(n26016), .ZN(n26018) );
  XNOR2HSV1 U28025 ( .A1(n26019), .A2(n26018), .ZN(n26020) );
  XOR2HSV0 U28026 ( .A1(n26021), .A2(n26020), .Z(n26022) );
  XOR2HSV0 U28027 ( .A1(n26023), .A2(n26022), .Z(n26024) );
  XOR2HSV0 U28028 ( .A1(n26025), .A2(n26024), .Z(n26026) );
  NAND2HSV0 U28029 ( .A1(n26082), .A2(n28593), .ZN(n26081) );
  CLKNAND2HSV1 U28030 ( .A1(n26031), .A2(\pe6/got [9]), .ZN(n26076) );
  NOR2HSV0 U28031 ( .A1(n25818), .A2(n26032), .ZN(n26074) );
  CLKNAND2HSV0 U28032 ( .A1(n28662), .A2(\pe6/got [7]), .ZN(n26072) );
  NAND2HSV0 U28033 ( .A1(\pe6/ti_7[7] ), .A2(\pe6/got [4]), .ZN(n26064) );
  NAND2HSV0 U28034 ( .A1(n26033), .A2(n14008), .ZN(n26062) );
  INAND2HSV0 U28035 ( .A1(n14029), .B1(\pe6/got [2]), .ZN(n26060) );
  NAND2HSV0 U28036 ( .A1(n28792), .A2(n26083), .ZN(n26058) );
  NAND2HSV0 U28037 ( .A1(\pe6/aot [11]), .A2(\pe6/bq[2] ), .ZN(n26036) );
  NAND2HSV0 U28038 ( .A1(\pe6/aot [6]), .A2(\pe6/bq[7] ), .ZN(n26035) );
  XOR2HSV0 U28039 ( .A1(n26036), .A2(n26035), .Z(n26040) );
  NAND2HSV0 U28040 ( .A1(\pe6/aot [4]), .A2(\pe6/bq[9] ), .ZN(n26038) );
  NAND2HSV0 U28041 ( .A1(\pe6/aot [1]), .A2(\pe6/bq[12] ), .ZN(n26037) );
  XOR2HSV0 U28042 ( .A1(n26038), .A2(n26037), .Z(n26039) );
  XOR2HSV0 U28043 ( .A1(n26040), .A2(n26039), .Z(n26050) );
  NAND2HSV0 U28044 ( .A1(\pe6/aot [9]), .A2(\pe6/bq[4] ), .ZN(n26042) );
  NAND2HSV0 U28045 ( .A1(\pe6/aot [3]), .A2(\pe6/bq[10] ), .ZN(n26041) );
  XOR2HSV0 U28046 ( .A1(n26042), .A2(n26041), .Z(n26048) );
  NOR2HSV0 U28047 ( .A1(n26044), .A2(n26043), .ZN(n26046) );
  AOI22HSV0 U28048 ( .A1(\pe6/aot [8]), .A2(\pe6/bq[5] ), .B1(\pe6/bq[11] ), 
        .B2(\pe6/aot [2]), .ZN(n26045) );
  NOR2HSV2 U28049 ( .A1(n26046), .A2(n26045), .ZN(n26047) );
  XNOR2HSV1 U28050 ( .A1(n26048), .A2(n26047), .ZN(n26049) );
  XNOR2HSV1 U28051 ( .A1(n26050), .A2(n26049), .ZN(n26056) );
  XNOR2HSV1 U28052 ( .A1(n26056), .A2(n26055), .ZN(n26057) );
  XNOR2HSV1 U28053 ( .A1(n26058), .A2(n26057), .ZN(n26059) );
  XNOR2HSV1 U28054 ( .A1(n26060), .A2(n26059), .ZN(n26061) );
  XNOR2HSV1 U28055 ( .A1(n26062), .A2(n26061), .ZN(n26063) );
  XNOR2HSV1 U28056 ( .A1(n26064), .A2(n26063), .ZN(n26067) );
  NAND2HSV0 U28057 ( .A1(n26065), .A2(n23041), .ZN(n26066) );
  XOR2HSV0 U28058 ( .A1(n26067), .A2(n26066), .Z(n26070) );
  NAND2HSV0 U28059 ( .A1(n26068), .A2(\pe6/got [6]), .ZN(n26069) );
  XNOR2HSV1 U28060 ( .A1(n26070), .A2(n26069), .ZN(n26071) );
  XNOR2HSV1 U28061 ( .A1(n26072), .A2(n26071), .ZN(n26073) );
  XOR2HSV0 U28062 ( .A1(n26074), .A2(n26073), .Z(n26075) );
  XOR2HSV0 U28063 ( .A1(n26076), .A2(n26075), .Z(n26077) );
  XOR2HSV0 U28064 ( .A1(n26081), .A2(n26080), .Z(\pe6/poht [4]) );
  NAND2HSV0 U28065 ( .A1(\pe6/got [2]), .A2(n26082), .ZN(n26090) );
  NAND2HSV0 U28066 ( .A1(\pe6/aot [2]), .A2(\pe6/bq[1] ), .ZN(n26086) );
  NAND2HSV0 U28067 ( .A1(\pe6/aot [1]), .A2(\pe6/bq[2] ), .ZN(n26085) );
  XOR2HSV0 U28068 ( .A1(n26086), .A2(n26085), .Z(n26087) );
  XOR2HSV0 U28069 ( .A1(n26090), .A2(n26089), .Z(\pe6/poht [14]) );
  NOR2HSV2 U28070 ( .A1(n27195), .A2(n26091), .ZN(n26150) );
  NOR2HSV2 U28071 ( .A1(n26093), .A2(n26092), .ZN(n26146) );
  NAND2HSV0 U28072 ( .A1(n28620), .A2(\pe10/got [7]), .ZN(n26140) );
  NAND2HSV0 U28073 ( .A1(\pe10/got [6]), .A2(n26094), .ZN(n26138) );
  NOR2HSV0 U28074 ( .A1(n26096), .A2(n26095), .ZN(n26136) );
  NAND2HSV0 U28075 ( .A1(n28794), .A2(\pe10/got [3]), .ZN(n26130) );
  NOR2HSV0 U28076 ( .A1(n26098), .A2(n26097), .ZN(n26100) );
  AOI22HSV0 U28077 ( .A1(\pe10/aot [13]), .A2(\pe10/bq[2] ), .B1(\pe10/bq[9] ), 
        .B2(\pe10/aot [6]), .ZN(n26099) );
  NOR2HSV2 U28078 ( .A1(n26100), .A2(n26099), .ZN(n26109) );
  NOR2HSV0 U28079 ( .A1(n26102), .A2(n26101), .ZN(n26104) );
  NAND2HSV0 U28080 ( .A1(\pe10/aot [9]), .A2(\pe10/bq[6] ), .ZN(n26103) );
  XOR2HSV0 U28081 ( .A1(n26104), .A2(n26103), .Z(n26108) );
  XOR2HSV0 U28082 ( .A1(n26106), .A2(n26105), .Z(n26107) );
  XOR3HSV2 U28083 ( .A1(n26109), .A2(n26108), .A3(n26107), .Z(n26126) );
  NAND2HSV0 U28084 ( .A1(\pe10/aot [1]), .A2(\pe10/bq[14] ), .ZN(n26111) );
  NAND2HSV0 U28085 ( .A1(\pe10/bq[1] ), .A2(\pe10/aot [14]), .ZN(n26110) );
  XOR2HSV0 U28086 ( .A1(n26111), .A2(n26110), .Z(n26115) );
  NAND2HSV0 U28087 ( .A1(\pe10/aot [8]), .A2(\pe10/bq[7] ), .ZN(n26113) );
  NAND2HSV0 U28088 ( .A1(\pe10/aot [4]), .A2(\pe10/bq[11] ), .ZN(n26112) );
  XOR2HSV0 U28089 ( .A1(n26113), .A2(n26112), .Z(n26114) );
  XOR2HSV0 U28090 ( .A1(n26115), .A2(n26114), .Z(n26123) );
  NAND2HSV0 U28091 ( .A1(\pe10/aot [11]), .A2(\pe10/bq[4] ), .ZN(n26117) );
  NAND2HSV0 U28092 ( .A1(\pe10/aot [12]), .A2(\pe10/bq[3] ), .ZN(n26116) );
  XOR2HSV0 U28093 ( .A1(n26117), .A2(n26116), .Z(n26121) );
  NAND2HSV0 U28094 ( .A1(\pe10/aot [10]), .A2(\pe10/bq[5] ), .ZN(n26119) );
  NAND2HSV0 U28095 ( .A1(\pe10/aot [5]), .A2(\pe10/bq[10] ), .ZN(n26118) );
  XOR2HSV0 U28096 ( .A1(n26119), .A2(n26118), .Z(n26120) );
  XOR2HSV0 U28097 ( .A1(n26121), .A2(n26120), .Z(n26122) );
  XOR2HSV0 U28098 ( .A1(n26123), .A2(n26122), .Z(n26125) );
  NAND2HSV0 U28099 ( .A1(n16850), .A2(n27196), .ZN(n26124) );
  XOR3HSV2 U28100 ( .A1(n26126), .A2(n26125), .A3(n26124), .Z(n26128) );
  NAND2HSV0 U28101 ( .A1(n28679), .A2(n14065), .ZN(n26127) );
  XNOR2HSV1 U28102 ( .A1(n26128), .A2(n26127), .ZN(n26129) );
  XNOR2HSV1 U28103 ( .A1(n26130), .A2(n26129), .ZN(n26134) );
  NAND2HSV0 U28104 ( .A1(n26132), .A2(n26131), .ZN(n26133) );
  XNOR2HSV1 U28105 ( .A1(n26134), .A2(n26133), .ZN(n26135) );
  XOR2HSV0 U28106 ( .A1(n26136), .A2(n26135), .Z(n26137) );
  XOR2HSV0 U28107 ( .A1(n26138), .A2(n26137), .Z(n26139) );
  XOR2HSV0 U28108 ( .A1(n26140), .A2(n26139), .Z(n26142) );
  NAND2HSV0 U28109 ( .A1(n28585), .A2(n28642), .ZN(n26141) );
  XOR2HSV0 U28110 ( .A1(n26142), .A2(n26141), .Z(n26144) );
  NAND2HSV0 U28111 ( .A1(n26209), .A2(\pe10/got [9]), .ZN(n26143) );
  XNOR2HSV1 U28112 ( .A1(n26144), .A2(n26143), .ZN(n26145) );
  XOR2HSV0 U28113 ( .A1(n26146), .A2(n26145), .Z(n26148) );
  NAND2HSV0 U28114 ( .A1(n28469), .A2(\pe10/got [11]), .ZN(n26147) );
  XOR2HSV0 U28115 ( .A1(n26148), .A2(n26147), .Z(n26149) );
  XOR2HSV2 U28116 ( .A1(n26150), .A2(n26149), .Z(n26152) );
  NAND2HSV0 U28117 ( .A1(n26221), .A2(n14070), .ZN(n26154) );
  XOR2HSV0 U28118 ( .A1(n26155), .A2(n26154), .Z(\pe10/poht [2]) );
  NOR2HSV2 U28119 ( .A1(n27195), .A2(n26156), .ZN(n26217) );
  NAND2HSV0 U28120 ( .A1(n28620), .A2(\pe10/got [9]), .ZN(n26208) );
  NAND2HSV0 U28121 ( .A1(n28642), .A2(n26157), .ZN(n26206) );
  NOR2HSV0 U28122 ( .A1(n26159), .A2(n26158), .ZN(n26204) );
  NAND2HSV0 U28123 ( .A1(n28794), .A2(\pe10/got [5]), .ZN(n26198) );
  NAND2HSV0 U28124 ( .A1(\pe10/aot [13]), .A2(\pe10/bq[4] ), .ZN(n26160) );
  XOR2HSV0 U28125 ( .A1(n26161), .A2(n26160), .Z(n26178) );
  XNOR2HSV1 U28126 ( .A1(n26169), .A2(n26168), .ZN(n26177) );
  NAND2HSV0 U28127 ( .A1(\pe10/aot [8]), .A2(\pe10/bq[9] ), .ZN(n26171) );
  NAND2HSV0 U28128 ( .A1(\pe10/bq[3] ), .A2(\pe10/aot [14]), .ZN(n26170) );
  XOR2HSV0 U28129 ( .A1(n26171), .A2(n26170), .Z(n26175) );
  NAND2HSV0 U28130 ( .A1(\pe10/aot [12]), .A2(\pe10/bq[5] ), .ZN(n26173) );
  NAND2HSV0 U28131 ( .A1(\pe10/aot [7]), .A2(\pe10/bq[10] ), .ZN(n26172) );
  XOR2HSV0 U28132 ( .A1(n26173), .A2(n26172), .Z(n26174) );
  XOR2HSV0 U28133 ( .A1(n26175), .A2(n26174), .Z(n26176) );
  XOR3HSV2 U28134 ( .A1(n26178), .A2(n26177), .A3(n26176), .Z(n26194) );
  NAND2HSV0 U28135 ( .A1(n28630), .A2(\pe10/got [3]), .ZN(n26193) );
  NAND2HSV0 U28136 ( .A1(n28811), .A2(\pe10/pq ), .ZN(n26180) );
  NAND2HSV0 U28137 ( .A1(\pe10/aot [4]), .A2(\pe10/bq[13] ), .ZN(n26179) );
  XOR2HSV0 U28138 ( .A1(n26180), .A2(n26179), .Z(n26184) );
  NAND2HSV0 U28139 ( .A1(\pe10/aot [10]), .A2(\pe10/bq[7] ), .ZN(n26182) );
  NAND2HSV0 U28140 ( .A1(\pe10/aot [6]), .A2(\pe10/bq[11] ), .ZN(n26181) );
  XOR2HSV0 U28141 ( .A1(n26182), .A2(n26181), .Z(n26183) );
  XOR2HSV0 U28142 ( .A1(n26184), .A2(n26183), .Z(n26188) );
  XOR2HSV0 U28143 ( .A1(n26188), .A2(n26187), .Z(n26191) );
  NAND2HSV0 U28144 ( .A1(n26189), .A2(n14065), .ZN(n26190) );
  XNOR2HSV1 U28145 ( .A1(n26191), .A2(n26190), .ZN(n26192) );
  XOR3HSV2 U28146 ( .A1(n26194), .A2(n26193), .A3(n26192), .Z(n26196) );
  NAND2HSV0 U28147 ( .A1(n28679), .A2(n26132), .ZN(n26195) );
  XNOR2HSV1 U28148 ( .A1(n26196), .A2(n26195), .ZN(n26197) );
  XNOR2HSV1 U28149 ( .A1(n26198), .A2(n26197), .ZN(n26202) );
  NOR2HSV0 U28150 ( .A1(n26200), .A2(n26199), .ZN(n26201) );
  XNOR2HSV1 U28151 ( .A1(n26202), .A2(n26201), .ZN(n26203) );
  XOR2HSV0 U28152 ( .A1(n26204), .A2(n26203), .Z(n26205) );
  XNOR2HSV1 U28153 ( .A1(n26206), .A2(n26205), .ZN(n26207) );
  NAND2HSV0 U28154 ( .A1(n26209), .A2(n16759), .ZN(n26210) );
  CLKAND2HSV0 U28155 ( .A1(n26210), .A2(n26212), .Z(n26214) );
  CLKNHSV1 U28156 ( .I(n26210), .ZN(n26211) );
  IOA21HSV2 U28157 ( .A1(n26215), .A2(\pe10/got [12]), .B(n26211), .ZN(n26213)
         );
  NAND2HSV0 U28158 ( .A1(n26229), .A2(n26230), .ZN(n26223) );
  XOR2HSV0 U28159 ( .A1(n26223), .A2(n26222), .Z(\pe8/poht [15]) );
  NAND2HSV0 U28160 ( .A1(n28426), .A2(n26230), .ZN(n26228) );
  NAND2HSV0 U28161 ( .A1(\pe8/aot [3]), .A2(\pe8/bq[1] ), .ZN(n26225) );
  NAND2HSV0 U28162 ( .A1(\pe8/aot [1]), .A2(\pe8/bq[3] ), .ZN(n26224) );
  XOR2HSV0 U28163 ( .A1(n26225), .A2(n26224), .Z(n26227) );
  NAND2HSV0 U28164 ( .A1(\pe8/aot [2]), .A2(\pe8/bq[1] ), .ZN(n26233) );
  NAND2HSV0 U28165 ( .A1(\pe8/aot [1]), .A2(\pe8/bq[2] ), .ZN(n26232) );
  XOR2HSV0 U28166 ( .A1(n26233), .A2(n26232), .Z(n26234) );
  XOR2HSV0 U28167 ( .A1(n26235), .A2(n26234), .Z(n26236) );
  XOR2HSV0 U28168 ( .A1(n26237), .A2(n26236), .Z(\pe8/poht [14]) );
  NAND2HSV2 U28169 ( .A1(n28461), .A2(\pe4/got [1]), .ZN(n26239) );
  NAND2HSV0 U28170 ( .A1(\pe4/aot [1]), .A2(\pe4/bq[1] ), .ZN(n26238) );
  XOR2HSV0 U28171 ( .A1(n26239), .A2(n26238), .Z(\pe4/poht [15]) );
  NOR2HSV2 U28172 ( .A1(n26602), .A2(n26241), .ZN(n26295) );
  NAND2HSV0 U28173 ( .A1(n26297), .A2(\pe3/got [9]), .ZN(n26288) );
  NAND2HSV0 U28174 ( .A1(n23327), .A2(n28648), .ZN(n26286) );
  CLKNAND2HSV0 U28175 ( .A1(n28588), .A2(\pe3/got [7]), .ZN(n26284) );
  NAND2HSV0 U28176 ( .A1(n26682), .A2(\pe3/got [6]), .ZN(n26280) );
  NAND2HSV0 U28177 ( .A1(n15240), .A2(\pe3/got [4]), .ZN(n26278) );
  NAND2HSV0 U28178 ( .A1(n26350), .A2(\pe3/got [2]), .ZN(n26276) );
  NAND2HSV0 U28179 ( .A1(n26242), .A2(n26751), .ZN(n26275) );
  NOR2HSV0 U28180 ( .A1(n26243), .A2(n26683), .ZN(n26245) );
  AOI22HSV0 U28181 ( .A1(\pe3/aot [14]), .A2(\pe3/bq[2] ), .B1(\pe3/bq[12] ), 
        .B2(\pe3/aot [4]), .ZN(n26244) );
  NOR2HSV2 U28182 ( .A1(n26245), .A2(n26244), .ZN(n26248) );
  NOR2HSV0 U28183 ( .A1(n26247), .A2(n26246), .ZN(n26308) );
  XNOR2HSV1 U28184 ( .A1(n26248), .A2(n26308), .ZN(n26258) );
  NAND2HSV0 U28185 ( .A1(\pe3/aot [11]), .A2(\pe3/bq[5] ), .ZN(n26250) );
  NAND2HSV0 U28186 ( .A1(\pe3/aot [10]), .A2(\pe3/bq[6] ), .ZN(n26249) );
  XOR2HSV0 U28187 ( .A1(n26250), .A2(n26249), .Z(n26254) );
  NAND2HSV0 U28188 ( .A1(\pe3/aot [5]), .A2(\pe3/bq[11] ), .ZN(n26252) );
  NAND2HSV0 U28189 ( .A1(\pe3/aot [12]), .A2(\pe3/bq[4] ), .ZN(n26251) );
  XOR2HSV0 U28190 ( .A1(n26252), .A2(n26251), .Z(n26253) );
  XOR2HSV0 U28191 ( .A1(n26254), .A2(n26253), .Z(n26257) );
  NAND2HSV0 U28192 ( .A1(n26255), .A2(\pe3/got [1]), .ZN(n26256) );
  XOR3HSV2 U28193 ( .A1(n26258), .A2(n26257), .A3(n26256), .Z(n26273) );
  NAND2HSV0 U28194 ( .A1(\pe3/aot [7]), .A2(\pe3/bq[9] ), .ZN(n26260) );
  NAND2HSV0 U28195 ( .A1(n11932), .A2(\pe3/bq[3] ), .ZN(n26259) );
  XOR2HSV0 U28196 ( .A1(n26260), .A2(n26259), .Z(n26264) );
  NAND2HSV0 U28197 ( .A1(\pe3/aot [1]), .A2(n26373), .ZN(n26262) );
  NAND2HSV0 U28198 ( .A1(\pe3/aot [2]), .A2(n14026), .ZN(n26261) );
  XOR2HSV0 U28199 ( .A1(n26262), .A2(n26261), .Z(n26263) );
  XOR2HSV0 U28200 ( .A1(n26264), .A2(n26263), .Z(n26271) );
  NAND2HSV0 U28201 ( .A1(\pe3/bq[8] ), .A2(\pe3/aot [8]), .ZN(n26740) );
  XOR2HSV0 U28202 ( .A1(n26740), .A2(n26265), .Z(n26269) );
  NAND2HSV0 U28203 ( .A1(\pe3/aot [6]), .A2(\pe3/bq[10] ), .ZN(n26267) );
  NAND2HSV0 U28204 ( .A1(\pe3/bq[1] ), .A2(\pe3/aot [15]), .ZN(n26266) );
  XOR2HSV0 U28205 ( .A1(n26267), .A2(n26266), .Z(n26268) );
  XOR2HSV0 U28206 ( .A1(n26269), .A2(n26268), .Z(n26270) );
  XOR2HSV0 U28207 ( .A1(n26271), .A2(n26270), .Z(n26272) );
  XNOR2HSV1 U28208 ( .A1(n26273), .A2(n26272), .ZN(n26274) );
  XOR3HSV1 U28209 ( .A1(n26276), .A2(n26275), .A3(n26274), .Z(n26277) );
  XNOR2HSV1 U28210 ( .A1(n26278), .A2(n26277), .ZN(n26279) );
  XNOR2HSV1 U28211 ( .A1(n26280), .A2(n26279), .ZN(n26282) );
  NOR2HSV0 U28212 ( .A1(n26714), .A2(n23329), .ZN(n26281) );
  XNOR2HSV1 U28213 ( .A1(n26282), .A2(n26281), .ZN(n26283) );
  XNOR2HSV1 U28214 ( .A1(n26284), .A2(n26283), .ZN(n26285) );
  XNOR2HSV1 U28215 ( .A1(n26286), .A2(n26285), .ZN(n26287) );
  XOR2HSV0 U28216 ( .A1(n26288), .A2(n26287), .Z(n26290) );
  NAND2HSV0 U28217 ( .A1(n26752), .A2(\pe3/got [10]), .ZN(n26289) );
  XOR2HSV0 U28218 ( .A1(n26290), .A2(n26289), .Z(n26293) );
  NAND2HSV0 U28219 ( .A1(\pe3/got [11]), .A2(n26291), .ZN(n26292) );
  XNOR2HSV1 U28220 ( .A1(n26293), .A2(n26292), .ZN(n26294) );
  NOR2HSV2 U28221 ( .A1(n26681), .A2(n26296), .ZN(n26347) );
  NAND2HSV0 U28222 ( .A1(n26297), .A2(n28648), .ZN(n26341) );
  NAND2HSV0 U28223 ( .A1(n23327), .A2(\pe3/got [7]), .ZN(n26339) );
  NAND2HSV0 U28224 ( .A1(n28588), .A2(\pe3/got [6]), .ZN(n26337) );
  NAND2HSV0 U28225 ( .A1(\pe3/got [5]), .A2(n26682), .ZN(n26332) );
  NAND2HSV0 U28226 ( .A1(n16112), .A2(n26751), .ZN(n26330) );
  NAND2HSV0 U28227 ( .A1(\pe3/aot [9]), .A2(\pe3/bq[6] ), .ZN(n26299) );
  NAND2HSV0 U28228 ( .A1(\pe3/aot [8]), .A2(\pe3/bq[7] ), .ZN(n26298) );
  XOR2HSV0 U28229 ( .A1(n26299), .A2(n26298), .Z(n26324) );
  NAND2HSV0 U28230 ( .A1(\pe3/aot [14]), .A2(\pe3/bq[1] ), .ZN(n26301) );
  NAND2HSV0 U28231 ( .A1(n11932), .A2(\pe3/bq[2] ), .ZN(n26300) );
  XOR2HSV0 U28232 ( .A1(n26301), .A2(n26300), .Z(n26305) );
  NAND2HSV0 U28233 ( .A1(\pe3/aot [10]), .A2(\pe3/bq[5] ), .ZN(n26303) );
  NAND2HSV0 U28234 ( .A1(\pe3/aot [7]), .A2(\pe3/bq[8] ), .ZN(n26302) );
  XOR2HSV0 U28235 ( .A1(n26303), .A2(n26302), .Z(n26304) );
  XNOR2HSV1 U28236 ( .A1(n26305), .A2(n26304), .ZN(n26323) );
  AOI22HSV0 U28237 ( .A1(\pe3/aot [3]), .A2(\pe3/bq[12] ), .B1(\pe3/bq[13] ), 
        .B2(\pe3/aot [2]), .ZN(n26306) );
  AOI21HSV1 U28238 ( .A1(n26308), .A2(n26307), .B(n26306), .ZN(n26314) );
  NOR2HSV0 U28239 ( .A1(n26310), .A2(n26309), .ZN(n26312) );
  AOI22HSV0 U28240 ( .A1(\pe3/aot [12]), .A2(\pe3/bq[3] ), .B1(n14026), .B2(
        \pe3/aot [1]), .ZN(n26311) );
  NOR2HSV1 U28241 ( .A1(n26312), .A2(n26311), .ZN(n26313) );
  XOR2HSV0 U28242 ( .A1(n26314), .A2(n26313), .Z(n26322) );
  NAND2HSV0 U28243 ( .A1(\pe3/aot [4]), .A2(\pe3/bq[11] ), .ZN(n26316) );
  NAND2HSV0 U28244 ( .A1(\pe3/aot [11]), .A2(\pe3/bq[4] ), .ZN(n26315) );
  XOR2HSV0 U28245 ( .A1(n26316), .A2(n26315), .Z(n26320) );
  NAND2HSV0 U28246 ( .A1(\pe3/aot [6]), .A2(\pe3/bq[9] ), .ZN(n26318) );
  NAND2HSV0 U28247 ( .A1(\pe3/aot [5]), .A2(\pe3/bq[10] ), .ZN(n26317) );
  XOR2HSV0 U28248 ( .A1(n26318), .A2(n26317), .Z(n26319) );
  XOR2HSV0 U28249 ( .A1(n26320), .A2(n26319), .Z(n26321) );
  XOR4HSV1 U28250 ( .A1(n26324), .A2(n26323), .A3(n26322), .A4(n26321), .Z(
        n26326) );
  NAND2HSV0 U28251 ( .A1(n26350), .A2(\pe3/got [1]), .ZN(n26325) );
  XOR2HSV0 U28252 ( .A1(n26326), .A2(n26325), .Z(n26328) );
  NAND2HSV0 U28253 ( .A1(n28920), .A2(\pe3/got [2]), .ZN(n26327) );
  XNOR2HSV1 U28254 ( .A1(n26328), .A2(n26327), .ZN(n26329) );
  XNOR2HSV1 U28255 ( .A1(n26330), .A2(n26329), .ZN(n26331) );
  XNOR2HSV1 U28256 ( .A1(n26332), .A2(n26331), .ZN(n26335) );
  NOR2HSV0 U28257 ( .A1(n26714), .A2(n26333), .ZN(n26334) );
  XNOR2HSV1 U28258 ( .A1(n26335), .A2(n26334), .ZN(n26336) );
  XNOR2HSV1 U28259 ( .A1(n26337), .A2(n26336), .ZN(n26338) );
  XNOR2HSV1 U28260 ( .A1(n26339), .A2(n26338), .ZN(n26340) );
  XOR2HSV0 U28261 ( .A1(n26341), .A2(n26340), .Z(n26343) );
  NAND2HSV0 U28262 ( .A1(n26752), .A2(\pe3/got [9]), .ZN(n26342) );
  XOR2HSV0 U28263 ( .A1(n26343), .A2(n26342), .Z(n26345) );
  NAND2HSV0 U28264 ( .A1(\pe3/got [10]), .A2(n28584), .ZN(n26344) );
  XOR2HSV0 U28265 ( .A1(n26345), .A2(n26344), .Z(n26346) );
  NAND2HSV0 U28266 ( .A1(n28438), .A2(\pe3/got [10]), .ZN(n26405) );
  NAND2HSV0 U28267 ( .A1(n23327), .A2(n26642), .ZN(n26403) );
  NAND2HSV0 U28268 ( .A1(n28588), .A2(n28648), .ZN(n26401) );
  NAND2HSV0 U28269 ( .A1(n26682), .A2(\pe3/got [7]), .ZN(n26396) );
  NAND2HSV0 U28270 ( .A1(n15240), .A2(n26603), .ZN(n26394) );
  NAND2HSV0 U28271 ( .A1(n26350), .A2(n26751), .ZN(n26392) );
  NAND2HSV0 U28272 ( .A1(n28920), .A2(\pe3/got [4]), .ZN(n26391) );
  NAND2HSV0 U28273 ( .A1(\pe3/aot [1]), .A2(n26351), .ZN(n26353) );
  NAND2HSV0 U28274 ( .A1(\pe3/aot [12]), .A2(\pe3/bq[5] ), .ZN(n26352) );
  XOR2HSV0 U28275 ( .A1(n26353), .A2(n26352), .Z(n26357) );
  NAND2HSV0 U28276 ( .A1(\pe3/aot [11]), .A2(\pe3/bq[6] ), .ZN(n26355) );
  NAND2HSV0 U28277 ( .A1(\pe3/aot [9]), .A2(\pe3/bq[8] ), .ZN(n26354) );
  XOR2HSV0 U28278 ( .A1(n26355), .A2(n26354), .Z(n26356) );
  XOR2HSV0 U28279 ( .A1(n26357), .A2(n26356), .Z(n26366) );
  NAND2HSV0 U28280 ( .A1(n26358), .A2(\pe3/bq[1] ), .ZN(n26360) );
  NAND2HSV0 U28281 ( .A1(\pe3/aot [15]), .A2(\pe3/bq[2] ), .ZN(n26359) );
  XOR2HSV0 U28282 ( .A1(n26360), .A2(n26359), .Z(n26364) );
  NAND2HSV0 U28283 ( .A1(\pe3/aot [3]), .A2(\pe3/bq[14] ), .ZN(n26362) );
  NAND2HSV0 U28284 ( .A1(\pe3/aot [4]), .A2(\pe3/bq[13] ), .ZN(n26361) );
  XOR2HSV0 U28285 ( .A1(n26362), .A2(n26361), .Z(n26363) );
  XOR2HSV0 U28286 ( .A1(n26364), .A2(n26363), .Z(n26365) );
  XOR2HSV0 U28287 ( .A1(n26366), .A2(n26365), .Z(n26369) );
  NAND2HSV0 U28288 ( .A1(n26367), .A2(\pe3/got [2]), .ZN(n26368) );
  XNOR2HSV1 U28289 ( .A1(n26369), .A2(n26368), .ZN(n26389) );
  NAND2HSV0 U28290 ( .A1(\pe3/bq[10] ), .A2(\pe3/aot [7]), .ZN(n26605) );
  XOR2HSV0 U28291 ( .A1(n26370), .A2(n26605), .Z(n26387) );
  NAND2HSV0 U28292 ( .A1(\pe3/aot [8]), .A2(\pe3/bq[9] ), .ZN(n26372) );
  NAND2HSV0 U28293 ( .A1(\pe3/aot [14]), .A2(\pe3/bq[3] ), .ZN(n26371) );
  XOR2HSV0 U28294 ( .A1(n26372), .A2(n26371), .Z(n26377) );
  NAND2HSV0 U28295 ( .A1(n11932), .A2(\pe3/bq[4] ), .ZN(n26375) );
  NAND2HSV0 U28296 ( .A1(\pe3/aot [2]), .A2(n26373), .ZN(n26374) );
  XOR2HSV0 U28297 ( .A1(n26375), .A2(n26374), .Z(n26376) );
  XNOR2HSV1 U28298 ( .A1(n26377), .A2(n26376), .ZN(n26386) );
  NAND2HSV2 U28299 ( .A1(n15937), .A2(\pe3/pq ), .ZN(n26379) );
  NAND2HSV0 U28300 ( .A1(\pe3/aot [10]), .A2(\pe3/bq[7] ), .ZN(n26378) );
  XOR2HSV0 U28301 ( .A1(n26379), .A2(n26378), .Z(n26384) );
  NAND2HSV0 U28302 ( .A1(\pe3/got [1]), .A2(n26380), .ZN(n26382) );
  NAND2HSV0 U28303 ( .A1(\pe3/aot [5]), .A2(\pe3/bq[12] ), .ZN(n26381) );
  XOR2HSV0 U28304 ( .A1(n26382), .A2(n26381), .Z(n26383) );
  XOR2HSV0 U28305 ( .A1(n26384), .A2(n26383), .Z(n26385) );
  XOR3HSV2 U28306 ( .A1(n26387), .A2(n26386), .A3(n26385), .Z(n26388) );
  XNOR2HSV1 U28307 ( .A1(n26389), .A2(n26388), .ZN(n26390) );
  XOR3HSV1 U28308 ( .A1(n26392), .A2(n26391), .A3(n26390), .Z(n26393) );
  XNOR2HSV1 U28309 ( .A1(n26394), .A2(n26393), .ZN(n26395) );
  XNOR2HSV1 U28310 ( .A1(n26396), .A2(n26395), .ZN(n26399) );
  NOR2HSV0 U28311 ( .A1(n26714), .A2(n26397), .ZN(n26398) );
  XNOR2HSV1 U28312 ( .A1(n26399), .A2(n26398), .ZN(n26400) );
  XNOR2HSV1 U28313 ( .A1(n26401), .A2(n26400), .ZN(n26402) );
  XNOR2HSV1 U28314 ( .A1(n26403), .A2(n26402), .ZN(n26404) );
  XOR2HSV0 U28315 ( .A1(n26405), .A2(n26404), .Z(n26407) );
  NAND2HSV0 U28316 ( .A1(n26634), .A2(\pe3/got [11]), .ZN(n26406) );
  XOR2HSV0 U28317 ( .A1(n26407), .A2(n26406), .Z(n26409) );
  NAND2HSV0 U28318 ( .A1(n11891), .A2(n26637), .ZN(n26408) );
  XOR2HSV0 U28319 ( .A1(n26409), .A2(n26408), .Z(n26410) );
  XOR2HSV0 U28320 ( .A1(n26411), .A2(n26410), .Z(n26412) );
  CLKNAND2HSV3 U28321 ( .A1(n26415), .A2(n26414), .ZN(n27136) );
  CLKNAND2HSV0 U28322 ( .A1(n27136), .A2(\pe1/got [14]), .ZN(n26476) );
  NAND2HSV0 U28323 ( .A1(n27137), .A2(\pe1/got [13]), .ZN(n26474) );
  INHSV2 U28324 ( .I(n26416), .ZN(n26888) );
  NOR2HSV1 U28325 ( .A1(n26888), .A2(n26417), .ZN(n26472) );
  CLKNHSV0 U28326 ( .I(\pe1/got [11]), .ZN(n26538) );
  NOR2HSV2 U28327 ( .A1(n26830), .A2(n26538), .ZN(n26470) );
  CLKNAND2HSV0 U28328 ( .A1(n26854), .A2(n28615), .ZN(n26468) );
  NAND2HSV0 U28329 ( .A1(n28609), .A2(\pe1/got [8]), .ZN(n26464) );
  NAND2HSV0 U28330 ( .A1(n27005), .A2(\pe1/got [4]), .ZN(n26457) );
  NAND2HSV0 U28331 ( .A1(\pe1/bq[1] ), .A2(\pe1/aot [13]), .ZN(n27024) );
  AO22HSV2 U28332 ( .A1(\pe1/bq[1] ), .A2(n28485), .B1(\pe1/aot [13]), .B2(
        \pe1/bq[4] ), .Z(n26419) );
  OAI21HSV0 U28333 ( .A1(n27024), .A2(n26420), .B(n26419), .ZN(n26425) );
  NAND2HSV0 U28334 ( .A1(\pe1/aot [14]), .A2(\pe1/bq[2] ), .ZN(n26557) );
  NOR2HSV0 U28335 ( .A1(n26421), .A2(n26557), .ZN(n26423) );
  AOI22HSV0 U28336 ( .A1(n28468), .A2(\pe1/bq[2] ), .B1(\pe1/aot [14]), .B2(
        \pe1/bq[3] ), .ZN(n26422) );
  NOR2HSV1 U28337 ( .A1(n26423), .A2(n26422), .ZN(n26424) );
  XOR2HSV0 U28338 ( .A1(n26425), .A2(n26424), .Z(n26428) );
  NAND2HSV0 U28339 ( .A1(n26426), .A2(\pe1/got [2]), .ZN(n26427) );
  XOR2HSV0 U28340 ( .A1(n26428), .A2(n26427), .Z(n26455) );
  NAND2HSV0 U28341 ( .A1(\pe1/aot [10]), .A2(\pe1/bq[7] ), .ZN(n26430) );
  NAND2HSV0 U28342 ( .A1(\pe1/aot [7]), .A2(\pe1/bq[10] ), .ZN(n26429) );
  XOR2HSV0 U28343 ( .A1(n26430), .A2(n26429), .Z(n26435) );
  NAND2HSV0 U28344 ( .A1(\pe1/aot [6]), .A2(\pe1/bq[11] ), .ZN(n26433) );
  NAND2HSV0 U28345 ( .A1(\pe1/aot [2]), .A2(n26431), .ZN(n26432) );
  XOR2HSV0 U28346 ( .A1(n26433), .A2(n26432), .Z(n26434) );
  XOR2HSV0 U28347 ( .A1(n26435), .A2(n26434), .Z(n26443) );
  NAND2HSV0 U28348 ( .A1(\pe1/aot [5]), .A2(\pe1/bq[12] ), .ZN(n26438) );
  NAND2HSV0 U28349 ( .A1(\pe1/aot [1]), .A2(n26436), .ZN(n26437) );
  XOR2HSV0 U28350 ( .A1(n26438), .A2(n26437), .Z(n26441) );
  NAND2HSV0 U28351 ( .A1(\pe1/aot [4]), .A2(\pe1/bq[5] ), .ZN(n26858) );
  XNOR2HSV1 U28352 ( .A1(n26441), .A2(n26440), .ZN(n26442) );
  XNOR2HSV1 U28353 ( .A1(n26443), .A2(n26442), .ZN(n26454) );
  NAND2HSV0 U28354 ( .A1(n26444), .A2(\pe1/got [3]), .ZN(n26452) );
  NAND2HSV0 U28355 ( .A1(\pe1/aot [9]), .A2(\pe1/bq[8] ), .ZN(n26446) );
  NAND2HSV0 U28356 ( .A1(\pe1/aot [11]), .A2(\pe1/bq[6] ), .ZN(n26445) );
  XOR2HSV0 U28357 ( .A1(n26446), .A2(n26445), .Z(n26450) );
  NAND2HSV0 U28358 ( .A1(\pe1/aot [8]), .A2(\pe1/bq[9] ), .ZN(n26448) );
  NAND2HSV0 U28359 ( .A1(\pe1/aot [3]), .A2(\pe1/bq[14] ), .ZN(n26447) );
  XOR2HSV0 U28360 ( .A1(n26448), .A2(n26447), .Z(n26449) );
  XOR2HSV0 U28361 ( .A1(n26450), .A2(n26449), .Z(n26451) );
  XOR2HSV0 U28362 ( .A1(n26452), .A2(n26451), .Z(n26453) );
  XOR3HSV2 U28363 ( .A1(n26455), .A2(n26454), .A3(n26453), .Z(n26456) );
  XNOR2HSV1 U28364 ( .A1(n26457), .A2(n26456), .ZN(n26459) );
  NAND2HSV0 U28365 ( .A1(n28635), .A2(\pe1/got [5]), .ZN(n26458) );
  XNOR2HSV1 U28366 ( .A1(n26459), .A2(n26458), .ZN(n26462) );
  NAND2HSV0 U28367 ( .A1(n28649), .A2(n28434), .ZN(n26461) );
  NAND2HSV0 U28368 ( .A1(n27166), .A2(\pe1/got [7]), .ZN(n26460) );
  XOR3HSV2 U28369 ( .A1(n26462), .A2(n26461), .A3(n26460), .Z(n26463) );
  XNOR2HSV1 U28370 ( .A1(n26464), .A2(n26463), .ZN(n26466) );
  NAND2HSV0 U28371 ( .A1(n28589), .A2(\pe1/got [9]), .ZN(n26465) );
  XNOR2HSV1 U28372 ( .A1(n26466), .A2(n26465), .ZN(n26467) );
  XNOR2HSV1 U28373 ( .A1(n26468), .A2(n26467), .ZN(n26469) );
  XOR2HSV0 U28374 ( .A1(n26470), .A2(n26469), .Z(n26471) );
  XOR2HSV0 U28375 ( .A1(n26472), .A2(n26471), .Z(n26473) );
  XNOR2HSV1 U28376 ( .A1(n26474), .A2(n26473), .ZN(n26475) );
  XNOR2HSV1 U28377 ( .A1(n26476), .A2(n26475), .ZN(n26478) );
  NAND2HSV0 U28378 ( .A1(\pe1/got [15]), .A2(n26909), .ZN(n26477) );
  XOR2HSV0 U28379 ( .A1(n26478), .A2(n26477), .Z(n26479) );
  XOR2HSV0 U28380 ( .A1(n26480), .A2(n26479), .Z(po1) );
  NAND2HSV0 U28381 ( .A1(n27000), .A2(n26595), .ZN(n26535) );
  NAND2HSV0 U28382 ( .A1(n27136), .A2(n28425), .ZN(n26531) );
  NAND2HSV0 U28383 ( .A1(n27137), .A2(\pe1/got [11]), .ZN(n26529) );
  NOR2HSV2 U28384 ( .A1(n26888), .A2(n26539), .ZN(n26527) );
  CLKNHSV0 U28385 ( .I(\pe1/got [9]), .ZN(n27001) );
  NOR2HSV2 U28386 ( .A1(n27004), .A2(n27001), .ZN(n26525) );
  NAND2HSV0 U28387 ( .A1(n26854), .A2(\pe1/got [8]), .ZN(n26523) );
  NAND2HSV0 U28388 ( .A1(n26541), .A2(\pe1/got [6]), .ZN(n26519) );
  NAND2HSV0 U28389 ( .A1(n27005), .A2(\pe1/got [2]), .ZN(n26512) );
  NAND2HSV0 U28390 ( .A1(n26562), .A2(\pe1/got [1]), .ZN(n26510) );
  NAND2HSV0 U28391 ( .A1(\pe1/aot [14]), .A2(\pe1/bq[1] ), .ZN(n26484) );
  NAND2HSV0 U28392 ( .A1(\pe1/bq[2] ), .A2(\pe1/aot [13]), .ZN(n26483) );
  XOR2HSV0 U28393 ( .A1(n26484), .A2(n26483), .Z(n26489) );
  NAND2HSV0 U28394 ( .A1(\pe1/aot [6]), .A2(\pe1/bq[6] ), .ZN(n27147) );
  OAI21HSV0 U28395 ( .A1(n26763), .A2(n27158), .B(n26485), .ZN(n26486) );
  OAI21HSV0 U28396 ( .A1(n26487), .A2(n27147), .B(n26486), .ZN(n26488) );
  XNOR2HSV1 U28397 ( .A1(n26489), .A2(n26488), .ZN(n26493) );
  NAND2HSV0 U28398 ( .A1(\pe1/aot [7]), .A2(\pe1/bq[8] ), .ZN(n26491) );
  NAND2HSV0 U28399 ( .A1(\pe1/aot [2]), .A2(\pe1/bq[13] ), .ZN(n26490) );
  XOR2HSV0 U28400 ( .A1(n26491), .A2(n26490), .Z(n26492) );
  XNOR2HSV1 U28401 ( .A1(n26493), .A2(n26492), .ZN(n26509) );
  NAND2HSV0 U28402 ( .A1(\pe1/aot [8]), .A2(\pe1/bq[7] ), .ZN(n26495) );
  NAND2HSV0 U28403 ( .A1(\pe1/aot [11]), .A2(\pe1/bq[4] ), .ZN(n26494) );
  XOR2HSV0 U28404 ( .A1(n26495), .A2(n26494), .Z(n26499) );
  NAND2HSV0 U28405 ( .A1(\pe1/aot [12]), .A2(\pe1/bq[3] ), .ZN(n26497) );
  NAND2HSV0 U28406 ( .A1(\pe1/aot [10]), .A2(\pe1/bq[5] ), .ZN(n26496) );
  XOR2HSV0 U28407 ( .A1(n26497), .A2(n26496), .Z(n26498) );
  XOR2HSV0 U28408 ( .A1(n26499), .A2(n26498), .Z(n26507) );
  NAND2HSV0 U28409 ( .A1(\pe1/aot [1]), .A2(\pe1/bq[14] ), .ZN(n26501) );
  NAND2HSV0 U28410 ( .A1(\pe1/aot [4]), .A2(\pe1/bq[11] ), .ZN(n26500) );
  XOR2HSV0 U28411 ( .A1(n26501), .A2(n26500), .Z(n26505) );
  NAND2HSV0 U28412 ( .A1(\pe1/aot [3]), .A2(\pe1/bq[12] ), .ZN(n26503) );
  NAND2HSV0 U28413 ( .A1(\pe1/aot [5]), .A2(\pe1/bq[10] ), .ZN(n26502) );
  XOR2HSV0 U28414 ( .A1(n26503), .A2(n26502), .Z(n26504) );
  XOR2HSV0 U28415 ( .A1(n26505), .A2(n26504), .Z(n26506) );
  XOR2HSV0 U28416 ( .A1(n26507), .A2(n26506), .Z(n26508) );
  XOR3HSV2 U28417 ( .A1(n26510), .A2(n26509), .A3(n26508), .Z(n26511) );
  XNOR2HSV1 U28418 ( .A1(n26512), .A2(n26511), .ZN(n26514) );
  NAND2HSV0 U28419 ( .A1(n28635), .A2(\pe1/got [3]), .ZN(n26513) );
  XNOR2HSV1 U28420 ( .A1(n26514), .A2(n26513), .ZN(n26517) );
  NAND2HSV0 U28421 ( .A1(n28649), .A2(\pe1/got [4]), .ZN(n26516) );
  NAND2HSV0 U28422 ( .A1(n27166), .A2(\pe1/got [5]), .ZN(n26515) );
  XOR3HSV2 U28423 ( .A1(n26517), .A2(n26516), .A3(n26515), .Z(n26518) );
  XNOR2HSV1 U28424 ( .A1(n26519), .A2(n26518), .ZN(n26521) );
  NAND2HSV0 U28425 ( .A1(n28589), .A2(\pe1/got [7]), .ZN(n26520) );
  XNOR2HSV1 U28426 ( .A1(n26521), .A2(n26520), .ZN(n26522) );
  XNOR2HSV1 U28427 ( .A1(n26523), .A2(n26522), .ZN(n26524) );
  XOR2HSV0 U28428 ( .A1(n26525), .A2(n26524), .Z(n26526) );
  XOR2HSV0 U28429 ( .A1(n26527), .A2(n26526), .Z(n26528) );
  XNOR2HSV1 U28430 ( .A1(n26529), .A2(n26528), .ZN(n26530) );
  XNOR2HSV1 U28431 ( .A1(n26531), .A2(n26530), .ZN(n26533) );
  NAND2HSV0 U28432 ( .A1(n26909), .A2(\pe1/got [13]), .ZN(n26532) );
  XOR2HSV0 U28433 ( .A1(n26533), .A2(n26532), .Z(n26534) );
  XOR2HSV0 U28434 ( .A1(n26535), .A2(n26534), .Z(\pe1/poht [2]) );
  NAND2HSV0 U28435 ( .A1(n27000), .A2(n17230), .ZN(n26599) );
  NAND2HSV0 U28436 ( .A1(n27136), .A2(\pe1/got [13]), .ZN(n26594) );
  NAND2HSV0 U28437 ( .A1(n28425), .A2(n26537), .ZN(n26592) );
  NOR2HSV2 U28438 ( .A1(n26888), .A2(n26538), .ZN(n26590) );
  NOR2HSV0 U28439 ( .A1(n26540), .A2(n26539), .ZN(n26588) );
  NAND2HSV0 U28440 ( .A1(n26854), .A2(\pe1/got [9]), .ZN(n26586) );
  NAND2HSV0 U28441 ( .A1(\pe1/got [7]), .A2(n26541), .ZN(n26582) );
  NAND2HSV0 U28442 ( .A1(n28481), .A2(\pe1/got [3]), .ZN(n26575) );
  NAND2HSV0 U28443 ( .A1(n28622), .A2(\pe1/got [1]), .ZN(n26545) );
  NAND2HSV0 U28444 ( .A1(\pe1/bq[1] ), .A2(\pe1/aot [11]), .ZN(n27150) );
  NAND2HSV0 U28445 ( .A1(\pe1/aot [6]), .A2(\pe1/bq[10] ), .ZN(n26770) );
  XNOR2HSV1 U28446 ( .A1(n26543), .A2(n26770), .ZN(n26544) );
  XNOR2HSV1 U28447 ( .A1(n26545), .A2(n26544), .ZN(n26573) );
  NAND2HSV0 U28448 ( .A1(\pe1/aot [8]), .A2(\pe1/bq[8] ), .ZN(n26547) );
  NAND2HSV0 U28449 ( .A1(\pe1/aot [3]), .A2(\pe1/bq[13] ), .ZN(n26546) );
  XOR2HSV0 U28450 ( .A1(n26547), .A2(n26546), .Z(n26552) );
  NAND2HSV0 U28451 ( .A1(\pe1/aot [1]), .A2(n26548), .ZN(n26550) );
  NAND2HSV0 U28452 ( .A1(\pe1/aot [2]), .A2(\pe1/bq[14] ), .ZN(n26549) );
  XOR2HSV0 U28453 ( .A1(n26550), .A2(n26549), .Z(n26551) );
  XNOR2HSV1 U28454 ( .A1(n26552), .A2(n26551), .ZN(n26561) );
  NAND2HSV0 U28455 ( .A1(\pe1/bq[6] ), .A2(\pe1/aot [10]), .ZN(n26554) );
  NAND2HSV0 U28456 ( .A1(\pe1/aot [7]), .A2(\pe1/bq[9] ), .ZN(n26553) );
  XOR2HSV0 U28457 ( .A1(n26554), .A2(n26553), .Z(n26559) );
  NOR2HSV0 U28458 ( .A1(n26555), .A2(n26652), .ZN(n27022) );
  XNOR2HSV1 U28459 ( .A1(n26559), .A2(n26558), .ZN(n26560) );
  XNOR2HSV1 U28460 ( .A1(n26561), .A2(n26560), .ZN(n26572) );
  NAND2HSV0 U28461 ( .A1(n26562), .A2(\pe1/got [2]), .ZN(n26570) );
  NAND2HSV0 U28462 ( .A1(\pe1/aot [13]), .A2(\pe1/bq[3] ), .ZN(n26564) );
  NAND2HSV0 U28463 ( .A1(\pe1/aot [9]), .A2(\pe1/bq[7] ), .ZN(n26563) );
  XOR2HSV0 U28464 ( .A1(n26564), .A2(n26563), .Z(n26568) );
  NAND2HSV0 U28465 ( .A1(\pe1/aot [4]), .A2(\pe1/bq[12] ), .ZN(n26566) );
  NAND2HSV0 U28466 ( .A1(\pe1/aot [5]), .A2(\pe1/bq[11] ), .ZN(n26565) );
  XOR2HSV0 U28467 ( .A1(n26566), .A2(n26565), .Z(n26567) );
  XOR2HSV0 U28468 ( .A1(n26568), .A2(n26567), .Z(n26569) );
  XOR2HSV0 U28469 ( .A1(n26570), .A2(n26569), .Z(n26571) );
  XOR3HSV2 U28470 ( .A1(n26573), .A2(n26572), .A3(n26571), .Z(n26574) );
  XNOR2HSV1 U28471 ( .A1(n26575), .A2(n26574), .ZN(n26577) );
  NAND2HSV0 U28472 ( .A1(n28635), .A2(\pe1/got [4]), .ZN(n26576) );
  XNOR2HSV1 U28473 ( .A1(n26577), .A2(n26576), .ZN(n26580) );
  NAND2HSV0 U28474 ( .A1(n28649), .A2(\pe1/got [5]), .ZN(n26579) );
  NAND2HSV0 U28475 ( .A1(n27166), .A2(n28434), .ZN(n26578) );
  XOR3HSV2 U28476 ( .A1(n26580), .A2(n26579), .A3(n26578), .Z(n26581) );
  XNOR2HSV1 U28477 ( .A1(n26582), .A2(n26581), .ZN(n26584) );
  NAND2HSV0 U28478 ( .A1(n28589), .A2(\pe1/got [8]), .ZN(n26583) );
  XNOR2HSV1 U28479 ( .A1(n26584), .A2(n26583), .ZN(n26585) );
  XNOR2HSV1 U28480 ( .A1(n26586), .A2(n26585), .ZN(n26587) );
  XOR2HSV0 U28481 ( .A1(n26588), .A2(n26587), .Z(n26589) );
  XOR2HSV0 U28482 ( .A1(n26590), .A2(n26589), .Z(n26591) );
  XNOR2HSV1 U28483 ( .A1(n26592), .A2(n26591), .ZN(n26593) );
  XNOR2HSV1 U28484 ( .A1(n26594), .A2(n26593), .ZN(n26597) );
  CLKNAND2HSV0 U28485 ( .A1(n27185), .A2(\pe1/got [14]), .ZN(n26596) );
  XOR2HSV0 U28486 ( .A1(n26597), .A2(n26596), .Z(n26598) );
  XOR2HSV0 U28487 ( .A1(n26599), .A2(n26598), .Z(\pe1/poht [1]) );
  NAND2HSV0 U28488 ( .A1(n26600), .A2(\pe3/got [11]), .ZN(n26649) );
  NAND2HSV0 U28489 ( .A1(n28438), .A2(n26603), .ZN(n26633) );
  NAND2HSV0 U28490 ( .A1(n23327), .A2(\pe3/got [4]), .ZN(n26631) );
  NAND2HSV0 U28491 ( .A1(n28588), .A2(n26751), .ZN(n26629) );
  NAND2HSV0 U28492 ( .A1(n26682), .A2(\pe3/got [2]), .ZN(n26623) );
  NAND2HSV0 U28493 ( .A1(\pe3/aot [8]), .A2(\pe3/bq[4] ), .ZN(n26606) );
  XOR2HSV0 U28494 ( .A1(n26607), .A2(n26606), .Z(n26621) );
  NAND2HSV0 U28495 ( .A1(\pe3/aot [11]), .A2(\pe3/bq[1] ), .ZN(n26609) );
  NAND2HSV0 U28496 ( .A1(\pe3/aot [9]), .A2(\pe3/bq[3] ), .ZN(n26608) );
  XOR2HSV0 U28497 ( .A1(n26609), .A2(n26608), .Z(n26612) );
  NAND2HSV0 U28498 ( .A1(\pe3/aot [5]), .A2(\pe3/bq[8] ), .ZN(n26700) );
  XNOR2HSV1 U28499 ( .A1(n26612), .A2(n26611), .ZN(n26620) );
  NAND2HSV0 U28500 ( .A1(\pe3/aot [1]), .A2(\pe3/bq[11] ), .ZN(n26614) );
  NAND2HSV0 U28501 ( .A1(\pe3/aot [3]), .A2(\pe3/bq[9] ), .ZN(n26613) );
  XOR2HSV0 U28502 ( .A1(n26614), .A2(n26613), .Z(n26618) );
  NAND2HSV0 U28503 ( .A1(\pe3/aot [10]), .A2(\pe3/bq[2] ), .ZN(n26616) );
  NAND2HSV0 U28504 ( .A1(\pe3/aot [6]), .A2(\pe3/bq[6] ), .ZN(n26615) );
  XOR2HSV0 U28505 ( .A1(n26616), .A2(n26615), .Z(n26617) );
  XOR2HSV0 U28506 ( .A1(n26618), .A2(n26617), .Z(n26619) );
  XOR3HSV2 U28507 ( .A1(n26621), .A2(n26620), .A3(n26619), .Z(n26622) );
  XNOR2HSV1 U28508 ( .A1(n26623), .A2(n26622), .ZN(n26627) );
  NOR2HSV0 U28509 ( .A1(n26625), .A2(n26624), .ZN(n26626) );
  XNOR2HSV1 U28510 ( .A1(n26627), .A2(n26626), .ZN(n26628) );
  XNOR2HSV1 U28511 ( .A1(n26629), .A2(n26628), .ZN(n26630) );
  XNOR2HSV1 U28512 ( .A1(n26631), .A2(n26630), .ZN(n26632) );
  XOR2HSV0 U28513 ( .A1(n26633), .A2(n26632), .Z(n26636) );
  NAND2HSV0 U28514 ( .A1(n26634), .A2(\pe3/got [6]), .ZN(n26635) );
  XOR2HSV0 U28515 ( .A1(n26636), .A2(n26635), .Z(n26639) );
  NAND2HSV0 U28516 ( .A1(n26637), .A2(\pe3/got [7]), .ZN(n26638) );
  XOR2HSV0 U28517 ( .A1(n26639), .A2(n26638), .Z(n26640) );
  NAND2HSV0 U28518 ( .A1(n26759), .A2(n26642), .ZN(n26643) );
  INAND2HSV2 U28519 ( .A1(n26645), .B1(n26729), .ZN(n26646) );
  XNOR2HSV1 U28520 ( .A1(n26647), .A2(n26646), .ZN(n26648) );
  XOR2HSV0 U28521 ( .A1(n26649), .A2(n26648), .Z(\pe3/poht [5]) );
  NAND2HSV0 U28522 ( .A1(n28700), .A2(\pe1/got [5]), .ZN(n26674) );
  NAND2HSV0 U28523 ( .A1(n28460), .A2(n28435), .ZN(n26672) );
  CLKNHSV0 U28524 ( .I(\pe1/got [3]), .ZN(n26853) );
  NOR2HSV2 U28525 ( .A1(n27002), .A2(n26853), .ZN(n26670) );
  CLKNHSV1 U28526 ( .I(\pe1/got [2]), .ZN(n26829) );
  NOR2HSV2 U28527 ( .A1(n26830), .A2(n26829), .ZN(n26668) );
  NAND2HSV0 U28528 ( .A1(n26854), .A2(\pe1/got [1]), .ZN(n26666) );
  NAND2HSV0 U28529 ( .A1(\pe1/aot [5]), .A2(\pe1/bq[3] ), .ZN(n26651) );
  NAND2HSV0 U28530 ( .A1(\pe1/aot [1]), .A2(\pe1/bq[7] ), .ZN(n26650) );
  XOR2HSV0 U28531 ( .A1(n26651), .A2(n26650), .Z(n26657) );
  NOR2HSV0 U28532 ( .A1(n26653), .A2(n26652), .ZN(n26655) );
  NAND2HSV0 U28533 ( .A1(\pe1/aot [4]), .A2(\pe1/bq[4] ), .ZN(n26654) );
  XOR2HSV0 U28534 ( .A1(n26655), .A2(n26654), .Z(n26656) );
  XNOR2HSV1 U28535 ( .A1(n26657), .A2(n26656), .ZN(n26664) );
  NAND2HSV0 U28536 ( .A1(\pe1/aot [7]), .A2(\pe1/bq[1] ), .ZN(n26864) );
  NAND2HSV0 U28537 ( .A1(\pe1/aot [3]), .A2(\pe1/bq[5] ), .ZN(n26660) );
  CLKNHSV0 U28538 ( .I(\pe1/aot [3]), .ZN(n26658) );
  NOR2HSV2 U28539 ( .A1(n26658), .A2(n27064), .ZN(n26821) );
  NOR2HSV0 U28540 ( .A1(n26764), .A2(n26659), .ZN(n27146) );
  AOI22HSV0 U28541 ( .A1(n26864), .A2(n26660), .B1(n26821), .B2(n27146), .ZN(
        n26662) );
  NAND2HSV0 U28542 ( .A1(\pe1/aot [2]), .A2(\pe1/bq[6] ), .ZN(n26661) );
  XOR2HSV0 U28543 ( .A1(n26662), .A2(n26661), .Z(n26663) );
  XNOR2HSV1 U28544 ( .A1(n26664), .A2(n26663), .ZN(n26665) );
  XNOR2HSV1 U28545 ( .A1(n26666), .A2(n26665), .ZN(n26667) );
  XOR2HSV0 U28546 ( .A1(n26668), .A2(n26667), .Z(n26669) );
  XOR2HSV0 U28547 ( .A1(n26670), .A2(n26669), .Z(n26671) );
  XNOR2HSV1 U28548 ( .A1(n26672), .A2(n26671), .ZN(n26673) );
  XNOR2HSV1 U28549 ( .A1(n26674), .A2(n26673), .ZN(n26676) );
  CLKNAND2HSV1 U28550 ( .A1(n26909), .A2(\pe1/got [6]), .ZN(n26675) );
  XOR2HSV0 U28551 ( .A1(n26676), .A2(n26675), .Z(n26677) );
  XOR2HSV0 U28552 ( .A1(n26678), .A2(n26677), .Z(\pe1/poht [9]) );
  NOR2HSV2 U28553 ( .A1(n26681), .A2(n26680), .ZN(n26728) );
  NAND2HSV0 U28554 ( .A1(n28438), .A2(\pe3/got [6]), .ZN(n26722) );
  NAND2HSV0 U28555 ( .A1(n23327), .A2(\pe3/got [5]), .ZN(n26720) );
  NAND2HSV0 U28556 ( .A1(n28588), .A2(\pe3/got [4]), .ZN(n26718) );
  NAND2HSV0 U28557 ( .A1(n26682), .A2(n26751), .ZN(n26712) );
  NAND2HSV0 U28558 ( .A1(n15240), .A2(\pe3/got [1]), .ZN(n26710) );
  NOR2HSV0 U28559 ( .A1(n26684), .A2(n26683), .ZN(n26686) );
  AOI22HSV0 U28560 ( .A1(\pe3/aot [11]), .A2(\pe3/bq[2] ), .B1(\pe3/bq[9] ), 
        .B2(\pe3/aot [4]), .ZN(n26685) );
  NOR2HSV2 U28561 ( .A1(n26686), .A2(n26685), .ZN(n26692) );
  NOR2HSV0 U28562 ( .A1(n26688), .A2(n26687), .ZN(n26690) );
  AOI22HSV0 U28563 ( .A1(\pe3/aot [7]), .A2(\pe3/bq[6] ), .B1(\pe3/bq[11] ), 
        .B2(\pe3/aot [2]), .ZN(n26689) );
  NOR2HSV1 U28564 ( .A1(n26690), .A2(n26689), .ZN(n26691) );
  XOR2HSV0 U28565 ( .A1(n26692), .A2(n26691), .Z(n26708) );
  NAND2HSV0 U28566 ( .A1(\pe3/aot [12]), .A2(\pe3/bq[1] ), .ZN(n26694) );
  NAND2HSV0 U28567 ( .A1(\pe3/aot [10]), .A2(\pe3/bq[3] ), .ZN(n26693) );
  XOR2HSV0 U28568 ( .A1(n26694), .A2(n26693), .Z(n26698) );
  NAND2HSV0 U28569 ( .A1(\pe3/aot [3]), .A2(\pe3/bq[10] ), .ZN(n26696) );
  NAND2HSV0 U28570 ( .A1(\pe3/aot [8]), .A2(\pe3/bq[5] ), .ZN(n26695) );
  XOR2HSV0 U28571 ( .A1(n26696), .A2(n26695), .Z(n26697) );
  XNOR2HSV1 U28572 ( .A1(n26698), .A2(n26697), .ZN(n26707) );
  NAND2HSV0 U28573 ( .A1(\pe3/aot [1]), .A2(\pe3/bq[12] ), .ZN(n26699) );
  XOR2HSV0 U28574 ( .A1(n26700), .A2(n26699), .Z(n26705) );
  NOR2HSV0 U28575 ( .A1(n26701), .A2(n23349), .ZN(n26703) );
  NAND2HSV0 U28576 ( .A1(\pe3/aot [6]), .A2(\pe3/bq[7] ), .ZN(n26702) );
  XOR2HSV0 U28577 ( .A1(n26703), .A2(n26702), .Z(n26704) );
  XOR2HSV0 U28578 ( .A1(n26705), .A2(n26704), .Z(n26706) );
  XOR3HSV2 U28579 ( .A1(n26708), .A2(n26707), .A3(n26706), .Z(n26709) );
  XNOR2HSV1 U28580 ( .A1(n26710), .A2(n26709), .ZN(n26711) );
  XNOR2HSV1 U28581 ( .A1(n26712), .A2(n26711), .ZN(n26716) );
  NOR2HSV0 U28582 ( .A1(n26714), .A2(n26713), .ZN(n26715) );
  XNOR2HSV1 U28583 ( .A1(n26716), .A2(n26715), .ZN(n26717) );
  XNOR2HSV1 U28584 ( .A1(n26718), .A2(n26717), .ZN(n26719) );
  XNOR2HSV1 U28585 ( .A1(n26720), .A2(n26719), .ZN(n26721) );
  XOR2HSV0 U28586 ( .A1(n26722), .A2(n26721), .Z(n26724) );
  NAND2HSV0 U28587 ( .A1(n26752), .A2(\pe3/got [7]), .ZN(n26723) );
  XOR2HSV0 U28588 ( .A1(n26724), .A2(n26723), .Z(n26726) );
  NAND2HSV0 U28589 ( .A1(n28584), .A2(n28648), .ZN(n26725) );
  XOR2HSV0 U28590 ( .A1(n26726), .A2(n26725), .Z(n26727) );
  NOR2HSV2 U28591 ( .A1(n26730), .A2(n23329), .ZN(n26758) );
  NAND2HSV0 U28592 ( .A1(n28438), .A2(\pe3/got [2]), .ZN(n26750) );
  NAND2HSV0 U28593 ( .A1(n23327), .A2(\pe3/got [1]), .ZN(n26748) );
  NAND2HSV0 U28594 ( .A1(\pe3/aot [7]), .A2(\pe3/bq[2] ), .ZN(n26732) );
  NAND2HSV0 U28595 ( .A1(\pe3/aot [2]), .A2(\pe3/bq[7] ), .ZN(n26731) );
  XOR2HSV0 U28596 ( .A1(n26732), .A2(n26731), .Z(n26736) );
  NAND2HSV0 U28597 ( .A1(\pe3/aot [3]), .A2(\pe3/bq[6] ), .ZN(n26734) );
  NAND2HSV0 U28598 ( .A1(\pe3/aot [6]), .A2(\pe3/bq[3] ), .ZN(n26733) );
  XOR2HSV0 U28599 ( .A1(n26734), .A2(n26733), .Z(n26735) );
  XOR2HSV0 U28600 ( .A1(n26736), .A2(n26735), .Z(n26746) );
  NAND2HSV0 U28601 ( .A1(\pe3/aot [4]), .A2(\pe3/bq[5] ), .ZN(n26738) );
  NAND2HSV0 U28602 ( .A1(\pe3/aot [5]), .A2(\pe3/bq[4] ), .ZN(n26737) );
  XOR2HSV0 U28603 ( .A1(n26738), .A2(n26737), .Z(n26744) );
  NOR2HSV0 U28604 ( .A1(n26740), .A2(n26739), .ZN(n26742) );
  AOI22HSV0 U28605 ( .A1(\pe3/aot [8]), .A2(\pe3/bq[1] ), .B1(\pe3/bq[8] ), 
        .B2(\pe3/aot [1]), .ZN(n26741) );
  NOR2HSV2 U28606 ( .A1(n26742), .A2(n26741), .ZN(n26743) );
  XNOR2HSV1 U28607 ( .A1(n26744), .A2(n26743), .ZN(n26745) );
  XNOR2HSV1 U28608 ( .A1(n26746), .A2(n26745), .ZN(n26747) );
  XNOR2HSV1 U28609 ( .A1(n26748), .A2(n26747), .ZN(n26749) );
  XOR2HSV0 U28610 ( .A1(n26750), .A2(n26749), .Z(n26754) );
  NAND2HSV0 U28611 ( .A1(n26634), .A2(n26751), .ZN(n26753) );
  XOR2HSV0 U28612 ( .A1(n26754), .A2(n26753), .Z(n26756) );
  NAND2HSV0 U28613 ( .A1(\pe3/got [4]), .A2(n28584), .ZN(n26755) );
  NAND2HSV0 U28614 ( .A1(n27000), .A2(\pe1/got [12]), .ZN(n26804) );
  CLKNAND2HSV0 U28615 ( .A1(n27184), .A2(n28700), .ZN(n26800) );
  NAND2HSV0 U28616 ( .A1(n28460), .A2(\pe1/got [9]), .ZN(n26798) );
  CLKNHSV0 U28617 ( .I(\pe1/got [8]), .ZN(n27003) );
  NOR2HSV2 U28618 ( .A1(n26888), .A2(n27003), .ZN(n26796) );
  CLKNHSV0 U28619 ( .I(\pe1/got [7]), .ZN(n27138) );
  NOR2HSV2 U28620 ( .A1(n27004), .A2(n27138), .ZN(n26794) );
  NAND2HSV0 U28621 ( .A1(n26854), .A2(\pe1/got [6]), .ZN(n26792) );
  NAND2HSV0 U28622 ( .A1(n28609), .A2(n28435), .ZN(n26788) );
  NAND2HSV0 U28623 ( .A1(n28635), .A2(\pe1/got [1]), .ZN(n26783) );
  NAND2HSV0 U28624 ( .A1(\pe1/aot [1]), .A2(\pe1/bq[12] ), .ZN(n26762) );
  NAND2HSV0 U28625 ( .A1(\pe1/aot [12]), .A2(\pe1/bq[1] ), .ZN(n26761) );
  XOR2HSV0 U28626 ( .A1(n26762), .A2(n26761), .Z(n26766) );
  XOR2HSV0 U28627 ( .A1(n26766), .A2(n26765), .Z(n26774) );
  NAND2HSV0 U28628 ( .A1(\pe1/aot [4]), .A2(\pe1/bq[9] ), .ZN(n26768) );
  NAND2HSV0 U28629 ( .A1(\pe1/aot [5]), .A2(\pe1/bq[8] ), .ZN(n26767) );
  XOR2HSV0 U28630 ( .A1(n26768), .A2(n26767), .Z(n26772) );
  XNOR2HSV1 U28631 ( .A1(n26772), .A2(n26771), .ZN(n26773) );
  XNOR2HSV1 U28632 ( .A1(n26774), .A2(n26773), .ZN(n26781) );
  NAND2HSV0 U28633 ( .A1(\pe1/aot [10]), .A2(\pe1/bq[3] ), .ZN(n26776) );
  NAND2HSV0 U28634 ( .A1(\pe1/aot [2]), .A2(\pe1/bq[11] ), .ZN(n26775) );
  XOR2HSV0 U28635 ( .A1(n26776), .A2(n26775), .Z(n26779) );
  NAND2HSV0 U28636 ( .A1(\pe1/aot [8]), .A2(\pe1/bq[5] ), .ZN(n27144) );
  NAND2HSV0 U28637 ( .A1(\pe1/aot [9]), .A2(\pe1/bq[4] ), .ZN(n26777) );
  XOR2HSV0 U28638 ( .A1(n27144), .A2(n26777), .Z(n26778) );
  XOR2HSV0 U28639 ( .A1(n26779), .A2(n26778), .Z(n26780) );
  XNOR2HSV1 U28640 ( .A1(n26781), .A2(n26780), .ZN(n26782) );
  XNOR2HSV1 U28641 ( .A1(n26783), .A2(n26782), .ZN(n26786) );
  NAND2HSV0 U28642 ( .A1(n28649), .A2(\pe1/got [2]), .ZN(n26785) );
  NAND2HSV0 U28643 ( .A1(n27166), .A2(\pe1/got [3]), .ZN(n26784) );
  XOR3HSV2 U28644 ( .A1(n26786), .A2(n26785), .A3(n26784), .Z(n26787) );
  XNOR2HSV1 U28645 ( .A1(n26788), .A2(n26787), .ZN(n26790) );
  NAND2HSV0 U28646 ( .A1(n28589), .A2(\pe1/got [5]), .ZN(n26789) );
  XNOR2HSV1 U28647 ( .A1(n26790), .A2(n26789), .ZN(n26791) );
  XNOR2HSV1 U28648 ( .A1(n26792), .A2(n26791), .ZN(n26793) );
  XOR2HSV0 U28649 ( .A1(n26794), .A2(n26793), .Z(n26795) );
  XOR2HSV0 U28650 ( .A1(n26796), .A2(n26795), .Z(n26797) );
  XNOR2HSV1 U28651 ( .A1(n26798), .A2(n26797), .ZN(n26799) );
  XNOR2HSV1 U28652 ( .A1(n26800), .A2(n26799), .ZN(n26802) );
  NAND2HSV0 U28653 ( .A1(n27185), .A2(\pe1/got [11]), .ZN(n26801) );
  XOR2HSV0 U28654 ( .A1(n26802), .A2(n26801), .Z(n26803) );
  XOR2HSV0 U28655 ( .A1(n26804), .A2(n26803), .Z(\pe1/poht [4]) );
  NAND2HSV0 U28656 ( .A1(n27000), .A2(\pe1/got [1]), .ZN(n26806) );
  XOR2HSV0 U28657 ( .A1(n26806), .A2(n26805), .Z(\pe1/poht [15]) );
  CLKNAND2HSV0 U28658 ( .A1(\pe1/got [4]), .A2(n27000), .ZN(n26818) );
  NAND2HSV0 U28659 ( .A1(n27136), .A2(\pe1/got [2]), .ZN(n26814) );
  NAND2HSV0 U28660 ( .A1(n28460), .A2(\pe1/got [1]), .ZN(n26813) );
  NAND2HSV0 U28661 ( .A1(\pe1/aot [4]), .A2(\pe1/bq[1] ), .ZN(n26808) );
  NAND2HSV0 U28662 ( .A1(\pe1/aot [1]), .A2(\pe1/bq[4] ), .ZN(n26807) );
  XOR2HSV0 U28663 ( .A1(n26808), .A2(n26807), .Z(n26811) );
  CLKNAND2HSV0 U28664 ( .A1(\pe1/bq[2] ), .A2(\pe1/aot [3]), .ZN(n26889) );
  NAND2HSV0 U28665 ( .A1(\pe1/aot [2]), .A2(\pe1/bq[3] ), .ZN(n26809) );
  XOR2HSV0 U28666 ( .A1(n26889), .A2(n26809), .Z(n26810) );
  XOR2HSV0 U28667 ( .A1(n26811), .A2(n26810), .Z(n26812) );
  NAND2HSV0 U28668 ( .A1(n26909), .A2(\pe1/got [3]), .ZN(n26815) );
  XOR2HSV0 U28669 ( .A1(n26816), .A2(n26815), .Z(n26817) );
  XOR2HSV0 U28670 ( .A1(n26818), .A2(n26817), .Z(\pe1/poht [12]) );
  NAND2HSV0 U28671 ( .A1(\pe1/aot [1]), .A2(\pe1/bq[3] ), .ZN(n26820) );
  NAND2HSV0 U28672 ( .A1(\pe1/aot [2]), .A2(\pe1/bq[2] ), .ZN(n26819) );
  CLKNHSV0 U28673 ( .I(n26822), .ZN(n26823) );
  CLKNAND2HSV0 U28674 ( .A1(n26824), .A2(n26823), .ZN(n26826) );
  NOR2HSV1 U28675 ( .A1(n26826), .A2(n26825), .ZN(n26828) );
  CLKNAND2HSV0 U28676 ( .A1(n28700), .A2(\pe1/got [4]), .ZN(n26847) );
  NAND2HSV0 U28677 ( .A1(n28460), .A2(\pe1/got [3]), .ZN(n26845) );
  NOR2HSV2 U28678 ( .A1(n27139), .A2(n26829), .ZN(n26843) );
  CLKNHSV0 U28679 ( .I(\pe1/got [1]), .ZN(n26887) );
  NOR2HSV2 U28680 ( .A1(n26830), .A2(n26887), .ZN(n26841) );
  NAND2HSV0 U28681 ( .A1(\pe1/aot [3]), .A2(\pe1/bq[4] ), .ZN(n26832) );
  NAND2HSV0 U28682 ( .A1(\pe1/aot [2]), .A2(\pe1/bq[5] ), .ZN(n26831) );
  XOR2HSV0 U28683 ( .A1(n26832), .A2(n26831), .Z(n26836) );
  NAND2HSV0 U28684 ( .A1(\pe1/aot [1]), .A2(\pe1/bq[6] ), .ZN(n26834) );
  NAND2HSV0 U28685 ( .A1(\pe1/aot [5]), .A2(\pe1/bq[2] ), .ZN(n26833) );
  XOR2HSV0 U28686 ( .A1(n26834), .A2(n26833), .Z(n26835) );
  XNOR2HSV1 U28687 ( .A1(n26836), .A2(n26835), .ZN(n26839) );
  CLKNAND2HSV0 U28688 ( .A1(\pe1/aot [4]), .A2(\pe1/bq[3] ), .ZN(n26890) );
  NAND2HSV0 U28689 ( .A1(\pe1/aot [6]), .A2(\pe1/bq[1] ), .ZN(n26837) );
  XOR2HSV0 U28690 ( .A1(n26890), .A2(n26837), .Z(n26838) );
  XNOR2HSV1 U28691 ( .A1(n26839), .A2(n26838), .ZN(n26840) );
  XOR2HSV0 U28692 ( .A1(n26841), .A2(n26840), .Z(n26842) );
  XOR2HSV0 U28693 ( .A1(n26843), .A2(n26842), .Z(n26844) );
  XNOR2HSV1 U28694 ( .A1(n26845), .A2(n26844), .ZN(n26846) );
  XNOR2HSV1 U28695 ( .A1(n26847), .A2(n26846), .ZN(n26849) );
  XOR2HSV0 U28696 ( .A1(n26849), .A2(n26848), .Z(n26850) );
  XOR2HSV0 U28697 ( .A1(n26851), .A2(n26850), .Z(\pe1/poht [10]) );
  CLKNAND2HSV0 U28698 ( .A1(n28700), .A2(\pe1/got [6]), .ZN(n26882) );
  NAND2HSV0 U28699 ( .A1(n27137), .A2(\pe1/got [5]), .ZN(n26880) );
  NOR2HSV2 U28700 ( .A1(n27002), .A2(n26852), .ZN(n26878) );
  NOR2HSV2 U28701 ( .A1(n27004), .A2(n26853), .ZN(n26876) );
  CLKNAND2HSV0 U28702 ( .A1(n26854), .A2(\pe1/got [2]), .ZN(n26874) );
  NAND2HSV0 U28703 ( .A1(n28589), .A2(\pe1/got [1]), .ZN(n26872) );
  NAND2HSV0 U28704 ( .A1(\pe1/aot [5]), .A2(\pe1/bq[4] ), .ZN(n26856) );
  NAND2HSV0 U28705 ( .A1(\pe1/aot [6]), .A2(\pe1/bq[3] ), .ZN(n26855) );
  XOR2HSV0 U28706 ( .A1(n26856), .A2(n26855), .Z(n26860) );
  NAND2HSV0 U28707 ( .A1(\pe1/aot [3]), .A2(\pe1/bq[6] ), .ZN(n26857) );
  XOR2HSV0 U28708 ( .A1(n26858), .A2(n26857), .Z(n26859) );
  XOR2HSV0 U28709 ( .A1(n26860), .A2(n26859), .Z(n26870) );
  NAND2HSV0 U28710 ( .A1(\pe1/aot [1]), .A2(\pe1/bq[8] ), .ZN(n26862) );
  NAND2HSV0 U28711 ( .A1(\pe1/aot [2]), .A2(\pe1/bq[7] ), .ZN(n26861) );
  XOR2HSV0 U28712 ( .A1(n26862), .A2(n26861), .Z(n26868) );
  NOR2HSV0 U28713 ( .A1(n26864), .A2(n26863), .ZN(n26866) );
  AOI22HSV0 U28714 ( .A1(\pe1/aot [8]), .A2(\pe1/bq[1] ), .B1(\pe1/aot [7]), 
        .B2(\pe1/bq[2] ), .ZN(n26865) );
  NOR2HSV2 U28715 ( .A1(n26866), .A2(n26865), .ZN(n26867) );
  XNOR2HSV1 U28716 ( .A1(n26868), .A2(n26867), .ZN(n26869) );
  XNOR2HSV1 U28717 ( .A1(n26870), .A2(n26869), .ZN(n26871) );
  XNOR2HSV1 U28718 ( .A1(n26872), .A2(n26871), .ZN(n26873) );
  XNOR2HSV1 U28719 ( .A1(n26874), .A2(n26873), .ZN(n26875) );
  XOR2HSV0 U28720 ( .A1(n26876), .A2(n26875), .Z(n26877) );
  XOR2HSV0 U28721 ( .A1(n26878), .A2(n26877), .Z(n26879) );
  XNOR2HSV1 U28722 ( .A1(n26880), .A2(n26879), .ZN(n26881) );
  XNOR2HSV1 U28723 ( .A1(n26882), .A2(n26881), .ZN(n26884) );
  CLKNAND2HSV0 U28724 ( .A1(n26909), .A2(\pe1/got [7]), .ZN(n26883) );
  XOR2HSV0 U28725 ( .A1(n26884), .A2(n26883), .Z(n26885) );
  XOR2HSV0 U28726 ( .A1(n26886), .A2(n26885), .Z(\pe1/poht [8]) );
  NAND2HSV0 U28727 ( .A1(n27000), .A2(\pe1/got [5]), .ZN(n26908) );
  NAND2HSV0 U28728 ( .A1(n27136), .A2(\pe1/got [3]), .ZN(n26904) );
  NAND2HSV0 U28729 ( .A1(n28460), .A2(\pe1/got [2]), .ZN(n26902) );
  NOR2HSV2 U28730 ( .A1(n26888), .A2(n26887), .ZN(n26900) );
  NAND2HSV0 U28731 ( .A1(\pe1/aot [5]), .A2(\pe1/bq[1] ), .ZN(n26898) );
  NOR2HSV0 U28732 ( .A1(n26890), .A2(n26889), .ZN(n26892) );
  AOI22HSV0 U28733 ( .A1(\pe1/aot [4]), .A2(\pe1/bq[2] ), .B1(\pe1/bq[3] ), 
        .B2(\pe1/aot [3]), .ZN(n26891) );
  NOR2HSV2 U28734 ( .A1(n26892), .A2(n26891), .ZN(n26897) );
  CLKNHSV0 U28735 ( .I(\pe1/aot [2]), .ZN(n26893) );
  NOR2HSV1 U28736 ( .A1(n26893), .A2(n27141), .ZN(n26895) );
  NAND2HSV0 U28737 ( .A1(\pe1/aot [1]), .A2(\pe1/bq[5] ), .ZN(n26894) );
  XOR2HSV0 U28738 ( .A1(n26895), .A2(n26894), .Z(n26896) );
  XOR3HSV2 U28739 ( .A1(n26898), .A2(n26897), .A3(n26896), .Z(n26899) );
  XOR2HSV0 U28740 ( .A1(n26900), .A2(n26899), .Z(n26901) );
  XNOR2HSV1 U28741 ( .A1(n26902), .A2(n26901), .ZN(n26903) );
  XNOR2HSV1 U28742 ( .A1(n26904), .A2(n26903), .ZN(n26906) );
  CLKNAND2HSV0 U28743 ( .A1(n26909), .A2(\pe1/got [4]), .ZN(n26905) );
  XOR2HSV0 U28744 ( .A1(n26906), .A2(n26905), .Z(n26907) );
  XOR2HSV0 U28745 ( .A1(n26908), .A2(n26907), .Z(\pe1/poht [11]) );
  NAND2HSV0 U28746 ( .A1(n27000), .A2(\pe1/got [2]), .ZN(n26915) );
  NAND2HSV2 U28747 ( .A1(n26909), .A2(\pe1/got [1]), .ZN(n26913) );
  NAND2HSV0 U28748 ( .A1(\pe1/aot [1]), .A2(\pe1/bq[2] ), .ZN(n26911) );
  NAND2HSV0 U28749 ( .A1(\pe1/aot [2]), .A2(\pe1/bq[1] ), .ZN(n26910) );
  XOR2HSV0 U28750 ( .A1(n26911), .A2(n26910), .Z(n26912) );
  XOR2HSV0 U28751 ( .A1(n26913), .A2(n26912), .Z(n26914) );
  XOR2HSV0 U28752 ( .A1(n26915), .A2(n26914), .Z(\pe1/poht [14]) );
  CLKNHSV0 U28753 ( .I(n26916), .ZN(n26918) );
  AND3HSV2 U28754 ( .A1(n26924), .A2(n28592), .A3(n26923), .Z(n26917) );
  CLKNAND2HSV1 U28755 ( .A1(n26918), .A2(n26917), .ZN(n26922) );
  NOR2HSV0 U28756 ( .A1(n27974), .A2(n26919), .ZN(n26920) );
  OAI21HSV2 U28757 ( .A1(n26928), .A2(n27976), .B(n26920), .ZN(n26921) );
  NOR2HSV0 U28758 ( .A1(n26930), .A2(n26926), .ZN(n26927) );
  CLKNAND2HSV0 U28759 ( .A1(n26930), .A2(n26929), .ZN(n26931) );
  NOR2HSV2 U28760 ( .A1(n25080), .A2(n26932), .ZN(n26997) );
  NAND2HSV0 U28761 ( .A1(n14038), .A2(n28428), .ZN(n26995) );
  NOR2HSV0 U28762 ( .A1(n27876), .A2(n27871), .ZN(n26993) );
  NAND2HSV0 U28763 ( .A1(\pe4/got [10]), .A2(n27784), .ZN(n26934) );
  NAND2HSV0 U28764 ( .A1(n28578), .A2(\pe4/got [9]), .ZN(n26933) );
  XNOR2HSV1 U28765 ( .A1(n26934), .A2(n26933), .ZN(n26991) );
  NAND2HSV0 U28766 ( .A1(\pe4/ti_7[7] ), .A2(\pe4/got [8]), .ZN(n26989) );
  NAND2HSV0 U28767 ( .A1(n22931), .A2(n13996), .ZN(n26987) );
  NAND2HSV0 U28768 ( .A1(n27739), .A2(\pe4/got [5]), .ZN(n26980) );
  NAND2HSV0 U28769 ( .A1(\pe4/aot [13]), .A2(\pe4/bq[4] ), .ZN(n26936) );
  NAND2HSV0 U28770 ( .A1(\pe4/aot [8]), .A2(\pe4/bq[9] ), .ZN(n26935) );
  XOR2HSV0 U28771 ( .A1(n26936), .A2(n26935), .Z(n26955) );
  NAND2HSV0 U28772 ( .A1(n27066), .A2(\pe4/pq ), .ZN(n26938) );
  NAND2HSV0 U28773 ( .A1(n28683), .A2(\pe4/bq[1] ), .ZN(n26937) );
  XOR2HSV0 U28774 ( .A1(n26938), .A2(n26937), .Z(n26945) );
  OAI21HSV0 U28775 ( .A1(n27088), .A2(n26940), .B(n26939), .ZN(n26941) );
  OAI21HSV0 U28776 ( .A1(n26943), .A2(n26942), .B(n26941), .ZN(n26944) );
  XNOR2HSV1 U28777 ( .A1(n26945), .A2(n26944), .ZN(n26954) );
  NAND2HSV0 U28778 ( .A1(\pe4/bq[3] ), .A2(n28660), .ZN(n26947) );
  NAND2HSV0 U28779 ( .A1(\pe4/aot [11]), .A2(\pe4/bq[6] ), .ZN(n26946) );
  XOR2HSV0 U28780 ( .A1(n26947), .A2(n26946), .Z(n26952) );
  NAND2HSV0 U28781 ( .A1(\pe4/aot [9]), .A2(\pe4/bq[8] ), .ZN(n26950) );
  NAND2HSV0 U28782 ( .A1(\pe4/aot [1]), .A2(n26948), .ZN(n26949) );
  XOR2HSV0 U28783 ( .A1(n26950), .A2(n26949), .Z(n26951) );
  XOR2HSV0 U28784 ( .A1(n26952), .A2(n26951), .Z(n26953) );
  XOR3HSV2 U28785 ( .A1(n26955), .A2(n26954), .A3(n26953), .Z(n26957) );
  NAND2HSV0 U28786 ( .A1(n28671), .A2(\pe4/got [3]), .ZN(n26956) );
  XOR2HSV0 U28787 ( .A1(n26957), .A2(n26956), .Z(n26978) );
  NAND2HSV0 U28788 ( .A1(\pe4/aot [2]), .A2(n26958), .ZN(n26960) );
  NAND2HSV0 U28789 ( .A1(\pe4/aot [3]), .A2(n27060), .ZN(n26959) );
  XOR2HSV0 U28790 ( .A1(n26960), .A2(n26959), .Z(n26965) );
  NAND2HSV0 U28791 ( .A1(\pe4/aot [10]), .A2(\pe4/bq[7] ), .ZN(n26963) );
  NAND2HSV0 U28792 ( .A1(\pe4/aot [4]), .A2(n26961), .ZN(n26962) );
  XOR2HSV0 U28793 ( .A1(n26963), .A2(n26962), .Z(n26964) );
  XOR2HSV0 U28794 ( .A1(n26965), .A2(n26964), .Z(n26974) );
  NAND2HSV0 U28795 ( .A1(\pe4/aot [7]), .A2(\pe4/bq[10] ), .ZN(n26967) );
  NAND2HSV0 U28796 ( .A1(\pe4/got [1]), .A2(n27128), .ZN(n26966) );
  XOR2HSV0 U28797 ( .A1(n26967), .A2(n26966), .Z(n26972) );
  CLKNHSV0 U28798 ( .I(\pe4/aot [6]), .ZN(n27847) );
  NOR2HSV0 U28799 ( .A1(n27847), .A2(n26968), .ZN(n26970) );
  NAND2HSV0 U28800 ( .A1(\pe4/aot [5]), .A2(\pe4/bq[12] ), .ZN(n26969) );
  XOR2HSV0 U28801 ( .A1(n26970), .A2(n26969), .Z(n26971) );
  XOR2HSV0 U28802 ( .A1(n26972), .A2(n26971), .Z(n26973) );
  XOR2HSV0 U28803 ( .A1(n26974), .A2(n26973), .Z(n26976) );
  NAND2HSV0 U28804 ( .A1(n28653), .A2(n28591), .ZN(n26975) );
  XNOR2HSV1 U28805 ( .A1(n26976), .A2(n26975), .ZN(n26977) );
  XNOR2HSV1 U28806 ( .A1(n26978), .A2(n26977), .ZN(n26979) );
  XNOR2HSV1 U28807 ( .A1(n26980), .A2(n26979), .ZN(n26983) );
  INHSV2 U28808 ( .I(\pe4/got [4]), .ZN(n27973) );
  NOR2HSV0 U28809 ( .A1(n26981), .A2(n27973), .ZN(n26982) );
  XNOR2HSV1 U28810 ( .A1(n26983), .A2(n26982), .ZN(n26985) );
  NAND2HSV0 U28811 ( .A1(n28696), .A2(n22826), .ZN(n26984) );
  XOR2HSV0 U28812 ( .A1(n26985), .A2(n26984), .Z(n26986) );
  XNOR2HSV1 U28813 ( .A1(n26987), .A2(n26986), .ZN(n26988) );
  XNOR2HSV1 U28814 ( .A1(n26989), .A2(n26988), .ZN(n26990) );
  XNOR2HSV1 U28815 ( .A1(n26991), .A2(n26990), .ZN(n26992) );
  XOR2HSV0 U28816 ( .A1(n26993), .A2(n26992), .Z(n26994) );
  XNOR2HSV1 U28817 ( .A1(n26995), .A2(n26994), .ZN(n26996) );
  XOR2HSV0 U28818 ( .A1(n26999), .A2(n26998), .Z(po4) );
  NAND2HSV0 U28819 ( .A1(n27000), .A2(\pe1/got [13]), .ZN(n27047) );
  NAND2HSV0 U28820 ( .A1(n27136), .A2(\pe1/got [11]), .ZN(n27043) );
  CLKNAND2HSV0 U28821 ( .A1(n27184), .A2(n27137), .ZN(n27041) );
  NAND2HSV0 U28822 ( .A1(n28609), .A2(\pe1/got [5]), .ZN(n27038) );
  NAND2HSV0 U28823 ( .A1(n27005), .A2(\pe1/got [1]), .ZN(n27031) );
  NAND2HSV0 U28824 ( .A1(\pe1/aot [3]), .A2(\pe1/bq[11] ), .ZN(n27007) );
  NAND2HSV0 U28825 ( .A1(\pe1/aot [8]), .A2(\pe1/bq[6] ), .ZN(n27006) );
  XOR2HSV0 U28826 ( .A1(n27007), .A2(n27006), .Z(n27011) );
  NAND2HSV0 U28827 ( .A1(\pe1/aot [11]), .A2(\pe1/bq[3] ), .ZN(n27009) );
  NAND2HSV0 U28828 ( .A1(\pe1/aot [2]), .A2(\pe1/bq[12] ), .ZN(n27008) );
  XOR2HSV0 U28829 ( .A1(n27009), .A2(n27008), .Z(n27010) );
  XOR2HSV0 U28830 ( .A1(n27011), .A2(n27010), .Z(n27019) );
  NAND2HSV0 U28831 ( .A1(\pe1/aot [4]), .A2(\pe1/bq[10] ), .ZN(n27013) );
  NAND2HSV0 U28832 ( .A1(\pe1/aot [6]), .A2(\pe1/bq[8] ), .ZN(n27012) );
  XOR2HSV0 U28833 ( .A1(n27013), .A2(n27012), .Z(n27017) );
  NAND2HSV0 U28834 ( .A1(\pe1/aot [10]), .A2(\pe1/bq[4] ), .ZN(n27015) );
  NAND2HSV0 U28835 ( .A1(\pe1/aot [9]), .A2(\pe1/bq[5] ), .ZN(n27014) );
  XOR2HSV0 U28836 ( .A1(n27015), .A2(n27014), .Z(n27016) );
  XOR2HSV0 U28837 ( .A1(n27017), .A2(n27016), .Z(n27018) );
  XOR2HSV0 U28838 ( .A1(n27019), .A2(n27018), .Z(n27029) );
  XOR2HSV0 U28839 ( .A1(n27023), .A2(n27022), .Z(n27027) );
  XOR2HSV0 U28840 ( .A1(n27025), .A2(n27024), .Z(n27026) );
  XOR2HSV0 U28841 ( .A1(n27027), .A2(n27026), .Z(n27028) );
  XNOR2HSV1 U28842 ( .A1(n27029), .A2(n27028), .ZN(n27030) );
  XNOR2HSV1 U28843 ( .A1(n27031), .A2(n27030), .ZN(n27033) );
  NAND2HSV0 U28844 ( .A1(n28635), .A2(\pe1/got [2]), .ZN(n27032) );
  XNOR2HSV1 U28845 ( .A1(n27033), .A2(n27032), .ZN(n27036) );
  NAND2HSV0 U28846 ( .A1(n28649), .A2(\pe1/got [3]), .ZN(n27035) );
  NAND2HSV0 U28847 ( .A1(n27166), .A2(n28435), .ZN(n27034) );
  XOR3HSV2 U28848 ( .A1(n27036), .A2(n27035), .A3(n27034), .Z(n27037) );
  NAND2HSV0 U28849 ( .A1(n28589), .A2(n28434), .ZN(n27039) );
  XNOR2HSV1 U28850 ( .A1(n27041), .A2(n27040), .ZN(n27042) );
  NAND2HSV0 U28851 ( .A1(n27185), .A2(n28425), .ZN(n27044) );
  XOR2HSV0 U28852 ( .A1(n27045), .A2(n27044), .Z(n27046) );
  XOR2HSV0 U28853 ( .A1(n27047), .A2(n27046), .Z(\pe1/poht [3]) );
  MUX2HSV2 U28854 ( .I0(\pe5/bq[10] ), .I1(bo5[10]), .S(n27048), .Z(n28712) );
  INHSV2 U28855 ( .I(n27050), .ZN(n27052) );
  MUX2HSV2 U28856 ( .I0(\pe5/bq[6] ), .I1(bo5[6]), .S(n27051), .Z(n28714) );
  MUX2HSV2 U28857 ( .I0(\pe5/bq[3] ), .I1(bo5[3]), .S(n27052), .Z(n28715) );
  MUX2HSV2 U28858 ( .I0(n27053), .I1(bo5[2]), .S(n27052), .Z(n28716) );
  CLKNHSV0 U28859 ( .I(\pe11/bq[13] ), .ZN(n27054) );
  INHSV2 U28860 ( .I(n27054), .ZN(n27056) );
  MUX2HSV2 U28861 ( .I0(bo11[13]), .I1(n27056), .S(n27055), .Z(n28726) );
  MUX2HSV2 U28862 ( .I0(bo11[16]), .I1(n27058), .S(n27057), .Z(n28729) );
  INHSV2 U28863 ( .I(n27692), .ZN(n27706) );
  MUX2HSV2 U28864 ( .I0(bo2[4]), .I1(n27706), .S(n27059), .Z(n28731) );
  MUX2HSV2 U28865 ( .I0(bo4[14]), .I1(n27060), .S(n23508), .Z(n28733) );
  CLKNHSV0 U28866 ( .I(\pe1/bq[10] ), .ZN(n27061) );
  INHSV2 U28867 ( .I(n27061), .ZN(n27063) );
  MUX2HSV2 U28868 ( .I0(bo1[10]), .I1(n27063), .S(n27062), .Z(n28735) );
  MUX2HSV2 U28869 ( .I0(bo1[5]), .I1(\pe1/bq[5] ), .S(n23534), .Z(n28737) );
  MUX2HSV2 U28870 ( .I0(bo4[3]), .I1(\pe4/bq[3] ), .S(n27066), .Z(n28739) );
  MUX2HSV2 U28871 ( .I0(bo1[16]), .I1(n27067), .S(n14005), .Z(n28740) );
  CLKNHSV0 U28872 ( .I(\pe1/bq[13] ), .ZN(n27068) );
  INHSV2 U28873 ( .I(n27068), .ZN(n27069) );
  MUX2HSV2 U28874 ( .I0(bo1[13]), .I1(n27069), .S(n14004), .Z(n28741) );
  MUX2HSV2 U28875 ( .I0(bo1[7]), .I1(\pe1/bq[7] ), .S(n14024), .Z(n28743) );
  MUX2HSV2 U28876 ( .I0(bo1[2]), .I1(\pe1/bq[2] ), .S(n14024), .Z(n28745) );
  MUX2HSV2 U28877 ( .I0(bo6[7]), .I1(\pe6/bq[7] ), .S(n27072), .Z(n28746) );
  MUX2HSV2 U28878 ( .I0(bo6[5]), .I1(\pe6/bq[5] ), .S(n27073), .Z(n28747) );
  MUX2HSV2 U28879 ( .I0(\pe6/bq[3] ), .I1(bo6[3]), .S(n27074), .Z(n28750) );
  CLKNHSV0 U28880 ( .I(\pe4/bq[1] ), .ZN(n27075) );
  INHSV2 U28881 ( .I(n27075), .ZN(n27077) );
  MUX2HSV2 U28882 ( .I0(bo4[1]), .I1(n27077), .S(n27076), .Z(n28751) );
  INHSV1 U28883 ( .I(n27078), .ZN(n27079) );
  MUX2HSV2 U28884 ( .I0(\pe9/bq[5] ), .I1(bo9[5]), .S(n27079), .Z(n28752) );
  CLKNHSV0 U28885 ( .I(\pe9/bq[13] ), .ZN(n27080) );
  INHSV2 U28886 ( .I(n27080), .ZN(n27081) );
  MUX2HSV2 U28887 ( .I0(bo9[13]), .I1(n27081), .S(n27093), .Z(n28754) );
  MUX2HSV2 U28888 ( .I0(bo7[15]), .I1(n27083), .S(n27082), .Z(n28756) );
  CLKNHSV0 U28889 ( .I(\pe7/bq[11] ), .ZN(n27084) );
  INHSV2 U28890 ( .I(n27084), .ZN(n27086) );
  INHSV1 U28891 ( .I(n27085), .ZN(n27094) );
  MUX2HSV2 U28892 ( .I0(bo7[11]), .I1(n27086), .S(n27094), .Z(n28757) );
  MUX2HSV2 U28893 ( .I0(bo7[7]), .I1(\pe7/bq[7] ), .S(n27087), .Z(n28758) );
  MUX2HSV2 U28894 ( .I0(bo7[2]), .I1(\pe7/bq[2] ), .S(n27087), .Z(n28759) );
  MUX2HSV2 U28895 ( .I0(bo4[10]), .I1(\pe4/bq[10] ), .S(n27089), .Z(n28761) );
  MUX2HSV2 U28896 ( .I0(bo4[7]), .I1(\pe4/bq[7] ), .S(n28924), .Z(n28762) );
  MUX2HSV2 U28897 ( .I0(bo4[2]), .I1(\pe4/bq[2] ), .S(n27089), .Z(n28763) );
  CLKNHSV0 U28898 ( .I(\pe9/bq[10] ), .ZN(n27090) );
  INHSV2 U28899 ( .I(n27090), .ZN(n27091) );
  MUX2HSV2 U28900 ( .I0(bo9[10]), .I1(n27091), .S(n27093), .Z(n28764) );
  MUX2HSV2 U28901 ( .I0(bo9[8]), .I1(\pe9/bq[8] ), .S(n27092), .Z(n28765) );
  MUX2HSV2 U28902 ( .I0(bo9[4]), .I1(\pe9/bq[4] ), .S(n27093), .Z(n28766) );
  MUX2HSV2 U28903 ( .I0(bo9[3]), .I1(\pe9/bq[3] ), .S(n27093), .Z(n28767) );
  MUX2HSV2 U28904 ( .I0(bo7[16]), .I1(n25273), .S(n27094), .Z(n28768) );
  MUX2HSV2 U28905 ( .I0(bo7[10]), .I1(\pe7/bq[10] ), .S(n12688), .Z(n28769) );
  MUX2HSV2 U28906 ( .I0(bo4[4]), .I1(\pe4/bq[4] ), .S(n28924), .Z(n28770) );
  MUX2HSV2 U28907 ( .I0(bo7[1]), .I1(\pe7/bq[1] ), .S(n27096), .Z(n28772) );
  MUX2HSV2 U28908 ( .I0(bo7[3]), .I1(\pe7/bq[3] ), .S(n27099), .Z(n28776) );
  MUX2HSV2 U28909 ( .I0(bo4[8]), .I1(\pe4/bq[8] ), .S(n27105), .Z(n28777) );
  MUX2HSV2 U28910 ( .I0(bo9[7]), .I1(\pe9/bq[7] ), .S(n27093), .Z(n28781) );
  MUX2HSV2 U28911 ( .I0(bo7[14]), .I1(n27103), .S(n27102), .Z(n28782) );
  MUX2HSV2 U28912 ( .I0(bo7[4]), .I1(\pe7/bq[4] ), .S(n27104), .Z(n28785) );
  MUX2HSV2 U28913 ( .I0(bo4[6]), .I1(\pe4/bq[6] ), .S(n27105), .Z(n28786) );
  NAND2HSV0 U28914 ( .A1(\pe5/aot [2]), .A2(\pe5/bq[1] ), .ZN(n27108) );
  NAND2HSV0 U28915 ( .A1(\pe5/aot [1]), .A2(\pe5/bq[2] ), .ZN(n27107) );
  XOR2HSV0 U28916 ( .A1(n27108), .A2(n27107), .Z(n27109) );
  NAND2HSV2 U28917 ( .A1(n27112), .A2(n28640), .ZN(n27114) );
  NAND2HSV0 U28918 ( .A1(\pe5/aot [1]), .A2(\pe5/bq[1] ), .ZN(n27113) );
  XOR2HSV0 U28919 ( .A1(n27114), .A2(n27113), .Z(\pe5/poht [15]) );
  NOR2HSV0 U28920 ( .A1(n27116), .A2(n27115), .ZN(n27118) );
  NAND2HSV0 U28921 ( .A1(n27118), .A2(n27117), .ZN(n27120) );
  XNOR2HSV1 U28922 ( .A1(n27120), .A2(n27119), .ZN(pov3[6]) );
  XNOR2HSV0 U28923 ( .A1(n27122), .A2(n27121), .ZN(n27124) );
  XOR2HSV0 U28924 ( .A1(n27124), .A2(n27123), .Z(n29040) );
  INHSV2 U28925 ( .I(\pe4/pq ), .ZN(n27130) );
  MUX2NHSV1 U28926 ( .I0(n27130), .I1(n15764), .S(n27129), .ZN(\pe4/ti_1t ) );
  NAND2HSV0 U28927 ( .A1(n27136), .A2(\pe1/got [9]), .ZN(n27183) );
  NAND2HSV0 U28928 ( .A1(n27137), .A2(\pe1/got [8]), .ZN(n27181) );
  NOR2HSV2 U28929 ( .A1(n27139), .A2(n27138), .ZN(n27179) );
  NOR2HSV2 U28930 ( .A1(n26830), .A2(n27140), .ZN(n27177) );
  NAND2HSV0 U28931 ( .A1(n26854), .A2(\pe1/got [5]), .ZN(n27175) );
  NAND2HSV0 U28932 ( .A1(n28609), .A2(\pe1/got [3]), .ZN(n27171) );
  CLKNHSV0 U28933 ( .I(\pe1/aot [8]), .ZN(n27142) );
  NOR2HSV0 U28934 ( .A1(n27142), .A2(n27141), .ZN(n27145) );
  OAI22HSV1 U28935 ( .A1(n27146), .A2(n27145), .B1(n27144), .B2(n27143), .ZN(
        n27148) );
  XOR2HSV0 U28936 ( .A1(n27148), .A2(n27147), .Z(n27165) );
  NAND2HSV0 U28937 ( .A1(\pe1/aot [4]), .A2(\pe1/bq[8] ), .ZN(n27149) );
  XOR2HSV0 U28938 ( .A1(n27150), .A2(n27149), .Z(n27154) );
  NAND2HSV0 U28939 ( .A1(\pe1/aot [5]), .A2(\pe1/bq[7] ), .ZN(n27152) );
  NAND2HSV0 U28940 ( .A1(\pe1/aot [1]), .A2(\pe1/bq[11] ), .ZN(n27151) );
  XOR2HSV0 U28941 ( .A1(n27152), .A2(n27151), .Z(n27153) );
  XNOR2HSV1 U28942 ( .A1(n27154), .A2(n27153), .ZN(n27164) );
  NAND2HSV0 U28943 ( .A1(\pe1/aot [10]), .A2(\pe1/bq[2] ), .ZN(n27156) );
  NAND2HSV0 U28944 ( .A1(\pe1/aot [2]), .A2(\pe1/bq[10] ), .ZN(n27155) );
  XOR2HSV0 U28945 ( .A1(n27156), .A2(n27155), .Z(n27162) );
  NOR2HSV0 U28946 ( .A1(n27158), .A2(n27157), .ZN(n27160) );
  NAND2HSV0 U28947 ( .A1(\pe1/aot [3]), .A2(\pe1/bq[9] ), .ZN(n27159) );
  XOR2HSV0 U28948 ( .A1(n27160), .A2(n27159), .Z(n27161) );
  XOR2HSV0 U28949 ( .A1(n27162), .A2(n27161), .Z(n27163) );
  XOR3HSV2 U28950 ( .A1(n27165), .A2(n27164), .A3(n27163), .Z(n27169) );
  NAND2HSV0 U28951 ( .A1(n28649), .A2(\pe1/got [1]), .ZN(n27168) );
  NAND2HSV0 U28952 ( .A1(n27166), .A2(\pe1/got [2]), .ZN(n27167) );
  XOR3HSV2 U28953 ( .A1(n27169), .A2(n27168), .A3(n27167), .Z(n27170) );
  XNOR2HSV1 U28954 ( .A1(n27171), .A2(n27170), .ZN(n27173) );
  NAND2HSV0 U28955 ( .A1(n28589), .A2(n28435), .ZN(n27172) );
  XNOR2HSV1 U28956 ( .A1(n27173), .A2(n27172), .ZN(n27174) );
  XNOR2HSV1 U28957 ( .A1(n27175), .A2(n27174), .ZN(n27176) );
  XOR2HSV0 U28958 ( .A1(n27177), .A2(n27176), .Z(n27178) );
  XOR2HSV0 U28959 ( .A1(n27179), .A2(n27178), .Z(n27180) );
  XNOR2HSV1 U28960 ( .A1(n27181), .A2(n27180), .ZN(n27182) );
  XNOR2HSV1 U28961 ( .A1(n27183), .A2(n27182), .ZN(n27187) );
  NAND2HSV0 U28962 ( .A1(n27185), .A2(n27184), .ZN(n27186) );
  XOR2HSV0 U28963 ( .A1(n27189), .A2(n27188), .Z(\pe1/poht [5]) );
  NOR2HSV0 U28964 ( .A1(n27191), .A2(n27190), .ZN(n27193) );
  XOR2HSV0 U28965 ( .A1(n27193), .A2(n27192), .Z(n29027) );
  NOR2HSV2 U28966 ( .A1(n27195), .A2(n27194), .ZN(n27207) );
  NAND2HSV0 U28967 ( .A1(n27197), .A2(n27196), .ZN(n27205) );
  XOR2HSV0 U28968 ( .A1(n27199), .A2(n27198), .Z(n27203) );
  NAND2HSV0 U28969 ( .A1(\pe10/aot [1]), .A2(\pe10/bq[4] ), .ZN(n27201) );
  NAND2HSV0 U28970 ( .A1(\pe10/aot [2]), .A2(\pe10/bq[3] ), .ZN(n27200) );
  XOR2HSV0 U28971 ( .A1(n27201), .A2(n27200), .Z(n27202) );
  XOR2HSV0 U28972 ( .A1(n27203), .A2(n27202), .Z(n27204) );
  XOR2HSV0 U28973 ( .A1(n27205), .A2(n27204), .Z(n27206) );
  INHSV2 U28974 ( .I(n27208), .ZN(n27209) );
  XNOR2HSV1 U28975 ( .A1(n27213), .A2(n27214), .ZN(n27216) );
  XNOR2HSV1 U28976 ( .A1(n27216), .A2(n27215), .ZN(n28985) );
  AOI21HSV1 U28977 ( .A1(n27219), .A2(n27218), .B(n27217), .ZN(n27222) );
  NAND2HSV2 U28978 ( .A1(n27222), .A2(n27221), .ZN(n27224) );
  XOR2HSV0 U28979 ( .A1(n27224), .A2(n27223), .Z(n28958) );
  NOR2HSV0 U28980 ( .A1(n27225), .A2(n28667), .ZN(n27227) );
  XOR2HSV0 U28981 ( .A1(n27227), .A2(n27226), .Z(n29011) );
  CLKNAND2HSV1 U28982 ( .A1(n27294), .A2(n27295), .ZN(n27230) );
  INHSV2 U28983 ( .I(n27230), .ZN(n27398) );
  INHSV2 U28984 ( .I(n27398), .ZN(n27691) );
  NAND2HSV2 U28985 ( .A1(n27231), .A2(n27691), .ZN(n27288) );
  NAND2HSV0 U28986 ( .A1(n27667), .A2(n27543), .ZN(n27282) );
  NAND2HSV0 U28987 ( .A1(n27614), .A2(\pe2/got [8]), .ZN(n27276) );
  NAND2HSV0 U28988 ( .A1(n28427), .A2(n28634), .ZN(n27268) );
  NOR2HSV0 U28989 ( .A1(n27452), .A2(n27633), .ZN(n27266) );
  INHSV2 U28990 ( .I(\pe2/got [2]), .ZN(n27735) );
  NOR2HSV0 U28991 ( .A1(n27423), .A2(n27735), .ZN(n27247) );
  NAND2HSV0 U28992 ( .A1(\pe2/aot [12]), .A2(\pe2/bq[4] ), .ZN(n27234) );
  NAND2HSV0 U28993 ( .A1(\pe2/aot [10]), .A2(\pe2/bq[6] ), .ZN(n27233) );
  XOR2HSV0 U28994 ( .A1(n27234), .A2(n27233), .Z(n27238) );
  NAND2HSV0 U28995 ( .A1(\pe2/aot [13]), .A2(\pe2/bq[3] ), .ZN(n27236) );
  NAND2HSV0 U28996 ( .A1(\pe2/aot [6]), .A2(\pe2/bq[10] ), .ZN(n27235) );
  XOR2HSV0 U28997 ( .A1(n27236), .A2(n27235), .Z(n27237) );
  XOR2HSV0 U28998 ( .A1(n27238), .A2(n27237), .Z(n27245) );
  NAND2HSV0 U28999 ( .A1(\pe2/aot [8]), .A2(\pe2/bq[8] ), .ZN(n27553) );
  NAND2HSV0 U29000 ( .A1(\pe2/aot [14]), .A2(\pe2/bq[2] ), .ZN(n27414) );
  XOR2HSV0 U29001 ( .A1(n27553), .A2(n27414), .Z(n27243) );
  NAND2HSV0 U29002 ( .A1(\pe2/aot [7]), .A2(\pe2/bq[9] ), .ZN(n27241) );
  NAND2HSV0 U29003 ( .A1(\pe2/aot [1]), .A2(\pe2/bq[15] ), .ZN(n27240) );
  XOR2HSV0 U29004 ( .A1(n27241), .A2(n27240), .Z(n27242) );
  XOR2HSV0 U29005 ( .A1(n27243), .A2(n27242), .Z(n27244) );
  XOR2HSV0 U29006 ( .A1(n27245), .A2(n27244), .Z(n27246) );
  XOR2HSV0 U29007 ( .A1(n27247), .A2(n27246), .Z(n27264) );
  NAND2HSV0 U29008 ( .A1(\pe2/aot [4]), .A2(\pe2/bq[12] ), .ZN(n27249) );
  NAND2HSV0 U29009 ( .A1(\pe2/aot [3]), .A2(\pe2/bq[13] ), .ZN(n27248) );
  XOR2HSV0 U29010 ( .A1(n27249), .A2(n27248), .Z(n27254) );
  NAND2HSV0 U29011 ( .A1(\pe2/aot [2]), .A2(n27312), .ZN(n27252) );
  NAND2HSV0 U29012 ( .A1(\pe2/aot [9]), .A2(\pe2/bq[7] ), .ZN(n27251) );
  XOR2HSV0 U29013 ( .A1(n27252), .A2(n27251), .Z(n27253) );
  XOR2HSV0 U29014 ( .A1(n27254), .A2(n27253), .Z(n27260) );
  NAND2HSV0 U29015 ( .A1(\pe2/aot [5]), .A2(\pe2/bq[1] ), .ZN(n27709) );
  NOR2HSV0 U29016 ( .A1(n27255), .A2(n27709), .ZN(n27257) );
  AOI22HSV0 U29017 ( .A1(\pe2/bq[1] ), .A2(\pe2/aot [15]), .B1(\pe2/bq[11] ), 
        .B2(\pe2/aot [5]), .ZN(n27256) );
  NOR2HSV2 U29018 ( .A1(n27257), .A2(n27256), .ZN(n27258) );
  NAND2HSV0 U29019 ( .A1(\pe2/aot [11]), .A2(\pe2/bq[5] ), .ZN(n27359) );
  XNOR2HSV1 U29020 ( .A1(n27258), .A2(n27359), .ZN(n27259) );
  XNOR2HSV1 U29021 ( .A1(n27260), .A2(n27259), .ZN(n27262) );
  NAND2HSV0 U29022 ( .A1(n28697), .A2(\pe2/got [1]), .ZN(n27261) );
  XOR2HSV0 U29023 ( .A1(n27262), .A2(n27261), .Z(n27263) );
  XNOR2HSV1 U29024 ( .A1(n27264), .A2(n27263), .ZN(n27265) );
  XOR2HSV0 U29025 ( .A1(n27266), .A2(n27265), .Z(n27267) );
  XNOR2HSV1 U29026 ( .A1(n27268), .A2(n27267), .ZN(n27270) );
  NAND2HSV0 U29027 ( .A1(n27485), .A2(n27719), .ZN(n27269) );
  XNOR2HSV1 U29028 ( .A1(n27270), .A2(n27269), .ZN(n27274) );
  CLKNHSV1 U29029 ( .I(n27271), .ZN(n27594) );
  NOR2HSV2 U29030 ( .A1(n27594), .A2(n27498), .ZN(n27273) );
  NAND2HSV0 U29031 ( .A1(n28617), .A2(n14046), .ZN(n27272) );
  XOR3HSV2 U29032 ( .A1(n27274), .A2(n27273), .A3(n27272), .Z(n27275) );
  XNOR2HSV1 U29033 ( .A1(n27276), .A2(n27275), .ZN(n27280) );
  BUFHSV2 U29034 ( .I(n27277), .Z(n27678) );
  NOR2HSV2 U29035 ( .A1(n27678), .A2(n27610), .ZN(n27279) );
  NAND2HSV0 U29036 ( .A1(\pe2/got [10]), .A2(n27344), .ZN(n27278) );
  XOR3HSV2 U29037 ( .A1(n27280), .A2(n27279), .A3(n27278), .Z(n27281) );
  XNOR2HSV1 U29038 ( .A1(n27282), .A2(n27281), .ZN(n27286) );
  NAND2HSV0 U29039 ( .A1(n27640), .A2(n27544), .ZN(n27285) );
  XOR2HSV0 U29040 ( .A1(n27286), .A2(n27285), .Z(n27287) );
  XNOR2HSV1 U29041 ( .A1(n27288), .A2(n27287), .ZN(n27293) );
  NAND2HSV2 U29042 ( .A1(n28456), .A2(n22085), .ZN(n27292) );
  CLKNAND2HSV3 U29043 ( .A1(n27290), .A2(n27289), .ZN(n27726) );
  CLKNAND2HSV1 U29044 ( .A1(n27726), .A2(\pe2/got [14]), .ZN(n27291) );
  XOR3HSV2 U29045 ( .A1(n27293), .A2(n27292), .A3(n27291), .Z(\pe2/poht [1])
         );
  CLKNAND2HSV0 U29046 ( .A1(n27731), .A2(n21144), .ZN(n27353) );
  NAND2HSV0 U29047 ( .A1(n27667), .A2(n27544), .ZN(n27349) );
  NAND2HSV0 U29048 ( .A1(n27614), .A2(n27647), .ZN(n27343) );
  NAND2HSV0 U29049 ( .A1(n28427), .A2(n27719), .ZN(n27336) );
  NOR2HSV0 U29050 ( .A1(n27452), .A2(n27718), .ZN(n27334) );
  NOR2HSV0 U29051 ( .A1(n27423), .A2(n27633), .ZN(n27310) );
  NAND2HSV0 U29052 ( .A1(\pe2/aot [13]), .A2(\pe2/bq[4] ), .ZN(n27469) );
  NAND2HSV0 U29053 ( .A1(\pe2/bq[7] ), .A2(\pe2/aot [10]), .ZN(n27364) );
  XOR2HSV0 U29054 ( .A1(n27469), .A2(n27364), .Z(n27308) );
  CLKNHSV0 U29055 ( .I(\pe2/aot [12]), .ZN(n27296) );
  NOR2HSV0 U29056 ( .A1(n27296), .A2(n27652), .ZN(n27501) );
  AOI22HSV0 U29057 ( .A1(n11953), .A2(n27723), .B1(\pe2/aot [12]), .B2(
        \pe2/bq[5] ), .ZN(n27297) );
  AOI21HSV0 U29058 ( .A1(n27501), .A2(n27298), .B(n27297), .ZN(n27301) );
  NAND2HSV0 U29059 ( .A1(\pe2/aot [2]), .A2(\pe2/bq[9] ), .ZN(n27576) );
  XOR2HSV0 U29060 ( .A1(n27301), .A2(n27300), .Z(n27307) );
  NAND2HSV0 U29061 ( .A1(\pe2/aot [4]), .A2(\pe2/bq[13] ), .ZN(n27303) );
  NAND2HSV0 U29062 ( .A1(\pe2/aot [7]), .A2(\pe2/bq[10] ), .ZN(n27302) );
  XOR2HSV0 U29063 ( .A1(n27303), .A2(n27302), .Z(n27305) );
  XOR2HSV0 U29064 ( .A1(n27305), .A2(n27304), .Z(n27306) );
  XOR3HSV2 U29065 ( .A1(n27308), .A2(n27307), .A3(n27306), .Z(n27309) );
  XNOR2HSV1 U29066 ( .A1(n27310), .A2(n27309), .ZN(n27332) );
  NAND2HSV0 U29067 ( .A1(n27311), .A2(\pe2/pq ), .ZN(n27314) );
  NAND2HSV0 U29068 ( .A1(\pe2/aot [3]), .A2(n27312), .ZN(n27313) );
  XOR2HSV0 U29069 ( .A1(n27314), .A2(n27313), .Z(n27318) );
  NAND2HSV0 U29070 ( .A1(n14020), .A2(\pe2/bq[3] ), .ZN(n27316) );
  NAND2HSV0 U29071 ( .A1(\pe2/aot [15]), .A2(\pe2/bq[2] ), .ZN(n27315) );
  XOR2HSV0 U29072 ( .A1(n27316), .A2(n27315), .Z(n27317) );
  XOR2HSV0 U29073 ( .A1(n27318), .A2(n27317), .Z(n27328) );
  NAND2HSV0 U29074 ( .A1(\pe2/aot [6]), .A2(\pe2/bq[11] ), .ZN(n27320) );
  NAND2HSV0 U29075 ( .A1(\pe2/aot [5]), .A2(\pe2/bq[12] ), .ZN(n27319) );
  XOR2HSV0 U29076 ( .A1(n27320), .A2(n27319), .Z(n27326) );
  NAND2HSV0 U29077 ( .A1(\pe2/got [1]), .A2(n27321), .ZN(n27324) );
  INAND2HSV0 U29078 ( .A1(n27322), .B1(\pe2/aot [1]), .ZN(n27323) );
  XOR2HSV0 U29079 ( .A1(n27324), .A2(n27323), .Z(n27325) );
  XOR2HSV0 U29080 ( .A1(n27326), .A2(n27325), .Z(n27327) );
  XOR2HSV0 U29081 ( .A1(n27328), .A2(n27327), .Z(n27330) );
  NAND2HSV0 U29082 ( .A1(n28697), .A2(\pe2/got [2]), .ZN(n27329) );
  XNOR2HSV1 U29083 ( .A1(n27330), .A2(n27329), .ZN(n27331) );
  XOR2HSV0 U29084 ( .A1(n27332), .A2(n27331), .Z(n27333) );
  XOR2HSV0 U29085 ( .A1(n27334), .A2(n27333), .Z(n27335) );
  XNOR2HSV1 U29086 ( .A1(n27336), .A2(n27335), .ZN(n27338) );
  NAND2HSV0 U29087 ( .A1(n27524), .A2(n14003), .ZN(n27337) );
  XNOR2HSV1 U29088 ( .A1(n27338), .A2(n27337), .ZN(n27341) );
  NOR2HSV2 U29089 ( .A1(n27594), .A2(n27572), .ZN(n27340) );
  CLKNHSV0 U29090 ( .I(n27432), .ZN(n27595) );
  NOR2HSV1 U29091 ( .A1(n27595), .A2(n27645), .ZN(n27339) );
  XOR3HSV2 U29092 ( .A1(n27341), .A2(n27340), .A3(n27339), .Z(n27342) );
  XNOR2HSV1 U29093 ( .A1(n27343), .A2(n27342), .ZN(n27347) );
  NOR2HSV0 U29094 ( .A1(n27438), .A2(n27394), .ZN(n27346) );
  NAND2HSV0 U29095 ( .A1(n27344), .A2(n27543), .ZN(n27345) );
  XOR3HSV2 U29096 ( .A1(n27347), .A2(n27346), .A3(n27345), .Z(n27348) );
  XNOR2HSV1 U29097 ( .A1(n27349), .A2(n27348), .ZN(n27351) );
  CLKNAND2HSV1 U29098 ( .A1(n27640), .A2(\pe2/got [13]), .ZN(n27350) );
  XNOR2HSV1 U29099 ( .A1(n27351), .A2(n27350), .ZN(n27352) );
  XNOR2HSV1 U29100 ( .A1(n27353), .A2(n27352), .ZN(n27357) );
  INHSV2 U29101 ( .I(n27354), .ZN(n27571) );
  NOR2HSV2 U29102 ( .A1(n27646), .A2(n21225), .ZN(n27356) );
  CLKNAND2HSV0 U29103 ( .A1(n27736), .A2(n28693), .ZN(n27355) );
  XOR3HSV2 U29104 ( .A1(n27357), .A2(n27356), .A3(n27355), .Z(po2) );
  CLKNAND2HSV0 U29105 ( .A1(n27731), .A2(n27647), .ZN(n27393) );
  NAND2HSV0 U29106 ( .A1(n27657), .A2(n14046), .ZN(n27389) );
  NAND2HSV0 U29107 ( .A1(n27614), .A2(n28634), .ZN(n27384) );
  NAND2HSV0 U29108 ( .A1(n14055), .A2(n27524), .ZN(n27379) );
  NAND2HSV0 U29109 ( .A1(\pe2/bq[1] ), .A2(\pe2/aot [7]), .ZN(n27675) );
  AO22HSV2 U29110 ( .A1(\pe2/aot [11]), .A2(\pe2/bq[1] ), .B1(\pe2/aot [7]), 
        .B2(\pe2/bq[5] ), .Z(n27358) );
  OAI21HSV1 U29111 ( .A1(n27675), .A2(n27359), .B(n27358), .ZN(n27361) );
  NAND2HSV0 U29112 ( .A1(\pe2/aot [4]), .A2(\pe2/bq[8] ), .ZN(n27360) );
  XNOR2HSV1 U29113 ( .A1(n27361), .A2(n27360), .ZN(n27377) );
  NAND2HSV0 U29114 ( .A1(\pe2/aot [8]), .A2(\pe2/bq[4] ), .ZN(n27363) );
  NAND2HSV0 U29115 ( .A1(\pe2/aot [9]), .A2(\pe2/bq[3] ), .ZN(n27362) );
  XOR2HSV0 U29116 ( .A1(n27363), .A2(n27362), .Z(n27368) );
  NAND2HSV0 U29117 ( .A1(\pe2/aot [5]), .A2(\pe2/bq[2] ), .ZN(n27651) );
  NOR2HSV0 U29118 ( .A1(n27364), .A2(n27651), .ZN(n27366) );
  AOI22HSV0 U29119 ( .A1(\pe2/aot [10]), .A2(\pe2/bq[2] ), .B1(\pe2/bq[7] ), 
        .B2(\pe2/aot [5]), .ZN(n27365) );
  NOR2HSV2 U29120 ( .A1(n27366), .A2(n27365), .ZN(n27367) );
  XNOR2HSV1 U29121 ( .A1(n27368), .A2(n27367), .ZN(n27376) );
  NAND2HSV0 U29122 ( .A1(\pe2/aot [2]), .A2(\pe2/bq[10] ), .ZN(n27370) );
  NAND2HSV0 U29123 ( .A1(\pe2/aot [1]), .A2(\pe2/bq[11] ), .ZN(n27369) );
  XOR2HSV0 U29124 ( .A1(n27370), .A2(n27369), .Z(n27374) );
  NAND2HSV0 U29125 ( .A1(\pe2/aot [3]), .A2(\pe2/bq[9] ), .ZN(n27372) );
  NAND2HSV0 U29126 ( .A1(\pe2/aot [6]), .A2(\pe2/bq[6] ), .ZN(n27371) );
  XOR2HSV0 U29127 ( .A1(n27372), .A2(n27371), .Z(n27373) );
  XOR2HSV0 U29128 ( .A1(n27374), .A2(n27373), .Z(n27375) );
  XOR3HSV2 U29129 ( .A1(n27377), .A2(n27376), .A3(n27375), .Z(n27378) );
  XNOR2HSV1 U29130 ( .A1(n27379), .A2(n27378), .ZN(n27382) );
  NOR2HSV2 U29131 ( .A1(n27594), .A2(n27735), .ZN(n27381) );
  NOR2HSV1 U29132 ( .A1(n27595), .A2(n27633), .ZN(n27380) );
  XOR3HSV2 U29133 ( .A1(n27382), .A2(n27381), .A3(n27380), .Z(n27383) );
  XNOR2HSV1 U29134 ( .A1(n27384), .A2(n27383), .ZN(n27387) );
  CLKNHSV0 U29135 ( .I(n28805), .ZN(n27634) );
  NOR2HSV2 U29136 ( .A1(n27634), .A2(n27663), .ZN(n27386) );
  BUFHSV2 U29137 ( .I(n27439), .Z(n27679) );
  CLKNAND2HSV1 U29138 ( .A1(n27679), .A2(n14003), .ZN(n27385) );
  XOR3HSV2 U29139 ( .A1(n27387), .A2(n27386), .A3(n27385), .Z(n27388) );
  XNOR2HSV1 U29140 ( .A1(n27389), .A2(n27388), .ZN(n27391) );
  NAND2HSV0 U29141 ( .A1(n28702), .A2(\pe2/got [8]), .ZN(n27390) );
  XOR2HSV0 U29142 ( .A1(n27391), .A2(n27390), .Z(n27392) );
  XOR2HSV0 U29143 ( .A1(n27393), .A2(n27392), .Z(n27397) );
  NOR2HSV2 U29144 ( .A1(n12302), .A2(n27394), .ZN(n27396) );
  XOR3HSV2 U29145 ( .A1(n27397), .A2(n27396), .A3(n27395), .Z(\pe2/poht [5])
         );
  INHSV4 U29146 ( .I(n27398), .ZN(n27705) );
  NAND2HSV2 U29147 ( .A1(n27705), .A2(n27544), .ZN(n27448) );
  NAND2HSV0 U29148 ( .A1(n27667), .A2(\pe2/got [10]), .ZN(n27444) );
  NAND2HSV0 U29149 ( .A1(n27614), .A2(n14046), .ZN(n27437) );
  NAND2HSV0 U29150 ( .A1(n28427), .A2(n14052), .ZN(n27429) );
  NOR2HSV0 U29151 ( .A1(n27452), .A2(n27735), .ZN(n27427) );
  NAND2HSV0 U29152 ( .A1(\pe2/aot [2]), .A2(\pe2/bq[13] ), .ZN(n27400) );
  NAND2HSV0 U29153 ( .A1(\pe2/aot [1]), .A2(n27312), .ZN(n27399) );
  XOR2HSV0 U29154 ( .A1(n27400), .A2(n27399), .Z(n27404) );
  NAND2HSV0 U29155 ( .A1(\pe2/aot [7]), .A2(\pe2/bq[8] ), .ZN(n27402) );
  NAND2HSV0 U29156 ( .A1(\pe2/aot [3]), .A2(\pe2/bq[12] ), .ZN(n27401) );
  XOR2HSV0 U29157 ( .A1(n27402), .A2(n27401), .Z(n27403) );
  XOR2HSV0 U29158 ( .A1(n27404), .A2(n27403), .Z(n27412) );
  NAND2HSV0 U29159 ( .A1(\pe2/aot [8]), .A2(\pe2/bq[7] ), .ZN(n27406) );
  NAND2HSV0 U29160 ( .A1(\pe2/aot [10]), .A2(\pe2/bq[5] ), .ZN(n27405) );
  XOR2HSV0 U29161 ( .A1(n27406), .A2(n27405), .Z(n27410) );
  NAND2HSV0 U29162 ( .A1(\pe2/aot [4]), .A2(\pe2/bq[11] ), .ZN(n27408) );
  NAND2HSV0 U29163 ( .A1(\pe2/aot [12]), .A2(\pe2/bq[3] ), .ZN(n27407) );
  XOR2HSV0 U29164 ( .A1(n27408), .A2(n27407), .Z(n27409) );
  XNOR2HSV1 U29165 ( .A1(n27410), .A2(n27409), .ZN(n27411) );
  XNOR2HSV1 U29166 ( .A1(n27412), .A2(n27411), .ZN(n27422) );
  NAND2HSV0 U29167 ( .A1(\pe2/aot [13]), .A2(\pe2/bq[1] ), .ZN(n27472) );
  AO22HSV2 U29168 ( .A1(n27723), .A2(n14020), .B1(\pe2/aot [13]), .B2(
        \pe2/bq[2] ), .Z(n27413) );
  OAI21HSV2 U29169 ( .A1(n27472), .A2(n27414), .B(n27413), .ZN(n27420) );
  NAND2HSV0 U29170 ( .A1(\pe2/aot [6]), .A2(\pe2/bq[9] ), .ZN(n27416) );
  NAND2HSV0 U29171 ( .A1(\pe2/aot [5]), .A2(\pe2/bq[10] ), .ZN(n27415) );
  XOR2HSV0 U29172 ( .A1(n27416), .A2(n27415), .Z(n27419) );
  NAND2HSV0 U29173 ( .A1(\pe2/bq[6] ), .A2(\pe2/aot [9]), .ZN(n27617) );
  XOR2HSV0 U29174 ( .A1(n27417), .A2(n27617), .Z(n27418) );
  XOR3HSV2 U29175 ( .A1(n27420), .A2(n27419), .A3(n27418), .Z(n27421) );
  XNOR2HSV1 U29176 ( .A1(n27422), .A2(n27421), .ZN(n27425) );
  NOR2HSV0 U29177 ( .A1(n27423), .A2(n27677), .ZN(n27424) );
  XNOR2HSV1 U29178 ( .A1(n27425), .A2(n27424), .ZN(n27426) );
  XOR2HSV0 U29179 ( .A1(n27427), .A2(n27426), .Z(n27428) );
  XNOR2HSV1 U29180 ( .A1(n27429), .A2(n27428), .ZN(n27431) );
  NAND2HSV0 U29181 ( .A1(n27485), .A2(n28634), .ZN(n27430) );
  XNOR2HSV1 U29182 ( .A1(n27431), .A2(n27430), .ZN(n27435) );
  NOR2HSV1 U29183 ( .A1(n27594), .A2(n27663), .ZN(n27434) );
  NAND2HSV0 U29184 ( .A1(n27432), .A2(n14003), .ZN(n27433) );
  XOR3HSV2 U29185 ( .A1(n27435), .A2(n27434), .A3(n27433), .Z(n27436) );
  XNOR2HSV1 U29186 ( .A1(n27437), .A2(n27436), .ZN(n27442) );
  NOR2HSV0 U29187 ( .A1(n27438), .A2(n27645), .ZN(n27441) );
  NAND2HSV0 U29188 ( .A1(n28474), .A2(n27647), .ZN(n27440) );
  XOR3HSV2 U29189 ( .A1(n27442), .A2(n27441), .A3(n27440), .Z(n27443) );
  XNOR2HSV1 U29190 ( .A1(n27444), .A2(n27443), .ZN(n27446) );
  NAND2HSV0 U29191 ( .A1(n27640), .A2(n27543), .ZN(n27445) );
  XOR2HSV0 U29192 ( .A1(n27446), .A2(n27445), .Z(n27447) );
  NAND2HSV2 U29193 ( .A1(n27726), .A2(n27231), .ZN(n27450) );
  CLKNAND2HSV0 U29194 ( .A1(n28456), .A2(n17767), .ZN(n27449) );
  XOR3HSV2 U29195 ( .A1(n27451), .A2(n27450), .A3(n27449), .Z(\pe2/poht [2])
         );
  NAND2HSV2 U29196 ( .A1(n27691), .A2(n27543), .ZN(n27493) );
  CLKNAND2HSV0 U29197 ( .A1(n27657), .A2(n27647), .ZN(n27489) );
  NAND2HSV0 U29198 ( .A1(n28427), .A2(\pe2/got [2]), .ZN(n27484) );
  NOR2HSV0 U29199 ( .A1(n27452), .A2(n27677), .ZN(n27482) );
  NAND2HSV0 U29200 ( .A1(\pe2/aot [8]), .A2(\pe2/bq[6] ), .ZN(n27454) );
  NAND2HSV0 U29201 ( .A1(\pe2/aot [6]), .A2(\pe2/bq[8] ), .ZN(n27453) );
  XOR2HSV0 U29202 ( .A1(n27454), .A2(n27453), .Z(n27458) );
  NAND2HSV0 U29203 ( .A1(\pe2/aot [3]), .A2(\pe2/bq[11] ), .ZN(n27456) );
  NAND2HSV0 U29204 ( .A1(\pe2/aot [1]), .A2(\pe2/bq[13] ), .ZN(n27455) );
  XOR2HSV0 U29205 ( .A1(n27456), .A2(n27455), .Z(n27457) );
  XOR2HSV0 U29206 ( .A1(n27458), .A2(n27457), .Z(n27468) );
  NAND2HSV0 U29207 ( .A1(\pe2/aot [4]), .A2(\pe2/bq[10] ), .ZN(n27460) );
  NAND2HSV0 U29208 ( .A1(\pe2/aot [5]), .A2(\pe2/bq[9] ), .ZN(n27459) );
  XOR2HSV0 U29209 ( .A1(n27460), .A2(n27459), .Z(n27466) );
  NOR2HSV0 U29210 ( .A1(n27580), .A2(n27461), .ZN(n27673) );
  CLKNHSV0 U29211 ( .I(\pe2/bq[3] ), .ZN(n27710) );
  NOR2HSV0 U29212 ( .A1(n27462), .A2(n27710), .ZN(n27464) );
  NAND2HSV0 U29213 ( .A1(\pe2/aot [7]), .A2(\pe2/bq[3] ), .ZN(n27618) );
  OAI22HSV0 U29214 ( .A1(n27673), .A2(n27464), .B1(n27463), .B2(n27618), .ZN(
        n27465) );
  XNOR2HSV1 U29215 ( .A1(n27466), .A2(n27465), .ZN(n27467) );
  XNOR2HSV1 U29216 ( .A1(n27468), .A2(n27467), .ZN(n27480) );
  NAND2HSV0 U29217 ( .A1(\pe2/aot [10]), .A2(\pe2/bq[4] ), .ZN(n27471) );
  NAND2HSV0 U29218 ( .A1(\pe2/bq[1] ), .A2(\pe2/aot [10]), .ZN(n27577) );
  NOR2HSV0 U29219 ( .A1(n27577), .A2(n27469), .ZN(n27470) );
  AOI21HSV2 U29220 ( .A1(n27472), .A2(n27471), .B(n27470), .ZN(n27474) );
  NAND2HSV0 U29221 ( .A1(\pe2/aot [9]), .A2(\pe2/bq[5] ), .ZN(n27473) );
  XNOR2HSV1 U29222 ( .A1(n27474), .A2(n27473), .ZN(n27478) );
  NAND2HSV0 U29223 ( .A1(\pe2/aot [12]), .A2(\pe2/bq[2] ), .ZN(n27476) );
  NAND2HSV0 U29224 ( .A1(\pe2/aot [2]), .A2(\pe2/bq[12] ), .ZN(n27475) );
  XOR2HSV0 U29225 ( .A1(n27476), .A2(n27475), .Z(n27477) );
  XOR2HSV0 U29226 ( .A1(n27478), .A2(n27477), .Z(n27479) );
  XNOR2HSV1 U29227 ( .A1(n27480), .A2(n27479), .ZN(n27481) );
  XOR2HSV0 U29228 ( .A1(n27482), .A2(n27481), .Z(n27483) );
  XNOR2HSV1 U29229 ( .A1(n27484), .A2(n27483), .ZN(n27487) );
  NAND2HSV0 U29230 ( .A1(n27485), .A2(n14052), .ZN(n27486) );
  NAND2HSV0 U29231 ( .A1(n27640), .A2(\pe2/got [10]), .ZN(n27490) );
  XOR2HSV0 U29232 ( .A1(n27491), .A2(n27490), .Z(n27492) );
  XNOR2HSV1 U29233 ( .A1(n27493), .A2(n27492), .ZN(n27497) );
  NAND2HSV2 U29234 ( .A1(n27726), .A2(n27544), .ZN(n27496) );
  CLKNAND2HSV1 U29235 ( .A1(n27727), .A2(n28429), .ZN(n27495) );
  XOR3HSV2 U29236 ( .A1(n27497), .A2(n27496), .A3(n27495), .Z(\pe2/poht [3])
         );
  NAND2HSV2 U29237 ( .A1(n27691), .A2(\pe2/got [10]), .ZN(n27542) );
  CLKNAND2HSV0 U29238 ( .A1(n27667), .A2(\pe2/got [8]), .ZN(n27538) );
  NOR2HSV2 U29239 ( .A1(n27678), .A2(n27498), .ZN(n27534) );
  NAND2HSV0 U29240 ( .A1(n27614), .A2(n27719), .ZN(n27532) );
  NAND2HSV0 U29241 ( .A1(n28427), .A2(n14055), .ZN(n27523) );
  NOR2HSV0 U29242 ( .A1(n27580), .A2(n27654), .ZN(n27500) );
  OAI22HSV0 U29243 ( .A1(n27501), .A2(n27500), .B1(n27499), .B2(n27675), .ZN(
        n27506) );
  NAND2HSV0 U29244 ( .A1(\pe2/aot [4]), .A2(\pe2/bq[2] ), .ZN(n27708) );
  NOR2HSV0 U29245 ( .A1(n27502), .A2(n27708), .ZN(n27504) );
  AOI22HSV0 U29246 ( .A1(\pe2/aot [11]), .A2(\pe2/bq[2] ), .B1(\pe2/bq[9] ), 
        .B2(\pe2/aot [4]), .ZN(n27503) );
  NOR2HSV1 U29247 ( .A1(n27504), .A2(n27503), .ZN(n27505) );
  XOR2HSV0 U29248 ( .A1(n27506), .A2(n27505), .Z(n27521) );
  NAND2HSV0 U29249 ( .A1(\pe2/aot [9]), .A2(\pe2/bq[4] ), .ZN(n27508) );
  NAND2HSV0 U29250 ( .A1(\pe2/aot [6]), .A2(\pe2/bq[7] ), .ZN(n27507) );
  XOR2HSV0 U29251 ( .A1(n27508), .A2(n27507), .Z(n27512) );
  NAND2HSV0 U29252 ( .A1(\pe2/aot [10]), .A2(\pe2/bq[3] ), .ZN(n27510) );
  NAND2HSV0 U29253 ( .A1(\pe2/aot [3]), .A2(\pe2/bq[10] ), .ZN(n27509) );
  XOR2HSV0 U29254 ( .A1(n27510), .A2(n27509), .Z(n27511) );
  XNOR2HSV1 U29255 ( .A1(n27512), .A2(n27511), .ZN(n27520) );
  NAND2HSV0 U29256 ( .A1(\pe2/aot [1]), .A2(\pe2/bq[12] ), .ZN(n27514) );
  NAND2HSV0 U29257 ( .A1(\pe2/aot [5]), .A2(\pe2/bq[8] ), .ZN(n27513) );
  XOR2HSV0 U29258 ( .A1(n27514), .A2(n27513), .Z(n27518) );
  NAND2HSV0 U29259 ( .A1(\pe2/aot [2]), .A2(\pe2/bq[11] ), .ZN(n27516) );
  NAND2HSV0 U29260 ( .A1(\pe2/aot [8]), .A2(\pe2/bq[5] ), .ZN(n27515) );
  XOR2HSV0 U29261 ( .A1(n27516), .A2(n27515), .Z(n27517) );
  XOR2HSV0 U29262 ( .A1(n27518), .A2(n27517), .Z(n27519) );
  XOR3HSV2 U29263 ( .A1(n27521), .A2(n27520), .A3(n27519), .Z(n27522) );
  XNOR2HSV1 U29264 ( .A1(n27523), .A2(n27522), .ZN(n27526) );
  NAND2HSV0 U29265 ( .A1(n27524), .A2(\pe2/got [2]), .ZN(n27525) );
  XNOR2HSV1 U29266 ( .A1(n27526), .A2(n27525), .ZN(n27530) );
  NOR2HSV1 U29267 ( .A1(n27527), .A2(n27633), .ZN(n27529) );
  NOR2HSV1 U29268 ( .A1(n27595), .A2(n27718), .ZN(n27528) );
  XOR3HSV2 U29269 ( .A1(n27530), .A2(n27529), .A3(n27528), .Z(n27531) );
  XNOR2HSV1 U29270 ( .A1(n27532), .A2(n27531), .ZN(n27533) );
  XNOR2HSV4 U29271 ( .A1(n27534), .A2(n27533), .ZN(n27536) );
  XOR2HSV2 U29272 ( .A1(n27536), .A2(n27535), .Z(n27537) );
  XNOR2HSV4 U29273 ( .A1(n27538), .A2(n27537), .ZN(n27540) );
  XNOR2HSV4 U29274 ( .A1(n27540), .A2(n27539), .ZN(n27541) );
  NAND2HSV2 U29275 ( .A1(n28701), .A2(n27543), .ZN(n27546) );
  NAND2HSV2 U29276 ( .A1(n27705), .A2(n14003), .ZN(n27570) );
  NAND2HSV0 U29277 ( .A1(n27657), .A2(n28634), .ZN(n27566) );
  NAND2HSV0 U29278 ( .A1(n14055), .A2(n21816), .ZN(n27561) );
  NAND2HSV0 U29279 ( .A1(\pe2/aot [3]), .A2(\pe2/bq[6] ), .ZN(n27548) );
  NAND2HSV0 U29280 ( .A1(\pe2/aot [5]), .A2(\pe2/bq[4] ), .ZN(n27547) );
  XOR2HSV0 U29281 ( .A1(n27548), .A2(n27547), .Z(n27552) );
  NAND2HSV0 U29282 ( .A1(\pe2/aot [4]), .A2(\pe2/bq[5] ), .ZN(n27550) );
  NAND2HSV0 U29283 ( .A1(\pe2/aot [6]), .A2(\pe2/bq[3] ), .ZN(n27549) );
  XOR2HSV0 U29284 ( .A1(n27550), .A2(n27549), .Z(n27551) );
  XOR2HSV0 U29285 ( .A1(n27552), .A2(n27551), .Z(n27559) );
  NOR2HSV2 U29286 ( .A1(n27554), .A2(n27250), .ZN(n27733) );
  AOI22HSV0 U29287 ( .A1(\pe2/aot [7]), .A2(\pe2/bq[2] ), .B1(\pe2/bq[7] ), 
        .B2(\pe2/aot [2]), .ZN(n27555) );
  AOI21HSV0 U29288 ( .A1(n27733), .A2(n27673), .B(n27555), .ZN(n27556) );
  XOR2HSV0 U29289 ( .A1(n27557), .A2(n27556), .Z(n27558) );
  XNOR2HSV1 U29290 ( .A1(n27559), .A2(n27558), .ZN(n27560) );
  XOR2HSV0 U29291 ( .A1(n27561), .A2(n27560), .Z(n27564) );
  NOR2HSV2 U29292 ( .A1(n27678), .A2(n27735), .ZN(n27563) );
  CLKNAND2HSV1 U29293 ( .A1(n27679), .A2(n14052), .ZN(n27562) );
  XOR3HSV2 U29294 ( .A1(n27564), .A2(n27563), .A3(n27562), .Z(n27565) );
  XNOR2HSV1 U29295 ( .A1(n27566), .A2(n27565), .ZN(n27568) );
  NAND2HSV0 U29296 ( .A1(n27719), .A2(n28702), .ZN(n27567) );
  XOR2HSV0 U29297 ( .A1(n27568), .A2(n27567), .Z(n27569) );
  XOR2HSV0 U29298 ( .A1(n27570), .A2(n27569), .Z(n27575) );
  NAND2HSV0 U29299 ( .A1(n27727), .A2(\pe2/got [8]), .ZN(n27573) );
  XOR3HSV2 U29300 ( .A1(n27575), .A2(n27574), .A3(n27573), .Z(\pe2/poht [8])
         );
  CLKNAND2HSV0 U29301 ( .A1(n28590), .A2(\pe2/got [8]), .ZN(n27609) );
  NAND2HSV0 U29302 ( .A1(n27657), .A2(n14003), .ZN(n27605) );
  NAND2HSV0 U29303 ( .A1(n27614), .A2(n14052), .ZN(n27600) );
  XOR2HSV0 U29304 ( .A1(n27577), .A2(n27576), .Z(n27593) );
  NAND2HSV0 U29305 ( .A1(\pe2/aot [9]), .A2(\pe2/bq[2] ), .ZN(n27579) );
  NAND2HSV0 U29306 ( .A1(\pe2/aot [1]), .A2(\pe2/bq[10] ), .ZN(n27578) );
  XOR2HSV0 U29307 ( .A1(n27579), .A2(n27578), .Z(n27584) );
  NOR2HSV0 U29308 ( .A1(n27580), .A2(n27692), .ZN(n27582) );
  NAND2HSV0 U29309 ( .A1(\pe2/aot [3]), .A2(\pe2/bq[8] ), .ZN(n27581) );
  XOR2HSV0 U29310 ( .A1(n27582), .A2(n27581), .Z(n27583) );
  XNOR2HSV1 U29311 ( .A1(n27584), .A2(n27583), .ZN(n27592) );
  NAND2HSV0 U29312 ( .A1(\pe2/aot [5]), .A2(\pe2/bq[6] ), .ZN(n27586) );
  NAND2HSV0 U29313 ( .A1(\pe2/aot [4]), .A2(\pe2/bq[7] ), .ZN(n27585) );
  XOR2HSV0 U29314 ( .A1(n27586), .A2(n27585), .Z(n27590) );
  NAND2HSV0 U29315 ( .A1(\pe2/aot [8]), .A2(\pe2/bq[3] ), .ZN(n27588) );
  NAND2HSV0 U29316 ( .A1(\pe2/aot [6]), .A2(\pe2/bq[5] ), .ZN(n27587) );
  XOR2HSV0 U29317 ( .A1(n27588), .A2(n27587), .Z(n27589) );
  XOR2HSV0 U29318 ( .A1(n27590), .A2(n27589), .Z(n27591) );
  XOR3HSV2 U29319 ( .A1(n27593), .A2(n27592), .A3(n27591), .Z(n27598) );
  NOR2HSV2 U29320 ( .A1(n27594), .A2(n27677), .ZN(n27597) );
  NOR2HSV1 U29321 ( .A1(n27595), .A2(n27735), .ZN(n27596) );
  XOR3HSV2 U29322 ( .A1(n27598), .A2(n27597), .A3(n27596), .Z(n27599) );
  XNOR2HSV1 U29323 ( .A1(n27600), .A2(n27599), .ZN(n27603) );
  NOR2HSV2 U29324 ( .A1(n27678), .A2(n27718), .ZN(n27602) );
  CLKNAND2HSV1 U29325 ( .A1(n27679), .A2(n27719), .ZN(n27601) );
  XOR3HSV2 U29326 ( .A1(n27603), .A2(n27602), .A3(n27601), .Z(n27604) );
  XNOR2HSV1 U29327 ( .A1(n27605), .A2(n27604), .ZN(n27607) );
  NAND2HSV0 U29328 ( .A1(n28702), .A2(n14046), .ZN(n27606) );
  XOR2HSV0 U29329 ( .A1(n27607), .A2(n27606), .Z(n27608) );
  XOR2HSV0 U29330 ( .A1(n27609), .A2(n27608), .Z(n27613) );
  NOR2HSV2 U29331 ( .A1(n27646), .A2(n27610), .ZN(n27612) );
  NAND2HSV0 U29332 ( .A1(n27727), .A2(\pe2/got [10]), .ZN(n27611) );
  XOR3HSV2 U29333 ( .A1(n27613), .A2(n27612), .A3(n27611), .Z(\pe2/poht [6])
         );
  NAND2HSV0 U29334 ( .A1(n28590), .A2(n14046), .ZN(n27644) );
  NAND2HSV0 U29335 ( .A1(n27667), .A2(n27719), .ZN(n27639) );
  NAND2HSV0 U29336 ( .A1(n27614), .A2(\pe2/got [2]), .ZN(n27632) );
  NAND2HSV0 U29337 ( .A1(n28617), .A2(n14055), .ZN(n27630) );
  NAND2HSV0 U29338 ( .A1(\pe2/aot [6]), .A2(\pe2/bq[4] ), .ZN(n27653) );
  NAND2HSV0 U29339 ( .A1(\pe2/aot [5]), .A2(\pe2/bq[5] ), .ZN(n27615) );
  XOR2HSV0 U29340 ( .A1(n27653), .A2(n27615), .Z(n27628) );
  CLKNAND2HSV0 U29341 ( .A1(\pe2/aot [4]), .A2(\pe2/bq[1] ), .ZN(n27695) );
  AO22HSV2 U29342 ( .A1(\pe2/aot [9]), .A2(\pe2/bq[1] ), .B1(\pe2/bq[6] ), 
        .B2(\pe2/aot [4]), .Z(n27616) );
  OAI21HSV0 U29343 ( .A1(n27695), .A2(n27617), .B(n27616), .ZN(n27619) );
  XOR2HSV0 U29344 ( .A1(n27619), .A2(n27618), .Z(n27627) );
  NAND2HSV0 U29345 ( .A1(\pe2/aot [1]), .A2(\pe2/bq[9] ), .ZN(n27621) );
  NAND2HSV0 U29346 ( .A1(\pe2/aot [3]), .A2(\pe2/bq[7] ), .ZN(n27620) );
  XOR2HSV0 U29347 ( .A1(n27621), .A2(n27620), .Z(n27625) );
  NAND2HSV0 U29348 ( .A1(\pe2/aot [2]), .A2(\pe2/bq[8] ), .ZN(n27623) );
  NAND2HSV0 U29349 ( .A1(\pe2/aot [8]), .A2(\pe2/bq[2] ), .ZN(n27622) );
  XOR2HSV0 U29350 ( .A1(n27623), .A2(n27622), .Z(n27624) );
  XOR2HSV0 U29351 ( .A1(n27625), .A2(n27624), .Z(n27626) );
  XOR3HSV2 U29352 ( .A1(n27628), .A2(n27627), .A3(n27626), .Z(n27629) );
  XNOR2HSV1 U29353 ( .A1(n27630), .A2(n27629), .ZN(n27631) );
  XNOR2HSV1 U29354 ( .A1(n27632), .A2(n27631), .ZN(n27637) );
  NOR2HSV2 U29355 ( .A1(n27634), .A2(n27633), .ZN(n27636) );
  CLKNAND2HSV0 U29356 ( .A1(n28474), .A2(n28634), .ZN(n27635) );
  XOR3HSV2 U29357 ( .A1(n27637), .A2(n27636), .A3(n27635), .Z(n27638) );
  XNOR2HSV1 U29358 ( .A1(n27639), .A2(n27638), .ZN(n27642) );
  NAND2HSV0 U29359 ( .A1(n27640), .A2(n14003), .ZN(n27641) );
  XOR2HSV0 U29360 ( .A1(n27642), .A2(n27641), .Z(n27643) );
  XOR2HSV0 U29361 ( .A1(n27644), .A2(n27643), .Z(n27650) );
  NOR2HSV2 U29362 ( .A1(n12302), .A2(n27645), .ZN(n27649) );
  CLKNAND2HSV1 U29363 ( .A1(n27736), .A2(n27647), .ZN(n27648) );
  XOR3HSV2 U29364 ( .A1(n27650), .A2(n27649), .A3(n27648), .Z(\pe2/poht [7])
         );
  NAND2HSV2 U29365 ( .A1(n27705), .A2(n28634), .ZN(n27662) );
  CLKNAND2HSV0 U29366 ( .A1(n28474), .A2(n14055), .ZN(n27656) );
  CLKNAND2HSV0 U29367 ( .A1(\pe2/aot [5]), .A2(\pe2/bq[3] ), .ZN(n27711) );
  NAND2HSV2 U29368 ( .A1(\pe2/aot [3]), .A2(\pe2/bq[1] ), .ZN(n27734) );
  XOR2HSV0 U29369 ( .A1(n27656), .A2(n27655), .Z(n27660) );
  CLKNAND2HSV1 U29370 ( .A1(n27657), .A2(\pe2/got [2]), .ZN(n27659) );
  XNOR3HSV1 U29371 ( .A1(n27660), .A2(n27659), .A3(n27658), .ZN(n27661) );
  XNOR2HSV1 U29372 ( .A1(n27662), .A2(n27661), .ZN(n27666) );
  NAND2HSV0 U29373 ( .A1(n27736), .A2(n14003), .ZN(n27664) );
  XOR3HSV2 U29374 ( .A1(n27666), .A2(n27665), .A3(n27664), .Z(\pe2/poht [10])
         );
  NAND2HSV2 U29375 ( .A1(n27691), .A2(n27719), .ZN(n27685) );
  NAND2HSV0 U29376 ( .A1(n27667), .A2(n14052), .ZN(n27681) );
  NAND2HSV0 U29377 ( .A1(\pe2/aot [2]), .A2(n27668), .ZN(n27670) );
  NAND2HSV0 U29378 ( .A1(\pe2/aot [6]), .A2(\pe2/bq[2] ), .ZN(n27669) );
  NAND2HSV0 U29379 ( .A1(\pe2/aot [4]), .A2(\pe2/bq[4] ), .ZN(n27707) );
  NAND2HSV0 U29380 ( .A1(\pe2/aot [3]), .A2(\pe2/bq[5] ), .ZN(n27671) );
  NAND2HSV0 U29381 ( .A1(\pe2/aot [1]), .A2(\pe2/bq[7] ), .ZN(n27674) );
  AOI22HSV0 U29382 ( .A1(n27675), .A2(n27674), .B1(n27673), .B2(n27672), .ZN(
        n27676) );
  XNOR2HSV1 U29383 ( .A1(n27681), .A2(n27680), .ZN(n27683) );
  NAND2HSV0 U29384 ( .A1(n28702), .A2(n28634), .ZN(n27682) );
  XOR2HSV0 U29385 ( .A1(n27683), .A2(n27682), .Z(n27684) );
  XNOR2HSV1 U29386 ( .A1(n27685), .A2(n27684), .ZN(n27690) );
  CLKNAND2HSV1 U29387 ( .A1(n28701), .A2(n14003), .ZN(n27688) );
  XOR3HSV2 U29388 ( .A1(n27690), .A2(n27689), .A3(n27688), .Z(\pe2/poht [9])
         );
  NAND2HSV2 U29389 ( .A1(n27705), .A2(\pe2/got [2]), .ZN(n27701) );
  CLKNAND2HSV1 U29390 ( .A1(n28702), .A2(n14055), .ZN(n27699) );
  NAND2HSV0 U29391 ( .A1(\pe2/aot [2]), .A2(\pe2/bq[3] ), .ZN(n27694) );
  XOR2HSV0 U29392 ( .A1(n27695), .A2(n27694), .Z(n27696) );
  XOR2HSV0 U29393 ( .A1(n27697), .A2(n27696), .Z(n27698) );
  XNOR2HSV1 U29394 ( .A1(n27699), .A2(n27698), .ZN(n27700) );
  XOR2HSV0 U29395 ( .A1(n27701), .A2(n27700), .Z(n27704) );
  NAND2HSV2 U29396 ( .A1(n28701), .A2(n14052), .ZN(n27703) );
  NAND2HSV0 U29397 ( .A1(n27736), .A2(n28634), .ZN(n27702) );
  XOR3HSV2 U29398 ( .A1(n27704), .A2(n27703), .A3(n27702), .Z(\pe2/poht [12])
         );
  NAND2HSV2 U29399 ( .A1(n27705), .A2(n14052), .ZN(n27717) );
  CLKNAND2HSV0 U29400 ( .A1(n27657), .A2(n14055), .ZN(n27712) );
  XOR2HSV0 U29401 ( .A1(n27713), .A2(n27712), .Z(n27715) );
  NAND2HSV0 U29402 ( .A1(n28702), .A2(\pe2/got [2]), .ZN(n27714) );
  XOR2HSV0 U29403 ( .A1(n27715), .A2(n27714), .Z(n27716) );
  XOR2HSV0 U29404 ( .A1(n27717), .A2(n27716), .Z(n27722) );
  NAND2HSV0 U29405 ( .A1(n27736), .A2(n27719), .ZN(n27720) );
  XOR3HSV2 U29406 ( .A1(n27722), .A2(n27721), .A3(n27720), .Z(\pe2/poht [11])
         );
  NAND2HSV0 U29407 ( .A1(\pe2/aot [1]), .A2(\pe2/bq[2] ), .ZN(n27725) );
  CLKNAND2HSV1 U29408 ( .A1(\pe2/aot [2]), .A2(n27723), .ZN(n27724) );
  XOR2HSV0 U29409 ( .A1(n27725), .A2(n27724), .Z(n27730) );
  NAND2HSV2 U29410 ( .A1(n27726), .A2(n14055), .ZN(n27729) );
  NAND2HSV0 U29411 ( .A1(n27736), .A2(\pe2/got [2]), .ZN(n27728) );
  XOR3HSV2 U29412 ( .A1(n27730), .A2(n27729), .A3(n27728), .Z(\pe2/poht [14])
         );
  NAND2HSV0 U29413 ( .A1(\pe2/aot [1]), .A2(\pe2/bq[3] ), .ZN(n27732) );
  NOR2HSV2 U29414 ( .A1(n27875), .A2(n27871), .ZN(n27783) );
  NOR2HSV2 U29415 ( .A1(n28001), .A2(n27826), .ZN(n27777) );
  NAND2HSV0 U29416 ( .A1(n28523), .A2(\pe4/got [8]), .ZN(n27775) );
  NOR2HSV0 U29417 ( .A1(n27942), .A2(n27969), .ZN(n27773) );
  NAND2HSV0 U29418 ( .A1(n22826), .A2(n27784), .ZN(n27738) );
  NAND2HSV0 U29419 ( .A1(n27957), .A2(\pe4/got [5]), .ZN(n27737) );
  XNOR2HSV1 U29420 ( .A1(n27738), .A2(n27737), .ZN(n27771) );
  NAND2HSV0 U29421 ( .A1(\pe4/ti_7[7] ), .A2(\pe4/got [4]), .ZN(n27769) );
  CLKNAND2HSV0 U29422 ( .A1(n28626), .A2(n22825), .ZN(n27767) );
  NAND2HSV0 U29423 ( .A1(n27830), .A2(n28591), .ZN(n27765) );
  NAND2HSV0 U29424 ( .A1(n27739), .A2(n28624), .ZN(n27763) );
  NAND2HSV0 U29425 ( .A1(\pe4/aot [3]), .A2(\pe4/bq[10] ), .ZN(n27741) );
  NAND2HSV0 U29426 ( .A1(\pe4/aot [2]), .A2(\pe4/bq[11] ), .ZN(n27740) );
  XOR2HSV0 U29427 ( .A1(n27741), .A2(n27740), .Z(n27745) );
  NAND2HSV0 U29428 ( .A1(\pe4/aot [8]), .A2(\pe4/bq[5] ), .ZN(n27743) );
  NAND2HSV0 U29429 ( .A1(\pe4/aot [9]), .A2(\pe4/bq[4] ), .ZN(n27742) );
  XOR2HSV0 U29430 ( .A1(n27743), .A2(n27742), .Z(n27744) );
  XOR2HSV0 U29431 ( .A1(n27745), .A2(n27744), .Z(n27754) );
  NAND2HSV0 U29432 ( .A1(\pe4/aot [1]), .A2(\pe4/bq[12] ), .ZN(n27747) );
  NAND2HSV0 U29433 ( .A1(\pe4/aot [7]), .A2(\pe4/bq[6] ), .ZN(n27746) );
  XOR2HSV0 U29434 ( .A1(n27747), .A2(n27746), .Z(n27752) );
  NOR2HSV0 U29435 ( .A1(n27748), .A2(n27886), .ZN(n27750) );
  AOI22HSV0 U29436 ( .A1(\pe4/aot [11]), .A2(\pe4/bq[2] ), .B1(\pe4/bq[7] ), 
        .B2(\pe4/aot [6]), .ZN(n27749) );
  NOR2HSV2 U29437 ( .A1(n27750), .A2(n27749), .ZN(n27751) );
  XNOR2HSV1 U29438 ( .A1(n27752), .A2(n27751), .ZN(n27753) );
  XNOR2HSV1 U29439 ( .A1(n27754), .A2(n27753), .ZN(n27761) );
  NAND2HSV0 U29440 ( .A1(\pe4/aot [5]), .A2(\pe4/bq[8] ), .ZN(n27756) );
  NAND2HSV0 U29441 ( .A1(\pe4/aot [12]), .A2(\pe4/bq[1] ), .ZN(n27755) );
  XOR2HSV0 U29442 ( .A1(n27756), .A2(n27755), .Z(n27759) );
  NAND2HSV0 U29443 ( .A1(\pe4/aot [10]), .A2(\pe4/bq[3] ), .ZN(n27840) );
  NAND2HSV0 U29444 ( .A1(\pe4/aot [4]), .A2(\pe4/bq[9] ), .ZN(n27757) );
  XOR2HSV0 U29445 ( .A1(n27840), .A2(n27757), .Z(n27758) );
  XOR2HSV0 U29446 ( .A1(n27759), .A2(n27758), .Z(n27760) );
  XNOR2HSV1 U29447 ( .A1(n27761), .A2(n27760), .ZN(n27762) );
  XNOR2HSV1 U29448 ( .A1(n27763), .A2(n27762), .ZN(n27764) );
  XNOR2HSV1 U29449 ( .A1(n27765), .A2(n27764), .ZN(n27766) );
  XNOR2HSV1 U29450 ( .A1(n27767), .A2(n27766), .ZN(n27768) );
  XNOR2HSV1 U29451 ( .A1(n27769), .A2(n27768), .ZN(n27770) );
  XNOR2HSV1 U29452 ( .A1(n27771), .A2(n27770), .ZN(n27772) );
  XOR2HSV0 U29453 ( .A1(n27773), .A2(n27772), .Z(n27774) );
  XNOR2HSV1 U29454 ( .A1(n27775), .A2(n27774), .ZN(n27776) );
  XOR2HSV0 U29455 ( .A1(n27777), .A2(n27776), .Z(n27778) );
  XOR2HSV0 U29456 ( .A1(n27779), .A2(n27778), .Z(n27782) );
  NOR2HSV0 U29457 ( .A1(n27900), .A2(n27780), .ZN(n27781) );
  XOR3HSV2 U29458 ( .A1(n27783), .A2(n27782), .A3(n27781), .Z(\pe4/poht [4])
         );
  NOR2HSV2 U29459 ( .A1(n27875), .A2(n27826), .ZN(n27824) );
  CLKAND2HSV2 U29460 ( .A1(n27940), .A2(\pe4/got [8]), .Z(n27821) );
  NOR2HSV2 U29461 ( .A1(n27979), .A2(n27969), .ZN(n27819) );
  NAND2HSV0 U29462 ( .A1(n27784), .A2(\pe4/got [4]), .ZN(n27786) );
  NAND2HSV0 U29463 ( .A1(n28578), .A2(n28626), .ZN(n27785) );
  XNOR2HSV1 U29464 ( .A1(n27786), .A2(n27785), .ZN(n27806) );
  NAND2HSV0 U29465 ( .A1(\pe4/ti_7[7] ), .A2(n28591), .ZN(n27804) );
  CLKNAND2HSV0 U29466 ( .A1(n22825), .A2(n28624), .ZN(n27802) );
  NAND2HSV0 U29467 ( .A1(\pe4/aot [5]), .A2(\pe4/bq[6] ), .ZN(n27788) );
  NAND2HSV0 U29468 ( .A1(\pe4/aot [8]), .A2(\pe4/bq[3] ), .ZN(n27787) );
  XOR2HSV0 U29469 ( .A1(n27788), .A2(n27787), .Z(n27792) );
  NAND2HSV0 U29470 ( .A1(\pe4/aot [1]), .A2(\pe4/bq[10] ), .ZN(n27790) );
  NAND2HSV0 U29471 ( .A1(\pe4/aot [4]), .A2(\pe4/bq[7] ), .ZN(n27789) );
  XOR2HSV0 U29472 ( .A1(n27790), .A2(n27789), .Z(n27791) );
  XOR2HSV0 U29473 ( .A1(n27792), .A2(n27791), .Z(n27800) );
  IOA22HSV1 U29474 ( .B1(n27847), .B2(n27793), .A1(\pe4/aot [2]), .A2(
        \pe4/bq[9] ), .ZN(n27794) );
  OAI21HSV1 U29475 ( .A1(n27796), .A2(n27795), .B(n27794), .ZN(n27798) );
  NAND2HSV0 U29476 ( .A1(\pe4/aot [3]), .A2(\pe4/bq[8] ), .ZN(n27797) );
  XNOR2HSV1 U29477 ( .A1(n27798), .A2(n27797), .ZN(n27799) );
  XNOR2HSV1 U29478 ( .A1(n27800), .A2(n27799), .ZN(n27801) );
  XOR2HSV0 U29479 ( .A1(n27802), .A2(n27801), .Z(n27803) );
  XOR2HSV0 U29480 ( .A1(n27804), .A2(n27803), .Z(n27805) );
  XNOR2HSV1 U29481 ( .A1(n27806), .A2(n27805), .ZN(n27808) );
  CLKNHSV0 U29482 ( .I(n27808), .ZN(n27807) );
  OAI21HSV0 U29483 ( .A1(n27876), .A2(n21997), .B(n27807), .ZN(n27810) );
  NAND3HSV0 U29484 ( .A1(n28583), .A2(\pe4/got [5]), .A3(n27808), .ZN(n27809)
         );
  CLKNAND2HSV1 U29485 ( .A1(n27810), .A2(n27809), .ZN(n27815) );
  NAND2HSV0 U29486 ( .A1(\pe4/aot [7]), .A2(\pe4/bq[4] ), .ZN(n27812) );
  NAND2HSV0 U29487 ( .A1(\pe4/aot [10]), .A2(\pe4/bq[1] ), .ZN(n27811) );
  XOR2HSV0 U29488 ( .A1(n27812), .A2(n27811), .Z(n27813) );
  XNOR2HSV1 U29489 ( .A1(n27813), .A2(n27841), .ZN(n27814) );
  NAND2HSV0 U29490 ( .A1(n22826), .A2(n14038), .ZN(n27816) );
  XNOR2HSV4 U29491 ( .A1(n27821), .A2(n27820), .ZN(n27823) );
  NOR2HSV0 U29492 ( .A1(n27900), .A2(n27825), .ZN(n27822) );
  XOR3HSV2 U29493 ( .A1(n27824), .A2(n27823), .A3(n27822), .Z(\pe4/poht [6])
         );
  NOR2HSV2 U29494 ( .A1(n27875), .A2(n27825), .ZN(n27874) );
  NOR2HSV2 U29495 ( .A1(n27977), .A2(n27826), .ZN(n27870) );
  NOR2HSV2 U29496 ( .A1(n27906), .A2(n27827), .ZN(n27868) );
  NAND2HSV0 U29497 ( .A1(n14038), .A2(n13996), .ZN(n27866) );
  NOR2HSV0 U29498 ( .A1(n27876), .A2(n27905), .ZN(n27864) );
  NAND2HSV0 U29499 ( .A1(\pe4/got [5]), .A2(n27877), .ZN(n27829) );
  NAND2HSV0 U29500 ( .A1(n28578), .A2(\pe4/got [4]), .ZN(n27828) );
  XNOR2HSV1 U29501 ( .A1(n27829), .A2(n27828), .ZN(n27862) );
  NAND2HSV0 U29502 ( .A1(\pe4/ti_7[7] ), .A2(n28626), .ZN(n27860) );
  NAND2HSV0 U29503 ( .A1(n22825), .A2(n28591), .ZN(n27858) );
  NAND2HSV0 U29504 ( .A1(n28624), .A2(n27830), .ZN(n27856) );
  NOR2HSV0 U29505 ( .A1(n27832), .A2(n27831), .ZN(n27834) );
  AOI22HSV0 U29506 ( .A1(\pe4/aot [11]), .A2(\pe4/bq[1] ), .B1(\pe4/bq[10] ), 
        .B2(\pe4/aot [2]), .ZN(n27833) );
  NOR2HSV2 U29507 ( .A1(n27834), .A2(n27833), .ZN(n27836) );
  NAND2HSV0 U29508 ( .A1(\pe4/aot [8]), .A2(\pe4/bq[4] ), .ZN(n27835) );
  XNOR2HSV1 U29509 ( .A1(n27836), .A2(n27835), .ZN(n27854) );
  NAND2HSV0 U29510 ( .A1(\pe4/aot [5]), .A2(\pe4/bq[7] ), .ZN(n27838) );
  NAND2HSV0 U29511 ( .A1(\pe4/aot [3]), .A2(\pe4/bq[9] ), .ZN(n27837) );
  XOR2HSV0 U29512 ( .A1(n27838), .A2(n27837), .Z(n27843) );
  AO22HSV2 U29513 ( .A1(\pe4/aot [10]), .A2(\pe4/bq[2] ), .B1(\pe4/aot [9]), 
        .B2(\pe4/bq[3] ), .Z(n27839) );
  OAI21HSV0 U29514 ( .A1(n27841), .A2(n27840), .B(n27839), .ZN(n27842) );
  XNOR2HSV1 U29515 ( .A1(n27843), .A2(n27842), .ZN(n27853) );
  NAND2HSV0 U29516 ( .A1(\pe4/aot [1]), .A2(\pe4/bq[11] ), .ZN(n27845) );
  NAND2HSV0 U29517 ( .A1(\pe4/aot [7]), .A2(\pe4/bq[5] ), .ZN(n27844) );
  XOR2HSV0 U29518 ( .A1(n27845), .A2(n27844), .Z(n27851) );
  NOR2HSV0 U29519 ( .A1(n27847), .A2(n27846), .ZN(n27849) );
  NAND2HSV0 U29520 ( .A1(\pe4/aot [4]), .A2(\pe4/bq[8] ), .ZN(n27848) );
  XOR2HSV0 U29521 ( .A1(n27849), .A2(n27848), .Z(n27850) );
  XOR2HSV0 U29522 ( .A1(n27851), .A2(n27850), .Z(n27852) );
  XOR3HSV2 U29523 ( .A1(n27854), .A2(n27853), .A3(n27852), .Z(n27855) );
  XNOR2HSV1 U29524 ( .A1(n27856), .A2(n27855), .ZN(n27857) );
  XNOR2HSV1 U29525 ( .A1(n27858), .A2(n27857), .ZN(n27859) );
  XNOR2HSV1 U29526 ( .A1(n27860), .A2(n27859), .ZN(n27861) );
  XNOR2HSV1 U29527 ( .A1(n27862), .A2(n27861), .ZN(n27863) );
  XOR2HSV0 U29528 ( .A1(n27864), .A2(n27863), .Z(n27865) );
  XNOR2HSV1 U29529 ( .A1(n27866), .A2(n27865), .ZN(n27867) );
  NOR2HSV0 U29530 ( .A1(n27900), .A2(n27871), .ZN(n27872) );
  XOR3HSV2 U29531 ( .A1(n27874), .A2(n27873), .A3(n27872), .Z(\pe4/poht [5])
         );
  NOR2HSV2 U29532 ( .A1(n27875), .A2(n27905), .ZN(n27903) );
  NOR2HSV2 U29533 ( .A1(n27977), .A2(n21997), .ZN(n27899) );
  NOR2HSV2 U29534 ( .A1(n27979), .A2(n27973), .ZN(n27897) );
  NAND2HSV0 U29535 ( .A1(n28626), .A2(n14038), .ZN(n27895) );
  NOR2HSV0 U29536 ( .A1(n27876), .A2(n27978), .ZN(n27893) );
  NAND2HSV0 U29537 ( .A1(n27877), .A2(n28624), .ZN(n27891) );
  NAND2HSV0 U29538 ( .A1(\pe4/aot [1]), .A2(\pe4/bq[7] ), .ZN(n27879) );
  NAND2HSV0 U29539 ( .A1(\pe4/aot [5]), .A2(\pe4/bq[3] ), .ZN(n27878) );
  XOR2HSV0 U29540 ( .A1(n27879), .A2(n27878), .Z(n27883) );
  NAND2HSV0 U29541 ( .A1(\pe4/aot [7]), .A2(\pe4/bq[1] ), .ZN(n27881) );
  NAND2HSV0 U29542 ( .A1(\pe4/aot [3]), .A2(\pe4/bq[5] ), .ZN(n27880) );
  XOR2HSV0 U29543 ( .A1(n27881), .A2(n27880), .Z(n27882) );
  XOR2HSV0 U29544 ( .A1(n27883), .A2(n27882), .Z(n27889) );
  NAND2HSV0 U29545 ( .A1(\pe4/aot [4]), .A2(\pe4/bq[4] ), .ZN(n27885) );
  NAND2HSV0 U29546 ( .A1(\pe4/aot [2]), .A2(\pe4/bq[6] ), .ZN(n27884) );
  XOR2HSV0 U29547 ( .A1(n27885), .A2(n27884), .Z(n27887) );
  XNOR2HSV1 U29548 ( .A1(n27887), .A2(n27886), .ZN(n27888) );
  XNOR2HSV1 U29549 ( .A1(n27889), .A2(n27888), .ZN(n27890) );
  XOR2HSV0 U29550 ( .A1(n27891), .A2(n27890), .Z(n27892) );
  XOR2HSV0 U29551 ( .A1(n27893), .A2(n27892), .Z(n27894) );
  XOR2HSV0 U29552 ( .A1(n27895), .A2(n27894), .Z(n27896) );
  NOR2HSV0 U29553 ( .A1(n27900), .A2(n27969), .ZN(n27901) );
  XOR3HSV2 U29554 ( .A1(n27903), .A2(n27902), .A3(n27901), .Z(\pe4/poht [9])
         );
  AND2HSV2 U29555 ( .A1(n27904), .A2(\pe4/got [8]), .Z(n27939) );
  NOR2HSV2 U29556 ( .A1(n27906), .A2(n27905), .ZN(n27934) );
  NAND2HSV0 U29557 ( .A1(n14038), .A2(\pe4/got [5]), .ZN(n27932) );
  NOR2HSV0 U29558 ( .A1(n27942), .A2(n27973), .ZN(n27930) );
  NAND2HSV0 U29559 ( .A1(n27784), .A2(n28626), .ZN(n27909) );
  NAND2HSV0 U29560 ( .A1(n28578), .A2(n28591), .ZN(n27908) );
  XNOR2HSV1 U29561 ( .A1(n27909), .A2(n27908), .ZN(n27928) );
  NAND2HSV0 U29562 ( .A1(\pe4/ti_7[7] ), .A2(n28624), .ZN(n27926) );
  NAND2HSV0 U29563 ( .A1(\pe4/aot [6]), .A2(\pe4/bq[4] ), .ZN(n27911) );
  NAND2HSV0 U29564 ( .A1(\pe4/aot [8]), .A2(\pe4/bq[2] ), .ZN(n27910) );
  XOR2HSV0 U29565 ( .A1(n27911), .A2(n27910), .Z(n27924) );
  NAND2HSV0 U29566 ( .A1(\pe4/aot [4]), .A2(\pe4/bq[6] ), .ZN(n27913) );
  NAND2HSV0 U29567 ( .A1(\pe4/aot [2]), .A2(\pe4/bq[8] ), .ZN(n27912) );
  XOR2HSV0 U29568 ( .A1(n27913), .A2(n27912), .Z(n27915) );
  NAND2HSV0 U29569 ( .A1(\pe4/aot [1]), .A2(\pe4/bq[9] ), .ZN(n27914) );
  XNOR2HSV1 U29570 ( .A1(n27915), .A2(n27914), .ZN(n27923) );
  NAND2HSV0 U29571 ( .A1(\pe4/aot [9]), .A2(\pe4/bq[1] ), .ZN(n27917) );
  NAND2HSV0 U29572 ( .A1(\pe4/aot [5]), .A2(\pe4/bq[5] ), .ZN(n27916) );
  XOR2HSV0 U29573 ( .A1(n27917), .A2(n27916), .Z(n27921) );
  NAND2HSV0 U29574 ( .A1(\pe4/aot [7]), .A2(\pe4/bq[3] ), .ZN(n27919) );
  NAND2HSV0 U29575 ( .A1(\pe4/aot [3]), .A2(\pe4/bq[7] ), .ZN(n27918) );
  XOR2HSV0 U29576 ( .A1(n27919), .A2(n27918), .Z(n27920) );
  XOR2HSV0 U29577 ( .A1(n27921), .A2(n27920), .Z(n27922) );
  XOR3HSV2 U29578 ( .A1(n27924), .A2(n27923), .A3(n27922), .Z(n27925) );
  XNOR2HSV1 U29579 ( .A1(n27926), .A2(n27925), .ZN(n27927) );
  XNOR2HSV1 U29580 ( .A1(n27928), .A2(n27927), .ZN(n27929) );
  XOR2HSV0 U29581 ( .A1(n27930), .A2(n27929), .Z(n27931) );
  XNOR2HSV1 U29582 ( .A1(n27932), .A2(n27931), .ZN(n27933) );
  XOR2HSV0 U29583 ( .A1(n27934), .A2(n27933), .Z(n27935) );
  XOR2HSV2 U29584 ( .A1(n27936), .A2(n27935), .Z(n27938) );
  NAND2HSV0 U29585 ( .A1(n28012), .A2(\pe4/got [9]), .ZN(n27937) );
  XOR3HSV2 U29586 ( .A1(n27939), .A2(n27938), .A3(n27937), .Z(\pe4/poht [7])
         );
  NAND2HSV2 U29587 ( .A1(\pe4/got [6]), .A2(n27940), .ZN(n27968) );
  NAND2HSV0 U29588 ( .A1(\pe4/got [4]), .A2(n14080), .ZN(n27964) );
  NOR2HSV0 U29589 ( .A1(n27942), .A2(n27998), .ZN(n27962) );
  NAND2HSV0 U29590 ( .A1(\pe4/aot [7]), .A2(\pe4/bq[2] ), .ZN(n27944) );
  NAND2HSV0 U29591 ( .A1(\pe4/aot [1]), .A2(\pe4/bq[8] ), .ZN(n27943) );
  XOR2HSV0 U29592 ( .A1(n27944), .A2(n27943), .Z(n27948) );
  NAND2HSV0 U29593 ( .A1(\pe4/aot [4]), .A2(\pe4/bq[5] ), .ZN(n27946) );
  NAND2HSV0 U29594 ( .A1(\pe4/aot [5]), .A2(\pe4/bq[4] ), .ZN(n27945) );
  XOR2HSV0 U29595 ( .A1(n27946), .A2(n27945), .Z(n27947) );
  XOR2HSV0 U29596 ( .A1(n27948), .A2(n27947), .Z(n27956) );
  NAND2HSV0 U29597 ( .A1(\pe4/aot [8]), .A2(\pe4/bq[1] ), .ZN(n27950) );
  NAND2HSV0 U29598 ( .A1(\pe4/aot [2]), .A2(\pe4/bq[7] ), .ZN(n27949) );
  XOR2HSV0 U29599 ( .A1(n27950), .A2(n27949), .Z(n27954) );
  NAND2HSV0 U29600 ( .A1(\pe4/aot [3]), .A2(\pe4/bq[6] ), .ZN(n27952) );
  NAND2HSV0 U29601 ( .A1(\pe4/aot [6]), .A2(\pe4/bq[3] ), .ZN(n27951) );
  XOR2HSV0 U29602 ( .A1(n27952), .A2(n27951), .Z(n27953) );
  XOR2HSV0 U29603 ( .A1(n27954), .A2(n27953), .Z(n27955) );
  XOR2HSV0 U29604 ( .A1(n27956), .A2(n27955), .Z(n27960) );
  NAND2HSV2 U29605 ( .A1(n27957), .A2(n28624), .ZN(n27959) );
  NAND2HSV0 U29606 ( .A1(n27784), .A2(\pe4/got [2]), .ZN(n27958) );
  XOR3HSV2 U29607 ( .A1(n27960), .A2(n27959), .A3(n27958), .Z(n27961) );
  XOR2HSV0 U29608 ( .A1(n27962), .A2(n27961), .Z(n27963) );
  XNOR2HSV1 U29609 ( .A1(n27964), .A2(n27963), .ZN(n27965) );
  XOR2HSV0 U29610 ( .A1(n27966), .A2(n27965), .Z(n27967) );
  OR2HSV1 U29611 ( .A1(n27999), .A2(n27969), .Z(n27971) );
  NAND2HSV0 U29612 ( .A1(n28012), .A2(\pe4/got [8]), .ZN(n27970) );
  XOR3HSV2 U29613 ( .A1(n27972), .A2(n27971), .A3(n27970), .Z(\pe4/poht [8])
         );
  NOR2HSV1 U29614 ( .A1(n27974), .A2(n27973), .ZN(n27975) );
  NOR2HSV2 U29615 ( .A1(n27977), .A2(n27998), .ZN(n27994) );
  NOR2HSV2 U29616 ( .A1(n27979), .A2(n27978), .ZN(n27992) );
  NAND2HSV0 U29617 ( .A1(n28624), .A2(n14038), .ZN(n27990) );
  NAND2HSV0 U29618 ( .A1(\pe4/aot [1]), .A2(\pe4/bq[5] ), .ZN(n27982) );
  NAND2HSV0 U29619 ( .A1(\pe4/aot [2]), .A2(\pe4/bq[4] ), .ZN(n27981) );
  XOR2HSV0 U29620 ( .A1(n27982), .A2(n27981), .Z(n27984) );
  XNOR2HSV1 U29621 ( .A1(n27984), .A2(n27983), .ZN(n27988) );
  NAND2HSV0 U29622 ( .A1(\pe4/aot [3]), .A2(\pe4/bq[3] ), .ZN(n27986) );
  NAND2HSV0 U29623 ( .A1(\pe4/aot [4]), .A2(\pe4/bq[2] ), .ZN(n27985) );
  XOR2HSV0 U29624 ( .A1(n27986), .A2(n27985), .Z(n27987) );
  XNOR2HSV1 U29625 ( .A1(n27988), .A2(n27987), .ZN(n27989) );
  XNOR2HSV1 U29626 ( .A1(n27990), .A2(n27989), .ZN(n27991) );
  XOR2HSV0 U29627 ( .A1(n27992), .A2(n27991), .Z(n27993) );
  XNOR2HSV4 U29628 ( .A1(n27994), .A2(n27993), .ZN(n27996) );
  NAND2HSV2 U29629 ( .A1(n28461), .A2(\pe4/got [5]), .ZN(n27995) );
  XOR3HSV2 U29630 ( .A1(n27997), .A2(n27996), .A3(n27995), .Z(\pe4/poht [11])
         );
  NOR2HSV2 U29631 ( .A1(n27999), .A2(n27998), .ZN(n28015) );
  CLKNAND2HSV1 U29632 ( .A1(n28480), .A2(\pe4/got [2]), .ZN(n28011) );
  NOR2HSV2 U29633 ( .A1(n28001), .A2(n28000), .ZN(n28009) );
  NAND2HSV0 U29634 ( .A1(\pe4/aot [1]), .A2(\pe4/bq[4] ), .ZN(n28003) );
  NAND2HSV0 U29635 ( .A1(\pe4/aot [4]), .A2(\pe4/bq[1] ), .ZN(n28002) );
  XOR2HSV0 U29636 ( .A1(n28003), .A2(n28002), .Z(n28007) );
  NAND2HSV0 U29637 ( .A1(\pe4/aot [3]), .A2(\pe4/bq[2] ), .ZN(n28005) );
  NAND2HSV0 U29638 ( .A1(\pe4/aot [2]), .A2(\pe4/bq[3] ), .ZN(n28004) );
  XOR2HSV0 U29639 ( .A1(n28005), .A2(n28004), .Z(n28006) );
  XOR2HSV0 U29640 ( .A1(n28007), .A2(n28006), .Z(n28008) );
  XOR2HSV0 U29641 ( .A1(n28009), .A2(n28008), .Z(n28010) );
  XOR2HSV0 U29642 ( .A1(n28011), .A2(n28010), .Z(n28014) );
  XOR3HSV2 U29643 ( .A1(n28015), .A2(n28014), .A3(n28013), .Z(\pe4/poht [12])
         );
  NOR2HSV0 U29644 ( .A1(n28146), .A2(n28016), .ZN(n28075) );
  CLKNAND2HSV0 U29645 ( .A1(n28231), .A2(n28423), .ZN(n28073) );
  NAND2HSV0 U29646 ( .A1(n19767), .A2(n28227), .ZN(n28071) );
  NAND2HSV0 U29647 ( .A1(n28264), .A2(\pe9/got [8]), .ZN(n28066) );
  NAND2HSV0 U29648 ( .A1(n28110), .A2(n28405), .ZN(n28058) );
  NAND2HSV0 U29649 ( .A1(\pe9/aot [12]), .A2(\pe9/bq[5] ), .ZN(n28018) );
  NAND2HSV0 U29650 ( .A1(\pe9/aot [10]), .A2(\pe9/bq[7] ), .ZN(n28017) );
  XOR2HSV0 U29651 ( .A1(n28018), .A2(n28017), .Z(n28023) );
  NAND2HSV0 U29652 ( .A1(\pe9/bq[4] ), .A2(\pe9/aot [13]), .ZN(n28021) );
  NAND2HSV0 U29653 ( .A1(n28019), .A2(\pe9/got [1]), .ZN(n28020) );
  XOR2HSV0 U29654 ( .A1(n28021), .A2(n28020), .Z(n28022) );
  XOR2HSV0 U29655 ( .A1(n28023), .A2(n28022), .Z(n28032) );
  NAND2HSV0 U29656 ( .A1(\pe9/aot [6]), .A2(\pe9/bq[11] ), .ZN(n28025) );
  NAND2HSV0 U29657 ( .A1(\pe9/aot [14]), .A2(\pe9/bq[3] ), .ZN(n28024) );
  XOR2HSV0 U29658 ( .A1(n28025), .A2(n28024), .Z(n28030) );
  NOR2HSV0 U29659 ( .A1(n28398), .A2(n28026), .ZN(n28028) );
  NAND2HSV0 U29660 ( .A1(\pe9/aot [9]), .A2(\pe9/bq[8] ), .ZN(n28027) );
  XOR2HSV0 U29661 ( .A1(n28028), .A2(n28027), .Z(n28029) );
  XOR2HSV0 U29662 ( .A1(n28030), .A2(n28029), .Z(n28031) );
  XOR2HSV0 U29663 ( .A1(n28032), .A2(n28031), .Z(n28034) );
  NAND2HSV0 U29664 ( .A1(n28688), .A2(\pe9/got [2]), .ZN(n28033) );
  XNOR2HSV1 U29665 ( .A1(n28034), .A2(n28033), .ZN(n28055) );
  NAND2HSV0 U29666 ( .A1(\pe9/aot [11]), .A2(\pe9/bq[6] ), .ZN(n28148) );
  NAND2HSV0 U29667 ( .A1(\pe9/aot [3]), .A2(n23822), .ZN(n28035) );
  XOR2HSV0 U29668 ( .A1(n28148), .A2(n28035), .Z(n28053) );
  NAND2HSV0 U29669 ( .A1(n27093), .A2(\pe9/pq ), .ZN(n28037) );
  XOR2HSV0 U29670 ( .A1(n28037), .A2(n28036), .Z(n28043) );
  CLKNHSV0 U29671 ( .I(\pe9/aot [15]), .ZN(n28038) );
  NOR2HSV0 U29672 ( .A1(n28038), .A2(n28397), .ZN(n28040) );
  NAND2HSV0 U29673 ( .A1(\pe9/aot [5]), .A2(\pe9/bq[2] ), .ZN(n28359) );
  OAI22HSV0 U29674 ( .A1(n28041), .A2(n28040), .B1(n28039), .B2(n28359), .ZN(
        n28042) );
  XNOR2HSV1 U29675 ( .A1(n28043), .A2(n28042), .ZN(n28052) );
  NAND2HSV0 U29676 ( .A1(\pe9/aot [1]), .A2(n28044), .ZN(n28046) );
  NAND2HSV0 U29677 ( .A1(\pe9/aot [8]), .A2(\pe9/bq[9] ), .ZN(n28045) );
  XOR2HSV0 U29678 ( .A1(n28046), .A2(n28045), .Z(n28050) );
  NAND2HSV0 U29679 ( .A1(\pe9/aot [7]), .A2(\pe9/bq[10] ), .ZN(n28048) );
  NAND2HSV0 U29680 ( .A1(\pe9/aot [4]), .A2(\pe9/bq[13] ), .ZN(n28047) );
  XOR2HSV0 U29681 ( .A1(n28048), .A2(n28047), .Z(n28049) );
  XOR2HSV0 U29682 ( .A1(n28050), .A2(n28049), .Z(n28051) );
  XOR3HSV2 U29683 ( .A1(n28053), .A2(n28052), .A3(n28051), .Z(n28054) );
  XNOR2HSV1 U29684 ( .A1(n28055), .A2(n28054), .ZN(n28057) );
  NAND2HSV0 U29685 ( .A1(n28804), .A2(\pe9/got [4]), .ZN(n28056) );
  XOR3HSV2 U29686 ( .A1(n28058), .A2(n28057), .A3(n28056), .Z(n28061) );
  NAND2HSV0 U29687 ( .A1(n28059), .A2(n28643), .ZN(n28060) );
  XOR2HSV0 U29688 ( .A1(n28061), .A2(n28060), .Z(n28064) );
  NAND2HSV0 U29689 ( .A1(n28689), .A2(\pe9/got [7]), .ZN(n28063) );
  NAND2HSV0 U29690 ( .A1(n28638), .A2(\pe9/got [6]), .ZN(n28062) );
  XOR3HSV1 U29691 ( .A1(n28064), .A2(n28063), .A3(n28062), .Z(n28065) );
  XNOR2HSV1 U29692 ( .A1(n28066), .A2(n28065), .ZN(n28069) );
  OR2HSV1 U29693 ( .A1(n28214), .A2(n28067), .Z(n28068) );
  XNOR2HSV1 U29694 ( .A1(n28069), .A2(n28068), .ZN(n28070) );
  XNOR2HSV1 U29695 ( .A1(n28071), .A2(n28070), .ZN(n28072) );
  XNOR2HSV1 U29696 ( .A1(n28073), .A2(n28072), .ZN(n28074) );
  XOR2HSV0 U29697 ( .A1(n28075), .A2(n28074), .Z(n28077) );
  NAND2HSV0 U29698 ( .A1(n28580), .A2(n28137), .ZN(n28076) );
  XOR2HSV0 U29699 ( .A1(n28077), .A2(n28076), .Z(n28079) );
  NAND2HSV0 U29700 ( .A1(n28394), .A2(n28928), .ZN(n28078) );
  XNOR2HSV1 U29701 ( .A1(n28079), .A2(n28078), .ZN(n28084) );
  INHSV4 U29702 ( .I(n28141), .ZN(n28413) );
  NAND3HSV2 U29703 ( .A1(n28413), .A2(n14039), .A3(n28412), .ZN(n28083) );
  NAND2HSV2 U29704 ( .A1(n28390), .A2(n28081), .ZN(n28082) );
  XOR3HSV2 U29705 ( .A1(n28084), .A2(n28083), .A3(n28082), .Z(po9) );
  NOR2HSV2 U29706 ( .A1(n28316), .A2(n28085), .ZN(n28132) );
  CLKNAND2HSV0 U29707 ( .A1(n28231), .A2(n28227), .ZN(n28130) );
  NAND2HSV0 U29708 ( .A1(n28437), .A2(n14073), .ZN(n28128) );
  NAND2HSV0 U29709 ( .A1(n28264), .A2(\pe9/got [7]), .ZN(n28123) );
  NAND2HSV0 U29710 ( .A1(n28949), .A2(n28389), .ZN(n28118) );
  NAND2HSV0 U29711 ( .A1(n28804), .A2(\pe9/got [3]), .ZN(n28116) );
  NAND2HSV0 U29712 ( .A1(\pe9/aot [1]), .A2(\pe9/bq[15] ), .ZN(n28087) );
  NAND2HSV0 U29713 ( .A1(\pe9/aot [10]), .A2(\pe9/bq[6] ), .ZN(n28086) );
  XOR2HSV0 U29714 ( .A1(n28087), .A2(n28086), .Z(n28094) );
  NAND2HSV0 U29715 ( .A1(\pe9/aot [4]), .A2(\pe9/bq[12] ), .ZN(n28091) );
  NAND2HSV0 U29716 ( .A1(\pe9/aot [5]), .A2(\pe9/bq[11] ), .ZN(n28090) );
  XOR2HSV0 U29717 ( .A1(n28091), .A2(n28090), .Z(n28092) );
  XOR4HSV1 U29718 ( .A1(n28095), .A2(n28094), .A3(n28093), .A4(n28092), .Z(
        n28114) );
  NAND2HSV0 U29719 ( .A1(\pe9/aot [8]), .A2(\pe9/bq[8] ), .ZN(n28097) );
  NAND2HSV0 U29720 ( .A1(\pe9/aot [6]), .A2(\pe9/bq[10] ), .ZN(n28096) );
  XOR2HSV0 U29721 ( .A1(n28097), .A2(n28096), .Z(n28101) );
  NAND2HSV0 U29722 ( .A1(\pe9/bq[3] ), .A2(\pe9/aot [13]), .ZN(n28099) );
  NAND2HSV0 U29723 ( .A1(\pe9/aot [7]), .A2(\pe9/bq[9] ), .ZN(n28098) );
  XOR2HSV0 U29724 ( .A1(n28099), .A2(n28098), .Z(n28100) );
  XOR2HSV0 U29725 ( .A1(n28101), .A2(n28100), .Z(n28109) );
  NAND2HSV0 U29726 ( .A1(n14079), .A2(\pe9/bq[1] ), .ZN(n28103) );
  NAND2HSV0 U29727 ( .A1(\pe9/aot [9]), .A2(\pe9/bq[7] ), .ZN(n28102) );
  XOR2HSV0 U29728 ( .A1(n28103), .A2(n28102), .Z(n28107) );
  NAND2HSV0 U29729 ( .A1(\pe9/aot [12]), .A2(\pe9/bq[4] ), .ZN(n28105) );
  NAND2HSV0 U29730 ( .A1(\pe9/aot [3]), .A2(\pe9/bq[13] ), .ZN(n28104) );
  XOR2HSV0 U29731 ( .A1(n28105), .A2(n28104), .Z(n28106) );
  XOR2HSV0 U29732 ( .A1(n28107), .A2(n28106), .Z(n28108) );
  XOR2HSV0 U29733 ( .A1(n28109), .A2(n28108), .Z(n28113) );
  NAND2HSV0 U29734 ( .A1(n28688), .A2(n28658), .ZN(n28112) );
  NAND2HSV0 U29735 ( .A1(\pe9/got [2]), .A2(n28110), .ZN(n28111) );
  XOR4HSV1 U29736 ( .A1(n28114), .A2(n28113), .A3(n28112), .A4(n28111), .Z(
        n28115) );
  XNOR2HSV1 U29737 ( .A1(n28116), .A2(n28115), .ZN(n28117) );
  XOR2HSV0 U29738 ( .A1(n28118), .A2(n28117), .Z(n28121) );
  NAND2HSV0 U29739 ( .A1(n28189), .A2(\pe9/got [6]), .ZN(n28120) );
  NAND2HSV0 U29740 ( .A1(n28166), .A2(n28643), .ZN(n28119) );
  XOR3HSV1 U29741 ( .A1(n28121), .A2(n28120), .A3(n28119), .Z(n28122) );
  XNOR2HSV1 U29742 ( .A1(n28123), .A2(n28122), .ZN(n28126) );
  OR2HSV1 U29743 ( .A1(n28287), .A2(n28124), .Z(n28125) );
  XNOR2HSV1 U29744 ( .A1(n28126), .A2(n28125), .ZN(n28127) );
  XNOR2HSV1 U29745 ( .A1(n28128), .A2(n28127), .ZN(n28129) );
  XNOR2HSV1 U29746 ( .A1(n28130), .A2(n28129), .ZN(n28131) );
  XOR2HSV0 U29747 ( .A1(n28132), .A2(n28131), .Z(n28136) );
  CLKBUFHSV4 U29748 ( .I(n28133), .Z(n28383) );
  NAND2HSV0 U29749 ( .A1(n28383), .A2(n28134), .ZN(n28135) );
  CLKNAND2HSV0 U29750 ( .A1(n28475), .A2(n28137), .ZN(n28138) );
  XNOR2HSV1 U29751 ( .A1(n28139), .A2(n28138), .ZN(n28145) );
  INHSV2 U29752 ( .I(n28140), .ZN(n28141) );
  INHSV2 U29753 ( .I(n28184), .ZN(n28403) );
  NAND3HSV2 U29754 ( .A1(n28373), .A2(n28928), .A3(n28403), .ZN(n28144) );
  XOR3HSV2 U29755 ( .A1(n28145), .A2(n28144), .A3(n28143), .Z(\pe9/poht [1])
         );
  NOR2HSV2 U29756 ( .A1(n28146), .A2(n28348), .ZN(n28179) );
  CLKNAND2HSV1 U29757 ( .A1(n28317), .A2(\pe9/got [6]), .ZN(n28177) );
  NAND2HSV0 U29758 ( .A1(n19767), .A2(n28643), .ZN(n28175) );
  INHSV2 U29759 ( .I(\pe9/got [3]), .ZN(n28315) );
  INHSV2 U29760 ( .I(n28315), .ZN(n28388) );
  NAND2HSV0 U29761 ( .A1(n28264), .A2(n28388), .ZN(n28171) );
  NAND2HSV0 U29762 ( .A1(\pe9/aot [6]), .A2(\pe9/bq[1] ), .ZN(n28361) );
  OAI21HSV0 U29763 ( .A1(n28361), .A2(n28148), .B(n28147), .ZN(n28150) );
  XOR2HSV0 U29764 ( .A1(n28150), .A2(n28149), .Z(n28165) );
  NAND2HSV0 U29765 ( .A1(\pe9/aot [3]), .A2(\pe9/bq[9] ), .ZN(n28152) );
  NAND2HSV0 U29766 ( .A1(\pe9/aot [2]), .A2(\pe9/bq[10] ), .ZN(n28151) );
  XOR2HSV0 U29767 ( .A1(n28152), .A2(n28151), .Z(n28156) );
  NAND2HSV0 U29768 ( .A1(\pe9/aot [1]), .A2(\pe9/bq[11] ), .ZN(n28154) );
  NAND2HSV0 U29769 ( .A1(\pe9/aot [5]), .A2(\pe9/bq[7] ), .ZN(n28153) );
  XOR2HSV0 U29770 ( .A1(n28154), .A2(n28153), .Z(n28155) );
  XNOR2HSV1 U29771 ( .A1(n28156), .A2(n28155), .ZN(n28164) );
  NAND2HSV0 U29772 ( .A1(\pe9/aot [4]), .A2(\pe9/bq[8] ), .ZN(n28158) );
  NAND2HSV0 U29773 ( .A1(\pe9/aot [7]), .A2(\pe9/bq[5] ), .ZN(n28157) );
  XOR2HSV0 U29774 ( .A1(n28158), .A2(n28157), .Z(n28162) );
  NAND2HSV0 U29775 ( .A1(\pe9/aot [9]), .A2(\pe9/bq[3] ), .ZN(n28160) );
  NAND2HSV0 U29776 ( .A1(\pe9/aot [8]), .A2(\pe9/bq[4] ), .ZN(n28159) );
  XOR2HSV0 U29777 ( .A1(n28160), .A2(n28159), .Z(n28161) );
  XOR2HSV0 U29778 ( .A1(n28162), .A2(n28161), .Z(n28163) );
  XOR3HSV2 U29779 ( .A1(n28165), .A2(n28164), .A3(n28163), .Z(n28169) );
  NAND2HSV0 U29780 ( .A1(n28689), .A2(\pe9/got [2]), .ZN(n28168) );
  NAND2HSV0 U29781 ( .A1(n28166), .A2(n28658), .ZN(n28167) );
  XOR3HSV1 U29782 ( .A1(n28169), .A2(n28168), .A3(n28167), .Z(n28170) );
  XNOR2HSV1 U29783 ( .A1(n28171), .A2(n28170), .ZN(n28173) );
  INHSV2 U29784 ( .I(\pe9/got [4]), .ZN(n28263) );
  OR2HSV1 U29785 ( .A1(n28214), .A2(n28263), .Z(n28172) );
  XNOR2HSV1 U29786 ( .A1(n28173), .A2(n28172), .ZN(n28174) );
  XNOR2HSV1 U29787 ( .A1(n28175), .A2(n28174), .ZN(n28176) );
  XNOR2HSV1 U29788 ( .A1(n28177), .A2(n28176), .ZN(n28178) );
  XOR2HSV0 U29789 ( .A1(n28179), .A2(n28178), .Z(n28181) );
  NAND2HSV0 U29790 ( .A1(n28383), .A2(\pe9/got [8]), .ZN(n28180) );
  NAND2HSV0 U29791 ( .A1(n28475), .A2(n14073), .ZN(n28182) );
  XNOR2HSV1 U29792 ( .A1(n28183), .A2(n28182), .ZN(n28187) );
  INHSV2 U29793 ( .I(n28184), .ZN(n28387) );
  NAND3HSV2 U29794 ( .A1(n28404), .A2(n28227), .A3(n28387), .ZN(n28186) );
  XOR3HSV2 U29795 ( .A1(n28187), .A2(n28186), .A3(n28185), .Z(\pe9/poht [5])
         );
  NOR2HSV1 U29796 ( .A1(n28368), .A2(n28188), .ZN(n28222) );
  CLKNAND2HSV1 U29797 ( .A1(n28317), .A2(n28643), .ZN(n28220) );
  NAND2HSV0 U29798 ( .A1(n28437), .A2(n28389), .ZN(n28218) );
  NAND2HSV0 U29799 ( .A1(n28264), .A2(n28654), .ZN(n28213) );
  NAND2HSV0 U29800 ( .A1(n28189), .A2(n28658), .ZN(n28211) );
  NAND2HSV0 U29801 ( .A1(\pe9/aot [7]), .A2(\pe9/bq[4] ), .ZN(n28190) );
  XOR2HSV0 U29802 ( .A1(n28191), .A2(n28190), .Z(n28209) );
  NAND2HSV0 U29803 ( .A1(\pe9/aot [3]), .A2(\pe9/bq[8] ), .ZN(n28193) );
  NAND2HSV0 U29804 ( .A1(\pe9/aot [10]), .A2(\pe9/bq[1] ), .ZN(n28192) );
  XOR2HSV0 U29805 ( .A1(n28193), .A2(n28192), .Z(n28198) );
  NOR2HSV0 U29806 ( .A1(n28194), .A2(n28240), .ZN(n28196) );
  NAND2HSV0 U29807 ( .A1(\pe9/aot [1]), .A2(\pe9/bq[10] ), .ZN(n28195) );
  XOR2HSV0 U29808 ( .A1(n28196), .A2(n28195), .Z(n28197) );
  XNOR2HSV1 U29809 ( .A1(n28198), .A2(n28197), .ZN(n28208) );
  NOR2HSV0 U29810 ( .A1(n28200), .A2(n28199), .ZN(n28202) );
  NAND2HSV0 U29811 ( .A1(\pe9/aot [6]), .A2(\pe9/bq[5] ), .ZN(n28201) );
  XOR2HSV0 U29812 ( .A1(n28202), .A2(n28201), .Z(n28206) );
  NAND2HSV0 U29813 ( .A1(\pe9/aot [9]), .A2(\pe9/bq[2] ), .ZN(n28204) );
  NAND2HSV0 U29814 ( .A1(\pe9/aot [8]), .A2(\pe9/bq[3] ), .ZN(n28203) );
  XOR2HSV0 U29815 ( .A1(n28204), .A2(n28203), .Z(n28205) );
  XOR2HSV0 U29816 ( .A1(n28206), .A2(n28205), .Z(n28207) );
  XOR3HSV2 U29817 ( .A1(n28209), .A2(n28208), .A3(n28207), .Z(n28210) );
  XOR2HSV0 U29818 ( .A1(n28211), .A2(n28210), .Z(n28212) );
  XNOR2HSV1 U29819 ( .A1(n28213), .A2(n28212), .ZN(n28216) );
  OR2HSV1 U29820 ( .A1(n28214), .A2(n28315), .Z(n28215) );
  XNOR2HSV1 U29821 ( .A1(n28216), .A2(n28215), .ZN(n28217) );
  XNOR2HSV1 U29822 ( .A1(n28218), .A2(n28217), .ZN(n28219) );
  XNOR2HSV1 U29823 ( .A1(n28220), .A2(n28219), .ZN(n28221) );
  XOR2HSV0 U29824 ( .A1(n28222), .A2(n28221), .Z(n28224) );
  CLKNAND2HSV0 U29825 ( .A1(n28383), .A2(\pe9/got [7]), .ZN(n28223) );
  XOR2HSV0 U29826 ( .A1(n28224), .A2(n28223), .Z(n28226) );
  NAND2HSV0 U29827 ( .A1(n28394), .A2(\pe9/got [8]), .ZN(n28225) );
  XNOR2HSV1 U29828 ( .A1(n28226), .A2(n28225), .ZN(n28230) );
  NAND3HSV2 U29829 ( .A1(n28413), .A2(\pe9/got [9]), .A3(n28387), .ZN(n28229)
         );
  XOR3HSV2 U29830 ( .A1(n28230), .A2(n28229), .A3(n28228), .Z(\pe9/poht [6])
         );
  NOR2HSV2 U29831 ( .A1(n28316), .A2(n28263), .ZN(n28254) );
  CLKNAND2HSV0 U29832 ( .A1(n28231), .A2(n28405), .ZN(n28252) );
  NAND2HSV0 U29833 ( .A1(n19767), .A2(n28654), .ZN(n28250) );
  OR2HSV1 U29834 ( .A1(n28287), .A2(n28303), .Z(n28248) );
  NAND2HSV0 U29835 ( .A1(\pe9/aot [7]), .A2(\pe9/bq[2] ), .ZN(n28233) );
  NAND2HSV0 U29836 ( .A1(\pe9/aot [1]), .A2(\pe9/bq[8] ), .ZN(n28232) );
  XOR2HSV0 U29837 ( .A1(n28233), .A2(n28232), .Z(n28237) );
  NAND2HSV0 U29838 ( .A1(\pe9/aot [3]), .A2(\pe9/bq[6] ), .ZN(n28235) );
  NAND2HSV0 U29839 ( .A1(\pe9/aot [5]), .A2(\pe9/bq[4] ), .ZN(n28234) );
  XOR2HSV0 U29840 ( .A1(n28235), .A2(n28234), .Z(n28236) );
  XOR2HSV0 U29841 ( .A1(n28237), .A2(n28236), .Z(n28246) );
  NAND2HSV0 U29842 ( .A1(\pe9/aot [6]), .A2(\pe9/bq[3] ), .ZN(n28239) );
  NAND2HSV0 U29843 ( .A1(\pe9/aot [8]), .A2(\pe9/bq[1] ), .ZN(n28238) );
  XOR2HSV0 U29844 ( .A1(n28239), .A2(n28238), .Z(n28244) );
  NOR2HSV0 U29845 ( .A1(n28398), .A2(n28240), .ZN(n28242) );
  NAND2HSV0 U29846 ( .A1(\pe9/aot [4]), .A2(\pe9/bq[5] ), .ZN(n28241) );
  XOR2HSV0 U29847 ( .A1(n28242), .A2(n28241), .Z(n28243) );
  XOR2HSV0 U29848 ( .A1(n28244), .A2(n28243), .Z(n28245) );
  XOR2HSV0 U29849 ( .A1(n28246), .A2(n28245), .Z(n28247) );
  XNOR2HSV1 U29850 ( .A1(n28248), .A2(n28247), .ZN(n28249) );
  XNOR2HSV1 U29851 ( .A1(n28250), .A2(n28249), .ZN(n28251) );
  XNOR2HSV1 U29852 ( .A1(n28252), .A2(n28251), .ZN(n28253) );
  XOR2HSV0 U29853 ( .A1(n28254), .A2(n28253), .Z(n28256) );
  NAND2HSV0 U29854 ( .A1(n28383), .A2(n28643), .ZN(n28255) );
  CLKNAND2HSV1 U29855 ( .A1(n28475), .A2(\pe9/got [6]), .ZN(n28257) );
  XNOR2HSV1 U29856 ( .A1(n28258), .A2(n28257), .ZN(n28261) );
  NAND3HSV2 U29857 ( .A1(n28413), .A2(\pe9/got [7]), .A3(n28387), .ZN(n28260)
         );
  XOR3HSV2 U29858 ( .A1(n28261), .A2(n28260), .A3(n28259), .Z(\pe9/poht [8])
         );
  NOR2HSV2 U29859 ( .A1(n28316), .A2(n28262), .ZN(n28295) );
  INHSV2 U29860 ( .I(n28263), .ZN(n28369) );
  CLKNAND2HSV1 U29861 ( .A1(n28317), .A2(n28369), .ZN(n28293) );
  NAND2HSV0 U29862 ( .A1(n28437), .A2(n28405), .ZN(n28291) );
  NAND2HSV0 U29863 ( .A1(n28264), .A2(n28658), .ZN(n28285) );
  CLKNHSV0 U29864 ( .I(\pe9/aot [1]), .ZN(n28267) );
  OAI21HSV0 U29865 ( .A1(n28267), .A2(n28266), .B(n28265), .ZN(n28268) );
  OAI21HSV0 U29866 ( .A1(n28270), .A2(n28269), .B(n28268), .ZN(n28271) );
  NAND2HSV0 U29867 ( .A1(\pe9/bq[7] ), .A2(\pe9/aot [3]), .ZN(n28324) );
  XNOR2HSV1 U29868 ( .A1(n28271), .A2(n28324), .ZN(n28275) );
  NAND2HSV0 U29869 ( .A1(\pe9/aot [7]), .A2(\pe9/bq[3] ), .ZN(n28273) );
  NAND2HSV0 U29870 ( .A1(\pe9/aot [2]), .A2(\pe9/bq[8] ), .ZN(n28272) );
  XOR2HSV0 U29871 ( .A1(n28273), .A2(n28272), .Z(n28274) );
  XNOR2HSV1 U29872 ( .A1(n28275), .A2(n28274), .ZN(n28283) );
  NAND2HSV0 U29873 ( .A1(\pe9/aot [6]), .A2(\pe9/bq[4] ), .ZN(n28277) );
  NAND2HSV0 U29874 ( .A1(\pe9/aot [8]), .A2(\pe9/bq[2] ), .ZN(n28276) );
  XOR2HSV0 U29875 ( .A1(n28277), .A2(n28276), .Z(n28281) );
  NAND2HSV0 U29876 ( .A1(\pe9/aot [4]), .A2(\pe9/bq[6] ), .ZN(n28279) );
  NAND2HSV0 U29877 ( .A1(\pe9/aot [5]), .A2(\pe9/bq[5] ), .ZN(n28278) );
  XOR2HSV0 U29878 ( .A1(n28279), .A2(n28278), .Z(n28280) );
  XOR2HSV0 U29879 ( .A1(n28281), .A2(n28280), .Z(n28282) );
  XNOR2HSV1 U29880 ( .A1(n28283), .A2(n28282), .ZN(n28284) );
  XNOR2HSV1 U29881 ( .A1(n28285), .A2(n28284), .ZN(n28289) );
  OR2HSV1 U29882 ( .A1(n28287), .A2(n28286), .Z(n28288) );
  XNOR2HSV1 U29883 ( .A1(n28289), .A2(n28288), .ZN(n28290) );
  XNOR2HSV1 U29884 ( .A1(n28291), .A2(n28290), .ZN(n28292) );
  XNOR2HSV1 U29885 ( .A1(n28293), .A2(n28292), .ZN(n28294) );
  XOR2HSV0 U29886 ( .A1(n28295), .A2(n28294), .Z(n28297) );
  CLKNAND2HSV0 U29887 ( .A1(n28580), .A2(\pe9/got [6]), .ZN(n28296) );
  XOR2HSV0 U29888 ( .A1(n28297), .A2(n28296), .Z(n28299) );
  CLKNAND2HSV0 U29889 ( .A1(n28475), .A2(\pe9/got [7]), .ZN(n28298) );
  XNOR2HSV1 U29890 ( .A1(n28299), .A2(n28298), .ZN(n28302) );
  NAND3HSV2 U29891 ( .A1(n28373), .A2(\pe9/got [8]), .A3(n28403), .ZN(n28301)
         );
  NAND2HSV2 U29892 ( .A1(n28390), .A2(\pe9/got [9]), .ZN(n28300) );
  XOR3HSV2 U29893 ( .A1(n28302), .A2(n28301), .A3(n28300), .Z(\pe9/poht [7])
         );
  NOR2HSV2 U29894 ( .A1(n28368), .A2(n28303), .ZN(n28312) );
  NAND2HSV0 U29895 ( .A1(\pe9/aot [3]), .A2(\pe9/bq[3] ), .ZN(n28305) );
  NAND2HSV0 U29896 ( .A1(\pe9/aot [2]), .A2(\pe9/bq[4] ), .ZN(n28304) );
  XOR2HSV0 U29897 ( .A1(n28305), .A2(n28304), .Z(n28306) );
  NAND2HSV0 U29898 ( .A1(\pe9/aot [1]), .A2(\pe9/bq[5] ), .ZN(n28325) );
  XNOR2HSV1 U29899 ( .A1(n28306), .A2(n28325), .ZN(n28310) );
  NAND2HSV0 U29900 ( .A1(\pe9/aot [5]), .A2(\pe9/bq[1] ), .ZN(n28307) );
  XOR2HSV0 U29901 ( .A1(n28308), .A2(n28307), .Z(n28309) );
  XNOR2HSV1 U29902 ( .A1(n28310), .A2(n28309), .ZN(n28311) );
  XOR2HSV0 U29903 ( .A1(n28312), .A2(n28311), .Z(n28314) );
  NAND2HSV0 U29904 ( .A1(n28383), .A2(n28654), .ZN(n28313) );
  NOR2HSV2 U29905 ( .A1(n28316), .A2(n28315), .ZN(n28335) );
  CLKNAND2HSV0 U29906 ( .A1(n28317), .A2(n28654), .ZN(n28333) );
  NAND2HSV0 U29907 ( .A1(n28437), .A2(n28658), .ZN(n28331) );
  NAND2HSV0 U29908 ( .A1(\pe9/aot [5]), .A2(\pe9/bq[3] ), .ZN(n28319) );
  NAND2HSV0 U29909 ( .A1(\pe9/aot [4]), .A2(\pe9/bq[4] ), .ZN(n28318) );
  XOR2HSV0 U29910 ( .A1(n28319), .A2(n28318), .Z(n28323) );
  NAND2HSV0 U29911 ( .A1(\pe9/aot [7]), .A2(\pe9/bq[1] ), .ZN(n28321) );
  NAND2HSV0 U29912 ( .A1(\pe9/aot [2]), .A2(\pe9/bq[6] ), .ZN(n28320) );
  XOR2HSV0 U29913 ( .A1(n28321), .A2(n28320), .Z(n28322) );
  XOR2HSV0 U29914 ( .A1(n28323), .A2(n28322), .Z(n28329) );
  XOR2HSV0 U29915 ( .A1(n28327), .A2(n28326), .Z(n28328) );
  XNOR2HSV1 U29916 ( .A1(n28329), .A2(n28328), .ZN(n28330) );
  XOR2HSV0 U29917 ( .A1(n28331), .A2(n28330), .Z(n28332) );
  XOR2HSV0 U29918 ( .A1(n28333), .A2(n28332), .Z(n28334) );
  XOR2HSV0 U29919 ( .A1(n28335), .A2(n28334), .Z(n28337) );
  CLKNAND2HSV0 U29920 ( .A1(n28580), .A2(n28389), .ZN(n28336) );
  XOR2HSV0 U29921 ( .A1(n28337), .A2(n28336), .Z(n28339) );
  NAND2HSV0 U29922 ( .A1(n28475), .A2(n28643), .ZN(n28338) );
  XNOR2HSV1 U29923 ( .A1(n28339), .A2(n28338), .ZN(n28355) );
  INHSV2 U29924 ( .I(n28373), .ZN(n28342) );
  NAND2HSV0 U29925 ( .A1(n28340), .A2(\pe9/got [6]), .ZN(n28341) );
  NOR2HSV4 U29926 ( .A1(n28342), .A2(n28341), .ZN(n28354) );
  INAND2HSV2 U29927 ( .A1(n28347), .B1(n28346), .ZN(n28351) );
  CLKNHSV0 U29928 ( .I(\pe9/ti_7t [15]), .ZN(n28349) );
  AOI21HSV0 U29929 ( .A1(n28349), .A2(n18641), .B(n28348), .ZN(n28350) );
  XOR3HSV2 U29930 ( .A1(n28355), .A2(n28354), .A3(n28353), .Z(\pe9/poht [9])
         );
  NAND2HSV2 U29931 ( .A1(\pe9/got [1]), .A2(n28231), .ZN(n28365) );
  NAND2HSV0 U29932 ( .A1(\pe9/aot [3]), .A2(\pe9/bq[4] ), .ZN(n28357) );
  NAND2HSV0 U29933 ( .A1(\pe9/aot [1]), .A2(\pe9/bq[6] ), .ZN(n28356) );
  XOR2HSV0 U29934 ( .A1(n28357), .A2(n28356), .Z(n28362) );
  NAND2HSV0 U29935 ( .A1(\pe9/aot [4]), .A2(\pe9/bq[3] ), .ZN(n28358) );
  XOR2HSV0 U29936 ( .A1(n28359), .A2(n28358), .Z(n28360) );
  XOR4HSV1 U29937 ( .A1(n28363), .A2(n28362), .A3(n28361), .A4(n28360), .Z(
        n28364) );
  XNOR2HSV1 U29938 ( .A1(n28365), .A2(n28364), .ZN(n28367) );
  OAI21HSV1 U29939 ( .A1(n28368), .A2(n28286), .B(n28367), .ZN(n28366) );
  NAND2HSV2 U29940 ( .A1(n28383), .A2(n28388), .ZN(n28371) );
  CLKNAND2HSV1 U29941 ( .A1(n28475), .A2(n28369), .ZN(n28370) );
  XOR3HSV2 U29942 ( .A1(n28372), .A2(n28371), .A3(n28370), .Z(n28376) );
  NAND3HSV2 U29943 ( .A1(n28373), .A2(n28643), .A3(n28412), .ZN(n28375) );
  XOR3HSV2 U29944 ( .A1(n28376), .A2(n28375), .A3(n28374), .Z(\pe9/poht [10])
         );
  NAND2HSV0 U29945 ( .A1(\pe9/aot [4]), .A2(\pe9/bq[1] ), .ZN(n28378) );
  NAND2HSV0 U29946 ( .A1(\pe9/aot [3]), .A2(\pe9/bq[2] ), .ZN(n28377) );
  XOR2HSV0 U29947 ( .A1(n28378), .A2(n28377), .Z(n28382) );
  NAND2HSV0 U29948 ( .A1(\pe9/aot [1]), .A2(\pe9/bq[4] ), .ZN(n28380) );
  NAND2HSV0 U29949 ( .A1(\pe9/aot [2]), .A2(\pe9/bq[3] ), .ZN(n28379) );
  XOR2HSV0 U29950 ( .A1(n28380), .A2(n28379), .Z(n28381) );
  XOR2HSV0 U29951 ( .A1(n28382), .A2(n28381), .Z(n28386) );
  NAND2HSV2 U29952 ( .A1(n28383), .A2(n28658), .ZN(n28385) );
  NAND2HSV0 U29953 ( .A1(n28475), .A2(n28654), .ZN(n28384) );
  XOR3HSV2 U29954 ( .A1(n28386), .A2(n28385), .A3(n28384), .Z(n28393) );
  NAND3HSV2 U29955 ( .A1(n28413), .A2(n28388), .A3(n28387), .ZN(n28392) );
  NAND2HSV2 U29956 ( .A1(n28390), .A2(n28389), .ZN(n28391) );
  XOR3HSV2 U29957 ( .A1(n28393), .A2(n28392), .A3(n28391), .Z(\pe9/poht [12])
         );
  NAND2HSV0 U29958 ( .A1(n28394), .A2(\pe9/got [1]), .ZN(n28402) );
  NAND2HSV0 U29959 ( .A1(\pe9/aot [1]), .A2(\pe9/bq[3] ), .ZN(n28396) );
  NAND2HSV0 U29960 ( .A1(\pe9/aot [3]), .A2(\pe9/bq[1] ), .ZN(n28395) );
  XOR2HSV0 U29961 ( .A1(n28396), .A2(n28395), .Z(n28400) );
  NOR2HSV2 U29962 ( .A1(n28398), .A2(n28397), .ZN(n28399) );
  XNOR2HSV1 U29963 ( .A1(n28400), .A2(n28399), .ZN(n28401) );
  XOR2HSV0 U29964 ( .A1(n28402), .A2(n28401), .Z(n28409) );
  NAND3HSV2 U29965 ( .A1(n28404), .A2(n28654), .A3(n28403), .ZN(n28408) );
  XOR3HSV2 U29966 ( .A1(n28409), .A2(n28408), .A3(n28407), .Z(\pe9/poht [13])
         );
  CLKNAND2HSV1 U29967 ( .A1(\pe9/aot [2]), .A2(\pe9/bq[1] ), .ZN(n28411) );
  NAND2HSV0 U29968 ( .A1(\pe9/aot [1]), .A2(\pe9/bq[2] ), .ZN(n28410) );
  XOR2HSV0 U29969 ( .A1(n28411), .A2(n28410), .Z(n28417) );
  NAND3HSV2 U29970 ( .A1(n28413), .A2(n28658), .A3(n28412), .ZN(n28416) );
  CLKNAND2HSV0 U29971 ( .A1(n28414), .A2(\pe9/got [2]), .ZN(n28415) );
  XOR3HSV2 U29972 ( .A1(n28417), .A2(n28416), .A3(n28415), .Z(\pe9/poht [14])
         );
endmodule

